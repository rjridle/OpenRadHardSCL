* SPICE3 file created from NAND3X1.ext - technology: sky130A

.subckt NAND3X1 Y A B VDD GND
X0 VDD.t11 B.t0 Y.t5 VDD.t10 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X1 Y a_599_989# a_372_210.t0 GND sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=0p ps=0u w=0u l=0u
X2 VDD.t7 a_599_989# Y.t3  DS sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X3 GND A.t1 a_91_103.t0 GND sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=0p ps=0u w=0u l=0u
X4 Y.t1 A.t0 VDD.t3 �DS sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X5 Y.t6 B.t1 VDD.t9  DS sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X6 Y.t4 a_599_989# VDD.t5 �DS sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X7 VDD.t1 A.t2 Y.t0  DS sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
C0 a_599_989# A 0.02fF
C1 VDD A 0.35fF
C2 B Y 0.12fF
C3 Y a_599_989# 0.26fF
C4 B a_599_989# 0.18fF
C5 VDD Y 2.50fF
C6 B VDD 0.30fF
C7 VDD a_599_989# 0.30fF
C8 Y A 0.02fF
C9 B A 0.18fF
R0 B.n0 B.t0 479.223
R1 B.n0 B.t1 375.52
R2 B.n1 B.t2 343.29
R3 B.n1 B.n0 140.752
R4 B.n2 B.n1 4.65
R5 B.n2 B 0.046
R6 Y.n9 Y.n8 280.357
R7 Y.n9 Y.n4 207.058
R8 Y.n3 Y.n2 161.352
R9 Y.n4 Y.n0 95.095
R10 Y.n3 Y.n1 95.095
R11 Y.n4 Y.n3 66.258
R12 Y.n8 Y.n7 30
R13 Y.n6 Y.n5 24.383
R14 Y.n8 Y.n6 23.684
R15 Y.n0 Y.t3 14.282
R16 Y.n0 Y.t4 14.282
R17 Y.n1 Y.t5 14.282
R18 Y.n1 Y.t6 14.282
R19 Y.n2 Y.t0 14.282
R20 Y.n2 Y.t1 14.282
R21 Y.n10 Y.n9 4.65
R22 Y.n10 Y 0.046
R23 VDD.n30 VDD.t7 143.754
R24 VDD.n74 VDD.t3 135.17
R25 VDD.n84 VDD.n83 129.472
R26 VDD.n39 VDD.n38 129.472
R27 VDD.n55 VDD.n54 92.5
R28 VDD.n53 VDD.n52 92.5
R29 VDD.n51 VDD.n50 92.5
R30 VDD.n49 VDD.n48 92.5
R31 VDD.n57 VDD.n56 92.5
R32 VDD.n14 VDD.n1 92.5
R33 VDD.n5 VDD.n4 92.5
R34 VDD.n7 VDD.n6 92.5
R35 VDD.n9 VDD.n8 92.5
R36 VDD.n11 VDD.n10 92.5
R37 VDD.n13 VDD.n12 92.5
R38 VDD.n21 VDD.n20 92.059
R39 VDD.n66 VDD.n65 92.059
R40 VDD.n20 VDD.n16 67.194
R41 VDD.n20 VDD.n17 67.194
R42 VDD.n20 VDD.n18 67.194
R43 VDD.n20 VDD.n19 67.194
R44 VDD.n5 VDD.n3 44.141
R45 VDD.n3 VDD.n2 44.107
R46 VDD.n20 VDD.n15 41.052
R47 VDD.n64 VDD.n62 39.742
R48 VDD.n64 VDD.n63 39.742
R49 VDD.n61 VDD.n60 39.742
R50 VDD.n32  DS 35.8
R51 VDD.n79 �DS 33.243
R52 VDD.n1 VDD.n0 30.923
R53 VDD.n65 VDD.n64 26.38
R54 VDD.n65 VDD.n61 26.38
R55 VDD.n65 VDD.n59 26.38
R56 VDD.n65 VDD.n58 26.38
R57 VDD.n68 VDD.n57 22.915
R58 VDD.n23 VDD.n14 22.915
R59 VDD.n36 �DS 15.343
R60 VDD.n57 VDD.n55 14.864
R61 VDD.n55 VDD.n53 14.864
R62 VDD.n53 VDD.n51 14.864
R63 VDD.n51 VDD.n49 14.864
R64 VDD.n49 VDD.n47 14.864
R65 VDD.n47 VDD.n46 14.864
R66 VDD.n14 VDD.n13 14.864
R67 VDD.n13 VDD.n11 14.864
R68 VDD.n11 VDD.n9 14.864
R69 VDD.n9 VDD.n7 14.864
R70 VDD.n7 VDD.n5 14.864
R71 VDD.n83 VDD.t9 14.282
R72 VDD.n83 VDD.t1 14.282
R73 VDD.n38 VDD.t5 14.282
R74 VDD.n38 VDD.t11 14.282
R75 VDD.n85  DS 12.786
R76 VDD.n23 VDD.n22 8.855
R77 VDD.n22 VDD.n21 8.855
R78 VDD.n26 VDD.n25 8.855
R79 VDD.n25 VDD.n24 8.855
R80 VDD.n30 VDD.n29 8.855
R81 VDD.n29 VDD.n28 8.855
R82 VDD.n34 VDD.n33 8.855
R83 VDD.n33 VDD.n32 8.855
R84 VDD.n40 VDD.n37 8.855
R85 VDD.n37 VDD.n36 8.855
R86 VDD.n44 VDD.n43 8.855
R87 VDD.n43 VDD.n42 8.855
R88 VDD.n91 VDD.n90 8.855
R89 VDD.n90 VDD.n89 8.855
R90 VDD.n87 VDD.n86 8.855
R91 VDD.n86 VDD.n85 8.855
R92 VDD.n81 VDD.n80 8.855
R93 VDD.n80 VDD.n79 8.855
R94 VDD.n77 VDD.n76 8.855
R95 VDD.n76 VDD.n75 8.855
R96 VDD.n72 VDD.n71 8.855
R97 VDD.n71 VDD.n70 8.855
R98 VDD.n68 VDD.n67 8.855
R99 VDD.n67 VDD.n66 8.855
R100 VDD.n89  DS 7.671
R101 VDD.n87 VDD.n84 7.019
R102 VDD.n40 VDD.n39 6.606
R103 VDD.n42 VDD.t10 5.114
R104 VDD.n31 VDD.n30 4.65
R105 VDD.n35 VDD.n34 4.65
R106 VDD.n41 VDD.n40 4.65
R107 VDD.n45 VDD.n44 4.65
R108 VDD.n92 VDD.n91 4.65
R109 VDD.n88 VDD.n87 4.65
R110 VDD.n82 VDD.n81 4.65
R111 VDD.n78 VDD.n77 4.65
R112 VDD.n73 VDD.n72 4.65
R113 VDD.n69 VDD.n68 4.65
R114 VDD.n27 VDD.n23 2.933
R115 VDD.n27 VDD.n26 2.844
R116 VDD.n31 VDD.n27 1.063
R117 VDD.n77 VDD.n74 0.412
R118 VDD.n69 VDD 0.207
R119 VDD.n35 VDD.n31 0.145
R120 VDD.n41 VDD.n35 0.145
R121 VDD.n45 VDD.n41 0.145
R122 VDD.n92 VDD.n88 0.145
R123 VDD.n88 VDD.n82 0.145
R124 VDD.n82 VDD.n78 0.145
R125 VDD.n78 VDD.n73 0.145
R126 VDD.n73 VDD.n69 0.145
R127 VDD VDD.n45 0.098
R128 VDD VDD.n92 0.098
R129 a_372_210.n9 a_372_210.n7 171.558
R130 a_372_210.t0 a_372_210.n9 75.765
R131 a_372_210.n3 a_372_210.n1 74.827
R132 a_372_210.n3 a_372_210.n2 27.476
R133 a_372_210.n7 a_372_210.n6 27.2
R134 a_372_210.n5 a_372_210.n4 23.498
R135 a_372_210.n7 a_372_210.n5 22.4
R136 a_372_210.t0 a_372_210.n11 20.241
R137 a_372_210.t0 a_372_210.n3 13.984
R138 a_372_210.n11 a_372_210.n10 13.494
R139 a_372_210.t0 a_372_210.n0 8.137
R140 a_372_210.n9 a_372_210.n8 1.505
R141 GND.n26 GND.n25 167.358
R142 GND.n25 GND.n23 23.03
R143 GND.n20 GND.n19 9.154
R144 GND.n27 GND.n22 9.154
R145 GND.n30 GND.n29 9.154
R146 GND.n33 GND.n32 9.154
R147 GND.n36 GND.n35 9.154
R148 GND.n14 GND.n13 9.154
R149 GND.n11 GND.n10 9.154
R150 GND.n8 GND.n7 9.154
R151 GND.n5 GND.n4 9.154
R152 GND.n2 GND.n1 9.154
R153 GND.n25 GND.n24 8.128
R154 GND.n18 GND.n17 4.65
R155 GND.n6 GND.n5 4.65
R156 GND.n9 GND.n8 4.65
R157 GND.n12 GND.n11 4.65
R158 GND.n15 GND.n14 4.65
R159 GND.n37 GND.n36 4.65
R160 GND.n34 GND.n33 4.65
R161 GND.n31 GND.n30 4.65
R162 GND.n28 GND.n27 4.65
R163 GND.n21 GND.n20 4.65
R164 GND.n3 GND.n0 3.407
R165 GND.n3 GND.n2 2.844
R166 GND.n6 GND.n3 1.063
R167 GND.n17 GND.n16 0.474
R168 GND.n18 GND 0.207
R169 GND.n27 GND.n26 0.206
R170 GND.n9 GND.n6 0.145
R171 GND.n12 GND.n9 0.145
R172 GND.n15 GND.n12 0.145
R173 GND.n37 GND.n34 0.145
R174 GND.n34 GND.n31 0.145
R175 GND.n31 GND.n28 0.145
R176 GND.n28 GND.n21 0.145
R177 GND.n21 GND.n18 0.145
R178 GND GND.n15 0.098
R179 GND GND.n37 0.098
R180 A.n0 A.t2 512.525
R181 A.n0 A.t0 371.139
R182 A.n1 A.t1 361.392
R183 A.n1 A.n0 235.554
R184 A.n2 A.n1 4.65
R185 A.n2 A 0.046
R186 a_91_103.n5 a_91_103.n4 66.708
R187 a_91_103.n2 a_91_103.n0 25.439
R188 a_91_103.n5 a_91_103.n3 19.496
R189 a_91_103.t0 a_91_103.n5 13.756
R190 a_91_103.n2 a_91_103.n1 2.455
R191 a_91_103.t0 a_91_103.n2 0.246
C10 VDD GND 1.92fF
C11 a_91_103.n0 GND 0.10fF
C12 a_91_103.n1 GND 0.03fF
C13 a_91_103.n2 GND 0.03fF
C14 a_91_103.n3 GND 0.07fF
C15 a_91_103.n4 GND 0.08fF
C16 a_91_103.n5 GND 0.03fF
C17 a_372_210.n0 GND 0.06fF
C18 a_372_210.n1 GND 0.09fF
C19 a_372_210.n2 GND 0.11fF
C20 a_372_210.n3 GND 0.08fF
C21 a_372_210.n4 GND 0.02fF
C22 a_372_210.n5 GND 0.03fF
C23 a_372_210.n6 GND 0.02fF
C24 a_372_210.n7 GND 0.03fF
C25 a_372_210.n8 GND 0.02fF
C26 a_372_210.n9 GND 0.13fF
C27 a_372_210.n10 GND 0.08fF
C28 a_372_210.n11 GND 0.02fF
C29 VDD.n1 GND 0.03fF
C30 VDD.n2 GND 0.14fF
C31 VDD.n3 GND 0.02fF
C32 VDD.n4 GND 0.02fF
C33 VDD.n5 GND 0.05fF
C34 VDD.n6 GND 0.02fF
C35 VDD.n7 GND 0.02fF
C36 VDD.n8 GND 0.02fF
C37 VDD.n9 GND 0.02fF
C38 VDD.n10 GND 0.02fF
C39 VDD.n11 GND 0.02fF
C40 VDD.n12 GND 0.02fF
C41 VDD.n13 GND 0.02fF
C42 VDD.n14 GND 0.03fF
C43 VDD.n15 GND 0.01fF
C44 VDD.n20 GND 0.35fF
C45 VDD.n21 GND 0.21fF
C46 VDD.n22 GND 0.01fF
C47 VDD.n23 GND 0.03fF
C48 VDD.n24 GND 0.21fF
C49 VDD.n25 GND 0.01fF
C50 VDD.n26 GND 0.02fF
C51 VDD.n27 GND 0.01fF
C52 VDD.n28 GND 0.17fF
C53 VDD.n29 GND 0.01fF
C54 VDD.n30 GND 0.05fF
C55 VDD.n31 GND 0.06fF
C56 VDD.n32 GND 0.13fF
C57 VDD.n33 GND 0.01fF
C58 VDD.n34 GND 0.02fF
C59 VDD.n35 GND 0.02fF
C60 VDD.n36 GND 0.12fF
C61 VDD.n37 GND 0.01fF
C62 VDD.n38 GND 0.06fF
C63 VDD.n39 GND 0.04fF
C64 VDD.n40 GND 0.01fF
C65 VDD.n41 GND 0.02fF
C66 VDD.n42 GND 0.11fF
C67 VDD.n43 GND 0.01fF
C68 VDD.n44 GND 0.02fF
C69 VDD.n45 GND 0.01fF
C70 VDD.n46 GND 0.04fF
C71 VDD.n47 GND 0.02fF
C72 VDD.n48 GND 0.02fF
C73 VDD.n49 GND 0.02fF
C74 VDD.n50 GND 0.02fF
C75 VDD.n51 GND 0.02fF
C76 VDD.n52 GND 0.02fF
C77 VDD.n53 GND 0.02fF
C78 VDD.n54 GND 0.02fF
C79 VDD.n55 GND 0.02fF
C80 VDD.n56 GND 0.03fF
C81 VDD.n57 GND 0.03fF
C82 VDD.n60 GND 0.02fF
C83 VDD.n62 GND 0.02fF
C84 VDD.n63 GND 0.14fF
C85 VDD.n65 GND 0.35fF
C86 VDD.n66 GND 0.21fF
C87 VDD.n67 GND 0.01fF
C88 VDD.n68 GND 0.03fF
C89 VDD.n69 GND 0.02fF
C90 VDD.n70 GND 0.21fF
C91 VDD.n71 GND 0.01fF
C92 VDD.n72 GND 0.02fF
C93 VDD.n73 GND 0.02fF
C94 VDD.n74 GND 0.05fF
C95 VDD.n75 GND 0.17fF
C96 VDD.n76 GND 0.01fF
C97 VDD.n77 GND 0.