** sch_path: /home/rjridle/OpenRadHardSCL/lib/xschem/LDO/LDO.sch
**.subckt LDO
V1 Vref GND 1.2
V2 VDD GND 1.68
R1 Vout Vfb 10k m=1
R2 net2 GND 20k m=1
C1 Vout GND 20p m=1
R3 net3 GND 70k m=1
x1 Vfb Vref Vg VDD GND opamp_2stage_V2
.save  v(vref)
.save  v(vout)
Vmeas net1 Vout 0
.save  i(vmeas)
.save  v(vg)
XM1 VDD Vg net1 GND sky130_fd_pr__nfet_01v8 L=0.15 W=7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.save  v(vfb)
Vmeas1 Vout net3 0
.save  i(vmeas1)
Vmeas2 Vfb net2 0
.save  i(vmeas2)
**** begin user architecture code

.lib /home/rjridle/OpenRadHardSCL/sky130A/libs.tech/ngspice/sky130.lib.spice tt


**** end user architecture code
**.ends

* expanding   symbol:  LDO/opamp_2stage_V2.sym # of pins=3
** sym_path: /home/rjridle/OpenRadHardSCL/lib/xschem/LDO/opamp_2stage_V2.sym
** sch_path: /home/rjridle/OpenRadHardSCL/lib/xschem/LDO/opamp_2stage_V2.sch
.subckt opamp_2stage_V2  MINUS PLUS Vout  VDD  GND
*.ipin PLUS
*.ipin MINUS
*.opin Vout
C3 net6 Vout 2p m=1
XM6 net3 net3 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 net5 net3 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 net2 PLUS net1 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM10 net4 MINUS net1 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM11 net1 Vbias VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM13 Vout net5 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM16 net7 Vbias VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.save  v(plus)
.save  v(minus)
.save  v(net2)
.save  v(net4)
.save  v(minus)
.save  v(vout)
.save  v(plus)
Vmeas1 net4 net3 0
.save  i(vmeas1)
Vmeas2 net2 net5 0
.save  i(vmeas2)
Vmeas3 net7 Vout 0
.save  i(vmeas3)
Vmeas5 net2 net8 0
.save  i(vmeas5)
x1 Vbias Vcs VDD GND casc_mirror
XM1 net6 Vcs net8 GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.save  v(net6)
.save  v(vbias)
.save  v(vbias)
.ends


* expanding   symbol:  LDO/casc_mirror.sym # of pins=2
** sym_path: /home/rjridle/OpenRadHardSCL/lib/xschem/LDO/casc_mirror.sym
** sch_path: /home/rjridle/OpenRadHardSCL/lib/xschem/LDO/casc_mirror.sch
.subckt casc_mirror  Vbias Vcs  VDD  GND
*.opin Vbias
*.opin Vcs
XM8 Vbias Vbias net3 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM9 net7 net1 net4 GND sky130_fd_pr__nfet_01v8 L=0.15 W=7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 Vcs Vbias net3 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 net9 net2 net8 GND sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 net2 net2 net6 GND sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 net1 net1 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
R1 net5 GND 1k m=1
Vmeas_ref2 net4 net5 0
.save  i(vmeas_ref2)
Vmeas1 net6 net1 0
.save  i(vmeas1)
Vmeas_ref1 net8 net7 0
.save  i(vmeas_ref1)
.save  v(net7)
.save  v(net5)
.save  v(net1)
Vmeas_ref3 Vbias net9 0
.save  i(vmeas_ref3)
Vmeas_ref4 Vcs net2 0
.save  i(vmeas_ref4)
Vmeas_ref5 VDD net10 0
.save  i(vmeas_ref5)
I0 net10 net3 0.25u
.save  v(vbias)
.save  v(vcs)
.ends

.GLOBAL VDD
.GLOBAL GND
**** begin user architecture code



.control
save all
op
write LDO.raw
*dc V2 1.62 1.98 0.005
*plot v(Vout) v(Vfb) v(Vg) vs v(VDD)
.endc


**** end user architecture code
.end
