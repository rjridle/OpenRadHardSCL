magic
tech sky130A
magscale 1 2
timestamp 1648751716
<< nwell >>
rect -84 832 4968 1575
<< nmos >>
rect 168 316 198 377
tri 198 316 214 332 sw
rect 362 324 392 377
tri 392 324 408 340 sw
rect 168 286 274 316
tri 274 286 304 316 sw
rect 362 294 468 324
tri 468 294 498 324 sw
rect 168 185 198 286
tri 198 270 214 286 nw
tri 258 270 274 286 ne
tri 198 185 214 201 sw
tri 258 185 274 201 se
rect 274 185 304 286
rect 362 193 392 294
tri 392 278 408 294 nw
tri 452 278 468 294 ne
tri 392 193 408 209 sw
tri 452 193 468 209 se
rect 468 193 498 294
tri 168 155 198 185 ne
rect 198 155 274 185
tri 274 155 304 185 nw
tri 362 163 392 193 ne
rect 392 163 468 193
tri 468 163 498 193 nw
rect 813 318 843 379
tri 843 318 859 334 sw
rect 1113 318 1143 379
rect 813 288 919 318
tri 919 288 949 318 sw
rect 813 187 843 288
tri 843 272 859 288 nw
tri 903 272 919 288 ne
tri 843 187 859 203 sw
tri 903 187 919 203 se
rect 919 187 949 288
tri 1008 288 1038 318 se
rect 1038 288 1143 318
rect 1008 194 1038 288
tri 1038 272 1054 288 nw
tri 1097 272 1113 288 ne
tri 1038 194 1054 210 sw
tri 1097 194 1113 210 se
rect 1113 194 1143 288
tri 813 157 843 187 ne
rect 843 157 919 187
tri 919 157 949 187 nw
tri 1008 164 1038 194 ne
rect 1038 164 1113 194
tri 1113 164 1143 194 nw
rect 1315 326 1345 379
tri 1345 326 1361 342 sw
rect 1315 296 1421 326
tri 1421 296 1451 326 sw
rect 1315 195 1345 296
tri 1345 280 1361 296 nw
tri 1405 280 1421 296 ne
tri 1345 195 1361 211 sw
tri 1405 195 1421 211 se
rect 1421 195 1451 296
tri 1315 165 1345 195 ne
rect 1345 165 1421 195
tri 1421 165 1451 195 nw
rect 1775 318 1805 379
tri 1805 318 1821 334 sw
rect 2075 318 2105 379
rect 1775 288 1881 318
tri 1881 288 1911 318 sw
rect 1775 187 1805 288
tri 1805 272 1821 288 nw
tri 1865 272 1881 288 ne
tri 1805 187 1821 203 sw
tri 1865 187 1881 203 se
rect 1881 187 1911 288
tri 1970 288 2000 318 se
rect 2000 288 2105 318
rect 1970 194 2000 288
tri 2000 272 2016 288 nw
tri 2059 272 2075 288 ne
tri 2000 194 2016 210 sw
tri 2059 194 2075 210 se
rect 2075 194 2105 288
tri 1775 157 1805 187 ne
rect 1805 157 1881 187
tri 1881 157 1911 187 nw
tri 1970 164 2000 194 ne
rect 2000 164 2075 194
tri 2075 164 2105 194 nw
rect 2277 326 2307 379
tri 2307 326 2323 342 sw
rect 2277 296 2383 326
tri 2383 296 2413 326 sw
rect 2277 195 2307 296
tri 2307 280 2323 296 nw
tri 2367 280 2383 296 ne
tri 2307 195 2323 211 sw
tri 2367 195 2383 211 se
rect 2383 195 2413 296
tri 2277 165 2307 195 ne
rect 2307 165 2383 195
tri 2383 165 2413 195 nw
rect 2758 316 2788 377
tri 2788 316 2804 332 sw
rect 2952 324 2982 377
tri 2982 324 2998 340 sw
rect 2758 286 2864 316
tri 2864 286 2894 316 sw
rect 2952 294 3058 324
tri 3058 294 3088 324 sw
rect 2758 185 2788 286
tri 2788 270 2804 286 nw
tri 2848 270 2864 286 ne
tri 2788 185 2804 201 sw
tri 2848 185 2864 201 se
rect 2864 185 2894 286
rect 2952 193 2982 294
tri 2982 278 2998 294 nw
tri 3042 278 3058 294 ne
tri 2982 193 2998 209 sw
tri 3042 193 3058 209 se
rect 3058 193 3088 294
tri 2758 155 2788 185 ne
rect 2788 155 2864 185
tri 2864 155 2894 185 nw
tri 2952 163 2982 193 ne
rect 2982 163 3058 193
tri 3058 163 3088 193 nw
rect 3424 316 3454 377
tri 3454 316 3470 332 sw
rect 3618 324 3648 377
tri 3648 324 3664 340 sw
rect 3424 286 3530 316
tri 3530 286 3560 316 sw
rect 3618 294 3724 324
tri 3724 294 3754 324 sw
rect 3424 185 3454 286
tri 3454 270 3470 286 nw
tri 3514 270 3530 286 ne
tri 3454 185 3470 201 sw
tri 3514 185 3530 201 se
rect 3530 185 3560 286
rect 3618 193 3648 294
tri 3648 278 3664 294 nw
tri 3708 278 3724 294 ne
tri 3648 193 3664 209 sw
tri 3708 193 3724 209 se
rect 3724 193 3754 294
tri 3424 155 3454 185 ne
rect 3454 155 3530 185
tri 3530 155 3560 185 nw
tri 3618 163 3648 193 ne
rect 3648 163 3724 193
tri 3724 163 3754 193 nw
rect 4069 318 4099 379
tri 4099 318 4115 334 sw
rect 4369 318 4399 379
rect 4069 288 4175 318
tri 4175 288 4205 318 sw
rect 4069 187 4099 288
tri 4099 272 4115 288 nw
tri 4159 272 4175 288 ne
tri 4099 187 4115 203 sw
tri 4159 187 4175 203 se
rect 4175 187 4205 288
tri 4264 288 4294 318 se
rect 4294 288 4399 318
rect 4264 194 4294 288
tri 4294 272 4310 288 nw
tri 4353 272 4369 288 ne
tri 4294 194 4310 210 sw
tri 4353 194 4369 210 se
rect 4369 194 4399 288
tri 4069 157 4099 187 ne
rect 4099 157 4175 187
tri 4175 157 4205 187 nw
tri 4264 164 4294 194 ne
rect 4294 164 4369 194
tri 4369 164 4399 194 nw
rect 4571 326 4601 379
tri 4601 326 4617 342 sw
rect 4571 296 4677 326
tri 4677 296 4707 326 sw
rect 4571 195 4601 296
tri 4601 280 4617 296 nw
tri 4661 280 4677 296 ne
tri 4601 195 4617 211 sw
tri 4661 195 4677 211 se
rect 4677 195 4707 296
tri 4571 165 4601 195 ne
rect 4601 165 4677 195
tri 4677 165 4707 195 nw
<< pmos >>
rect 187 1050 217 1450
rect 275 1050 305 1450
rect 363 1050 393 1450
rect 451 1050 481 1450
rect 913 1050 943 1450
rect 1001 1050 1031 1450
rect 1089 1050 1119 1450
rect 1177 1050 1207 1450
rect 1265 1050 1295 1450
rect 1353 1050 1383 1450
rect 1875 1050 1905 1450
rect 1963 1050 1993 1450
rect 2051 1050 2081 1450
rect 2139 1050 2169 1450
rect 2227 1050 2257 1450
rect 2315 1050 2345 1450
rect 2777 1050 2807 1450
rect 2865 1050 2895 1450
rect 2953 1050 2983 1450
rect 3041 1050 3071 1450
rect 3443 1050 3473 1450
rect 3531 1050 3561 1450
rect 3619 1050 3649 1450
rect 3707 1050 3737 1450
rect 4169 1050 4199 1450
rect 4257 1050 4287 1450
rect 4345 1050 4375 1450
rect 4433 1050 4463 1450
rect 4521 1050 4551 1450
rect 4609 1050 4639 1450
<< ndiff >>
rect 112 361 168 377
rect 112 327 122 361
rect 156 327 168 361
rect 112 289 168 327
rect 198 361 362 377
rect 198 332 219 361
tri 198 316 214 332 ne
rect 214 327 219 332
rect 253 327 316 361
rect 350 327 362 361
rect 214 316 362 327
rect 392 340 554 377
tri 392 324 408 340 ne
rect 408 324 554 340
rect 112 255 122 289
rect 156 255 168 289
tri 274 286 304 316 ne
rect 304 289 362 316
tri 468 294 498 324 ne
rect 112 221 168 255
rect 112 187 122 221
rect 156 187 168 221
rect 112 155 168 187
tri 198 270 214 286 se
rect 214 270 258 286
tri 258 270 274 286 sw
rect 198 236 274 270
rect 198 202 219 236
rect 253 202 274 236
rect 198 201 274 202
tri 198 185 214 201 ne
rect 214 185 258 201
tri 258 185 274 201 nw
rect 304 255 316 289
rect 350 255 362 289
rect 304 221 362 255
rect 304 187 316 221
rect 350 187 362 221
tri 392 278 408 294 se
rect 408 278 452 294
tri 452 278 468 294 sw
rect 392 245 468 278
rect 392 211 413 245
rect 447 211 468 245
rect 392 209 468 211
tri 392 193 408 209 ne
rect 408 193 452 209
tri 452 193 468 209 nw
rect 498 289 554 324
rect 498 255 510 289
rect 544 255 554 289
rect 498 221 554 255
tri 168 155 198 185 sw
tri 274 155 304 185 se
rect 304 163 362 187
tri 362 163 392 193 sw
tri 468 163 498 193 se
rect 498 187 510 221
rect 544 187 554 221
rect 498 163 554 187
rect 304 155 554 163
rect 112 151 554 155
rect 112 117 122 151
rect 156 117 316 151
rect 350 117 413 151
rect 447 117 510 151
rect 544 117 554 151
rect 112 101 554 117
rect 757 363 813 379
rect 757 329 767 363
rect 801 329 813 363
rect 757 291 813 329
rect 843 363 1113 379
rect 843 334 864 363
tri 843 318 859 334 ne
rect 859 329 864 334
rect 898 329 961 363
rect 995 329 1058 363
rect 1092 329 1113 363
rect 859 318 1113 329
rect 1143 363 1199 379
rect 1143 329 1155 363
rect 1189 329 1199 363
rect 757 257 767 291
rect 801 257 813 291
tri 919 288 949 318 ne
rect 949 291 1008 318
rect 757 223 813 257
rect 757 189 767 223
rect 801 189 813 223
rect 757 157 813 189
tri 843 272 859 288 se
rect 859 272 903 288
tri 903 272 919 288 sw
rect 843 238 919 272
rect 843 204 864 238
rect 898 204 919 238
rect 843 203 919 204
tri 843 187 859 203 ne
rect 859 187 903 203
tri 903 187 919 203 nw
rect 949 257 961 291
rect 995 257 1008 291
tri 1008 288 1038 318 nw
rect 949 223 1008 257
rect 949 189 961 223
rect 995 189 1008 223
tri 1038 272 1054 288 se
rect 1054 272 1097 288
tri 1097 272 1113 288 sw
rect 1038 244 1113 272
rect 1038 210 1059 244
rect 1093 210 1113 244
tri 1038 194 1054 210 ne
rect 1054 194 1097 210
tri 1097 194 1113 210 nw
tri 813 157 843 187 sw
tri 919 157 949 187 se
rect 949 164 1008 189
tri 1008 164 1038 194 sw
tri 1113 164 1143 194 se
rect 1143 164 1199 329
rect 949 157 1199 164
rect 757 153 1199 157
rect 757 119 767 153
rect 801 119 961 153
rect 995 119 1058 153
rect 1092 119 1155 153
rect 1189 119 1199 153
rect 757 103 1199 119
rect 1259 363 1315 379
rect 1259 329 1269 363
rect 1303 329 1315 363
rect 1259 291 1315 329
rect 1345 342 1507 379
tri 1345 326 1361 342 ne
rect 1361 326 1507 342
tri 1421 296 1451 326 ne
rect 1259 257 1269 291
rect 1303 257 1315 291
rect 1259 223 1315 257
rect 1259 189 1269 223
rect 1303 189 1315 223
tri 1345 280 1361 296 se
rect 1361 280 1405 296
tri 1405 280 1421 296 sw
rect 1345 247 1421 280
rect 1345 213 1366 247
rect 1400 213 1421 247
rect 1345 211 1421 213
tri 1345 195 1361 211 ne
rect 1361 195 1405 211
tri 1405 195 1421 211 nw
rect 1451 291 1507 326
rect 1451 257 1463 291
rect 1497 257 1507 291
rect 1451 223 1507 257
rect 1259 165 1315 189
tri 1315 165 1345 195 sw
tri 1421 165 1451 195 se
rect 1451 189 1463 223
rect 1497 189 1507 223
rect 1451 165 1507 189
rect 1259 153 1507 165
rect 1259 119 1269 153
rect 1303 119 1366 153
rect 1400 119 1463 153
rect 1497 119 1507 153
rect 1259 103 1507 119
rect 1719 363 1775 379
rect 1719 329 1729 363
rect 1763 329 1775 363
rect 1719 291 1775 329
rect 1805 363 2075 379
rect 1805 334 1826 363
tri 1805 318 1821 334 ne
rect 1821 329 1826 334
rect 1860 329 1923 363
rect 1957 329 2020 363
rect 2054 329 2075 363
rect 1821 318 2075 329
rect 2105 363 2161 379
rect 2105 329 2117 363
rect 2151 329 2161 363
rect 1719 257 1729 291
rect 1763 257 1775 291
tri 1881 288 1911 318 ne
rect 1911 291 1970 318
rect 1719 223 1775 257
rect 1719 189 1729 223
rect 1763 189 1775 223
rect 1719 157 1775 189
tri 1805 272 1821 288 se
rect 1821 272 1865 288
tri 1865 272 1881 288 sw
rect 1805 238 1881 272
rect 1805 204 1826 238
rect 1860 204 1881 238
rect 1805 203 1881 204
tri 1805 187 1821 203 ne
rect 1821 187 1865 203
tri 1865 187 1881 203 nw
rect 1911 257 1923 291
rect 1957 257 1970 291
tri 1970 288 2000 318 nw
rect 1911 223 1970 257
rect 1911 189 1923 223
rect 1957 189 1970 223
tri 2000 272 2016 288 se
rect 2016 272 2059 288
tri 2059 272 2075 288 sw
rect 2000 244 2075 272
rect 2000 210 2021 244
rect 2055 210 2075 244
tri 2000 194 2016 210 ne
rect 2016 194 2059 210
tri 2059 194 2075 210 nw
tri 1775 157 1805 187 sw
tri 1881 157 1911 187 se
rect 1911 164 1970 189
tri 1970 164 2000 194 sw
tri 2075 164 2105 194 se
rect 2105 164 2161 329
rect 1911 157 2161 164
rect 1719 153 2161 157
rect 1719 119 1729 153
rect 1763 119 1923 153
rect 1957 119 2020 153
rect 2054 119 2117 153
rect 2151 119 2161 153
rect 1719 103 2161 119
rect 2221 363 2277 379
rect 2221 329 2231 363
rect 2265 329 2277 363
rect 2221 291 2277 329
rect 2307 342 2469 379
tri 2307 326 2323 342 ne
rect 2323 326 2469 342
tri 2383 296 2413 326 ne
rect 2221 257 2231 291
rect 2265 257 2277 291
rect 2221 223 2277 257
rect 2221 189 2231 223
rect 2265 189 2277 223
tri 2307 280 2323 296 se
rect 2323 280 2367 296
tri 2367 280 2383 296 sw
rect 2307 247 2383 280
rect 2307 213 2328 247
rect 2362 213 2383 247
rect 2307 211 2383 213
tri 2307 195 2323 211 ne
rect 2323 195 2367 211
tri 2367 195 2383 211 nw
rect 2413 291 2469 326
rect 2413 257 2425 291
rect 2459 257 2469 291
rect 2413 223 2469 257
rect 2221 165 2277 189
tri 2277 165 2307 195 sw
tri 2383 165 2413 195 se
rect 2413 189 2425 223
rect 2459 189 2469 223
rect 2413 165 2469 189
rect 2221 153 2469 165
rect 2221 119 2231 153
rect 2265 119 2328 153
rect 2362 119 2425 153
rect 2459 119 2469 153
rect 2221 103 2469 119
rect 2702 361 2758 377
rect 2702 327 2712 361
rect 2746 327 2758 361
rect 2702 289 2758 327
rect 2788 361 2952 377
rect 2788 332 2809 361
tri 2788 316 2804 332 ne
rect 2804 327 2809 332
rect 2843 327 2906 361
rect 2940 327 2952 361
rect 2804 316 2952 327
rect 2982 340 3144 377
tri 2982 324 2998 340 ne
rect 2998 324 3144 340
rect 2702 255 2712 289
rect 2746 255 2758 289
tri 2864 286 2894 316 ne
rect 2894 289 2952 316
tri 3058 294 3088 324 ne
rect 2702 221 2758 255
rect 2702 187 2712 221
rect 2746 187 2758 221
rect 2702 155 2758 187
tri 2788 270 2804 286 se
rect 2804 270 2848 286
tri 2848 270 2864 286 sw
rect 2788 236 2864 270
rect 2788 202 2809 236
rect 2843 202 2864 236
rect 2788 201 2864 202
tri 2788 185 2804 201 ne
rect 2804 185 2848 201
tri 2848 185 2864 201 nw
rect 2894 255 2906 289
rect 2940 255 2952 289
rect 2894 221 2952 255
rect 2894 187 2906 221
rect 2940 187 2952 221
tri 2982 278 2998 294 se
rect 2998 278 3042 294
tri 3042 278 3058 294 sw
rect 2982 245 3058 278
rect 2982 211 3003 245
rect 3037 211 3058 245
rect 2982 209 3058 211
tri 2982 193 2998 209 ne
rect 2998 193 3042 209
tri 3042 193 3058 209 nw
rect 3088 289 3144 324
rect 3088 255 3100 289
rect 3134 255 3144 289
rect 3088 221 3144 255
tri 2758 155 2788 185 sw
tri 2864 155 2894 185 se
rect 2894 163 2952 187
tri 2952 163 2982 193 sw
tri 3058 163 3088 193 se
rect 3088 187 3100 221
rect 3134 187 3144 221
rect 3088 163 3144 187
rect 2894 155 3144 163
rect 2702 151 3144 155
rect 2702 117 2712 151
rect 2746 117 2906 151
rect 2940 117 3003 151
rect 3037 117 3100 151
rect 3134 117 3144 151
rect 2702 101 3144 117
rect 3368 361 3424 377
rect 3368 327 3378 361
rect 3412 327 3424 361
rect 3368 289 3424 327
rect 3454 361 3618 377
rect 3454 332 3475 361
tri 3454 316 3470 332 ne
rect 3470 327 3475 332
rect 3509 327 3572 361
rect 3606 327 3618 361
rect 3470 316 3618 327
rect 3648 340 3810 377
tri 3648 324 3664 340 ne
rect 3664 324 3810 340
rect 3368 255 3378 289
rect 3412 255 3424 289
tri 3530 286 3560 316 ne
rect 3560 289 3618 316
tri 3724 294 3754 324 ne
rect 3368 221 3424 255
rect 3368 187 3378 221
rect 3412 187 3424 221
rect 3368 155 3424 187
tri 3454 270 3470 286 se
rect 3470 270 3514 286
tri 3514 270 3530 286 sw
rect 3454 236 3530 270
rect 3454 202 3475 236
rect 3509 202 3530 236
rect 3454 201 3530 202
tri 3454 185 3470 201 ne
rect 3470 185 3514 201
tri 3514 185 3530 201 nw
rect 3560 255 3572 289
rect 3606 255 3618 289
rect 3560 221 3618 255
rect 3560 187 3572 221
rect 3606 187 3618 221
tri 3648 278 3664 294 se
rect 3664 278 3708 294
tri 3708 278 3724 294 sw
rect 3648 245 3724 278
rect 3648 211 3669 245
rect 3703 211 3724 245
rect 3648 209 3724 211
tri 3648 193 3664 209 ne
rect 3664 193 3708 209
tri 3708 193 3724 209 nw
rect 3754 289 3810 324
rect 3754 255 3766 289
rect 3800 255 3810 289
rect 3754 221 3810 255
tri 3424 155 3454 185 sw
tri 3530 155 3560 185 se
rect 3560 163 3618 187
tri 3618 163 3648 193 sw
tri 3724 163 3754 193 se
rect 3754 187 3766 221
rect 3800 187 3810 221
rect 3754 163 3810 187
rect 3560 155 3810 163
rect 3368 151 3810 155
rect 3368 117 3378 151
rect 3412 117 3572 151
rect 3606 117 3669 151
rect 3703 117 3766 151
rect 3800 117 3810 151
rect 3368 101 3810 117
rect 4013 363 4069 379
rect 4013 329 4023 363
rect 4057 329 4069 363
rect 4013 291 4069 329
rect 4099 363 4369 379
rect 4099 334 4120 363
tri 4099 318 4115 334 ne
rect 4115 329 4120 334
rect 4154 329 4217 363
rect 4251 329 4314 363
rect 4348 329 4369 363
rect 4115 318 4369 329
rect 4399 363 4455 379
rect 4399 329 4411 363
rect 4445 329 4455 363
rect 4013 257 4023 291
rect 4057 257 4069 291
tri 4175 288 4205 318 ne
rect 4205 291 4264 318
rect 4013 223 4069 257
rect 4013 189 4023 223
rect 4057 189 4069 223
rect 4013 157 4069 189
tri 4099 272 4115 288 se
rect 4115 272 4159 288
tri 4159 272 4175 288 sw
rect 4099 238 4175 272
rect 4099 204 4120 238
rect 4154 204 4175 238
rect 4099 203 4175 204
tri 4099 187 4115 203 ne
rect 4115 187 4159 203
tri 4159 187 4175 203 nw
rect 4205 257 4217 291
rect 4251 257 4264 291
tri 4264 288 4294 318 nw
rect 4205 223 4264 257
rect 4205 189 4217 223
rect 4251 189 4264 223
tri 4294 272 4310 288 se
rect 4310 272 4353 288
tri 4353 272 4369 288 sw
rect 4294 244 4369 272
rect 4294 210 4315 244
rect 4349 210 4369 244
tri 4294 194 4310 210 ne
rect 4310 194 4353 210
tri 4353 194 4369 210 nw
tri 4069 157 4099 187 sw
tri 4175 157 4205 187 se
rect 4205 164 4264 189
tri 4264 164 4294 194 sw
tri 4369 164 4399 194 se
rect 4399 164 4455 329
rect 4205 157 4455 164
rect 4013 153 4455 157
rect 4013 119 4023 153
rect 4057 119 4217 153
rect 4251 119 4314 153
rect 4348 119 4411 153
rect 4445 119 4455 153
rect 4013 103 4455 119
rect 4515 363 4571 379
rect 4515 329 4525 363
rect 4559 329 4571 363
rect 4515 291 4571 329
rect 4601 342 4763 379
tri 4601 326 4617 342 ne
rect 4617 326 4763 342
tri 4677 296 4707 326 ne
rect 4515 257 4525 291
rect 4559 257 4571 291
rect 4515 223 4571 257
rect 4515 189 4525 223
rect 4559 189 4571 223
tri 4601 280 4617 296 se
rect 4617 280 4661 296
tri 4661 280 4677 296 sw
rect 4601 247 4677 280
rect 4601 213 4622 247
rect 4656 213 4677 247
rect 4601 211 4677 213
tri 4601 195 4617 211 ne
rect 4617 195 4661 211
tri 4661 195 4677 211 nw
rect 4707 291 4763 326
rect 4707 257 4719 291
rect 4753 257 4763 291
rect 4707 223 4763 257
rect 4515 165 4571 189
tri 4571 165 4601 195 sw
tri 4677 165 4707 195 se
rect 4707 189 4719 223
rect 4753 189 4763 223
rect 4707 165 4763 189
rect 4515 153 4763 165
rect 4515 119 4525 153
rect 4559 119 4622 153
rect 4656 119 4719 153
rect 4753 119 4763 153
rect 4515 103 4763 119
<< pdiff >>
rect 131 1412 187 1450
rect 131 1378 141 1412
rect 175 1378 187 1412
rect 131 1344 187 1378
rect 131 1310 141 1344
rect 175 1310 187 1344
rect 131 1276 187 1310
rect 131 1242 141 1276
rect 175 1242 187 1276
rect 131 1208 187 1242
rect 131 1174 141 1208
rect 175 1174 187 1208
rect 131 1139 187 1174
rect 131 1105 141 1139
rect 175 1105 187 1139
rect 131 1050 187 1105
rect 217 1412 275 1450
rect 217 1378 229 1412
rect 263 1378 275 1412
rect 217 1344 275 1378
rect 217 1310 229 1344
rect 263 1310 275 1344
rect 217 1276 275 1310
rect 217 1242 229 1276
rect 263 1242 275 1276
rect 217 1208 275 1242
rect 217 1174 229 1208
rect 263 1174 275 1208
rect 217 1139 275 1174
rect 217 1105 229 1139
rect 263 1105 275 1139
rect 217 1050 275 1105
rect 305 1412 363 1450
rect 305 1378 317 1412
rect 351 1378 363 1412
rect 305 1344 363 1378
rect 305 1310 317 1344
rect 351 1310 363 1344
rect 305 1276 363 1310
rect 305 1242 317 1276
rect 351 1242 363 1276
rect 305 1208 363 1242
rect 305 1174 317 1208
rect 351 1174 363 1208
rect 305 1050 363 1174
rect 393 1412 451 1450
rect 393 1378 405 1412
rect 439 1378 451 1412
rect 393 1344 451 1378
rect 393 1310 405 1344
rect 439 1310 451 1344
rect 393 1276 451 1310
rect 393 1242 405 1276
rect 439 1242 451 1276
rect 393 1208 451 1242
rect 393 1174 405 1208
rect 439 1174 451 1208
rect 393 1139 451 1174
rect 393 1105 405 1139
rect 439 1105 451 1139
rect 393 1050 451 1105
rect 481 1412 535 1450
rect 481 1378 493 1412
rect 527 1378 535 1412
rect 481 1344 535 1378
rect 481 1310 493 1344
rect 527 1310 535 1344
rect 481 1276 535 1310
rect 481 1242 493 1276
rect 527 1242 535 1276
rect 481 1208 535 1242
rect 481 1174 493 1208
rect 527 1174 535 1208
rect 481 1050 535 1174
rect 857 1412 913 1450
rect 857 1378 867 1412
rect 901 1378 913 1412
rect 857 1344 913 1378
rect 857 1310 867 1344
rect 901 1310 913 1344
rect 857 1276 913 1310
rect 857 1242 867 1276
rect 901 1242 913 1276
rect 857 1208 913 1242
rect 857 1174 867 1208
rect 901 1174 913 1208
rect 857 1139 913 1174
rect 857 1105 867 1139
rect 901 1105 913 1139
rect 857 1050 913 1105
rect 943 1412 1001 1450
rect 943 1378 955 1412
rect 989 1378 1001 1412
rect 943 1344 1001 1378
rect 943 1310 955 1344
rect 989 1310 1001 1344
rect 943 1276 1001 1310
rect 943 1242 955 1276
rect 989 1242 1001 1276
rect 943 1208 1001 1242
rect 943 1174 955 1208
rect 989 1174 1001 1208
rect 943 1139 1001 1174
rect 943 1105 955 1139
rect 989 1105 1001 1139
rect 943 1050 1001 1105
rect 1031 1412 1089 1450
rect 1031 1378 1043 1412
rect 1077 1378 1089 1412
rect 1031 1344 1089 1378
rect 1031 1310 1043 1344
rect 1077 1310 1089 1344
rect 1031 1276 1089 1310
rect 1031 1242 1043 1276
rect 1077 1242 1089 1276
rect 1031 1208 1089 1242
rect 1031 1174 1043 1208
rect 1077 1174 1089 1208
rect 1031 1050 1089 1174
rect 1119 1412 1177 1450
rect 1119 1378 1131 1412
rect 1165 1378 1177 1412
rect 1119 1344 1177 1378
rect 1119 1310 1131 1344
rect 1165 1310 1177 1344
rect 1119 1276 1177 1310
rect 1119 1242 1131 1276
rect 1165 1242 1177 1276
rect 1119 1208 1177 1242
rect 1119 1174 1131 1208
rect 1165 1174 1177 1208
rect 1119 1139 1177 1174
rect 1119 1105 1131 1139
rect 1165 1105 1177 1139
rect 1119 1050 1177 1105
rect 1207 1412 1265 1450
rect 1207 1378 1219 1412
rect 1253 1378 1265 1412
rect 1207 1344 1265 1378
rect 1207 1310 1219 1344
rect 1253 1310 1265 1344
rect 1207 1276 1265 1310
rect 1207 1242 1219 1276
rect 1253 1242 1265 1276
rect 1207 1208 1265 1242
rect 1207 1174 1219 1208
rect 1253 1174 1265 1208
rect 1207 1050 1265 1174
rect 1295 1412 1353 1450
rect 1295 1378 1307 1412
rect 1341 1378 1353 1412
rect 1295 1344 1353 1378
rect 1295 1310 1307 1344
rect 1341 1310 1353 1344
rect 1295 1276 1353 1310
rect 1295 1242 1307 1276
rect 1341 1242 1353 1276
rect 1295 1208 1353 1242
rect 1295 1174 1307 1208
rect 1341 1174 1353 1208
rect 1295 1139 1353 1174
rect 1295 1105 1307 1139
rect 1341 1105 1353 1139
rect 1295 1050 1353 1105
rect 1383 1412 1437 1450
rect 1383 1378 1395 1412
rect 1429 1378 1437 1412
rect 1383 1344 1437 1378
rect 1383 1310 1395 1344
rect 1429 1310 1437 1344
rect 1383 1276 1437 1310
rect 1383 1242 1395 1276
rect 1429 1242 1437 1276
rect 1383 1208 1437 1242
rect 1383 1174 1395 1208
rect 1429 1174 1437 1208
rect 1383 1050 1437 1174
rect 1819 1412 1875 1450
rect 1819 1378 1829 1412
rect 1863 1378 1875 1412
rect 1819 1344 1875 1378
rect 1819 1310 1829 1344
rect 1863 1310 1875 1344
rect 1819 1276 1875 1310
rect 1819 1242 1829 1276
rect 1863 1242 1875 1276
rect 1819 1208 1875 1242
rect 1819 1174 1829 1208
rect 1863 1174 1875 1208
rect 1819 1139 1875 1174
rect 1819 1105 1829 1139
rect 1863 1105 1875 1139
rect 1819 1050 1875 1105
rect 1905 1412 1963 1450
rect 1905 1378 1917 1412
rect 1951 1378 1963 1412
rect 1905 1344 1963 1378
rect 1905 1310 1917 1344
rect 1951 1310 1963 1344
rect 1905 1276 1963 1310
rect 1905 1242 1917 1276
rect 1951 1242 1963 1276
rect 1905 1208 1963 1242
rect 1905 1174 1917 1208
rect 1951 1174 1963 1208
rect 1905 1139 1963 1174
rect 1905 1105 1917 1139
rect 1951 1105 1963 1139
rect 1905 1050 1963 1105
rect 1993 1412 2051 1450
rect 1993 1378 2005 1412
rect 2039 1378 2051 1412
rect 1993 1344 2051 1378
rect 1993 1310 2005 1344
rect 2039 1310 2051 1344
rect 1993 1276 2051 1310
rect 1993 1242 2005 1276
rect 2039 1242 2051 1276
rect 1993 1208 2051 1242
rect 1993 1174 2005 1208
rect 2039 1174 2051 1208
rect 1993 1050 2051 1174
rect 2081 1412 2139 1450
rect 2081 1378 2093 1412
rect 2127 1378 2139 1412
rect 2081 1344 2139 1378
rect 2081 1310 2093 1344
rect 2127 1310 2139 1344
rect 2081 1276 2139 1310
rect 2081 1242 2093 1276
rect 2127 1242 2139 1276
rect 2081 1208 2139 1242
rect 2081 1174 2093 1208
rect 2127 1174 2139 1208
rect 2081 1139 2139 1174
rect 2081 1105 2093 1139
rect 2127 1105 2139 1139
rect 2081 1050 2139 1105
rect 2169 1412 2227 1450
rect 2169 1378 2181 1412
rect 2215 1378 2227 1412
rect 2169 1344 2227 1378
rect 2169 1310 2181 1344
rect 2215 1310 2227 1344
rect 2169 1276 2227 1310
rect 2169 1242 2181 1276
rect 2215 1242 2227 1276
rect 2169 1208 2227 1242
rect 2169 1174 2181 1208
rect 2215 1174 2227 1208
rect 2169 1050 2227 1174
rect 2257 1412 2315 1450
rect 2257 1378 2269 1412
rect 2303 1378 2315 1412
rect 2257 1344 2315 1378
rect 2257 1310 2269 1344
rect 2303 1310 2315 1344
rect 2257 1276 2315 1310
rect 2257 1242 2269 1276
rect 2303 1242 2315 1276
rect 2257 1208 2315 1242
rect 2257 1174 2269 1208
rect 2303 1174 2315 1208
rect 2257 1139 2315 1174
rect 2257 1105 2269 1139
rect 2303 1105 2315 1139
rect 2257 1050 2315 1105
rect 2345 1412 2399 1450
rect 2345 1378 2357 1412
rect 2391 1378 2399 1412
rect 2345 1344 2399 1378
rect 2345 1310 2357 1344
rect 2391 1310 2399 1344
rect 2345 1276 2399 1310
rect 2345 1242 2357 1276
rect 2391 1242 2399 1276
rect 2345 1208 2399 1242
rect 2345 1174 2357 1208
rect 2391 1174 2399 1208
rect 2345 1050 2399 1174
rect 2721 1412 2777 1450
rect 2721 1378 2731 1412
rect 2765 1378 2777 1412
rect 2721 1344 2777 1378
rect 2721 1310 2731 1344
rect 2765 1310 2777 1344
rect 2721 1276 2777 1310
rect 2721 1242 2731 1276
rect 2765 1242 2777 1276
rect 2721 1208 2777 1242
rect 2721 1174 2731 1208
rect 2765 1174 2777 1208
rect 2721 1139 2777 1174
rect 2721 1105 2731 1139
rect 2765 1105 2777 1139
rect 2721 1050 2777 1105
rect 2807 1412 2865 1450
rect 2807 1378 2819 1412
rect 2853 1378 2865 1412
rect 2807 1344 2865 1378
rect 2807 1310 2819 1344
rect 2853 1310 2865 1344
rect 2807 1276 2865 1310
rect 2807 1242 2819 1276
rect 2853 1242 2865 1276
rect 2807 1208 2865 1242
rect 2807 1174 2819 1208
rect 2853 1174 2865 1208
rect 2807 1139 2865 1174
rect 2807 1105 2819 1139
rect 2853 1105 2865 1139
rect 2807 1050 2865 1105
rect 2895 1412 2953 1450
rect 2895 1378 2907 1412
rect 2941 1378 2953 1412
rect 2895 1344 2953 1378
rect 2895 1310 2907 1344
rect 2941 1310 2953 1344
rect 2895 1276 2953 1310
rect 2895 1242 2907 1276
rect 2941 1242 2953 1276
rect 2895 1208 2953 1242
rect 2895 1174 2907 1208
rect 2941 1174 2953 1208
rect 2895 1050 2953 1174
rect 2983 1412 3041 1450
rect 2983 1378 2995 1412
rect 3029 1378 3041 1412
rect 2983 1344 3041 1378
rect 2983 1310 2995 1344
rect 3029 1310 3041 1344
rect 2983 1276 3041 1310
rect 2983 1242 2995 1276
rect 3029 1242 3041 1276
rect 2983 1208 3041 1242
rect 2983 1174 2995 1208
rect 3029 1174 3041 1208
rect 2983 1139 3041 1174
rect 2983 1105 2995 1139
rect 3029 1105 3041 1139
rect 2983 1050 3041 1105
rect 3071 1412 3125 1450
rect 3071 1378 3083 1412
rect 3117 1378 3125 1412
rect 3071 1344 3125 1378
rect 3071 1310 3083 1344
rect 3117 1310 3125 1344
rect 3071 1276 3125 1310
rect 3071 1242 3083 1276
rect 3117 1242 3125 1276
rect 3071 1208 3125 1242
rect 3071 1174 3083 1208
rect 3117 1174 3125 1208
rect 3071 1050 3125 1174
rect 3387 1412 3443 1450
rect 3387 1378 3397 1412
rect 3431 1378 3443 1412
rect 3387 1344 3443 1378
rect 3387 1310 3397 1344
rect 3431 1310 3443 1344
rect 3387 1276 3443 1310
rect 3387 1242 3397 1276
rect 3431 1242 3443 1276
rect 3387 1208 3443 1242
rect 3387 1174 3397 1208
rect 3431 1174 3443 1208
rect 3387 1139 3443 1174
rect 3387 1105 3397 1139
rect 3431 1105 3443 1139
rect 3387 1050 3443 1105
rect 3473 1412 3531 1450
rect 3473 1378 3485 1412
rect 3519 1378 3531 1412
rect 3473 1344 3531 1378
rect 3473 1310 3485 1344
rect 3519 1310 3531 1344
rect 3473 1276 3531 1310
rect 3473 1242 3485 1276
rect 3519 1242 3531 1276
rect 3473 1208 3531 1242
rect 3473 1174 3485 1208
rect 3519 1174 3531 1208
rect 3473 1139 3531 1174
rect 3473 1105 3485 1139
rect 3519 1105 3531 1139
rect 3473 1050 3531 1105
rect 3561 1412 3619 1450
rect 3561 1378 3573 1412
rect 3607 1378 3619 1412
rect 3561 1344 3619 1378
rect 3561 1310 3573 1344
rect 3607 1310 3619 1344
rect 3561 1276 3619 1310
rect 3561 1242 3573 1276
rect 3607 1242 3619 1276
rect 3561 1208 3619 1242
rect 3561 1174 3573 1208
rect 3607 1174 3619 1208
rect 3561 1050 3619 1174
rect 3649 1412 3707 1450
rect 3649 1378 3661 1412
rect 3695 1378 3707 1412
rect 3649 1344 3707 1378
rect 3649 1310 3661 1344
rect 3695 1310 3707 1344
rect 3649 1276 3707 1310
rect 3649 1242 3661 1276
rect 3695 1242 3707 1276
rect 3649 1208 3707 1242
rect 3649 1174 3661 1208
rect 3695 1174 3707 1208
rect 3649 1139 3707 1174
rect 3649 1105 3661 1139
rect 3695 1105 3707 1139
rect 3649 1050 3707 1105
rect 3737 1412 3791 1450
rect 3737 1378 3749 1412
rect 3783 1378 3791 1412
rect 3737 1344 3791 1378
rect 3737 1310 3749 1344
rect 3783 1310 3791 1344
rect 3737 1276 3791 1310
rect 3737 1242 3749 1276
rect 3783 1242 3791 1276
rect 3737 1208 3791 1242
rect 3737 1174 3749 1208
rect 3783 1174 3791 1208
rect 3737 1050 3791 1174
rect 4113 1412 4169 1450
rect 4113 1378 4123 1412
rect 4157 1378 4169 1412
rect 4113 1344 4169 1378
rect 4113 1310 4123 1344
rect 4157 1310 4169 1344
rect 4113 1276 4169 1310
rect 4113 1242 4123 1276
rect 4157 1242 4169 1276
rect 4113 1208 4169 1242
rect 4113 1174 4123 1208
rect 4157 1174 4169 1208
rect 4113 1139 4169 1174
rect 4113 1105 4123 1139
rect 4157 1105 4169 1139
rect 4113 1050 4169 1105
rect 4199 1412 4257 1450
rect 4199 1378 4211 1412
rect 4245 1378 4257 1412
rect 4199 1344 4257 1378
rect 4199 1310 4211 1344
rect 4245 1310 4257 1344
rect 4199 1276 4257 1310
rect 4199 1242 4211 1276
rect 4245 1242 4257 1276
rect 4199 1208 4257 1242
rect 4199 1174 4211 1208
rect 4245 1174 4257 1208
rect 4199 1139 4257 1174
rect 4199 1105 4211 1139
rect 4245 1105 4257 1139
rect 4199 1050 4257 1105
rect 4287 1412 4345 1450
rect 4287 1378 4299 1412
rect 4333 1378 4345 1412
rect 4287 1344 4345 1378
rect 4287 1310 4299 1344
rect 4333 1310 4345 1344
rect 4287 1276 4345 1310
rect 4287 1242 4299 1276
rect 4333 1242 4345 1276
rect 4287 1208 4345 1242
rect 4287 1174 4299 1208
rect 4333 1174 4345 1208
rect 4287 1050 4345 1174
rect 4375 1412 4433 1450
rect 4375 1378 4387 1412
rect 4421 1378 4433 1412
rect 4375 1344 4433 1378
rect 4375 1310 4387 1344
rect 4421 1310 4433 1344
rect 4375 1276 4433 1310
rect 4375 1242 4387 1276
rect 4421 1242 4433 1276
rect 4375 1208 4433 1242
rect 4375 1174 4387 1208
rect 4421 1174 4433 1208
rect 4375 1139 4433 1174
rect 4375 1105 4387 1139
rect 4421 1105 4433 1139
rect 4375 1050 4433 1105
rect 4463 1412 4521 1450
rect 4463 1378 4475 1412
rect 4509 1378 4521 1412
rect 4463 1344 4521 1378
rect 4463 1310 4475 1344
rect 4509 1310 4521 1344
rect 4463 1276 4521 1310
rect 4463 1242 4475 1276
rect 4509 1242 4521 1276
rect 4463 1208 4521 1242
rect 4463 1174 4475 1208
rect 4509 1174 4521 1208
rect 4463 1050 4521 1174
rect 4551 1412 4609 1450
rect 4551 1378 4563 1412
rect 4597 1378 4609 1412
rect 4551 1344 4609 1378
rect 4551 1310 4563 1344
rect 4597 1310 4609 1344
rect 4551 1276 4609 1310
rect 4551 1242 4563 1276
rect 4597 1242 4609 1276
rect 4551 1208 4609 1242
rect 4551 1174 4563 1208
rect 4597 1174 4609 1208
rect 4551 1139 4609 1174
rect 4551 1105 4563 1139
rect 4597 1105 4609 1139
rect 4551 1050 4609 1105
rect 4639 1412 4693 1450
rect 4639 1378 4651 1412
rect 4685 1378 4693 1412
rect 4639 1344 4693 1378
rect 4639 1310 4651 1344
rect 4685 1310 4693 1344
rect 4639 1276 4693 1310
rect 4639 1242 4651 1276
rect 4685 1242 4693 1276
rect 4639 1208 4693 1242
rect 4639 1174 4651 1208
rect 4685 1174 4693 1208
rect 4639 1050 4693 1174
<< ndiffc >>
rect 122 327 156 361
rect 219 327 253 361
rect 316 327 350 361
rect 122 255 156 289
rect 122 187 156 221
rect 219 202 253 236
rect 316 255 350 289
rect 316 187 350 221
rect 413 211 447 245
rect 510 255 544 289
rect 510 187 544 221
rect 122 117 156 151
rect 316 117 350 151
rect 413 117 447 151
rect 510 117 544 151
rect 767 329 801 363
rect 864 329 898 363
rect 961 329 995 363
rect 1058 329 1092 363
rect 1155 329 1189 363
rect 767 257 801 291
rect 767 189 801 223
rect 864 204 898 238
rect 961 257 995 291
rect 961 189 995 223
rect 1059 210 1093 244
rect 767 119 801 153
rect 961 119 995 153
rect 1058 119 1092 153
rect 1155 119 1189 153
rect 1269 329 1303 363
rect 1269 257 1303 291
rect 1269 189 1303 223
rect 1366 213 1400 247
rect 1463 257 1497 291
rect 1463 189 1497 223
rect 1269 119 1303 153
rect 1366 119 1400 153
rect 1463 119 1497 153
rect 1729 329 1763 363
rect 1826 329 1860 363
rect 1923 329 1957 363
rect 2020 329 2054 363
rect 2117 329 2151 363
rect 1729 257 1763 291
rect 1729 189 1763 223
rect 1826 204 1860 238
rect 1923 257 1957 291
rect 1923 189 1957 223
rect 2021 210 2055 244
rect 1729 119 1763 153
rect 1923 119 1957 153
rect 2020 119 2054 153
rect 2117 119 2151 153
rect 2231 329 2265 363
rect 2231 257 2265 291
rect 2231 189 2265 223
rect 2328 213 2362 247
rect 2425 257 2459 291
rect 2425 189 2459 223
rect 2231 119 2265 153
rect 2328 119 2362 153
rect 2425 119 2459 153
rect 2712 327 2746 361
rect 2809 327 2843 361
rect 2906 327 2940 361
rect 2712 255 2746 289
rect 2712 187 2746 221
rect 2809 202 2843 236
rect 2906 255 2940 289
rect 2906 187 2940 221
rect 3003 211 3037 245
rect 3100 255 3134 289
rect 3100 187 3134 221
rect 2712 117 2746 151
rect 2906 117 2940 151
rect 3003 117 3037 151
rect 3100 117 3134 151
rect 3378 327 3412 361
rect 3475 327 3509 361
rect 3572 327 3606 361
rect 3378 255 3412 289
rect 3378 187 3412 221
rect 3475 202 3509 236
rect 3572 255 3606 289
rect 3572 187 3606 221
rect 3669 211 3703 245
rect 3766 255 3800 289
rect 3766 187 3800 221
rect 3378 117 3412 151
rect 3572 117 3606 151
rect 3669 117 3703 151
rect 3766 117 3800 151
rect 4023 329 4057 363
rect 4120 329 4154 363
rect 4217 329 4251 363
rect 4314 329 4348 363
rect 4411 329 4445 363
rect 4023 257 4057 291
rect 4023 189 4057 223
rect 4120 204 4154 238
rect 4217 257 4251 291
rect 4217 189 4251 223
rect 4315 210 4349 244
rect 4023 119 4057 153
rect 4217 119 4251 153
rect 4314 119 4348 153
rect 4411 119 4445 153
rect 4525 329 4559 363
rect 4525 257 4559 291
rect 4525 189 4559 223
rect 4622 213 4656 247
rect 4719 257 4753 291
rect 4719 189 4753 223
rect 4525 119 4559 153
rect 4622 119 4656 153
rect 4719 119 4753 153
<< pdiffc >>
rect 141 1378 175 1412
rect 141 1310 175 1344
rect 141 1242 175 1276
rect 141 1174 175 1208
rect 141 1105 175 1139
rect 229 1378 263 1412
rect 229 1310 263 1344
rect 229 1242 263 1276
rect 229 1174 263 1208
rect 229 1105 263 1139
rect 317 1378 351 1412
rect 317 1310 351 1344
rect 317 1242 351 1276
rect 317 1174 351 1208
rect 405 1378 439 1412
rect 405 1310 439 1344
rect 405 1242 439 1276
rect 405 1174 439 1208
rect 405 1105 439 1139
rect 493 1378 527 1412
rect 493 1310 527 1344
rect 493 1242 527 1276
rect 493 1174 527 1208
rect 867 1378 901 1412
rect 867 1310 901 1344
rect 867 1242 901 1276
rect 867 1174 901 1208
rect 867 1105 901 1139
rect 955 1378 989 1412
rect 955 1310 989 1344
rect 955 1242 989 1276
rect 955 1174 989 1208
rect 955 1105 989 1139
rect 1043 1378 1077 1412
rect 1043 1310 1077 1344
rect 1043 1242 1077 1276
rect 1043 1174 1077 1208
rect 1131 1378 1165 1412
rect 1131 1310 1165 1344
rect 1131 1242 1165 1276
rect 1131 1174 1165 1208
rect 1131 1105 1165 1139
rect 1219 1378 1253 1412
rect 1219 1310 1253 1344
rect 1219 1242 1253 1276
rect 1219 1174 1253 1208
rect 1307 1378 1341 1412
rect 1307 1310 1341 1344
rect 1307 1242 1341 1276
rect 1307 1174 1341 1208
rect 1307 1105 1341 1139
rect 1395 1378 1429 1412
rect 1395 1310 1429 1344
rect 1395 1242 1429 1276
rect 1395 1174 1429 1208
rect 1829 1378 1863 1412
rect 1829 1310 1863 1344
rect 1829 1242 1863 1276
rect 1829 1174 1863 1208
rect 1829 1105 1863 1139
rect 1917 1378 1951 1412
rect 1917 1310 1951 1344
rect 1917 1242 1951 1276
rect 1917 1174 1951 1208
rect 1917 1105 1951 1139
rect 2005 1378 2039 1412
rect 2005 1310 2039 1344
rect 2005 1242 2039 1276
rect 2005 1174 2039 1208
rect 2093 1378 2127 1412
rect 2093 1310 2127 1344
rect 2093 1242 2127 1276
rect 2093 1174 2127 1208
rect 2093 1105 2127 1139
rect 2181 1378 2215 1412
rect 2181 1310 2215 1344
rect 2181 1242 2215 1276
rect 2181 1174 2215 1208
rect 2269 1378 2303 1412
rect 2269 1310 2303 1344
rect 2269 1242 2303 1276
rect 2269 1174 2303 1208
rect 2269 1105 2303 1139
rect 2357 1378 2391 1412
rect 2357 1310 2391 1344
rect 2357 1242 2391 1276
rect 2357 1174 2391 1208
rect 2731 1378 2765 1412
rect 2731 1310 2765 1344
rect 2731 1242 2765 1276
rect 2731 1174 2765 1208
rect 2731 1105 2765 1139
rect 2819 1378 2853 1412
rect 2819 1310 2853 1344
rect 2819 1242 2853 1276
rect 2819 1174 2853 1208
rect 2819 1105 2853 1139
rect 2907 1378 2941 1412
rect 2907 1310 2941 1344
rect 2907 1242 2941 1276
rect 2907 1174 2941 1208
rect 2995 1378 3029 1412
rect 2995 1310 3029 1344
rect 2995 1242 3029 1276
rect 2995 1174 3029 1208
rect 2995 1105 3029 1139
rect 3083 1378 3117 1412
rect 3083 1310 3117 1344
rect 3083 1242 3117 1276
rect 3083 1174 3117 1208
rect 3397 1378 3431 1412
rect 3397 1310 3431 1344
rect 3397 1242 3431 1276
rect 3397 1174 3431 1208
rect 3397 1105 3431 1139
rect 3485 1378 3519 1412
rect 3485 1310 3519 1344
rect 3485 1242 3519 1276
rect 3485 1174 3519 1208
rect 3485 1105 3519 1139
rect 3573 1378 3607 1412
rect 3573 1310 3607 1344
rect 3573 1242 3607 1276
rect 3573 1174 3607 1208
rect 3661 1378 3695 1412
rect 3661 1310 3695 1344
rect 3661 1242 3695 1276
rect 3661 1174 3695 1208
rect 3661 1105 3695 1139
rect 3749 1378 3783 1412
rect 3749 1310 3783 1344
rect 3749 1242 3783 1276
rect 3749 1174 3783 1208
rect 4123 1378 4157 1412
rect 4123 1310 4157 1344
rect 4123 1242 4157 1276
rect 4123 1174 4157 1208
rect 4123 1105 4157 1139
rect 4211 1378 4245 1412
rect 4211 1310 4245 1344
rect 4211 1242 4245 1276
rect 4211 1174 4245 1208
rect 4211 1105 4245 1139
rect 4299 1378 4333 1412
rect 4299 1310 4333 1344
rect 4299 1242 4333 1276
rect 4299 1174 4333 1208
rect 4387 1378 4421 1412
rect 4387 1310 4421 1344
rect 4387 1242 4421 1276
rect 4387 1174 4421 1208
rect 4387 1105 4421 1139
rect 4475 1378 4509 1412
rect 4475 1310 4509 1344
rect 4475 1242 4509 1276
rect 4475 1174 4509 1208
rect 4563 1378 4597 1412
rect 4563 1310 4597 1344
rect 4563 1242 4597 1276
rect 4563 1174 4597 1208
rect 4563 1105 4597 1139
rect 4651 1378 4685 1412
rect 4651 1310 4685 1344
rect 4651 1242 4685 1276
rect 4651 1174 4685 1208
<< psubdiff >>
rect -31 546 4915 572
rect -31 512 -17 546
rect 17 512 649 546
rect 683 512 1611 546
rect 1645 512 2573 546
rect 2607 512 3239 546
rect 3273 512 3905 546
rect 3939 512 4867 546
rect 4901 512 4915 546
rect -31 510 4915 512
rect -31 474 31 510
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect -31 368 -17 402
rect 17 368 31 402
rect 635 474 697 510
rect 635 440 649 474
rect 683 440 697 474
rect 635 402 697 440
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect 635 368 649 402
rect 683 368 697 402
rect 1597 474 1659 510
rect 1597 440 1611 474
rect 1645 440 1659 474
rect 1597 402 1659 440
rect 635 330 697 368
rect 635 296 649 330
rect 683 296 697 330
rect 635 258 697 296
rect 635 224 649 258
rect 683 224 697 258
rect 635 186 697 224
rect 635 152 649 186
rect 683 152 697 186
rect 635 114 697 152
rect -31 47 31 80
rect 635 80 649 114
rect 683 80 697 114
rect 1597 368 1611 402
rect 1645 368 1659 402
rect 2559 474 2621 510
rect 2559 440 2573 474
rect 2607 440 2621 474
rect 2559 402 2621 440
rect 1597 330 1659 368
rect 1597 296 1611 330
rect 1645 296 1659 330
rect 1597 258 1659 296
rect 1597 224 1611 258
rect 1645 224 1659 258
rect 1597 186 1659 224
rect 1597 152 1611 186
rect 1645 152 1659 186
rect 1597 114 1659 152
rect 635 47 697 80
rect 1597 80 1611 114
rect 1645 80 1659 114
rect 2559 368 2573 402
rect 2607 368 2621 402
rect 3225 474 3287 510
rect 3225 440 3239 474
rect 3273 440 3287 474
rect 3225 402 3287 440
rect 2559 330 2621 368
rect 2559 296 2573 330
rect 2607 296 2621 330
rect 2559 258 2621 296
rect 2559 224 2573 258
rect 2607 224 2621 258
rect 2559 186 2621 224
rect 2559 152 2573 186
rect 2607 152 2621 186
rect 2559 114 2621 152
rect 1597 47 1659 80
rect 2559 80 2573 114
rect 2607 80 2621 114
rect 3225 368 3239 402
rect 3273 368 3287 402
rect 3891 474 3953 510
rect 3891 440 3905 474
rect 3939 440 3953 474
rect 3891 402 3953 440
rect 3225 330 3287 368
rect 3225 296 3239 330
rect 3273 296 3287 330
rect 3225 258 3287 296
rect 3225 224 3239 258
rect 3273 224 3287 258
rect 3225 186 3287 224
rect 3225 152 3239 186
rect 3273 152 3287 186
rect 3225 114 3287 152
rect 2559 47 2621 80
rect 3225 80 3239 114
rect 3273 80 3287 114
rect 3891 368 3905 402
rect 3939 368 3953 402
rect 4853 474 4915 510
rect 4853 440 4867 474
rect 4901 440 4915 474
rect 4853 402 4915 440
rect 3891 330 3953 368
rect 3891 296 3905 330
rect 3939 296 3953 330
rect 3891 258 3953 296
rect 3891 224 3905 258
rect 3939 224 3953 258
rect 3891 186 3953 224
rect 3891 152 3905 186
rect 3939 152 3953 186
rect 3891 114 3953 152
rect 3225 47 3287 80
rect 3891 80 3905 114
rect 3939 80 3953 114
rect 4853 368 4867 402
rect 4901 368 4915 402
rect 4853 330 4915 368
rect 4853 296 4867 330
rect 4901 296 4915 330
rect 4853 258 4915 296
rect 4853 224 4867 258
rect 4901 224 4915 258
rect 4853 186 4915 224
rect 4853 152 4867 186
rect 4901 152 4915 186
rect 4853 114 4915 152
rect 3891 47 3953 80
rect 4853 80 4867 114
rect 4901 80 4915 114
rect 4853 47 4915 80
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 361 47
rect 395 13 433 47
rect 467 13 505 47
rect 539 13 577 47
rect 611 13 721 47
rect 755 13 793 47
rect 827 13 865 47
rect 899 13 937 47
rect 971 13 1009 47
rect 1043 13 1081 47
rect 1115 13 1179 47
rect 1213 13 1251 47
rect 1285 13 1323 47
rect 1357 13 1395 47
rect 1429 13 1467 47
rect 1501 13 1539 47
rect 1573 13 1683 47
rect 1717 13 1755 47
rect 1789 13 1827 47
rect 1861 13 1899 47
rect 1933 13 1971 47
rect 2005 13 2043 47
rect 2077 13 2141 47
rect 2175 13 2213 47
rect 2247 13 2285 47
rect 2319 13 2357 47
rect 2391 13 2429 47
rect 2463 13 2501 47
rect 2535 13 2645 47
rect 2679 13 2717 47
rect 2751 13 2789 47
rect 2823 13 2861 47
rect 2895 13 2951 47
rect 2985 13 3023 47
rect 3057 13 3095 47
rect 3129 13 3167 47
rect 3201 13 3311 47
rect 3345 13 3383 47
rect 3417 13 3455 47
rect 3489 13 3527 47
rect 3561 13 3617 47
rect 3651 13 3689 47
rect 3723 13 3761 47
rect 3795 13 3833 47
rect 3867 13 3977 47
rect 4011 13 4049 47
rect 4083 13 4121 47
rect 4155 13 4193 47
rect 4227 13 4265 47
rect 4299 13 4337 47
rect 4371 13 4435 47
rect 4469 13 4507 47
rect 4541 13 4579 47
rect 4613 13 4651 47
rect 4685 13 4723 47
rect 4757 13 4795 47
rect 4829 13 4915 47
rect -31 11 31 13
rect 635 11 697 13
rect 1597 11 1659 13
rect 2559 11 2621 13
rect 3225 11 3287 13
rect 3891 11 3953 13
rect 4853 11 4915 13
<< nsubdiff >>
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 361 1539
rect 395 1505 433 1539
rect 467 1505 505 1539
rect 539 1505 577 1539
rect 611 1505 721 1539
rect 755 1505 793 1539
rect 827 1505 865 1539
rect 899 1505 937 1539
rect 971 1505 1009 1539
rect 1043 1505 1081 1539
rect 1115 1505 1179 1539
rect 1213 1505 1251 1539
rect 1285 1505 1323 1539
rect 1357 1505 1395 1539
rect 1429 1505 1467 1539
rect 1501 1505 1539 1539
rect 1573 1505 1683 1539
rect 1717 1505 1755 1539
rect 1789 1505 1827 1539
rect 1861 1505 1899 1539
rect 1933 1505 1971 1539
rect 2005 1505 2043 1539
rect 2077 1505 2141 1539
rect 2175 1505 2213 1539
rect 2247 1505 2285 1539
rect 2319 1505 2357 1539
rect 2391 1505 2429 1539
rect 2463 1505 2501 1539
rect 2535 1505 2645 1539
rect 2679 1505 2717 1539
rect 2751 1505 2789 1539
rect 2823 1505 2861 1539
rect 2895 1505 2951 1539
rect 2985 1505 3023 1539
rect 3057 1505 3095 1539
rect 3129 1505 3167 1539
rect 3201 1505 3311 1539
rect 3345 1505 3383 1539
rect 3417 1505 3455 1539
rect 3489 1505 3527 1539
rect 3561 1505 3617 1539
rect 3651 1505 3689 1539
rect 3723 1505 3761 1539
rect 3795 1505 3833 1539
rect 3867 1505 3977 1539
rect 4011 1505 4049 1539
rect 4083 1505 4121 1539
rect 4155 1505 4193 1539
rect 4227 1505 4265 1539
rect 4299 1505 4337 1539
rect 4371 1505 4435 1539
rect 4469 1505 4507 1539
rect 4541 1505 4579 1539
rect 4613 1505 4651 1539
rect 4685 1505 4723 1539
rect 4757 1505 4795 1539
rect 4829 1505 4915 1539
rect -31 1470 31 1505
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect 635 1470 697 1505
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect -31 1038 31 1076
rect 635 1436 649 1470
rect 683 1436 697 1470
rect 1597 1470 1659 1505
rect 635 1398 697 1436
rect 635 1364 649 1398
rect 683 1364 697 1398
rect 635 1326 697 1364
rect 635 1292 649 1326
rect 683 1292 697 1326
rect 635 1254 697 1292
rect 635 1220 649 1254
rect 683 1220 697 1254
rect 635 1182 697 1220
rect 635 1148 649 1182
rect 683 1148 697 1182
rect 635 1110 697 1148
rect 635 1076 649 1110
rect 683 1076 697 1110
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect 635 1038 697 1076
rect 1597 1436 1611 1470
rect 1645 1436 1659 1470
rect 2559 1470 2621 1505
rect 1597 1398 1659 1436
rect 1597 1364 1611 1398
rect 1645 1364 1659 1398
rect 1597 1326 1659 1364
rect 1597 1292 1611 1326
rect 1645 1292 1659 1326
rect 1597 1254 1659 1292
rect 1597 1220 1611 1254
rect 1645 1220 1659 1254
rect 1597 1182 1659 1220
rect 1597 1148 1611 1182
rect 1645 1148 1659 1182
rect 1597 1110 1659 1148
rect 1597 1076 1611 1110
rect 1645 1076 1659 1110
rect 635 1004 649 1038
rect 683 1004 697 1038
rect 635 966 697 1004
rect -31 930 31 932
rect 635 932 649 966
rect 683 932 697 966
rect 1597 1038 1659 1076
rect 2559 1436 2573 1470
rect 2607 1436 2621 1470
rect 3225 1470 3287 1505
rect 2559 1398 2621 1436
rect 2559 1364 2573 1398
rect 2607 1364 2621 1398
rect 2559 1326 2621 1364
rect 2559 1292 2573 1326
rect 2607 1292 2621 1326
rect 2559 1254 2621 1292
rect 2559 1220 2573 1254
rect 2607 1220 2621 1254
rect 2559 1182 2621 1220
rect 2559 1148 2573 1182
rect 2607 1148 2621 1182
rect 2559 1110 2621 1148
rect 2559 1076 2573 1110
rect 2607 1076 2621 1110
rect 1597 1004 1611 1038
rect 1645 1004 1659 1038
rect 1597 966 1659 1004
rect 635 930 697 932
rect 1597 932 1611 966
rect 1645 932 1659 966
rect 2559 1038 2621 1076
rect 3225 1436 3239 1470
rect 3273 1436 3287 1470
rect 3891 1470 3953 1505
rect 3225 1398 3287 1436
rect 3225 1364 3239 1398
rect 3273 1364 3287 1398
rect 3225 1326 3287 1364
rect 3225 1292 3239 1326
rect 3273 1292 3287 1326
rect 3225 1254 3287 1292
rect 3225 1220 3239 1254
rect 3273 1220 3287 1254
rect 3225 1182 3287 1220
rect 3225 1148 3239 1182
rect 3273 1148 3287 1182
rect 3225 1110 3287 1148
rect 3225 1076 3239 1110
rect 3273 1076 3287 1110
rect 2559 1004 2573 1038
rect 2607 1004 2621 1038
rect 2559 966 2621 1004
rect 1597 930 1659 932
rect 2559 932 2573 966
rect 2607 932 2621 966
rect 3225 1038 3287 1076
rect 3891 1436 3905 1470
rect 3939 1436 3953 1470
rect 4853 1470 4915 1505
rect 3891 1398 3953 1436
rect 3891 1364 3905 1398
rect 3939 1364 3953 1398
rect 3891 1326 3953 1364
rect 3891 1292 3905 1326
rect 3939 1292 3953 1326
rect 3891 1254 3953 1292
rect 3891 1220 3905 1254
rect 3939 1220 3953 1254
rect 3891 1182 3953 1220
rect 3891 1148 3905 1182
rect 3939 1148 3953 1182
rect 3891 1110 3953 1148
rect 3891 1076 3905 1110
rect 3939 1076 3953 1110
rect 3225 1004 3239 1038
rect 3273 1004 3287 1038
rect 3225 966 3287 1004
rect 2559 930 2621 932
rect 3225 932 3239 966
rect 3273 932 3287 966
rect 3891 1038 3953 1076
rect 4853 1436 4867 1470
rect 4901 1436 4915 1470
rect 4853 1398 4915 1436
rect 4853 1364 4867 1398
rect 4901 1364 4915 1398
rect 4853 1326 4915 1364
rect 4853 1292 4867 1326
rect 4901 1292 4915 1326
rect 4853 1254 4915 1292
rect 4853 1220 4867 1254
rect 4901 1220 4915 1254
rect 4853 1182 4915 1220
rect 4853 1148 4867 1182
rect 4901 1148 4915 1182
rect 4853 1110 4915 1148
rect 4853 1076 4867 1110
rect 4901 1076 4915 1110
rect 3891 1004 3905 1038
rect 3939 1004 3953 1038
rect 3891 966 3953 1004
rect 3225 930 3287 932
rect 3891 932 3905 966
rect 3939 932 3953 966
rect 4853 1038 4915 1076
rect 4853 1004 4867 1038
rect 4901 1004 4915 1038
rect 4853 966 4915 1004
rect 3891 930 3953 932
rect 4853 932 4867 966
rect 4901 932 4915 966
rect 4853 930 4915 932
rect -31 868 4915 930
<< psubdiffcont >>
rect -17 512 17 546
rect 649 512 683 546
rect 1611 512 1645 546
rect 2573 512 2607 546
rect 3239 512 3273 546
rect 3905 512 3939 546
rect 4867 512 4901 546
rect -17 440 17 474
rect -17 368 17 402
rect 649 440 683 474
rect -17 296 17 330
rect -17 224 17 258
rect -17 152 17 186
rect -17 80 17 114
rect 649 368 683 402
rect 1611 440 1645 474
rect 649 296 683 330
rect 649 224 683 258
rect 649 152 683 186
rect 649 80 683 114
rect 1611 368 1645 402
rect 2573 440 2607 474
rect 1611 296 1645 330
rect 1611 224 1645 258
rect 1611 152 1645 186
rect 1611 80 1645 114
rect 2573 368 2607 402
rect 3239 440 3273 474
rect 2573 296 2607 330
rect 2573 224 2607 258
rect 2573 152 2607 186
rect 2573 80 2607 114
rect 3239 368 3273 402
rect 3905 440 3939 474
rect 3239 296 3273 330
rect 3239 224 3273 258
rect 3239 152 3273 186
rect 3239 80 3273 114
rect 3905 368 3939 402
rect 4867 440 4901 474
rect 3905 296 3939 330
rect 3905 224 3939 258
rect 3905 152 3939 186
rect 3905 80 3939 114
rect 4867 368 4901 402
rect 4867 296 4901 330
rect 4867 224 4901 258
rect 4867 152 4901 186
rect 4867 80 4901 114
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 361 13 395 47
rect 433 13 467 47
rect 505 13 539 47
rect 577 13 611 47
rect 721 13 755 47
rect 793 13 827 47
rect 865 13 899 47
rect 937 13 971 47
rect 1009 13 1043 47
rect 1081 13 1115 47
rect 1179 13 1213 47
rect 1251 13 1285 47
rect 1323 13 1357 47
rect 1395 13 1429 47
rect 1467 13 1501 47
rect 1539 13 1573 47
rect 1683 13 1717 47
rect 1755 13 1789 47
rect 1827 13 1861 47
rect 1899 13 1933 47
rect 1971 13 2005 47
rect 2043 13 2077 47
rect 2141 13 2175 47
rect 2213 13 2247 47
rect 2285 13 2319 47
rect 2357 13 2391 47
rect 2429 13 2463 47
rect 2501 13 2535 47
rect 2645 13 2679 47
rect 2717 13 2751 47
rect 2789 13 2823 47
rect 2861 13 2895 47
rect 2951 13 2985 47
rect 3023 13 3057 47
rect 3095 13 3129 47
rect 3167 13 3201 47
rect 3311 13 3345 47
rect 3383 13 3417 47
rect 3455 13 3489 47
rect 3527 13 3561 47
rect 3617 13 3651 47
rect 3689 13 3723 47
rect 3761 13 3795 47
rect 3833 13 3867 47
rect 3977 13 4011 47
rect 4049 13 4083 47
rect 4121 13 4155 47
rect 4193 13 4227 47
rect 4265 13 4299 47
rect 4337 13 4371 47
rect 4435 13 4469 47
rect 4507 13 4541 47
rect 4579 13 4613 47
rect 4651 13 4685 47
rect 4723 13 4757 47
rect 4795 13 4829 47
<< nsubdiffcont >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 361 1505 395 1539
rect 433 1505 467 1539
rect 505 1505 539 1539
rect 577 1505 611 1539
rect 721 1505 755 1539
rect 793 1505 827 1539
rect 865 1505 899 1539
rect 937 1505 971 1539
rect 1009 1505 1043 1539
rect 1081 1505 1115 1539
rect 1179 1505 1213 1539
rect 1251 1505 1285 1539
rect 1323 1505 1357 1539
rect 1395 1505 1429 1539
rect 1467 1505 1501 1539
rect 1539 1505 1573 1539
rect 1683 1505 1717 1539
rect 1755 1505 1789 1539
rect 1827 1505 1861 1539
rect 1899 1505 1933 1539
rect 1971 1505 2005 1539
rect 2043 1505 2077 1539
rect 2141 1505 2175 1539
rect 2213 1505 2247 1539
rect 2285 1505 2319 1539
rect 2357 1505 2391 1539
rect 2429 1505 2463 1539
rect 2501 1505 2535 1539
rect 2645 1505 2679 1539
rect 2717 1505 2751 1539
rect 2789 1505 2823 1539
rect 2861 1505 2895 1539
rect 2951 1505 2985 1539
rect 3023 1505 3057 1539
rect 3095 1505 3129 1539
rect 3167 1505 3201 1539
rect 3311 1505 3345 1539
rect 3383 1505 3417 1539
rect 3455 1505 3489 1539
rect 3527 1505 3561 1539
rect 3617 1505 3651 1539
rect 3689 1505 3723 1539
rect 3761 1505 3795 1539
rect 3833 1505 3867 1539
rect 3977 1505 4011 1539
rect 4049 1505 4083 1539
rect 4121 1505 4155 1539
rect 4193 1505 4227 1539
rect 4265 1505 4299 1539
rect 4337 1505 4371 1539
rect 4435 1505 4469 1539
rect 4507 1505 4541 1539
rect 4579 1505 4613 1539
rect 4651 1505 4685 1539
rect 4723 1505 4757 1539
rect 4795 1505 4829 1539
rect -17 1436 17 1470
rect -17 1364 17 1398
rect -17 1292 17 1326
rect -17 1220 17 1254
rect -17 1148 17 1182
rect -17 1076 17 1110
rect 649 1436 683 1470
rect 649 1364 683 1398
rect 649 1292 683 1326
rect 649 1220 683 1254
rect 649 1148 683 1182
rect 649 1076 683 1110
rect -17 1004 17 1038
rect -17 932 17 966
rect 1611 1436 1645 1470
rect 1611 1364 1645 1398
rect 1611 1292 1645 1326
rect 1611 1220 1645 1254
rect 1611 1148 1645 1182
rect 1611 1076 1645 1110
rect 649 1004 683 1038
rect 649 932 683 966
rect 2573 1436 2607 1470
rect 2573 1364 2607 1398
rect 2573 1292 2607 1326
rect 2573 1220 2607 1254
rect 2573 1148 2607 1182
rect 2573 1076 2607 1110
rect 1611 1004 1645 1038
rect 1611 932 1645 966
rect 3239 1436 3273 1470
rect 3239 1364 3273 1398
rect 3239 1292 3273 1326
rect 3239 1220 3273 1254
rect 3239 1148 3273 1182
rect 3239 1076 3273 1110
rect 2573 1004 2607 1038
rect 2573 932 2607 966
rect 3905 1436 3939 1470
rect 3905 1364 3939 1398
rect 3905 1292 3939 1326
rect 3905 1220 3939 1254
rect 3905 1148 3939 1182
rect 3905 1076 3939 1110
rect 3239 1004 3273 1038
rect 3239 932 3273 966
rect 4867 1436 4901 1470
rect 4867 1364 4901 1398
rect 4867 1292 4901 1326
rect 4867 1220 4901 1254
rect 4867 1148 4901 1182
rect 4867 1076 4901 1110
rect 3905 1004 3939 1038
rect 3905 932 3939 966
rect 4867 1004 4901 1038
rect 4867 932 4901 966
<< poly >>
rect 187 1450 217 1476
rect 275 1450 305 1476
rect 363 1450 393 1476
rect 451 1450 481 1476
rect 913 1450 943 1476
rect 1001 1450 1031 1476
rect 1089 1450 1119 1476
rect 1177 1450 1207 1476
rect 1265 1450 1295 1476
rect 1353 1450 1383 1476
rect 187 1019 217 1050
rect 275 1019 305 1050
rect 363 1019 393 1050
rect 451 1019 481 1050
rect 187 1003 305 1019
rect 187 989 205 1003
rect 195 969 205 989
rect 239 989 305 1003
rect 349 1003 481 1019
rect 239 969 249 989
rect 195 953 249 969
rect 349 969 359 1003
rect 393 989 481 1003
rect 1875 1450 1905 1476
rect 1963 1450 1993 1476
rect 2051 1450 2081 1476
rect 2139 1450 2169 1476
rect 2227 1450 2257 1476
rect 2315 1450 2345 1476
rect 913 1019 943 1050
rect 1001 1019 1031 1050
rect 1089 1019 1119 1050
rect 1177 1019 1207 1050
rect 393 969 403 989
rect 349 953 403 969
rect 861 1003 1031 1019
rect 861 969 871 1003
rect 905 989 1031 1003
rect 1083 1003 1207 1019
rect 905 969 915 989
rect 861 953 915 969
rect 1083 969 1093 1003
rect 1127 989 1207 1003
rect 1265 1019 1295 1050
rect 1353 1019 1383 1050
rect 1265 1003 1383 1019
rect 1265 989 1315 1003
rect 1127 969 1137 989
rect 1083 953 1137 969
rect 1305 969 1315 989
rect 1349 989 1383 1003
rect 2777 1450 2807 1476
rect 2865 1450 2895 1476
rect 2953 1450 2983 1476
rect 3041 1450 3071 1476
rect 1875 1019 1905 1050
rect 1963 1019 1993 1050
rect 2051 1019 2081 1050
rect 2139 1019 2169 1050
rect 1349 969 1359 989
rect 1305 953 1359 969
rect 1823 1003 1993 1019
rect 1823 969 1833 1003
rect 1867 989 1993 1003
rect 2045 1003 2169 1019
rect 1867 969 1877 989
rect 1823 953 1877 969
rect 2045 969 2055 1003
rect 2089 989 2169 1003
rect 2227 1019 2257 1050
rect 2315 1019 2345 1050
rect 2227 1003 2345 1019
rect 2227 989 2277 1003
rect 2089 969 2099 989
rect 2045 953 2099 969
rect 2267 969 2277 989
rect 2311 989 2345 1003
rect 3443 1450 3473 1476
rect 3531 1450 3561 1476
rect 3619 1450 3649 1476
rect 3707 1450 3737 1476
rect 2311 969 2321 989
rect 2267 953 2321 969
rect 2777 1019 2807 1050
rect 2865 1019 2895 1050
rect 2953 1019 2983 1050
rect 3041 1019 3071 1050
rect 2777 1003 2895 1019
rect 2777 989 2795 1003
rect 2785 969 2795 989
rect 2829 989 2895 1003
rect 2939 1003 3071 1019
rect 2829 969 2839 989
rect 2785 953 2839 969
rect 2939 969 2949 1003
rect 2983 989 3071 1003
rect 4169 1450 4199 1476
rect 4257 1450 4287 1476
rect 4345 1450 4375 1476
rect 4433 1450 4463 1476
rect 4521 1450 4551 1476
rect 4609 1450 4639 1476
rect 2983 969 2993 989
rect 2939 953 2993 969
rect 3443 1019 3473 1050
rect 3531 1019 3561 1050
rect 3619 1019 3649 1050
rect 3707 1019 3737 1050
rect 3443 1003 3561 1019
rect 3443 989 3461 1003
rect 3451 969 3461 989
rect 3495 989 3561 1003
rect 3605 1003 3737 1019
rect 3495 969 3505 989
rect 3451 953 3505 969
rect 3605 969 3615 1003
rect 3649 989 3737 1003
rect 4169 1019 4199 1050
rect 4257 1019 4287 1050
rect 4345 1019 4375 1050
rect 4433 1019 4463 1050
rect 3649 969 3659 989
rect 3605 953 3659 969
rect 4117 1003 4287 1019
rect 4117 969 4127 1003
rect 4161 989 4287 1003
rect 4339 1003 4463 1019
rect 4161 969 4171 989
rect 4117 953 4171 969
rect 4339 969 4349 1003
rect 4383 989 4463 1003
rect 4521 1019 4551 1050
rect 4609 1019 4639 1050
rect 4521 1003 4639 1019
rect 4521 989 4571 1003
rect 4383 969 4393 989
rect 4339 953 4393 969
rect 4561 969 4571 989
rect 4605 989 4639 1003
rect 4605 969 4615 989
rect 4561 953 4615 969
rect 195 461 249 477
rect 195 441 205 461
rect 168 427 205 441
rect 239 427 249 461
rect 168 411 249 427
rect 343 461 397 477
rect 343 427 353 461
rect 387 427 397 461
rect 343 411 397 427
rect 861 461 915 477
rect 861 441 871 461
rect 168 377 198 411
rect 362 377 392 411
rect 813 427 871 441
rect 905 427 915 461
rect 813 411 915 427
rect 1083 461 1137 477
rect 1083 427 1093 461
rect 1127 441 1137 461
rect 1305 461 1359 477
rect 1127 427 1143 441
rect 1083 411 1143 427
rect 1305 427 1315 461
rect 1349 427 1359 461
rect 1305 411 1359 427
rect 1823 461 1877 477
rect 1823 441 1833 461
rect 813 379 843 411
rect 1113 379 1143 411
rect 1315 379 1345 411
rect 1775 427 1833 441
rect 1867 427 1877 461
rect 1775 411 1877 427
rect 2045 461 2099 477
rect 2045 427 2055 461
rect 2089 441 2099 461
rect 2267 461 2321 477
rect 2089 427 2105 441
rect 2045 411 2105 427
rect 2267 427 2277 461
rect 2311 427 2321 461
rect 2267 411 2321 427
rect 2785 461 2839 477
rect 2785 441 2795 461
rect 1775 379 1805 411
rect 2075 379 2105 411
rect 2277 379 2307 411
rect 2758 427 2795 441
rect 2829 427 2839 461
rect 2758 411 2839 427
rect 2933 461 2987 477
rect 2933 427 2943 461
rect 2977 427 2987 461
rect 2933 411 2987 427
rect 3451 461 3505 477
rect 3451 441 3461 461
rect 2758 377 2788 411
rect 2952 377 2982 411
rect 3424 427 3461 441
rect 3495 427 3505 461
rect 3424 411 3505 427
rect 3599 461 3653 477
rect 3599 427 3609 461
rect 3643 427 3653 461
rect 3599 411 3653 427
rect 4117 461 4171 477
rect 4117 441 4127 461
rect 3424 377 3454 411
rect 3618 377 3648 411
rect 4069 427 4127 441
rect 4161 427 4171 461
rect 4069 411 4171 427
rect 4339 461 4393 477
rect 4339 427 4349 461
rect 4383 441 4393 461
rect 4561 461 4615 477
rect 4383 427 4399 441
rect 4339 411 4399 427
rect 4561 427 4571 461
rect 4605 427 4615 461
rect 4561 411 4615 427
rect 4069 379 4099 411
rect 4369 379 4399 411
rect 4571 379 4601 411
<< polycont >>
rect 205 969 239 1003
rect 359 969 393 1003
rect 871 969 905 1003
rect 1093 969 1127 1003
rect 1315 969 1349 1003
rect 1833 969 1867 1003
rect 2055 969 2089 1003
rect 2277 969 2311 1003
rect 2795 969 2829 1003
rect 2949 969 2983 1003
rect 3461 969 3495 1003
rect 3615 969 3649 1003
rect 4127 969 4161 1003
rect 4349 969 4383 1003
rect 4571 969 4605 1003
rect 205 427 239 461
rect 353 427 387 461
rect 871 427 905 461
rect 1093 427 1127 461
rect 1315 427 1349 461
rect 1833 427 1867 461
rect 2055 427 2089 461
rect 2277 427 2311 461
rect 2795 427 2829 461
rect 2943 427 2977 461
rect 3461 427 3495 461
rect 3609 427 3643 461
rect 4127 427 4161 461
rect 4349 427 4383 461
rect 4571 427 4605 461
<< locali >>
rect -31 1539 4915 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 361 1539
rect 395 1505 433 1539
rect 467 1505 505 1539
rect 539 1505 577 1539
rect 611 1505 721 1539
rect 755 1505 793 1539
rect 827 1505 865 1539
rect 899 1505 937 1539
rect 971 1505 1009 1539
rect 1043 1505 1081 1539
rect 1115 1505 1179 1539
rect 1213 1505 1251 1539
rect 1285 1505 1323 1539
rect 1357 1505 1395 1539
rect 1429 1505 1467 1539
rect 1501 1505 1539 1539
rect 1573 1505 1683 1539
rect 1717 1505 1755 1539
rect 1789 1505 1827 1539
rect 1861 1505 1899 1539
rect 1933 1505 1971 1539
rect 2005 1505 2043 1539
rect 2077 1505 2141 1539
rect 2175 1505 2213 1539
rect 2247 1505 2285 1539
rect 2319 1505 2357 1539
rect 2391 1505 2429 1539
rect 2463 1505 2501 1539
rect 2535 1505 2645 1539
rect 2679 1505 2717 1539
rect 2751 1505 2789 1539
rect 2823 1505 2861 1539
rect 2895 1505 2951 1539
rect 2985 1505 3023 1539
rect 3057 1505 3095 1539
rect 3129 1505 3167 1539
rect 3201 1505 3311 1539
rect 3345 1505 3383 1539
rect 3417 1505 3455 1539
rect 3489 1505 3527 1539
rect 3561 1505 3617 1539
rect 3651 1505 3689 1539
rect 3723 1505 3761 1539
rect 3795 1505 3833 1539
rect 3867 1505 3977 1539
rect 4011 1505 4049 1539
rect 4083 1505 4121 1539
rect 4155 1505 4193 1539
rect 4227 1505 4265 1539
rect 4299 1505 4337 1539
rect 4371 1505 4435 1539
rect 4469 1505 4507 1539
rect 4541 1505 4579 1539
rect 4613 1505 4651 1539
rect 4685 1505 4723 1539
rect 4757 1505 4795 1539
rect 4829 1505 4915 1539
rect -31 1492 4915 1505
rect -31 1470 31 1492
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect -31 1038 31 1076
rect 141 1412 175 1492
rect 141 1344 175 1378
rect 141 1276 175 1310
rect 141 1208 175 1242
rect 141 1139 175 1174
rect 141 1073 175 1105
rect 229 1412 263 1450
rect 229 1344 263 1378
rect 229 1276 263 1310
rect 229 1208 263 1242
rect 229 1139 263 1174
rect 317 1412 351 1492
rect 317 1344 351 1378
rect 317 1276 351 1310
rect 317 1208 351 1242
rect 317 1157 351 1174
rect 405 1412 439 1450
rect 405 1344 439 1378
rect 405 1276 439 1310
rect 405 1208 439 1242
rect 229 1103 263 1105
rect 405 1139 439 1174
rect 493 1412 527 1492
rect 493 1344 527 1378
rect 493 1276 527 1310
rect 493 1208 527 1242
rect 493 1157 527 1174
rect 635 1470 697 1492
rect 635 1436 649 1470
rect 683 1436 697 1470
rect 635 1398 697 1436
rect 635 1364 649 1398
rect 683 1364 697 1398
rect 635 1326 697 1364
rect 635 1292 649 1326
rect 683 1292 697 1326
rect 635 1254 697 1292
rect 635 1220 649 1254
rect 683 1220 697 1254
rect 635 1182 697 1220
rect 405 1103 439 1105
rect 635 1148 649 1182
rect 683 1148 697 1182
rect 635 1110 697 1148
rect 229 1069 535 1103
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect -31 868 31 932
rect 205 1003 239 1019
rect 359 1003 393 1019
rect 205 831 239 969
rect -31 546 31 572
rect -31 512 -17 546
rect 17 512 31 546
rect -31 474 31 512
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect 205 461 239 797
rect 205 411 239 427
rect 353 969 359 988
rect 353 953 393 969
rect 353 905 387 953
rect 353 461 387 871
rect 353 411 387 427
rect 501 609 535 1069
rect 635 1076 649 1110
rect 683 1076 697 1110
rect 867 1412 901 1492
rect 867 1344 901 1378
rect 867 1276 901 1310
rect 867 1208 901 1242
rect 867 1139 901 1174
rect 867 1089 901 1105
rect 955 1412 989 1450
rect 955 1344 989 1378
rect 955 1276 989 1310
rect 955 1208 989 1242
rect 955 1139 989 1174
rect 1043 1412 1077 1492
rect 1043 1344 1077 1378
rect 1043 1276 1077 1310
rect 1043 1208 1077 1242
rect 1043 1157 1077 1174
rect 1131 1412 1165 1450
rect 1131 1344 1165 1378
rect 1131 1276 1165 1310
rect 1131 1208 1165 1242
rect 955 1094 989 1105
rect 1131 1139 1165 1174
rect 1219 1412 1253 1492
rect 1219 1344 1253 1378
rect 1219 1276 1253 1310
rect 1219 1208 1253 1242
rect 1219 1157 1253 1174
rect 1307 1412 1341 1450
rect 1307 1344 1341 1378
rect 1307 1276 1341 1310
rect 1307 1208 1341 1242
rect 1131 1094 1165 1105
rect 1307 1139 1341 1174
rect 1395 1412 1429 1492
rect 1395 1344 1429 1378
rect 1395 1276 1429 1310
rect 1395 1208 1429 1242
rect 1395 1157 1429 1174
rect 1597 1470 1659 1492
rect 1597 1436 1611 1470
rect 1645 1436 1659 1470
rect 1597 1398 1659 1436
rect 1597 1364 1611 1398
rect 1645 1364 1659 1398
rect 1597 1326 1659 1364
rect 1597 1292 1611 1326
rect 1645 1292 1659 1326
rect 1597 1254 1659 1292
rect 1597 1220 1611 1254
rect 1645 1220 1659 1254
rect 1597 1182 1659 1220
rect 1307 1094 1341 1105
rect 1597 1148 1611 1182
rect 1645 1148 1659 1182
rect 1597 1110 1659 1148
rect 635 1038 697 1076
rect 955 1060 1497 1094
rect 635 1004 649 1038
rect 683 1004 697 1038
rect 635 966 697 1004
rect 635 932 649 966
rect 683 932 697 966
rect 635 868 697 932
rect 871 1003 905 1019
rect -31 368 -17 402
rect 17 368 31 402
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect 122 361 156 377
rect 316 361 350 377
rect 501 376 535 575
rect 871 608 905 969
rect 156 327 219 361
rect 253 327 316 361
rect 122 289 156 327
rect 122 221 156 255
rect 316 289 350 327
rect 122 151 156 187
rect 122 101 156 117
rect 219 236 253 252
rect -31 62 31 80
rect 219 62 253 202
rect 316 221 350 255
rect 413 342 535 376
rect 635 546 697 572
rect 635 512 649 546
rect 683 512 697 546
rect 635 474 697 512
rect 635 440 649 474
rect 683 440 697 474
rect 635 402 697 440
rect 871 461 905 574
rect 871 411 905 427
rect 1093 1003 1127 1019
rect 1093 461 1127 945
rect 1093 411 1127 427
rect 1315 1003 1349 1019
rect 1315 831 1349 969
rect 1463 921 1497 1060
rect 1462 905 1497 921
rect 1496 871 1497 905
rect 1462 855 1497 871
rect 1597 1076 1611 1110
rect 1645 1076 1659 1110
rect 1829 1412 1863 1492
rect 1829 1344 1863 1378
rect 1829 1276 1863 1310
rect 1829 1208 1863 1242
rect 1829 1139 1863 1174
rect 1829 1089 1863 1105
rect 1917 1412 1951 1450
rect 1917 1344 1951 1378
rect 1917 1276 1951 1310
rect 1917 1208 1951 1242
rect 1917 1139 1951 1174
rect 2005 1412 2039 1492
rect 2005 1344 2039 1378
rect 2005 1276 2039 1310
rect 2005 1208 2039 1242
rect 2005 1157 2039 1174
rect 2093 1412 2127 1450
rect 2093 1344 2127 1378
rect 2093 1276 2127 1310
rect 2093 1208 2127 1242
rect 1917 1094 1951 1105
rect 2093 1139 2127 1174
rect 2181 1412 2215 1492
rect 2181 1344 2215 1378
rect 2181 1276 2215 1310
rect 2181 1208 2215 1242
rect 2181 1157 2215 1174
rect 2269 1412 2303 1450
rect 2269 1344 2303 1378
rect 2269 1276 2303 1310
rect 2269 1208 2303 1242
rect 2093 1094 2127 1105
rect 2269 1139 2303 1174
rect 2357 1412 2391 1492
rect 2357 1344 2391 1378
rect 2357 1276 2391 1310
rect 2357 1208 2391 1242
rect 2357 1157 2391 1174
rect 2559 1470 2621 1492
rect 2559 1436 2573 1470
rect 2607 1436 2621 1470
rect 2559 1398 2621 1436
rect 2559 1364 2573 1398
rect 2607 1364 2621 1398
rect 2559 1326 2621 1364
rect 2559 1292 2573 1326
rect 2607 1292 2621 1326
rect 2559 1254 2621 1292
rect 2559 1220 2573 1254
rect 2607 1220 2621 1254
rect 2559 1182 2621 1220
rect 2269 1094 2303 1105
rect 2559 1148 2573 1182
rect 2607 1148 2621 1182
rect 2559 1110 2621 1148
rect 1597 1038 1659 1076
rect 1917 1060 2459 1094
rect 1597 1004 1611 1038
rect 1645 1004 1659 1038
rect 1597 966 1659 1004
rect 1597 932 1611 966
rect 1645 932 1659 966
rect 1597 868 1659 932
rect 1833 1003 1867 1019
rect 1315 461 1349 797
rect 1315 411 1349 427
rect 635 368 649 402
rect 683 368 697 402
rect 413 245 447 342
rect 635 330 697 368
rect 413 195 447 211
rect 510 289 544 305
rect 510 221 544 255
rect 316 151 350 187
rect 510 151 544 187
rect 350 117 413 151
rect 447 117 510 151
rect 316 101 350 117
rect 510 101 544 117
rect 635 296 649 330
rect 683 296 697 330
rect 635 258 697 296
rect 635 224 649 258
rect 683 224 697 258
rect 635 186 697 224
rect 635 152 649 186
rect 683 152 697 186
rect 635 114 697 152
rect 635 80 649 114
rect 683 80 697 114
rect 767 363 801 379
rect 961 363 995 379
rect 1155 363 1189 379
rect 801 329 864 363
rect 898 329 961 363
rect 995 329 1058 363
rect 1092 329 1155 363
rect 767 291 801 329
rect 767 223 801 257
rect 961 291 995 329
rect 1155 313 1189 329
rect 1269 363 1303 379
rect 1463 378 1497 855
rect 1833 609 1867 969
rect 1269 291 1303 329
rect 767 153 801 189
rect 767 103 801 119
rect 864 238 898 254
rect 635 62 697 80
rect 864 62 898 204
rect 961 223 995 257
rect 1059 244 1093 260
rect 1269 244 1303 257
rect 1093 223 1303 244
rect 1093 210 1269 223
rect 1059 194 1093 210
rect 961 153 995 189
rect 1366 344 1497 378
rect 1597 546 1659 572
rect 1597 512 1611 546
rect 1645 512 1659 546
rect 1597 474 1659 512
rect 1597 440 1611 474
rect 1645 440 1659 474
rect 1597 402 1659 440
rect 1833 461 1867 575
rect 1833 411 1867 427
rect 2055 1003 2089 1019
rect 2055 535 2089 969
rect 2055 461 2089 501
rect 2055 411 2089 427
rect 2277 1003 2311 1019
rect 2277 831 2311 969
rect 2277 461 2311 797
rect 2277 411 2311 427
rect 2425 609 2459 1060
rect 2559 1076 2573 1110
rect 2607 1076 2621 1110
rect 2559 1038 2621 1076
rect 2731 1412 2765 1492
rect 2731 1344 2765 1378
rect 2731 1276 2765 1310
rect 2731 1208 2765 1242
rect 2731 1139 2765 1174
rect 2731 1073 2765 1105
rect 2819 1412 2853 1450
rect 2819 1344 2853 1378
rect 2819 1276 2853 1310
rect 2819 1208 2853 1242
rect 2819 1139 2853 1174
rect 2907 1412 2941 1492
rect 2907 1344 2941 1378
rect 2907 1276 2941 1310
rect 2907 1208 2941 1242
rect 2907 1157 2941 1174
rect 2995 1412 3029 1450
rect 2995 1344 3029 1378
rect 2995 1276 3029 1310
rect 2995 1208 3029 1242
rect 2819 1103 2853 1105
rect 2995 1139 3029 1174
rect 3083 1412 3117 1492
rect 3083 1344 3117 1378
rect 3083 1276 3117 1310
rect 3083 1208 3117 1242
rect 3083 1157 3117 1174
rect 3225 1470 3287 1492
rect 3225 1436 3239 1470
rect 3273 1436 3287 1470
rect 3225 1398 3287 1436
rect 3225 1364 3239 1398
rect 3273 1364 3287 1398
rect 3225 1326 3287 1364
rect 3225 1292 3239 1326
rect 3273 1292 3287 1326
rect 3225 1254 3287 1292
rect 3225 1220 3239 1254
rect 3273 1220 3287 1254
rect 3225 1182 3287 1220
rect 2995 1103 3029 1105
rect 3225 1148 3239 1182
rect 3273 1148 3287 1182
rect 3225 1110 3287 1148
rect 2819 1069 3125 1103
rect 2559 1004 2573 1038
rect 2607 1004 2621 1038
rect 2559 966 2621 1004
rect 2559 932 2573 966
rect 2607 932 2621 966
rect 2559 868 2621 932
rect 2795 1003 2829 1019
rect 2949 1003 2983 1019
rect 1597 368 1611 402
rect 1645 368 1659 402
rect 1366 247 1400 344
rect 1597 330 1659 368
rect 1366 197 1400 213
rect 1463 291 1497 307
rect 1463 223 1497 257
rect 1155 153 1189 169
rect 995 119 1058 153
rect 1092 119 1155 153
rect 961 103 995 119
rect 1155 103 1189 119
rect 1269 153 1303 189
rect 1463 153 1497 189
rect 1303 119 1366 153
rect 1400 119 1463 153
rect 1269 103 1303 119
rect 1463 103 1497 119
rect 1597 296 1611 330
rect 1645 296 1659 330
rect 1597 258 1659 296
rect 1597 224 1611 258
rect 1645 224 1659 258
rect 1597 186 1659 224
rect 1597 152 1611 186
rect 1645 152 1659 186
rect 1597 114 1659 152
rect 1597 80 1611 114
rect 1645 80 1659 114
rect 1729 363 1763 379
rect 1923 363 1957 379
rect 2117 363 2151 379
rect 1763 329 1826 363
rect 1860 329 1923 363
rect 1957 329 2020 363
rect 2054 329 2117 363
rect 1729 291 1763 329
rect 1729 223 1763 257
rect 1923 291 1957 329
rect 2117 313 2151 329
rect 2231 363 2265 379
rect 2425 378 2459 575
rect 2795 609 2829 969
rect 2231 291 2265 329
rect 1729 153 1763 189
rect 1729 103 1763 119
rect 1826 238 1860 254
rect 1597 62 1659 80
rect 1826 62 1860 204
rect 1923 223 1957 257
rect 2021 244 2055 260
rect 2231 244 2265 257
rect 2055 223 2265 244
rect 2055 210 2231 223
rect 2021 194 2055 210
rect 1923 153 1957 189
rect 2328 344 2459 378
rect 2559 546 2621 572
rect 2559 512 2573 546
rect 2607 512 2621 546
rect 2559 474 2621 512
rect 2559 440 2573 474
rect 2607 440 2621 474
rect 2559 402 2621 440
rect 2795 461 2829 575
rect 2795 411 2829 427
rect 2943 979 2949 995
rect 2977 953 2983 969
rect 2943 461 2977 945
rect 2943 411 2977 427
rect 3091 831 3125 1069
rect 3225 1076 3239 1110
rect 3273 1076 3287 1110
rect 3225 1038 3287 1076
rect 3397 1412 3431 1492
rect 3397 1344 3431 1378
rect 3397 1276 3431 1310
rect 3397 1208 3431 1242
rect 3397 1139 3431 1174
rect 3397 1073 3431 1105
rect 3485 1412 3519 1450
rect 3485 1344 3519 1378
rect 3485 1276 3519 1310
rect 3485 1208 3519 1242
rect 3485 1139 3519 1174
rect 3573 1412 3607 1492
rect 3573 1344 3607 1378
rect 3573 1276 3607 1310
rect 3573 1208 3607 1242
rect 3573 1157 3607 1174
rect 3661 1412 3695 1450
rect 3661 1344 3695 1378
rect 3661 1276 3695 1310
rect 3661 1208 3695 1242
rect 3485 1103 3519 1105
rect 3661 1139 3695 1174
rect 3749 1412 3783 1492
rect 3749 1344 3783 1378
rect 3749 1276 3783 1310
rect 3749 1208 3783 1242
rect 3749 1157 3783 1174
rect 3891 1470 3953 1492
rect 3891 1436 3905 1470
rect 3939 1436 3953 1470
rect 3891 1398 3953 1436
rect 3891 1364 3905 1398
rect 3939 1364 3953 1398
rect 3891 1326 3953 1364
rect 3891 1292 3905 1326
rect 3939 1292 3953 1326
rect 3891 1254 3953 1292
rect 3891 1220 3905 1254
rect 3939 1220 3953 1254
rect 3891 1182 3953 1220
rect 3661 1103 3695 1105
rect 3891 1148 3905 1182
rect 3939 1148 3953 1182
rect 3891 1110 3953 1148
rect 3485 1069 3791 1103
rect 3225 1004 3239 1038
rect 3273 1004 3287 1038
rect 3225 966 3287 1004
rect 3225 932 3239 966
rect 3273 932 3287 966
rect 3225 868 3287 932
rect 3461 1003 3495 1019
rect 3615 1003 3649 1019
rect 3461 905 3495 969
rect 2559 368 2573 402
rect 2607 368 2621 402
rect 2328 247 2362 344
rect 2559 330 2621 368
rect 2328 197 2362 213
rect 2425 291 2459 307
rect 2425 223 2459 257
rect 2117 153 2151 169
rect 1957 119 2020 153
rect 2054 119 2117 153
rect 1923 103 1957 119
rect 2117 103 2151 119
rect 2231 153 2265 189
rect 2425 153 2459 189
rect 2265 119 2328 153
rect 2362 119 2425 153
rect 2231 103 2265 119
rect 2425 103 2459 119
rect 2559 296 2573 330
rect 2607 296 2621 330
rect 2559 258 2621 296
rect 2559 224 2573 258
rect 2607 224 2621 258
rect 2559 186 2621 224
rect 2559 152 2573 186
rect 2607 152 2621 186
rect 2559 114 2621 152
rect 2559 80 2573 114
rect 2607 80 2621 114
rect 2712 361 2746 377
rect 2906 361 2940 377
rect 3091 376 3125 797
rect 2746 327 2809 361
rect 2843 327 2906 361
rect 2712 289 2746 327
rect 2712 221 2746 255
rect 2906 289 2940 327
rect 2712 151 2746 187
rect 2712 101 2746 117
rect 2809 236 2843 252
rect 2559 62 2621 80
rect 2809 62 2843 202
rect 2906 221 2940 255
rect 3003 342 3125 376
rect 3225 546 3287 572
rect 3225 512 3239 546
rect 3273 512 3287 546
rect 3225 474 3287 512
rect 3225 440 3239 474
rect 3273 440 3287 474
rect 3225 402 3287 440
rect 3461 461 3495 871
rect 3461 411 3495 427
rect 3609 969 3615 988
rect 3609 953 3649 969
rect 3609 757 3643 953
rect 3609 461 3643 723
rect 3609 411 3643 427
rect 3757 683 3791 1069
rect 3891 1076 3905 1110
rect 3939 1076 3953 1110
rect 4123 1412 4157 1492
rect 4123 1344 4157 1378
rect 4123 1276 4157 1310
rect 4123 1208 4157 1242
rect 4123 1139 4157 1174
rect 4123 1089 4157 1105
rect 4211 1412 4245 1450
rect 4211 1344 4245 1378
rect 4211 1276 4245 1310
rect 4211 1208 4245 1242
rect 4211 1139 4245 1174
rect 4299 1412 4333 1492
rect 4299 1344 4333 1378
rect 4299 1276 4333 1310
rect 4299 1208 4333 1242
rect 4299 1157 4333 1174
rect 4387 1412 4421 1450
rect 4387 1344 4421 1378
rect 4387 1276 4421 1310
rect 4387 1208 4421 1242
rect 4211 1094 4245 1105
rect 4387 1139 4421 1174
rect 4475 1412 4509 1492
rect 4475 1344 4509 1378
rect 4475 1276 4509 1310
rect 4475 1208 4509 1242
rect 4475 1157 4509 1174
rect 4563 1412 4597 1450
rect 4563 1344 4597 1378
rect 4563 1276 4597 1310
rect 4563 1208 4597 1242
rect 4387 1094 4421 1105
rect 4563 1139 4597 1174
rect 4651 1412 4685 1492
rect 4651 1344 4685 1378
rect 4651 1276 4685 1310
rect 4651 1208 4685 1242
rect 4651 1157 4685 1174
rect 4853 1470 4915 1492
rect 4853 1436 4867 1470
rect 4901 1436 4915 1470
rect 4853 1398 4915 1436
rect 4853 1364 4867 1398
rect 4901 1364 4915 1398
rect 4853 1326 4915 1364
rect 4853 1292 4867 1326
rect 4901 1292 4915 1326
rect 4853 1254 4915 1292
rect 4853 1220 4867 1254
rect 4901 1220 4915 1254
rect 4853 1182 4915 1220
rect 4563 1094 4597 1105
rect 4853 1148 4867 1182
rect 4901 1148 4915 1182
rect 4853 1110 4915 1148
rect 3891 1038 3953 1076
rect 4211 1060 4753 1094
rect 3891 1004 3905 1038
rect 3939 1004 3953 1038
rect 3891 966 3953 1004
rect 3891 932 3905 966
rect 3939 932 3953 966
rect 3891 868 3953 932
rect 4127 1003 4161 1019
rect 3225 368 3239 402
rect 3273 368 3287 402
rect 3003 245 3037 342
rect 3225 330 3287 368
rect 3003 195 3037 211
rect 3100 289 3134 305
rect 3100 221 3134 255
rect 2906 151 2940 187
rect 3100 151 3134 187
rect 2940 117 3003 151
rect 3037 117 3100 151
rect 2906 101 2940 117
rect 3100 101 3134 117
rect 3225 296 3239 330
rect 3273 296 3287 330
rect 3225 258 3287 296
rect 3225 224 3239 258
rect 3273 224 3287 258
rect 3225 186 3287 224
rect 3225 152 3239 186
rect 3273 152 3287 186
rect 3225 114 3287 152
rect 3225 80 3239 114
rect 3273 80 3287 114
rect 3378 361 3412 377
rect 3572 361 3606 377
rect 3757 376 3791 649
rect 4127 683 4161 969
rect 3412 327 3475 361
rect 3509 327 3572 361
rect 3378 289 3412 327
rect 3378 221 3412 255
rect 3572 289 3606 327
rect 3378 151 3412 187
rect 3378 101 3412 117
rect 3475 236 3509 252
rect 3225 62 3287 80
rect 3475 62 3509 202
rect 3572 221 3606 255
rect 3669 342 3791 376
rect 3891 546 3953 572
rect 3891 512 3905 546
rect 3939 512 3953 546
rect 3891 474 3953 512
rect 3891 440 3905 474
rect 3939 440 3953 474
rect 3891 402 3953 440
rect 4127 461 4161 649
rect 4127 411 4161 427
rect 4349 1003 4383 1019
rect 4349 535 4383 969
rect 4349 461 4383 501
rect 4349 411 4383 427
rect 4571 1003 4605 1019
rect 4571 831 4605 969
rect 4571 461 4605 797
rect 4571 411 4605 427
rect 4719 757 4753 1060
rect 4853 1076 4867 1110
rect 4901 1076 4915 1110
rect 4853 1038 4915 1076
rect 4853 1004 4867 1038
rect 4901 1004 4915 1038
rect 4853 966 4915 1004
rect 4853 932 4867 966
rect 4901 932 4915 966
rect 4853 868 4915 932
rect 3891 368 3905 402
rect 3939 368 3953 402
rect 3669 245 3703 342
rect 3891 330 3953 368
rect 3669 195 3703 211
rect 3766 289 3800 305
rect 3766 221 3800 255
rect 3572 151 3606 187
rect 3766 151 3800 187
rect 3606 117 3669 151
rect 3703 117 3766 151
rect 3572 101 3606 117
rect 3766 101 3800 117
rect 3891 296 3905 330
rect 3939 296 3953 330
rect 3891 258 3953 296
rect 3891 224 3905 258
rect 3939 224 3953 258
rect 3891 186 3953 224
rect 3891 152 3905 186
rect 3939 152 3953 186
rect 3891 114 3953 152
rect 3891 80 3905 114
rect 3939 80 3953 114
rect 4023 363 4057 379
rect 4217 363 4251 379
rect 4411 363 4445 379
rect 4057 329 4120 363
rect 4154 329 4217 363
rect 4251 329 4314 363
rect 4348 329 4411 363
rect 4023 291 4057 329
rect 4023 223 4057 257
rect 4217 291 4251 329
rect 4411 313 4445 329
rect 4525 363 4559 379
rect 4719 378 4753 723
rect 4525 291 4559 329
rect 4023 153 4057 189
rect 4023 103 4057 119
rect 4120 238 4154 254
rect 3891 62 3953 80
rect 4120 62 4154 204
rect 4217 223 4251 257
rect 4315 244 4349 260
rect 4525 244 4559 257
rect 4349 223 4559 244
rect 4349 210 4525 223
rect 4315 194 4349 210
rect 4217 153 4251 189
rect 4622 344 4753 378
rect 4853 546 4915 572
rect 4853 512 4867 546
rect 4901 512 4915 546
rect 4853 474 4915 512
rect 4853 440 4867 474
rect 4901 440 4915 474
rect 4853 402 4915 440
rect 4853 368 4867 402
rect 4901 368 4915 402
rect 4622 247 4656 344
rect 4853 330 4915 368
rect 4622 197 4656 213
rect 4719 291 4753 307
rect 4719 223 4753 257
rect 4411 153 4445 169
rect 4251 119 4314 153
rect 4348 119 4411 153
rect 4217 103 4251 119
rect 4411 103 4445 119
rect 4525 153 4559 189
rect 4719 153 4753 189
rect 4559 119 4622 153
rect 4656 119 4719 153
rect 4525 103 4559 119
rect 4719 103 4753 119
rect 4853 296 4867 330
rect 4901 296 4915 330
rect 4853 258 4915 296
rect 4853 224 4867 258
rect 4901 224 4915 258
rect 4853 186 4915 224
rect 4853 152 4867 186
rect 4901 152 4915 186
rect 4853 114 4915 152
rect 4853 80 4867 114
rect 4901 80 4915 114
rect 4853 62 4915 80
rect -31 47 4915 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 361 47
rect 395 13 433 47
rect 467 13 505 47
rect 539 13 577 47
rect 611 13 721 47
rect 755 13 793 47
rect 827 13 865 47
rect 899 13 937 47
rect 971 13 1009 47
rect 1043 13 1081 47
rect 1115 13 1179 47
rect 1213 13 1251 47
rect 1285 13 1323 47
rect 1357 13 1395 47
rect 1429 13 1467 47
rect 1501 13 1539 47
rect 1573 13 1683 47
rect 1717 13 1755 47
rect 1789 13 1827 47
rect 1861 13 1899 47
rect 1933 13 1971 47
rect 2005 13 2043 47
rect 2077 13 2141 47
rect 2175 13 2213 47
rect 2247 13 2285 47
rect 2319 13 2357 47
rect 2391 13 2429 47
rect 2463 13 2501 47
rect 2535 13 2645 47
rect 2679 13 2717 47
rect 2751 13 2789 47
rect 2823 13 2861 47
rect 2895 13 2951 47
rect 2985 13 3023 47
rect 3057 13 3095 47
rect 3129 13 3167 47
rect 3201 13 3311 47
rect 3345 13 3383 47
rect 3417 13 3455 47
rect 3489 13 3527 47
rect 3561 13 3617 47
rect 3651 13 3689 47
rect 3723 13 3761 47
rect 3795 13 3833 47
rect 3867 13 3977 47
rect 4011 13 4049 47
rect 4083 13 4121 47
rect 4155 13 4193 47
rect 4227 13 4265 47
rect 4299 13 4337 47
rect 4371 13 4435 47
rect 4469 13 4507 47
rect 4541 13 4579 47
rect 4613 13 4651 47
rect 4685 13 4723 47
rect 4757 13 4795 47
rect 4829 13 4915 47
rect -31 0 4915 13
<< viali >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 361 1505 395 1539
rect 433 1505 467 1539
rect 505 1505 539 1539
rect 577 1505 611 1539
rect 721 1505 755 1539
rect 793 1505 827 1539
rect 865 1505 899 1539
rect 937 1505 971 1539
rect 1009 1505 1043 1539
rect 1081 1505 1115 1539
rect 1179 1505 1213 1539
rect 1251 1505 1285 1539
rect 1323 1505 1357 1539
rect 1395 1505 1429 1539
rect 1467 1505 1501 1539
rect 1539 1505 1573 1539
rect 1683 1505 1717 1539
rect 1755 1505 1789 1539
rect 1827 1505 1861 1539
rect 1899 1505 1933 1539
rect 1971 1505 2005 1539
rect 2043 1505 2077 1539
rect 2141 1505 2175 1539
rect 2213 1505 2247 1539
rect 2285 1505 2319 1539
rect 2357 1505 2391 1539
rect 2429 1505 2463 1539
rect 2501 1505 2535 1539
rect 2645 1505 2679 1539
rect 2717 1505 2751 1539
rect 2789 1505 2823 1539
rect 2861 1505 2895 1539
rect 2951 1505 2985 1539
rect 3023 1505 3057 1539
rect 3095 1505 3129 1539
rect 3167 1505 3201 1539
rect 3311 1505 3345 1539
rect 3383 1505 3417 1539
rect 3455 1505 3489 1539
rect 3527 1505 3561 1539
rect 3617 1505 3651 1539
rect 3689 1505 3723 1539
rect 3761 1505 3795 1539
rect 3833 1505 3867 1539
rect 3977 1505 4011 1539
rect 4049 1505 4083 1539
rect 4121 1505 4155 1539
rect 4193 1505 4227 1539
rect 4265 1505 4299 1539
rect 4337 1505 4371 1539
rect 4435 1505 4469 1539
rect 4507 1505 4541 1539
rect 4579 1505 4613 1539
rect 4651 1505 4685 1539
rect 4723 1505 4757 1539
rect 4795 1505 4829 1539
rect 205 797 239 831
rect 353 871 387 905
rect 501 575 535 609
rect 871 574 905 608
rect 1093 969 1127 979
rect 1093 945 1127 969
rect 1462 871 1496 905
rect 1315 797 1349 831
rect 1833 575 1867 609
rect 2055 501 2089 535
rect 2277 797 2311 831
rect 2425 575 2459 609
rect 2795 575 2829 609
rect 2943 969 2949 979
rect 2949 969 2977 979
rect 2943 945 2977 969
rect 3461 871 3495 905
rect 3091 797 3125 831
rect 3609 723 3643 757
rect 3757 649 3791 683
rect 4127 649 4161 683
rect 4349 501 4383 535
rect 4571 797 4605 831
rect 4719 723 4753 757
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 361 13 395 47
rect 433 13 467 47
rect 505 13 539 47
rect 577 13 611 47
rect 721 13 755 47
rect 793 13 827 47
rect 865 13 899 47
rect 937 13 971 47
rect 1009 13 1043 47
rect 1081 13 1115 47
rect 1179 13 1213 47
rect 1251 13 1285 47
rect 1323 13 1357 47
rect 1395 13 1429 47
rect 1467 13 1501 47
rect 1539 13 1573 47
rect 1683 13 1717 47
rect 1755 13 1789 47
rect 1827 13 1861 47
rect 1899 13 1933 47
rect 1971 13 2005 47
rect 2043 13 2077 47
rect 2141 13 2175 47
rect 2213 13 2247 47
rect 2285 13 2319 47
rect 2357 13 2391 47
rect 2429 13 2463 47
rect 2501 13 2535 47
rect 2645 13 2679 47
rect 2717 13 2751 47
rect 2789 13 2823 47
rect 2861 13 2895 47
rect 2951 13 2985 47
rect 3023 13 3057 47
rect 3095 13 3129 47
rect 3167 13 3201 47
rect 3311 13 3345 47
rect 3383 13 3417 47
rect 3455 13 3489 47
rect 3527 13 3561 47
rect 3617 13 3651 47
rect 3689 13 3723 47
rect 3761 13 3795 47
rect 3833 13 3867 47
rect 3977 13 4011 47
rect 4049 13 4083 47
rect 4121 13 4155 47
rect 4193 13 4227 47
rect 4265 13 4299 47
rect 4337 13 4371 47
rect 4435 13 4469 47
rect 4507 13 4541 47
rect 4579 13 4613 47
rect 4651 13 4685 47
rect 4723 13 4757 47
rect 4795 13 4829 47
<< metal1 >>
rect -31 1539 4915 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 361 1539
rect 395 1505 433 1539
rect 467 1505 505 1539
rect 539 1505 577 1539
rect 611 1505 721 1539
rect 755 1505 793 1539
rect 827 1505 865 1539
rect 899 1505 937 1539
rect 971 1505 1009 1539
rect 1043 1505 1081 1539
rect 1115 1505 1179 1539
rect 1213 1505 1251 1539
rect 1285 1505 1323 1539
rect 1357 1505 1395 1539
rect 1429 1505 1467 1539
rect 1501 1505 1539 1539
rect 1573 1505 1683 1539
rect 1717 1505 1755 1539
rect 1789 1505 1827 1539
rect 1861 1505 1899 1539
rect 1933 1505 1971 1539
rect 2005 1505 2043 1539
rect 2077 1505 2141 1539
rect 2175 1505 2213 1539
rect 2247 1505 2285 1539
rect 2319 1505 2357 1539
rect 2391 1505 2429 1539
rect 2463 1505 2501 1539
rect 2535 1505 2645 1539
rect 2679 1505 2717 1539
rect 2751 1505 2789 1539
rect 2823 1505 2861 1539
rect 2895 1505 2951 1539
rect 2985 1505 3023 1539
rect 3057 1505 3095 1539
rect 3129 1505 3167 1539
rect 3201 1505 3311 1539
rect 3345 1505 3383 1539
rect 3417 1505 3455 1539
rect 3489 1505 3527 1539
rect 3561 1505 3617 1539
rect 3651 1505 3689 1539
rect 3723 1505 3761 1539
rect 3795 1505 3833 1539
rect 3867 1505 3977 1539
rect 4011 1505 4049 1539
rect 4083 1505 4121 1539
rect 4155 1505 4193 1539
rect 4227 1505 4265 1539
rect 4299 1505 4337 1539
rect 4371 1505 4435 1539
rect 4469 1505 4507 1539
rect 4541 1505 4579 1539
rect 4613 1505 4651 1539
rect 4685 1505 4723 1539
rect 4757 1505 4795 1539
rect 4829 1505 4915 1539
rect -31 1492 4915 1505
rect 1087 979 1133 985
rect 2937 979 2983 985
rect 1081 945 1093 979
rect 1127 945 2943 979
rect 2977 945 2989 979
rect 1087 939 1133 945
rect 2937 939 2983 945
rect 347 905 393 911
rect 1456 905 1502 911
rect 3455 905 3501 911
rect 341 871 353 905
rect 387 871 1462 905
rect 1496 871 3461 905
rect 3495 871 3507 905
rect 347 865 393 871
rect 1456 865 1502 871
rect 3455 865 3501 871
rect 199 831 245 837
rect 1309 831 1355 837
rect 2271 831 2317 837
rect 3085 831 3131 837
rect 4565 831 4611 837
rect 169 797 205 831
rect 239 797 251 831
rect 1303 797 1315 831
rect 1349 797 2277 831
rect 2311 797 3091 831
rect 3125 797 4571 831
rect 4605 797 4617 831
rect 199 791 245 797
rect 1309 791 1355 797
rect 2271 791 2317 797
rect 3085 791 3131 797
rect 4565 791 4611 797
rect 3603 757 3649 763
rect 4713 757 4759 763
rect 3597 723 3609 757
rect 3643 723 4719 757
rect 4753 723 4765 757
rect 3603 717 3649 723
rect 4713 717 4759 723
rect 3751 683 3797 689
rect 4121 683 4167 689
rect 3745 649 3757 683
rect 3791 649 4127 683
rect 4161 649 4173 683
rect 3751 643 3797 649
rect 4121 643 4167 649
rect 495 609 541 615
rect 865 609 911 614
rect 1827 609 1873 615
rect 2419 609 2465 615
rect 2789 609 2835 615
rect 489 575 501 609
rect 535 608 1833 609
rect 535 575 871 608
rect 495 569 541 575
rect 859 574 871 575
rect 905 575 1833 608
rect 1867 575 1879 609
rect 2413 575 2425 609
rect 2459 575 2795 609
rect 2829 575 2841 609
rect 905 574 941 575
rect 865 568 911 574
rect 1827 569 1873 575
rect 2419 569 2465 575
rect 2789 569 2835 575
rect 2049 535 2095 541
rect 4343 535 4389 541
rect 2043 501 2055 535
rect 2089 501 4349 535
rect 4383 501 4395 535
rect 2049 495 2095 501
rect 4343 495 4389 501
rect -31 47 4915 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 361 47
rect 395 13 433 47
rect 467 13 505 47
rect 539 13 577 47
rect 611 13 721 47
rect 755 13 793 47
rect 827 13 865 47
rect 899 13 937 47
rect 971 13 1009 47
rect 1043 13 1081 47
rect 1115 13 1179 47
rect 1213 13 1251 47
rect 1285 13 1323 47
rect 1357 13 1395 47
rect 1429 13 1467 47
rect 1501 13 1539 47
rect 1573 13 1683 47
rect 1717 13 1755 47
rect 1789 13 1827 47
rect 1861 13 1899 47
rect 1933 13 1971 47
rect 2005 13 2043 47
rect 2077 13 2141 47
rect 2175 13 2213 47
rect 2247 13 2285 47
rect 2319 13 2357 47
rect 2391 13 2429 47
rect 2463 13 2501 47
rect 2535 13 2645 47
rect 2679 13 2717 47
rect 2751 13 2789 47
rect 2823 13 2861 47
rect 2895 13 2951 47
rect 2985 13 3023 47
rect 3057 13 3095 47
rect 3129 13 3167 47
rect 3201 13 3311 47
rect 3345 13 3383 47
rect 3417 13 3455 47
rect 3489 13 3527 47
rect 3561 13 3617 47
rect 3651 13 3689 47
rect 3723 13 3761 47
rect 3795 13 3833 47
rect 3867 13 3977 47
rect 4011 13 4049 47
rect 4083 13 4121 47
rect 4155 13 4193 47
rect 4227 13 4265 47
rect 4299 13 4337 47
rect 4371 13 4435 47
rect 4469 13 4507 47
rect 4541 13 4579 47
rect 4613 13 4651 47
rect 4685 13 4723 47
rect 4757 13 4795 47
rect 4829 13 4915 47
rect -31 0 4915 13
<< labels >>
rlabel metal1 4719 723 4753 757 1 Q
port 1 n
rlabel metal1 205 797 239 831 1 D
port 2 n
rlabel metal1 1093 945 1127 979 1 CLK
port 3 n
rlabel metal1 2055 501 2089 535 1 SN
port 4 n
rlabel metal1 55 1505 89 1539 1 VDD
port 5 n
rlabel metal1 55 13 89 47 1 VSS
port 6 n
rlabel space 205 461 239 969 1 dffsnx1_pcell_0/D
rlabel space 1081 945 2952 979 1 dffsnx1_pcell_0/CLK
rlabel space 2043 501 4381 535 1 dffsnx1_pcell_0/SN
rlabel space 4719 344 4753 1094 1 dffsnx1_pcell_0/Q
rlabel space 4127 461 4161 969 1 dffsnx1_pcell_0/QN
rlabel space 3757 342 3791 1103 1 dffsnx1_pcell_0/QN
rlabel space 3609 461 3643 969 1 dffsnx1_pcell_0/Q
<< end >>
