magic
tech sky130A
magscale 1 2
timestamp 1651077792
<< nwell >>
rect -84 832 7854 1575
<< nmos >>
rect 155 324 185 377
tri 185 324 201 340 sw
rect 155 294 261 324
tri 261 294 291 324 sw
rect 155 193 185 294
tri 185 278 201 294 nw
tri 245 278 261 294 ne
tri 185 193 201 209 sw
tri 245 193 261 209 se
rect 261 193 291 294
tri 155 163 185 193 ne
rect 185 163 261 193
tri 261 163 291 193 nw
rect 612 316 642 377
tri 642 316 658 332 sw
rect 806 324 836 377
tri 836 324 852 340 sw
rect 612 286 718 316
tri 718 286 748 316 sw
rect 806 294 912 324
tri 912 294 942 324 sw
rect 612 185 642 286
tri 642 270 658 286 nw
tri 702 270 718 286 ne
tri 642 185 658 201 sw
tri 702 185 718 201 se
rect 718 185 748 286
rect 806 193 836 294
tri 836 278 852 294 nw
tri 896 278 912 294 ne
tri 836 193 852 209 sw
tri 896 193 912 209 se
rect 912 193 942 294
tri 612 155 642 185 ne
rect 642 155 718 185
tri 718 155 748 185 nw
tri 806 163 836 193 ne
rect 836 163 912 193
tri 912 163 942 193 nw
rect 1278 316 1308 377
tri 1308 316 1324 332 sw
rect 1472 324 1502 377
tri 1502 324 1518 340 sw
rect 1278 286 1384 316
tri 1384 286 1414 316 sw
rect 1472 294 1578 324
tri 1578 294 1608 324 sw
rect 1278 185 1308 286
tri 1308 270 1324 286 nw
tri 1368 270 1384 286 ne
tri 1308 185 1324 201 sw
tri 1368 185 1384 201 se
rect 1384 185 1414 286
rect 1472 193 1502 294
tri 1502 278 1518 294 nw
tri 1562 278 1578 294 ne
tri 1502 193 1518 209 sw
tri 1562 193 1578 209 se
rect 1578 193 1608 294
tri 1278 155 1308 185 ne
rect 1308 155 1384 185
tri 1384 155 1414 185 nw
tri 1472 163 1502 193 ne
rect 1502 163 1578 193
tri 1578 163 1608 193 nw
tri 2019 324 2035 340 se
rect 2035 324 2065 377
tri 1929 294 1959 324 se
rect 1959 294 2065 324
rect 1929 193 1959 294
tri 1959 278 1975 294 nw
tri 2019 278 2035 294 ne
tri 1959 193 1975 209 sw
tri 2019 193 2035 209 se
rect 2035 193 2065 294
tri 1929 163 1959 193 ne
rect 1959 163 2035 193
tri 2035 163 2065 193 nw
rect 2375 324 2405 377
tri 2405 324 2421 340 sw
rect 2375 294 2481 324
tri 2481 294 2511 324 sw
rect 2375 193 2405 294
tri 2405 278 2421 294 nw
tri 2465 278 2481 294 ne
tri 2405 193 2421 209 sw
tri 2465 193 2481 209 se
rect 2481 193 2511 294
tri 2375 163 2405 193 ne
rect 2405 163 2481 193
tri 2481 163 2511 193 nw
rect 2832 316 2862 377
tri 2862 316 2878 332 sw
rect 3026 324 3056 377
tri 3056 324 3072 340 sw
rect 2832 286 2938 316
tri 2938 286 2968 316 sw
rect 3026 294 3132 324
tri 3132 294 3162 324 sw
rect 2832 185 2862 286
tri 2862 270 2878 286 nw
tri 2922 270 2938 286 ne
tri 2862 185 2878 201 sw
tri 2922 185 2938 201 se
rect 2938 185 2968 286
rect 3026 193 3056 294
tri 3056 278 3072 294 nw
tri 3116 278 3132 294 ne
tri 3056 193 3072 209 sw
tri 3116 193 3132 209 se
rect 3132 193 3162 294
tri 2832 155 2862 185 ne
rect 2862 155 2938 185
tri 2938 155 2968 185 nw
tri 3026 163 3056 193 ne
rect 3056 163 3132 193
tri 3132 163 3162 193 nw
rect 3498 316 3528 377
tri 3528 316 3544 332 sw
rect 3692 324 3722 377
tri 3722 324 3738 340 sw
rect 3498 286 3604 316
tri 3604 286 3634 316 sw
rect 3692 294 3798 324
tri 3798 294 3828 324 sw
rect 3498 185 3528 286
tri 3528 270 3544 286 nw
tri 3588 270 3604 286 ne
tri 3528 185 3544 201 sw
tri 3588 185 3604 201 se
rect 3604 185 3634 286
rect 3692 193 3722 294
tri 3722 278 3738 294 nw
tri 3782 278 3798 294 ne
tri 3722 193 3738 209 sw
tri 3782 193 3798 209 se
rect 3798 193 3828 294
tri 3498 155 3528 185 ne
rect 3528 155 3604 185
tri 3604 155 3634 185 nw
tri 3692 163 3722 193 ne
rect 3722 163 3798 193
tri 3798 163 3828 193 nw
tri 4239 324 4255 340 se
rect 4255 324 4285 377
tri 4149 294 4179 324 se
rect 4179 294 4285 324
rect 4149 193 4179 294
tri 4179 278 4195 294 nw
tri 4239 278 4255 294 ne
tri 4179 193 4195 209 sw
tri 4239 193 4255 209 se
rect 4255 193 4285 294
tri 4149 163 4179 193 ne
rect 4179 163 4255 193
tri 4255 163 4285 193 nw
rect 4608 316 4638 377
tri 4638 316 4654 332 sw
rect 4802 324 4832 377
tri 4832 324 4848 340 sw
rect 4608 286 4714 316
tri 4714 286 4744 316 sw
rect 4802 294 4908 324
tri 4908 294 4938 324 sw
rect 4608 185 4638 286
tri 4638 270 4654 286 nw
tri 4698 270 4714 286 ne
tri 4638 185 4654 201 sw
tri 4698 185 4714 201 se
rect 4714 185 4744 286
rect 4802 193 4832 294
tri 4832 278 4848 294 nw
tri 4892 278 4908 294 ne
tri 4832 193 4848 209 sw
tri 4892 193 4908 209 se
rect 4908 193 4938 294
tri 4608 155 4638 185 ne
rect 4638 155 4714 185
tri 4714 155 4744 185 nw
tri 4802 163 4832 193 ne
rect 4832 163 4908 193
tri 4908 163 4938 193 nw
rect 5261 324 5291 377
tri 5291 324 5307 340 sw
rect 5261 294 5367 324
tri 5367 294 5397 324 sw
rect 5261 193 5291 294
tri 5291 278 5307 294 nw
tri 5351 278 5367 294 ne
tri 5291 193 5307 209 sw
tri 5351 193 5367 209 se
rect 5367 193 5397 294
tri 5261 163 5291 193 ne
rect 5291 163 5367 193
tri 5367 163 5397 193 nw
rect 5718 316 5748 377
tri 5748 316 5764 332 sw
rect 5912 324 5942 377
tri 5942 324 5958 340 sw
rect 5718 286 5824 316
tri 5824 286 5854 316 sw
rect 5912 294 6018 324
tri 6018 294 6048 324 sw
rect 5718 185 5748 286
tri 5748 270 5764 286 nw
tri 5808 270 5824 286 ne
tri 5748 185 5764 201 sw
tri 5808 185 5824 201 se
rect 5824 185 5854 286
rect 5912 193 5942 294
tri 5942 278 5958 294 nw
tri 6002 278 6018 294 ne
tri 5942 193 5958 209 sw
tri 6002 193 6018 209 se
rect 6018 193 6048 294
tri 5718 155 5748 185 ne
rect 5748 155 5824 185
tri 5824 155 5854 185 nw
tri 5912 163 5942 193 ne
rect 5942 163 6018 193
tri 6018 163 6048 193 nw
rect 6371 324 6401 377
tri 6401 324 6417 340 sw
rect 6371 294 6477 324
tri 6477 294 6507 324 sw
rect 6371 193 6401 294
tri 6401 278 6417 294 nw
tri 6461 278 6477 294 ne
tri 6401 193 6417 209 sw
tri 6461 193 6477 209 se
rect 6477 193 6507 294
tri 6371 163 6401 193 ne
rect 6401 163 6477 193
tri 6477 163 6507 193 nw
rect 6828 324 6858 377
tri 6858 324 6874 340 sw
rect 7022 324 7052 377
tri 7052 324 7068 340 sw
rect 6828 294 6934 324
tri 6934 294 6964 324 sw
rect 6828 193 6858 294
tri 6858 278 6874 294 nw
tri 6918 278 6934 294 ne
tri 6858 193 6874 209 sw
tri 6918 193 6934 209 se
rect 6934 193 6964 294
rect 7022 294 7128 324
tri 7128 294 7158 324 sw
rect 7022 279 7053 294
tri 7053 279 7068 294 nw
tri 7112 279 7127 294 ne
rect 7127 279 7158 294
tri 6828 163 6858 193 ne
rect 6858 163 6934 193
tri 6934 163 6964 193 nw
rect 7022 193 7052 279
tri 7052 193 7068 209 sw
tri 7112 193 7128 209 se
rect 7128 193 7158 279
tri 7022 163 7052 193 ne
rect 7052 163 7128 193
tri 7128 163 7158 193 nw
rect 7481 324 7511 377
tri 7511 324 7527 340 sw
rect 7481 294 7587 324
tri 7587 294 7617 324 sw
rect 7481 193 7511 294
tri 7511 278 7527 294 nw
tri 7571 278 7587 294 ne
tri 7511 193 7527 209 sw
tri 7571 193 7587 209 se
rect 7587 193 7617 294
tri 7481 163 7511 193 ne
rect 7511 163 7587 193
tri 7587 163 7617 193 nw
<< pmos >>
rect 163 1050 193 1450
rect 251 1050 281 1450
rect 631 1051 661 1451
rect 719 1051 749 1451
rect 807 1051 837 1451
rect 895 1051 925 1451
rect 1297 1051 1327 1451
rect 1385 1051 1415 1451
rect 1473 1051 1503 1451
rect 1561 1051 1591 1451
rect 1939 1050 1969 1450
rect 2027 1050 2057 1450
rect 2383 1050 2413 1450
rect 2471 1050 2501 1450
rect 2851 1051 2881 1451
rect 2939 1051 2969 1451
rect 3027 1051 3057 1451
rect 3115 1051 3145 1451
rect 3517 1051 3547 1451
rect 3605 1051 3635 1451
rect 3693 1051 3723 1451
rect 3781 1051 3811 1451
rect 4159 1050 4189 1450
rect 4247 1050 4277 1450
rect 4627 1050 4657 1450
rect 4715 1050 4745 1450
rect 4803 1050 4833 1450
rect 4891 1050 4921 1450
rect 5269 1050 5299 1450
rect 5357 1050 5387 1450
rect 5737 1050 5767 1450
rect 5825 1050 5855 1450
rect 5913 1050 5943 1450
rect 6001 1050 6031 1450
rect 6379 1050 6409 1450
rect 6467 1050 6497 1450
rect 6847 1051 6877 1451
rect 6935 1051 6965 1451
rect 7023 1051 7053 1451
rect 7111 1051 7141 1451
rect 7489 1050 7519 1450
rect 7577 1050 7607 1450
<< ndiff >>
rect 99 361 155 377
rect 99 327 109 361
rect 143 327 155 361
rect 99 289 155 327
rect 185 361 345 377
rect 185 340 303 361
tri 185 324 201 340 ne
rect 201 327 303 340
rect 337 327 345 361
rect 201 324 345 327
tri 261 294 291 324 ne
rect 99 255 109 289
rect 143 255 155 289
rect 99 221 155 255
rect 99 187 109 221
rect 143 187 155 221
tri 185 278 201 294 se
rect 201 278 245 294
tri 245 278 261 294 sw
rect 185 245 261 278
rect 185 211 205 245
rect 239 211 261 245
rect 185 209 261 211
tri 185 193 201 209 ne
rect 201 193 245 209
tri 245 193 261 209 nw
rect 291 289 345 324
rect 291 255 303 289
rect 337 255 345 289
rect 291 221 345 255
rect 99 163 155 187
tri 155 163 185 193 sw
tri 261 163 291 193 se
rect 291 187 303 221
rect 337 187 345 221
rect 291 163 345 187
rect 99 151 345 163
rect 99 117 109 151
rect 143 117 205 151
rect 239 117 303 151
rect 337 117 345 151
rect 99 101 345 117
rect 556 361 612 377
rect 556 327 566 361
rect 600 327 612 361
rect 556 289 612 327
rect 642 361 806 377
rect 642 332 663 361
tri 642 316 658 332 ne
rect 658 327 663 332
rect 697 327 760 361
rect 794 327 806 361
rect 658 316 806 327
rect 836 340 998 377
tri 836 324 852 340 ne
rect 852 324 998 340
rect 556 255 566 289
rect 600 255 612 289
tri 718 286 748 316 ne
rect 748 289 806 316
tri 912 294 942 324 ne
rect 556 221 612 255
rect 556 187 566 221
rect 600 187 612 221
rect 556 155 612 187
tri 642 270 658 286 se
rect 658 270 702 286
tri 702 270 718 286 sw
rect 642 236 718 270
rect 642 202 663 236
rect 697 202 718 236
rect 642 201 718 202
tri 642 185 658 201 ne
rect 658 185 702 201
tri 702 185 718 201 nw
rect 748 255 760 289
rect 794 255 806 289
rect 748 221 806 255
rect 748 187 760 221
rect 794 187 806 221
tri 836 278 852 294 se
rect 852 278 896 294
tri 896 278 912 294 sw
rect 836 245 912 278
rect 836 211 857 245
rect 891 211 912 245
rect 836 209 912 211
tri 836 193 852 209 ne
rect 852 193 896 209
tri 896 193 912 209 nw
rect 942 289 998 324
rect 942 255 954 289
rect 988 255 998 289
rect 942 221 998 255
tri 612 155 642 185 sw
tri 718 155 748 185 se
rect 748 163 806 187
tri 806 163 836 193 sw
tri 912 163 942 193 se
rect 942 187 954 221
rect 988 187 998 221
rect 942 163 998 187
rect 748 155 998 163
rect 556 151 998 155
rect 556 117 566 151
rect 600 117 760 151
rect 794 117 857 151
rect 891 117 954 151
rect 988 117 998 151
rect 556 101 998 117
rect 1222 361 1278 377
rect 1222 327 1232 361
rect 1266 327 1278 361
rect 1222 289 1278 327
rect 1308 361 1472 377
rect 1308 332 1329 361
tri 1308 316 1324 332 ne
rect 1324 327 1329 332
rect 1363 327 1426 361
rect 1460 327 1472 361
rect 1324 316 1472 327
rect 1502 340 1664 377
tri 1502 324 1518 340 ne
rect 1518 324 1664 340
rect 1222 255 1232 289
rect 1266 255 1278 289
tri 1384 286 1414 316 ne
rect 1414 289 1472 316
tri 1578 294 1608 324 ne
rect 1222 221 1278 255
rect 1222 187 1232 221
rect 1266 187 1278 221
rect 1222 155 1278 187
tri 1308 270 1324 286 se
rect 1324 270 1368 286
tri 1368 270 1384 286 sw
rect 1308 236 1384 270
rect 1308 202 1329 236
rect 1363 202 1384 236
rect 1308 201 1384 202
tri 1308 185 1324 201 ne
rect 1324 185 1368 201
tri 1368 185 1384 201 nw
rect 1414 255 1426 289
rect 1460 255 1472 289
rect 1414 221 1472 255
rect 1414 187 1426 221
rect 1460 187 1472 221
tri 1502 278 1518 294 se
rect 1518 278 1562 294
tri 1562 278 1578 294 sw
rect 1502 245 1578 278
rect 1502 211 1523 245
rect 1557 211 1578 245
rect 1502 209 1578 211
tri 1502 193 1518 209 ne
rect 1518 193 1562 209
tri 1562 193 1578 209 nw
rect 1608 289 1664 324
rect 1608 255 1620 289
rect 1654 255 1664 289
rect 1608 221 1664 255
tri 1278 155 1308 185 sw
tri 1384 155 1414 185 se
rect 1414 163 1472 187
tri 1472 163 1502 193 sw
tri 1578 163 1608 193 se
rect 1608 187 1620 221
rect 1654 187 1664 221
rect 1608 163 1664 187
rect 1414 155 1664 163
rect 1222 151 1664 155
rect 1222 117 1232 151
rect 1266 117 1426 151
rect 1460 117 1523 151
rect 1557 117 1620 151
rect 1654 117 1664 151
rect 1222 101 1664 117
rect 1875 361 2035 377
rect 1875 327 1883 361
rect 1917 340 2035 361
rect 1917 327 2019 340
rect 1875 324 2019 327
tri 2019 324 2035 340 nw
rect 2065 361 2121 377
rect 2065 327 2077 361
rect 2111 327 2121 361
rect 1875 289 1929 324
tri 1929 294 1959 324 nw
rect 1875 255 1883 289
rect 1917 255 1929 289
rect 1875 221 1929 255
rect 1875 187 1883 221
rect 1917 187 1929 221
tri 1959 278 1975 294 se
rect 1975 278 2019 294
tri 2019 278 2035 294 sw
rect 1959 245 2035 278
rect 1959 211 1981 245
rect 2015 211 2035 245
rect 1959 209 2035 211
tri 1959 193 1975 209 ne
rect 1975 193 2019 209
tri 2019 193 2035 209 nw
rect 2065 289 2121 327
rect 2065 255 2077 289
rect 2111 255 2121 289
rect 2065 221 2121 255
rect 1875 163 1929 187
tri 1929 163 1959 193 sw
tri 2035 163 2065 193 se
rect 2065 187 2077 221
rect 2111 187 2121 221
rect 2065 163 2121 187
rect 1875 151 2121 163
rect 1875 117 1883 151
rect 1917 117 1981 151
rect 2015 117 2077 151
rect 2111 117 2121 151
rect 1875 101 2121 117
rect 2319 361 2375 377
rect 2319 327 2329 361
rect 2363 327 2375 361
rect 2319 289 2375 327
rect 2405 361 2565 377
rect 2405 340 2523 361
tri 2405 324 2421 340 ne
rect 2421 327 2523 340
rect 2557 327 2565 361
rect 2421 324 2565 327
tri 2481 294 2511 324 ne
rect 2319 255 2329 289
rect 2363 255 2375 289
rect 2319 221 2375 255
rect 2319 187 2329 221
rect 2363 187 2375 221
tri 2405 278 2421 294 se
rect 2421 278 2465 294
tri 2465 278 2481 294 sw
rect 2405 245 2481 278
rect 2405 211 2425 245
rect 2459 211 2481 245
rect 2405 209 2481 211
tri 2405 193 2421 209 ne
rect 2421 193 2465 209
tri 2465 193 2481 209 nw
rect 2511 289 2565 324
rect 2511 255 2523 289
rect 2557 255 2565 289
rect 2511 221 2565 255
rect 2319 163 2375 187
tri 2375 163 2405 193 sw
tri 2481 163 2511 193 se
rect 2511 187 2523 221
rect 2557 187 2565 221
rect 2511 163 2565 187
rect 2319 151 2565 163
rect 2319 117 2329 151
rect 2363 117 2425 151
rect 2459 117 2523 151
rect 2557 117 2565 151
rect 2319 101 2565 117
rect 2776 361 2832 377
rect 2776 327 2786 361
rect 2820 327 2832 361
rect 2776 289 2832 327
rect 2862 361 3026 377
rect 2862 332 2883 361
tri 2862 316 2878 332 ne
rect 2878 327 2883 332
rect 2917 327 2980 361
rect 3014 327 3026 361
rect 2878 316 3026 327
rect 3056 340 3218 377
tri 3056 324 3072 340 ne
rect 3072 324 3218 340
rect 2776 255 2786 289
rect 2820 255 2832 289
tri 2938 286 2968 316 ne
rect 2968 289 3026 316
tri 3132 294 3162 324 ne
rect 2776 221 2832 255
rect 2776 187 2786 221
rect 2820 187 2832 221
rect 2776 155 2832 187
tri 2862 270 2878 286 se
rect 2878 270 2922 286
tri 2922 270 2938 286 sw
rect 2862 236 2938 270
rect 2862 202 2883 236
rect 2917 202 2938 236
rect 2862 201 2938 202
tri 2862 185 2878 201 ne
rect 2878 185 2922 201
tri 2922 185 2938 201 nw
rect 2968 255 2980 289
rect 3014 255 3026 289
rect 2968 221 3026 255
rect 2968 187 2980 221
rect 3014 187 3026 221
tri 3056 278 3072 294 se
rect 3072 278 3116 294
tri 3116 278 3132 294 sw
rect 3056 245 3132 278
rect 3056 211 3077 245
rect 3111 211 3132 245
rect 3056 209 3132 211
tri 3056 193 3072 209 ne
rect 3072 193 3116 209
tri 3116 193 3132 209 nw
rect 3162 289 3218 324
rect 3162 255 3174 289
rect 3208 255 3218 289
rect 3162 221 3218 255
tri 2832 155 2862 185 sw
tri 2938 155 2968 185 se
rect 2968 163 3026 187
tri 3026 163 3056 193 sw
tri 3132 163 3162 193 se
rect 3162 187 3174 221
rect 3208 187 3218 221
rect 3162 163 3218 187
rect 2968 155 3218 163
rect 2776 151 3218 155
rect 2776 117 2786 151
rect 2820 117 2980 151
rect 3014 117 3077 151
rect 3111 117 3174 151
rect 3208 117 3218 151
rect 2776 101 3218 117
rect 3442 361 3498 377
rect 3442 327 3452 361
rect 3486 327 3498 361
rect 3442 289 3498 327
rect 3528 361 3692 377
rect 3528 332 3549 361
tri 3528 316 3544 332 ne
rect 3544 327 3549 332
rect 3583 327 3646 361
rect 3680 327 3692 361
rect 3544 316 3692 327
rect 3722 340 3884 377
tri 3722 324 3738 340 ne
rect 3738 324 3884 340
rect 3442 255 3452 289
rect 3486 255 3498 289
tri 3604 286 3634 316 ne
rect 3634 289 3692 316
tri 3798 294 3828 324 ne
rect 3442 221 3498 255
rect 3442 187 3452 221
rect 3486 187 3498 221
rect 3442 155 3498 187
tri 3528 270 3544 286 se
rect 3544 270 3588 286
tri 3588 270 3604 286 sw
rect 3528 236 3604 270
rect 3528 202 3549 236
rect 3583 202 3604 236
rect 3528 201 3604 202
tri 3528 185 3544 201 ne
rect 3544 185 3588 201
tri 3588 185 3604 201 nw
rect 3634 255 3646 289
rect 3680 255 3692 289
rect 3634 221 3692 255
rect 3634 187 3646 221
rect 3680 187 3692 221
tri 3722 278 3738 294 se
rect 3738 278 3782 294
tri 3782 278 3798 294 sw
rect 3722 245 3798 278
rect 3722 211 3743 245
rect 3777 211 3798 245
rect 3722 209 3798 211
tri 3722 193 3738 209 ne
rect 3738 193 3782 209
tri 3782 193 3798 209 nw
rect 3828 289 3884 324
rect 3828 255 3840 289
rect 3874 255 3884 289
rect 3828 221 3884 255
tri 3498 155 3528 185 sw
tri 3604 155 3634 185 se
rect 3634 163 3692 187
tri 3692 163 3722 193 sw
tri 3798 163 3828 193 se
rect 3828 187 3840 221
rect 3874 187 3884 221
rect 3828 163 3884 187
rect 3634 155 3884 163
rect 3442 151 3884 155
rect 3442 117 3452 151
rect 3486 117 3646 151
rect 3680 117 3743 151
rect 3777 117 3840 151
rect 3874 117 3884 151
rect 3442 101 3884 117
rect 4095 361 4255 377
rect 4095 327 4103 361
rect 4137 340 4255 361
rect 4137 327 4239 340
rect 4095 324 4239 327
tri 4239 324 4255 340 nw
rect 4285 361 4341 377
rect 4285 327 4297 361
rect 4331 327 4341 361
rect 4095 289 4149 324
tri 4149 294 4179 324 nw
rect 4095 255 4103 289
rect 4137 255 4149 289
rect 4095 221 4149 255
rect 4095 187 4103 221
rect 4137 187 4149 221
tri 4179 278 4195 294 se
rect 4195 278 4239 294
tri 4239 278 4255 294 sw
rect 4179 245 4255 278
rect 4179 211 4201 245
rect 4235 211 4255 245
rect 4179 209 4255 211
tri 4179 193 4195 209 ne
rect 4195 193 4239 209
tri 4239 193 4255 209 nw
rect 4285 289 4341 327
rect 4285 255 4297 289
rect 4331 255 4341 289
rect 4285 221 4341 255
rect 4095 163 4149 187
tri 4149 163 4179 193 sw
tri 4255 163 4285 193 se
rect 4285 187 4297 221
rect 4331 187 4341 221
rect 4285 163 4341 187
rect 4095 151 4341 163
rect 4095 117 4103 151
rect 4137 117 4201 151
rect 4235 117 4297 151
rect 4331 117 4341 151
rect 4095 101 4341 117
rect 4552 361 4608 377
rect 4552 327 4562 361
rect 4596 327 4608 361
rect 4552 289 4608 327
rect 4638 361 4802 377
rect 4638 332 4659 361
tri 4638 316 4654 332 ne
rect 4654 327 4659 332
rect 4693 327 4756 361
rect 4790 327 4802 361
rect 4654 316 4802 327
rect 4832 340 4994 377
tri 4832 324 4848 340 ne
rect 4848 324 4994 340
rect 4552 255 4562 289
rect 4596 255 4608 289
tri 4714 286 4744 316 ne
rect 4744 289 4802 316
tri 4908 294 4938 324 ne
rect 4552 221 4608 255
rect 4552 187 4562 221
rect 4596 187 4608 221
rect 4552 155 4608 187
tri 4638 270 4654 286 se
rect 4654 270 4698 286
tri 4698 270 4714 286 sw
rect 4638 236 4714 270
rect 4638 202 4659 236
rect 4693 202 4714 236
rect 4638 201 4714 202
tri 4638 185 4654 201 ne
rect 4654 185 4698 201
tri 4698 185 4714 201 nw
rect 4744 255 4756 289
rect 4790 255 4802 289
rect 4744 221 4802 255
rect 4744 187 4756 221
rect 4790 187 4802 221
tri 4832 278 4848 294 se
rect 4848 278 4892 294
tri 4892 278 4908 294 sw
rect 4832 245 4908 278
rect 4832 211 4853 245
rect 4887 211 4908 245
rect 4832 209 4908 211
tri 4832 193 4848 209 ne
rect 4848 193 4892 209
tri 4892 193 4908 209 nw
rect 4938 289 4994 324
rect 4938 255 4950 289
rect 4984 255 4994 289
rect 4938 221 4994 255
tri 4608 155 4638 185 sw
tri 4714 155 4744 185 se
rect 4744 163 4802 187
tri 4802 163 4832 193 sw
tri 4908 163 4938 193 se
rect 4938 187 4950 221
rect 4984 187 4994 221
rect 4938 163 4994 187
rect 4744 155 4994 163
rect 4552 151 4994 155
rect 4552 117 4562 151
rect 4596 117 4756 151
rect 4790 117 4853 151
rect 4887 117 4950 151
rect 4984 117 4994 151
rect 4552 101 4994 117
rect 5205 361 5261 377
rect 5205 327 5215 361
rect 5249 327 5261 361
rect 5205 289 5261 327
rect 5291 361 5451 377
rect 5291 340 5409 361
tri 5291 324 5307 340 ne
rect 5307 327 5409 340
rect 5443 327 5451 361
rect 5307 324 5451 327
tri 5367 294 5397 324 ne
rect 5205 255 5215 289
rect 5249 255 5261 289
rect 5205 221 5261 255
rect 5205 187 5215 221
rect 5249 187 5261 221
tri 5291 278 5307 294 se
rect 5307 278 5351 294
tri 5351 278 5367 294 sw
rect 5291 245 5367 278
rect 5291 211 5311 245
rect 5345 211 5367 245
rect 5291 209 5367 211
tri 5291 193 5307 209 ne
rect 5307 193 5351 209
tri 5351 193 5367 209 nw
rect 5397 289 5451 324
rect 5397 255 5409 289
rect 5443 255 5451 289
rect 5397 221 5451 255
rect 5205 163 5261 187
tri 5261 163 5291 193 sw
tri 5367 163 5397 193 se
rect 5397 187 5409 221
rect 5443 187 5451 221
rect 5397 163 5451 187
rect 5205 151 5451 163
rect 5205 117 5215 151
rect 5249 117 5311 151
rect 5345 117 5409 151
rect 5443 117 5451 151
rect 5205 101 5451 117
rect 5662 361 5718 377
rect 5662 327 5672 361
rect 5706 327 5718 361
rect 5662 289 5718 327
rect 5748 361 5912 377
rect 5748 332 5769 361
tri 5748 316 5764 332 ne
rect 5764 327 5769 332
rect 5803 327 5866 361
rect 5900 327 5912 361
rect 5764 316 5912 327
rect 5942 340 6104 377
tri 5942 324 5958 340 ne
rect 5958 324 6104 340
rect 5662 255 5672 289
rect 5706 255 5718 289
tri 5824 286 5854 316 ne
rect 5854 289 5912 316
tri 6018 294 6048 324 ne
rect 5662 221 5718 255
rect 5662 187 5672 221
rect 5706 187 5718 221
rect 5662 155 5718 187
tri 5748 270 5764 286 se
rect 5764 270 5808 286
tri 5808 270 5824 286 sw
rect 5748 236 5824 270
rect 5748 202 5769 236
rect 5803 202 5824 236
rect 5748 201 5824 202
tri 5748 185 5764 201 ne
rect 5764 185 5808 201
tri 5808 185 5824 201 nw
rect 5854 255 5866 289
rect 5900 255 5912 289
rect 5854 221 5912 255
rect 5854 187 5866 221
rect 5900 187 5912 221
tri 5942 278 5958 294 se
rect 5958 278 6002 294
tri 6002 278 6018 294 sw
rect 5942 245 6018 278
rect 5942 211 5963 245
rect 5997 211 6018 245
rect 5942 209 6018 211
tri 5942 193 5958 209 ne
rect 5958 193 6002 209
tri 6002 193 6018 209 nw
rect 6048 289 6104 324
rect 6048 255 6060 289
rect 6094 255 6104 289
rect 6048 221 6104 255
tri 5718 155 5748 185 sw
tri 5824 155 5854 185 se
rect 5854 163 5912 187
tri 5912 163 5942 193 sw
tri 6018 163 6048 193 se
rect 6048 187 6060 221
rect 6094 187 6104 221
rect 6048 163 6104 187
rect 5854 155 6104 163
rect 5662 151 6104 155
rect 5662 117 5672 151
rect 5706 117 5866 151
rect 5900 117 5963 151
rect 5997 117 6060 151
rect 6094 117 6104 151
rect 5662 101 6104 117
rect 6315 361 6371 377
rect 6315 327 6325 361
rect 6359 327 6371 361
rect 6315 289 6371 327
rect 6401 361 6561 377
rect 6401 340 6519 361
tri 6401 324 6417 340 ne
rect 6417 327 6519 340
rect 6553 327 6561 361
rect 6417 324 6561 327
tri 6477 294 6507 324 ne
rect 6315 255 6325 289
rect 6359 255 6371 289
rect 6315 221 6371 255
rect 6315 187 6325 221
rect 6359 187 6371 221
tri 6401 278 6417 294 se
rect 6417 278 6461 294
tri 6461 278 6477 294 sw
rect 6401 245 6477 278
rect 6401 211 6421 245
rect 6455 211 6477 245
rect 6401 209 6477 211
tri 6401 193 6417 209 ne
rect 6417 193 6461 209
tri 6461 193 6477 209 nw
rect 6507 289 6561 324
rect 6507 255 6519 289
rect 6553 255 6561 289
rect 6507 221 6561 255
rect 6315 163 6371 187
tri 6371 163 6401 193 sw
tri 6477 163 6507 193 se
rect 6507 187 6519 221
rect 6553 187 6561 221
rect 6507 163 6561 187
rect 6315 151 6561 163
rect 6315 117 6325 151
rect 6359 117 6421 151
rect 6455 117 6519 151
rect 6553 117 6561 151
rect 6315 101 6561 117
rect 6772 361 6828 377
rect 6772 327 6782 361
rect 6816 327 6828 361
rect 6772 289 6828 327
rect 6858 340 7022 377
tri 6858 324 6874 340 ne
rect 6874 324 7022 340
rect 7052 340 7214 377
tri 7052 324 7068 340 ne
rect 7068 324 7214 340
tri 6934 294 6964 324 ne
rect 6772 255 6782 289
rect 6816 255 6828 289
rect 6772 221 6828 255
rect 6772 187 6782 221
rect 6816 187 6828 221
tri 6858 278 6874 294 se
rect 6874 278 6918 294
tri 6918 278 6934 294 sw
rect 6858 245 6934 278
rect 6858 211 6879 245
rect 6913 211 6934 245
rect 6858 209 6934 211
tri 6858 193 6874 209 ne
rect 6874 193 6918 209
tri 6918 193 6934 209 nw
rect 6964 289 7022 324
tri 7128 294 7158 324 ne
rect 6964 255 6976 289
rect 7010 255 7022 289
tri 7053 279 7068 294 se
rect 7068 279 7112 294
tri 7112 279 7127 294 sw
rect 7158 289 7214 324
rect 6964 221 7022 255
rect 6772 163 6828 187
tri 6828 163 6858 193 sw
tri 6934 163 6964 193 se
rect 6964 187 6976 221
rect 7010 187 7022 221
rect 7052 245 7128 279
rect 7052 211 7073 245
rect 7107 211 7128 245
rect 7052 209 7128 211
tri 7052 193 7068 209 ne
rect 7068 193 7112 209
tri 7112 193 7128 209 nw
rect 7158 255 7170 289
rect 7204 255 7214 289
rect 7158 221 7214 255
rect 6964 163 7022 187
tri 7022 163 7052 193 sw
tri 7128 163 7158 193 se
rect 7158 187 7170 221
rect 7204 187 7214 221
rect 7158 163 7214 187
rect 6772 151 7214 163
rect 6772 117 6782 151
rect 6816 117 6879 151
rect 6913 117 6976 151
rect 7010 117 7073 151
rect 7107 117 7170 151
rect 7204 117 7214 151
rect 6772 101 7214 117
rect 7425 361 7481 377
rect 7425 327 7435 361
rect 7469 327 7481 361
rect 7425 289 7481 327
rect 7511 361 7671 377
rect 7511 340 7629 361
tri 7511 324 7527 340 ne
rect 7527 327 7629 340
rect 7663 327 7671 361
rect 7527 324 7671 327
tri 7587 294 7617 324 ne
rect 7425 255 7435 289
rect 7469 255 7481 289
rect 7425 221 7481 255
rect 7425 187 7435 221
rect 7469 187 7481 221
tri 7511 278 7527 294 se
rect 7527 278 7571 294
tri 7571 278 7587 294 sw
rect 7511 245 7587 278
rect 7511 211 7531 245
rect 7565 211 7587 245
rect 7511 209 7587 211
tri 7511 193 7527 209 ne
rect 7527 193 7571 209
tri 7571 193 7587 209 nw
rect 7617 289 7671 324
rect 7617 255 7629 289
rect 7663 255 7671 289
rect 7617 221 7671 255
rect 7425 163 7481 187
tri 7481 163 7511 193 sw
tri 7587 163 7617 193 se
rect 7617 187 7629 221
rect 7663 187 7671 221
rect 7617 163 7671 187
rect 7425 151 7671 163
rect 7425 117 7435 151
rect 7469 117 7531 151
rect 7565 117 7629 151
rect 7663 117 7671 151
rect 7425 101 7671 117
<< pdiff >>
rect 107 1412 163 1450
rect 107 1378 117 1412
rect 151 1378 163 1412
rect 107 1344 163 1378
rect 107 1310 117 1344
rect 151 1310 163 1344
rect 107 1276 163 1310
rect 107 1242 117 1276
rect 151 1242 163 1276
rect 107 1208 163 1242
rect 107 1174 117 1208
rect 151 1174 163 1208
rect 107 1139 163 1174
rect 107 1105 117 1139
rect 151 1105 163 1139
rect 107 1050 163 1105
rect 193 1412 251 1450
rect 193 1378 205 1412
rect 239 1378 251 1412
rect 193 1344 251 1378
rect 193 1310 205 1344
rect 239 1310 251 1344
rect 193 1276 251 1310
rect 193 1242 205 1276
rect 239 1242 251 1276
rect 193 1208 251 1242
rect 193 1174 205 1208
rect 239 1174 251 1208
rect 193 1139 251 1174
rect 193 1105 205 1139
rect 239 1105 251 1139
rect 193 1050 251 1105
rect 281 1412 335 1450
rect 281 1378 293 1412
rect 327 1378 335 1412
rect 281 1344 335 1378
rect 281 1310 293 1344
rect 327 1310 335 1344
rect 281 1276 335 1310
rect 281 1242 293 1276
rect 327 1242 335 1276
rect 281 1208 335 1242
rect 281 1174 293 1208
rect 327 1174 335 1208
rect 281 1139 335 1174
rect 281 1105 293 1139
rect 327 1105 335 1139
rect 281 1050 335 1105
rect 575 1411 631 1451
rect 575 1377 585 1411
rect 619 1377 631 1411
rect 575 1343 631 1377
rect 575 1309 585 1343
rect 619 1309 631 1343
rect 575 1275 631 1309
rect 575 1241 585 1275
rect 619 1241 631 1275
rect 575 1207 631 1241
rect 575 1173 585 1207
rect 619 1173 631 1207
rect 575 1139 631 1173
rect 575 1105 585 1139
rect 619 1105 631 1139
rect 575 1051 631 1105
rect 661 1343 719 1451
rect 661 1309 673 1343
rect 707 1309 719 1343
rect 661 1275 719 1309
rect 661 1241 673 1275
rect 707 1241 719 1275
rect 661 1207 719 1241
rect 661 1173 673 1207
rect 707 1173 719 1207
rect 661 1051 719 1173
rect 749 1411 807 1451
rect 749 1377 761 1411
rect 795 1377 807 1411
rect 749 1343 807 1377
rect 749 1309 761 1343
rect 795 1309 807 1343
rect 749 1275 807 1309
rect 749 1241 761 1275
rect 795 1241 807 1275
rect 749 1207 807 1241
rect 749 1173 761 1207
rect 795 1173 807 1207
rect 749 1139 807 1173
rect 749 1105 761 1139
rect 795 1105 807 1139
rect 749 1051 807 1105
rect 837 1343 895 1451
rect 837 1309 849 1343
rect 883 1309 895 1343
rect 837 1275 895 1309
rect 837 1241 849 1275
rect 883 1241 895 1275
rect 837 1207 895 1241
rect 837 1173 849 1207
rect 883 1173 895 1207
rect 837 1139 895 1173
rect 837 1105 849 1139
rect 883 1105 895 1139
rect 837 1051 895 1105
rect 925 1411 979 1451
rect 925 1377 937 1411
rect 971 1377 979 1411
rect 925 1343 979 1377
rect 925 1309 937 1343
rect 971 1309 979 1343
rect 925 1275 979 1309
rect 925 1241 937 1275
rect 971 1241 979 1275
rect 925 1207 979 1241
rect 925 1173 937 1207
rect 971 1173 979 1207
rect 925 1051 979 1173
rect 1241 1411 1297 1451
rect 1241 1377 1251 1411
rect 1285 1377 1297 1411
rect 1241 1343 1297 1377
rect 1241 1309 1251 1343
rect 1285 1309 1297 1343
rect 1241 1275 1297 1309
rect 1241 1241 1251 1275
rect 1285 1241 1297 1275
rect 1241 1207 1297 1241
rect 1241 1173 1251 1207
rect 1285 1173 1297 1207
rect 1241 1139 1297 1173
rect 1241 1105 1251 1139
rect 1285 1105 1297 1139
rect 1241 1051 1297 1105
rect 1327 1343 1385 1451
rect 1327 1309 1339 1343
rect 1373 1309 1385 1343
rect 1327 1275 1385 1309
rect 1327 1241 1339 1275
rect 1373 1241 1385 1275
rect 1327 1207 1385 1241
rect 1327 1173 1339 1207
rect 1373 1173 1385 1207
rect 1327 1051 1385 1173
rect 1415 1411 1473 1451
rect 1415 1377 1427 1411
rect 1461 1377 1473 1411
rect 1415 1343 1473 1377
rect 1415 1309 1427 1343
rect 1461 1309 1473 1343
rect 1415 1275 1473 1309
rect 1415 1241 1427 1275
rect 1461 1241 1473 1275
rect 1415 1207 1473 1241
rect 1415 1173 1427 1207
rect 1461 1173 1473 1207
rect 1415 1139 1473 1173
rect 1415 1105 1427 1139
rect 1461 1105 1473 1139
rect 1415 1051 1473 1105
rect 1503 1343 1561 1451
rect 1503 1309 1515 1343
rect 1549 1309 1561 1343
rect 1503 1275 1561 1309
rect 1503 1241 1515 1275
rect 1549 1241 1561 1275
rect 1503 1207 1561 1241
rect 1503 1173 1515 1207
rect 1549 1173 1561 1207
rect 1503 1139 1561 1173
rect 1503 1105 1515 1139
rect 1549 1105 1561 1139
rect 1503 1051 1561 1105
rect 1591 1411 1645 1451
rect 1591 1377 1603 1411
rect 1637 1377 1645 1411
rect 1591 1343 1645 1377
rect 1591 1309 1603 1343
rect 1637 1309 1645 1343
rect 1591 1275 1645 1309
rect 1591 1241 1603 1275
rect 1637 1241 1645 1275
rect 1591 1207 1645 1241
rect 1591 1173 1603 1207
rect 1637 1173 1645 1207
rect 1591 1051 1645 1173
rect 1885 1412 1939 1450
rect 1885 1378 1893 1412
rect 1927 1378 1939 1412
rect 1885 1344 1939 1378
rect 1885 1310 1893 1344
rect 1927 1310 1939 1344
rect 1885 1276 1939 1310
rect 1885 1242 1893 1276
rect 1927 1242 1939 1276
rect 1885 1208 1939 1242
rect 1885 1174 1893 1208
rect 1927 1174 1939 1208
rect 1885 1139 1939 1174
rect 1885 1105 1893 1139
rect 1927 1105 1939 1139
rect 1885 1050 1939 1105
rect 1969 1412 2027 1450
rect 1969 1378 1981 1412
rect 2015 1378 2027 1412
rect 1969 1344 2027 1378
rect 1969 1310 1981 1344
rect 2015 1310 2027 1344
rect 1969 1276 2027 1310
rect 1969 1242 1981 1276
rect 2015 1242 2027 1276
rect 1969 1208 2027 1242
rect 1969 1174 1981 1208
rect 2015 1174 2027 1208
rect 1969 1139 2027 1174
rect 1969 1105 1981 1139
rect 2015 1105 2027 1139
rect 1969 1050 2027 1105
rect 2057 1412 2113 1450
rect 2057 1378 2069 1412
rect 2103 1378 2113 1412
rect 2057 1344 2113 1378
rect 2057 1310 2069 1344
rect 2103 1310 2113 1344
rect 2057 1276 2113 1310
rect 2057 1242 2069 1276
rect 2103 1242 2113 1276
rect 2057 1208 2113 1242
rect 2057 1174 2069 1208
rect 2103 1174 2113 1208
rect 2057 1139 2113 1174
rect 2057 1105 2069 1139
rect 2103 1105 2113 1139
rect 2057 1050 2113 1105
rect 2327 1412 2383 1450
rect 2327 1378 2337 1412
rect 2371 1378 2383 1412
rect 2327 1344 2383 1378
rect 2327 1310 2337 1344
rect 2371 1310 2383 1344
rect 2327 1276 2383 1310
rect 2327 1242 2337 1276
rect 2371 1242 2383 1276
rect 2327 1208 2383 1242
rect 2327 1174 2337 1208
rect 2371 1174 2383 1208
rect 2327 1139 2383 1174
rect 2327 1105 2337 1139
rect 2371 1105 2383 1139
rect 2327 1050 2383 1105
rect 2413 1412 2471 1450
rect 2413 1378 2425 1412
rect 2459 1378 2471 1412
rect 2413 1344 2471 1378
rect 2413 1310 2425 1344
rect 2459 1310 2471 1344
rect 2413 1276 2471 1310
rect 2413 1242 2425 1276
rect 2459 1242 2471 1276
rect 2413 1208 2471 1242
rect 2413 1174 2425 1208
rect 2459 1174 2471 1208
rect 2413 1139 2471 1174
rect 2413 1105 2425 1139
rect 2459 1105 2471 1139
rect 2413 1050 2471 1105
rect 2501 1412 2555 1450
rect 2501 1378 2513 1412
rect 2547 1378 2555 1412
rect 2501 1344 2555 1378
rect 2501 1310 2513 1344
rect 2547 1310 2555 1344
rect 2501 1276 2555 1310
rect 2501 1242 2513 1276
rect 2547 1242 2555 1276
rect 2501 1208 2555 1242
rect 2501 1174 2513 1208
rect 2547 1174 2555 1208
rect 2501 1139 2555 1174
rect 2501 1105 2513 1139
rect 2547 1105 2555 1139
rect 2501 1050 2555 1105
rect 2795 1411 2851 1451
rect 2795 1377 2805 1411
rect 2839 1377 2851 1411
rect 2795 1343 2851 1377
rect 2795 1309 2805 1343
rect 2839 1309 2851 1343
rect 2795 1275 2851 1309
rect 2795 1241 2805 1275
rect 2839 1241 2851 1275
rect 2795 1207 2851 1241
rect 2795 1173 2805 1207
rect 2839 1173 2851 1207
rect 2795 1139 2851 1173
rect 2795 1105 2805 1139
rect 2839 1105 2851 1139
rect 2795 1051 2851 1105
rect 2881 1343 2939 1451
rect 2881 1309 2893 1343
rect 2927 1309 2939 1343
rect 2881 1275 2939 1309
rect 2881 1241 2893 1275
rect 2927 1241 2939 1275
rect 2881 1207 2939 1241
rect 2881 1173 2893 1207
rect 2927 1173 2939 1207
rect 2881 1051 2939 1173
rect 2969 1411 3027 1451
rect 2969 1377 2981 1411
rect 3015 1377 3027 1411
rect 2969 1343 3027 1377
rect 2969 1309 2981 1343
rect 3015 1309 3027 1343
rect 2969 1275 3027 1309
rect 2969 1241 2981 1275
rect 3015 1241 3027 1275
rect 2969 1207 3027 1241
rect 2969 1173 2981 1207
rect 3015 1173 3027 1207
rect 2969 1139 3027 1173
rect 2969 1105 2981 1139
rect 3015 1105 3027 1139
rect 2969 1051 3027 1105
rect 3057 1343 3115 1451
rect 3057 1309 3069 1343
rect 3103 1309 3115 1343
rect 3057 1275 3115 1309
rect 3057 1241 3069 1275
rect 3103 1241 3115 1275
rect 3057 1207 3115 1241
rect 3057 1173 3069 1207
rect 3103 1173 3115 1207
rect 3057 1139 3115 1173
rect 3057 1105 3069 1139
rect 3103 1105 3115 1139
rect 3057 1051 3115 1105
rect 3145 1411 3199 1451
rect 3145 1377 3157 1411
rect 3191 1377 3199 1411
rect 3145 1343 3199 1377
rect 3145 1309 3157 1343
rect 3191 1309 3199 1343
rect 3145 1275 3199 1309
rect 3145 1241 3157 1275
rect 3191 1241 3199 1275
rect 3145 1207 3199 1241
rect 3145 1173 3157 1207
rect 3191 1173 3199 1207
rect 3145 1051 3199 1173
rect 3461 1411 3517 1451
rect 3461 1377 3471 1411
rect 3505 1377 3517 1411
rect 3461 1343 3517 1377
rect 3461 1309 3471 1343
rect 3505 1309 3517 1343
rect 3461 1275 3517 1309
rect 3461 1241 3471 1275
rect 3505 1241 3517 1275
rect 3461 1207 3517 1241
rect 3461 1173 3471 1207
rect 3505 1173 3517 1207
rect 3461 1139 3517 1173
rect 3461 1105 3471 1139
rect 3505 1105 3517 1139
rect 3461 1051 3517 1105
rect 3547 1343 3605 1451
rect 3547 1309 3559 1343
rect 3593 1309 3605 1343
rect 3547 1275 3605 1309
rect 3547 1241 3559 1275
rect 3593 1241 3605 1275
rect 3547 1207 3605 1241
rect 3547 1173 3559 1207
rect 3593 1173 3605 1207
rect 3547 1051 3605 1173
rect 3635 1411 3693 1451
rect 3635 1377 3647 1411
rect 3681 1377 3693 1411
rect 3635 1343 3693 1377
rect 3635 1309 3647 1343
rect 3681 1309 3693 1343
rect 3635 1275 3693 1309
rect 3635 1241 3647 1275
rect 3681 1241 3693 1275
rect 3635 1207 3693 1241
rect 3635 1173 3647 1207
rect 3681 1173 3693 1207
rect 3635 1139 3693 1173
rect 3635 1105 3647 1139
rect 3681 1105 3693 1139
rect 3635 1051 3693 1105
rect 3723 1343 3781 1451
rect 3723 1309 3735 1343
rect 3769 1309 3781 1343
rect 3723 1275 3781 1309
rect 3723 1241 3735 1275
rect 3769 1241 3781 1275
rect 3723 1207 3781 1241
rect 3723 1173 3735 1207
rect 3769 1173 3781 1207
rect 3723 1139 3781 1173
rect 3723 1105 3735 1139
rect 3769 1105 3781 1139
rect 3723 1051 3781 1105
rect 3811 1411 3865 1451
rect 3811 1377 3823 1411
rect 3857 1377 3865 1411
rect 3811 1343 3865 1377
rect 3811 1309 3823 1343
rect 3857 1309 3865 1343
rect 3811 1275 3865 1309
rect 3811 1241 3823 1275
rect 3857 1241 3865 1275
rect 3811 1207 3865 1241
rect 3811 1173 3823 1207
rect 3857 1173 3865 1207
rect 3811 1051 3865 1173
rect 4105 1412 4159 1450
rect 4105 1378 4113 1412
rect 4147 1378 4159 1412
rect 4105 1344 4159 1378
rect 4105 1310 4113 1344
rect 4147 1310 4159 1344
rect 4105 1276 4159 1310
rect 4105 1242 4113 1276
rect 4147 1242 4159 1276
rect 4105 1208 4159 1242
rect 4105 1174 4113 1208
rect 4147 1174 4159 1208
rect 4105 1139 4159 1174
rect 4105 1105 4113 1139
rect 4147 1105 4159 1139
rect 4105 1050 4159 1105
rect 4189 1412 4247 1450
rect 4189 1378 4201 1412
rect 4235 1378 4247 1412
rect 4189 1344 4247 1378
rect 4189 1310 4201 1344
rect 4235 1310 4247 1344
rect 4189 1276 4247 1310
rect 4189 1242 4201 1276
rect 4235 1242 4247 1276
rect 4189 1208 4247 1242
rect 4189 1174 4201 1208
rect 4235 1174 4247 1208
rect 4189 1139 4247 1174
rect 4189 1105 4201 1139
rect 4235 1105 4247 1139
rect 4189 1050 4247 1105
rect 4277 1412 4333 1450
rect 4277 1378 4289 1412
rect 4323 1378 4333 1412
rect 4277 1344 4333 1378
rect 4277 1310 4289 1344
rect 4323 1310 4333 1344
rect 4277 1276 4333 1310
rect 4277 1242 4289 1276
rect 4323 1242 4333 1276
rect 4277 1208 4333 1242
rect 4277 1174 4289 1208
rect 4323 1174 4333 1208
rect 4277 1139 4333 1174
rect 4277 1105 4289 1139
rect 4323 1105 4333 1139
rect 4277 1050 4333 1105
rect 4571 1412 4627 1450
rect 4571 1378 4581 1412
rect 4615 1378 4627 1412
rect 4571 1344 4627 1378
rect 4571 1310 4581 1344
rect 4615 1310 4627 1344
rect 4571 1276 4627 1310
rect 4571 1242 4581 1276
rect 4615 1242 4627 1276
rect 4571 1208 4627 1242
rect 4571 1174 4581 1208
rect 4615 1174 4627 1208
rect 4571 1139 4627 1174
rect 4571 1105 4581 1139
rect 4615 1105 4627 1139
rect 4571 1050 4627 1105
rect 4657 1412 4715 1450
rect 4657 1378 4669 1412
rect 4703 1378 4715 1412
rect 4657 1344 4715 1378
rect 4657 1310 4669 1344
rect 4703 1310 4715 1344
rect 4657 1276 4715 1310
rect 4657 1242 4669 1276
rect 4703 1242 4715 1276
rect 4657 1208 4715 1242
rect 4657 1174 4669 1208
rect 4703 1174 4715 1208
rect 4657 1139 4715 1174
rect 4657 1105 4669 1139
rect 4703 1105 4715 1139
rect 4657 1050 4715 1105
rect 4745 1412 4803 1450
rect 4745 1378 4757 1412
rect 4791 1378 4803 1412
rect 4745 1344 4803 1378
rect 4745 1310 4757 1344
rect 4791 1310 4803 1344
rect 4745 1276 4803 1310
rect 4745 1242 4757 1276
rect 4791 1242 4803 1276
rect 4745 1208 4803 1242
rect 4745 1174 4757 1208
rect 4791 1174 4803 1208
rect 4745 1050 4803 1174
rect 4833 1412 4891 1450
rect 4833 1378 4845 1412
rect 4879 1378 4891 1412
rect 4833 1344 4891 1378
rect 4833 1310 4845 1344
rect 4879 1310 4891 1344
rect 4833 1276 4891 1310
rect 4833 1242 4845 1276
rect 4879 1242 4891 1276
rect 4833 1208 4891 1242
rect 4833 1174 4845 1208
rect 4879 1174 4891 1208
rect 4833 1139 4891 1174
rect 4833 1105 4845 1139
rect 4879 1105 4891 1139
rect 4833 1050 4891 1105
rect 4921 1412 4975 1450
rect 4921 1378 4933 1412
rect 4967 1378 4975 1412
rect 4921 1344 4975 1378
rect 4921 1310 4933 1344
rect 4967 1310 4975 1344
rect 4921 1276 4975 1310
rect 4921 1242 4933 1276
rect 4967 1242 4975 1276
rect 4921 1208 4975 1242
rect 4921 1174 4933 1208
rect 4967 1174 4975 1208
rect 4921 1050 4975 1174
rect 5213 1412 5269 1450
rect 5213 1378 5223 1412
rect 5257 1378 5269 1412
rect 5213 1344 5269 1378
rect 5213 1310 5223 1344
rect 5257 1310 5269 1344
rect 5213 1276 5269 1310
rect 5213 1242 5223 1276
rect 5257 1242 5269 1276
rect 5213 1208 5269 1242
rect 5213 1174 5223 1208
rect 5257 1174 5269 1208
rect 5213 1139 5269 1174
rect 5213 1105 5223 1139
rect 5257 1105 5269 1139
rect 5213 1050 5269 1105
rect 5299 1412 5357 1450
rect 5299 1378 5311 1412
rect 5345 1378 5357 1412
rect 5299 1344 5357 1378
rect 5299 1310 5311 1344
rect 5345 1310 5357 1344
rect 5299 1276 5357 1310
rect 5299 1242 5311 1276
rect 5345 1242 5357 1276
rect 5299 1208 5357 1242
rect 5299 1174 5311 1208
rect 5345 1174 5357 1208
rect 5299 1139 5357 1174
rect 5299 1105 5311 1139
rect 5345 1105 5357 1139
rect 5299 1050 5357 1105
rect 5387 1412 5441 1450
rect 5387 1378 5399 1412
rect 5433 1378 5441 1412
rect 5387 1344 5441 1378
rect 5387 1310 5399 1344
rect 5433 1310 5441 1344
rect 5387 1276 5441 1310
rect 5387 1242 5399 1276
rect 5433 1242 5441 1276
rect 5387 1208 5441 1242
rect 5387 1174 5399 1208
rect 5433 1174 5441 1208
rect 5387 1139 5441 1174
rect 5387 1105 5399 1139
rect 5433 1105 5441 1139
rect 5387 1050 5441 1105
rect 5681 1412 5737 1450
rect 5681 1378 5691 1412
rect 5725 1378 5737 1412
rect 5681 1344 5737 1378
rect 5681 1310 5691 1344
rect 5725 1310 5737 1344
rect 5681 1276 5737 1310
rect 5681 1242 5691 1276
rect 5725 1242 5737 1276
rect 5681 1208 5737 1242
rect 5681 1174 5691 1208
rect 5725 1174 5737 1208
rect 5681 1139 5737 1174
rect 5681 1105 5691 1139
rect 5725 1105 5737 1139
rect 5681 1050 5737 1105
rect 5767 1412 5825 1450
rect 5767 1378 5779 1412
rect 5813 1378 5825 1412
rect 5767 1344 5825 1378
rect 5767 1310 5779 1344
rect 5813 1310 5825 1344
rect 5767 1276 5825 1310
rect 5767 1242 5779 1276
rect 5813 1242 5825 1276
rect 5767 1208 5825 1242
rect 5767 1174 5779 1208
rect 5813 1174 5825 1208
rect 5767 1139 5825 1174
rect 5767 1105 5779 1139
rect 5813 1105 5825 1139
rect 5767 1050 5825 1105
rect 5855 1412 5913 1450
rect 5855 1378 5867 1412
rect 5901 1378 5913 1412
rect 5855 1344 5913 1378
rect 5855 1310 5867 1344
rect 5901 1310 5913 1344
rect 5855 1276 5913 1310
rect 5855 1242 5867 1276
rect 5901 1242 5913 1276
rect 5855 1208 5913 1242
rect 5855 1174 5867 1208
rect 5901 1174 5913 1208
rect 5855 1050 5913 1174
rect 5943 1412 6001 1450
rect 5943 1378 5955 1412
rect 5989 1378 6001 1412
rect 5943 1344 6001 1378
rect 5943 1310 5955 1344
rect 5989 1310 6001 1344
rect 5943 1276 6001 1310
rect 5943 1242 5955 1276
rect 5989 1242 6001 1276
rect 5943 1208 6001 1242
rect 5943 1174 5955 1208
rect 5989 1174 6001 1208
rect 5943 1139 6001 1174
rect 5943 1105 5955 1139
rect 5989 1105 6001 1139
rect 5943 1050 6001 1105
rect 6031 1412 6085 1450
rect 6031 1378 6043 1412
rect 6077 1378 6085 1412
rect 6031 1344 6085 1378
rect 6031 1310 6043 1344
rect 6077 1310 6085 1344
rect 6031 1276 6085 1310
rect 6031 1242 6043 1276
rect 6077 1242 6085 1276
rect 6031 1208 6085 1242
rect 6031 1174 6043 1208
rect 6077 1174 6085 1208
rect 6031 1050 6085 1174
rect 6323 1412 6379 1450
rect 6323 1378 6333 1412
rect 6367 1378 6379 1412
rect 6323 1344 6379 1378
rect 6323 1310 6333 1344
rect 6367 1310 6379 1344
rect 6323 1276 6379 1310
rect 6323 1242 6333 1276
rect 6367 1242 6379 1276
rect 6323 1208 6379 1242
rect 6323 1174 6333 1208
rect 6367 1174 6379 1208
rect 6323 1139 6379 1174
rect 6323 1105 6333 1139
rect 6367 1105 6379 1139
rect 6323 1050 6379 1105
rect 6409 1412 6467 1450
rect 6409 1378 6421 1412
rect 6455 1378 6467 1412
rect 6409 1344 6467 1378
rect 6409 1310 6421 1344
rect 6455 1310 6467 1344
rect 6409 1276 6467 1310
rect 6409 1242 6421 1276
rect 6455 1242 6467 1276
rect 6409 1208 6467 1242
rect 6409 1174 6421 1208
rect 6455 1174 6467 1208
rect 6409 1139 6467 1174
rect 6409 1105 6421 1139
rect 6455 1105 6467 1139
rect 6409 1050 6467 1105
rect 6497 1412 6551 1450
rect 6497 1378 6509 1412
rect 6543 1378 6551 1412
rect 6497 1344 6551 1378
rect 6497 1310 6509 1344
rect 6543 1310 6551 1344
rect 6497 1276 6551 1310
rect 6497 1242 6509 1276
rect 6543 1242 6551 1276
rect 6497 1208 6551 1242
rect 6497 1174 6509 1208
rect 6543 1174 6551 1208
rect 6497 1139 6551 1174
rect 6497 1105 6509 1139
rect 6543 1105 6551 1139
rect 6497 1050 6551 1105
rect 6791 1411 6847 1451
rect 6791 1377 6801 1411
rect 6835 1377 6847 1411
rect 6791 1343 6847 1377
rect 6791 1309 6801 1343
rect 6835 1309 6847 1343
rect 6791 1275 6847 1309
rect 6791 1241 6801 1275
rect 6835 1241 6847 1275
rect 6791 1207 6847 1241
rect 6791 1173 6801 1207
rect 6835 1173 6847 1207
rect 6791 1139 6847 1173
rect 6791 1105 6801 1139
rect 6835 1105 6847 1139
rect 6791 1051 6847 1105
rect 6877 1411 6935 1451
rect 6877 1377 6889 1411
rect 6923 1377 6935 1411
rect 6877 1343 6935 1377
rect 6877 1309 6889 1343
rect 6923 1309 6935 1343
rect 6877 1275 6935 1309
rect 6877 1241 6889 1275
rect 6923 1241 6935 1275
rect 6877 1207 6935 1241
rect 6877 1173 6889 1207
rect 6923 1173 6935 1207
rect 6877 1051 6935 1173
rect 6965 1411 7023 1451
rect 6965 1377 6977 1411
rect 7011 1377 7023 1411
rect 6965 1343 7023 1377
rect 6965 1309 6977 1343
rect 7011 1309 7023 1343
rect 6965 1275 7023 1309
rect 6965 1241 6977 1275
rect 7011 1241 7023 1275
rect 6965 1207 7023 1241
rect 6965 1173 6977 1207
rect 7011 1173 7023 1207
rect 6965 1139 7023 1173
rect 6965 1105 6977 1139
rect 7011 1105 7023 1139
rect 6965 1051 7023 1105
rect 7053 1343 7111 1451
rect 7053 1309 7065 1343
rect 7099 1309 7111 1343
rect 7053 1275 7111 1309
rect 7053 1241 7065 1275
rect 7099 1241 7111 1275
rect 7053 1207 7111 1241
rect 7053 1173 7065 1207
rect 7099 1173 7111 1207
rect 7053 1139 7111 1173
rect 7053 1105 7065 1139
rect 7099 1105 7111 1139
rect 7053 1051 7111 1105
rect 7141 1411 7195 1451
rect 7141 1377 7153 1411
rect 7187 1377 7195 1411
rect 7141 1343 7195 1377
rect 7141 1309 7153 1343
rect 7187 1309 7195 1343
rect 7141 1275 7195 1309
rect 7141 1241 7153 1275
rect 7187 1241 7195 1275
rect 7141 1207 7195 1241
rect 7141 1173 7153 1207
rect 7187 1173 7195 1207
rect 7141 1051 7195 1173
rect 7433 1412 7489 1450
rect 7433 1378 7443 1412
rect 7477 1378 7489 1412
rect 7433 1344 7489 1378
rect 7433 1310 7443 1344
rect 7477 1310 7489 1344
rect 7433 1276 7489 1310
rect 7433 1242 7443 1276
rect 7477 1242 7489 1276
rect 7433 1208 7489 1242
rect 7433 1174 7443 1208
rect 7477 1174 7489 1208
rect 7433 1139 7489 1174
rect 7433 1105 7443 1139
rect 7477 1105 7489 1139
rect 7433 1050 7489 1105
rect 7519 1412 7577 1450
rect 7519 1378 7531 1412
rect 7565 1378 7577 1412
rect 7519 1344 7577 1378
rect 7519 1310 7531 1344
rect 7565 1310 7577 1344
rect 7519 1276 7577 1310
rect 7519 1242 7531 1276
rect 7565 1242 7577 1276
rect 7519 1208 7577 1242
rect 7519 1174 7531 1208
rect 7565 1174 7577 1208
rect 7519 1139 7577 1174
rect 7519 1105 7531 1139
rect 7565 1105 7577 1139
rect 7519 1050 7577 1105
rect 7607 1412 7661 1450
rect 7607 1378 7619 1412
rect 7653 1378 7661 1412
rect 7607 1344 7661 1378
rect 7607 1310 7619 1344
rect 7653 1310 7661 1344
rect 7607 1276 7661 1310
rect 7607 1242 7619 1276
rect 7653 1242 7661 1276
rect 7607 1208 7661 1242
rect 7607 1174 7619 1208
rect 7653 1174 7661 1208
rect 7607 1139 7661 1174
rect 7607 1105 7619 1139
rect 7653 1105 7661 1139
rect 7607 1050 7661 1105
<< ndiffc >>
rect 109 327 143 361
rect 303 327 337 361
rect 109 255 143 289
rect 109 187 143 221
rect 205 211 239 245
rect 303 255 337 289
rect 303 187 337 221
rect 109 117 143 151
rect 205 117 239 151
rect 303 117 337 151
rect 566 327 600 361
rect 663 327 697 361
rect 760 327 794 361
rect 566 255 600 289
rect 566 187 600 221
rect 663 202 697 236
rect 760 255 794 289
rect 760 187 794 221
rect 857 211 891 245
rect 954 255 988 289
rect 954 187 988 221
rect 566 117 600 151
rect 760 117 794 151
rect 857 117 891 151
rect 954 117 988 151
rect 1232 327 1266 361
rect 1329 327 1363 361
rect 1426 327 1460 361
rect 1232 255 1266 289
rect 1232 187 1266 221
rect 1329 202 1363 236
rect 1426 255 1460 289
rect 1426 187 1460 221
rect 1523 211 1557 245
rect 1620 255 1654 289
rect 1620 187 1654 221
rect 1232 117 1266 151
rect 1426 117 1460 151
rect 1523 117 1557 151
rect 1620 117 1654 151
rect 1883 327 1917 361
rect 2077 327 2111 361
rect 1883 255 1917 289
rect 1883 187 1917 221
rect 1981 211 2015 245
rect 2077 255 2111 289
rect 2077 187 2111 221
rect 1883 117 1917 151
rect 1981 117 2015 151
rect 2077 117 2111 151
rect 2329 327 2363 361
rect 2523 327 2557 361
rect 2329 255 2363 289
rect 2329 187 2363 221
rect 2425 211 2459 245
rect 2523 255 2557 289
rect 2523 187 2557 221
rect 2329 117 2363 151
rect 2425 117 2459 151
rect 2523 117 2557 151
rect 2786 327 2820 361
rect 2883 327 2917 361
rect 2980 327 3014 361
rect 2786 255 2820 289
rect 2786 187 2820 221
rect 2883 202 2917 236
rect 2980 255 3014 289
rect 2980 187 3014 221
rect 3077 211 3111 245
rect 3174 255 3208 289
rect 3174 187 3208 221
rect 2786 117 2820 151
rect 2980 117 3014 151
rect 3077 117 3111 151
rect 3174 117 3208 151
rect 3452 327 3486 361
rect 3549 327 3583 361
rect 3646 327 3680 361
rect 3452 255 3486 289
rect 3452 187 3486 221
rect 3549 202 3583 236
rect 3646 255 3680 289
rect 3646 187 3680 221
rect 3743 211 3777 245
rect 3840 255 3874 289
rect 3840 187 3874 221
rect 3452 117 3486 151
rect 3646 117 3680 151
rect 3743 117 3777 151
rect 3840 117 3874 151
rect 4103 327 4137 361
rect 4297 327 4331 361
rect 4103 255 4137 289
rect 4103 187 4137 221
rect 4201 211 4235 245
rect 4297 255 4331 289
rect 4297 187 4331 221
rect 4103 117 4137 151
rect 4201 117 4235 151
rect 4297 117 4331 151
rect 4562 327 4596 361
rect 4659 327 4693 361
rect 4756 327 4790 361
rect 4562 255 4596 289
rect 4562 187 4596 221
rect 4659 202 4693 236
rect 4756 255 4790 289
rect 4756 187 4790 221
rect 4853 211 4887 245
rect 4950 255 4984 289
rect 4950 187 4984 221
rect 4562 117 4596 151
rect 4756 117 4790 151
rect 4853 117 4887 151
rect 4950 117 4984 151
rect 5215 327 5249 361
rect 5409 327 5443 361
rect 5215 255 5249 289
rect 5215 187 5249 221
rect 5311 211 5345 245
rect 5409 255 5443 289
rect 5409 187 5443 221
rect 5215 117 5249 151
rect 5311 117 5345 151
rect 5409 117 5443 151
rect 5672 327 5706 361
rect 5769 327 5803 361
rect 5866 327 5900 361
rect 5672 255 5706 289
rect 5672 187 5706 221
rect 5769 202 5803 236
rect 5866 255 5900 289
rect 5866 187 5900 221
rect 5963 211 5997 245
rect 6060 255 6094 289
rect 6060 187 6094 221
rect 5672 117 5706 151
rect 5866 117 5900 151
rect 5963 117 5997 151
rect 6060 117 6094 151
rect 6325 327 6359 361
rect 6519 327 6553 361
rect 6325 255 6359 289
rect 6325 187 6359 221
rect 6421 211 6455 245
rect 6519 255 6553 289
rect 6519 187 6553 221
rect 6325 117 6359 151
rect 6421 117 6455 151
rect 6519 117 6553 151
rect 6782 327 6816 361
rect 6782 255 6816 289
rect 6782 187 6816 221
rect 6879 211 6913 245
rect 6976 255 7010 289
rect 6976 187 7010 221
rect 7073 211 7107 245
rect 7170 255 7204 289
rect 7170 187 7204 221
rect 6782 117 6816 151
rect 6879 117 6913 151
rect 6976 117 7010 151
rect 7073 117 7107 151
rect 7170 117 7204 151
rect 7435 327 7469 361
rect 7629 327 7663 361
rect 7435 255 7469 289
rect 7435 187 7469 221
rect 7531 211 7565 245
rect 7629 255 7663 289
rect 7629 187 7663 221
rect 7435 117 7469 151
rect 7531 117 7565 151
rect 7629 117 7663 151
<< pdiffc >>
rect 117 1378 151 1412
rect 117 1310 151 1344
rect 117 1242 151 1276
rect 117 1174 151 1208
rect 117 1105 151 1139
rect 205 1378 239 1412
rect 205 1310 239 1344
rect 205 1242 239 1276
rect 205 1174 239 1208
rect 205 1105 239 1139
rect 293 1378 327 1412
rect 293 1310 327 1344
rect 293 1242 327 1276
rect 293 1174 327 1208
rect 293 1105 327 1139
rect 585 1377 619 1411
rect 585 1309 619 1343
rect 585 1241 619 1275
rect 585 1173 619 1207
rect 585 1105 619 1139
rect 673 1309 707 1343
rect 673 1241 707 1275
rect 673 1173 707 1207
rect 761 1377 795 1411
rect 761 1309 795 1343
rect 761 1241 795 1275
rect 761 1173 795 1207
rect 761 1105 795 1139
rect 849 1309 883 1343
rect 849 1241 883 1275
rect 849 1173 883 1207
rect 849 1105 883 1139
rect 937 1377 971 1411
rect 937 1309 971 1343
rect 937 1241 971 1275
rect 937 1173 971 1207
rect 1251 1377 1285 1411
rect 1251 1309 1285 1343
rect 1251 1241 1285 1275
rect 1251 1173 1285 1207
rect 1251 1105 1285 1139
rect 1339 1309 1373 1343
rect 1339 1241 1373 1275
rect 1339 1173 1373 1207
rect 1427 1377 1461 1411
rect 1427 1309 1461 1343
rect 1427 1241 1461 1275
rect 1427 1173 1461 1207
rect 1427 1105 1461 1139
rect 1515 1309 1549 1343
rect 1515 1241 1549 1275
rect 1515 1173 1549 1207
rect 1515 1105 1549 1139
rect 1603 1377 1637 1411
rect 1603 1309 1637 1343
rect 1603 1241 1637 1275
rect 1603 1173 1637 1207
rect 1893 1378 1927 1412
rect 1893 1310 1927 1344
rect 1893 1242 1927 1276
rect 1893 1174 1927 1208
rect 1893 1105 1927 1139
rect 1981 1378 2015 1412
rect 1981 1310 2015 1344
rect 1981 1242 2015 1276
rect 1981 1174 2015 1208
rect 1981 1105 2015 1139
rect 2069 1378 2103 1412
rect 2069 1310 2103 1344
rect 2069 1242 2103 1276
rect 2069 1174 2103 1208
rect 2069 1105 2103 1139
rect 2337 1378 2371 1412
rect 2337 1310 2371 1344
rect 2337 1242 2371 1276
rect 2337 1174 2371 1208
rect 2337 1105 2371 1139
rect 2425 1378 2459 1412
rect 2425 1310 2459 1344
rect 2425 1242 2459 1276
rect 2425 1174 2459 1208
rect 2425 1105 2459 1139
rect 2513 1378 2547 1412
rect 2513 1310 2547 1344
rect 2513 1242 2547 1276
rect 2513 1174 2547 1208
rect 2513 1105 2547 1139
rect 2805 1377 2839 1411
rect 2805 1309 2839 1343
rect 2805 1241 2839 1275
rect 2805 1173 2839 1207
rect 2805 1105 2839 1139
rect 2893 1309 2927 1343
rect 2893 1241 2927 1275
rect 2893 1173 2927 1207
rect 2981 1377 3015 1411
rect 2981 1309 3015 1343
rect 2981 1241 3015 1275
rect 2981 1173 3015 1207
rect 2981 1105 3015 1139
rect 3069 1309 3103 1343
rect 3069 1241 3103 1275
rect 3069 1173 3103 1207
rect 3069 1105 3103 1139
rect 3157 1377 3191 1411
rect 3157 1309 3191 1343
rect 3157 1241 3191 1275
rect 3157 1173 3191 1207
rect 3471 1377 3505 1411
rect 3471 1309 3505 1343
rect 3471 1241 3505 1275
rect 3471 1173 3505 1207
rect 3471 1105 3505 1139
rect 3559 1309 3593 1343
rect 3559 1241 3593 1275
rect 3559 1173 3593 1207
rect 3647 1377 3681 1411
rect 3647 1309 3681 1343
rect 3647 1241 3681 1275
rect 3647 1173 3681 1207
rect 3647 1105 3681 1139
rect 3735 1309 3769 1343
rect 3735 1241 3769 1275
rect 3735 1173 3769 1207
rect 3735 1105 3769 1139
rect 3823 1377 3857 1411
rect 3823 1309 3857 1343
rect 3823 1241 3857 1275
rect 3823 1173 3857 1207
rect 4113 1378 4147 1412
rect 4113 1310 4147 1344
rect 4113 1242 4147 1276
rect 4113 1174 4147 1208
rect 4113 1105 4147 1139
rect 4201 1378 4235 1412
rect 4201 1310 4235 1344
rect 4201 1242 4235 1276
rect 4201 1174 4235 1208
rect 4201 1105 4235 1139
rect 4289 1378 4323 1412
rect 4289 1310 4323 1344
rect 4289 1242 4323 1276
rect 4289 1174 4323 1208
rect 4289 1105 4323 1139
rect 4581 1378 4615 1412
rect 4581 1310 4615 1344
rect 4581 1242 4615 1276
rect 4581 1174 4615 1208
rect 4581 1105 4615 1139
rect 4669 1378 4703 1412
rect 4669 1310 4703 1344
rect 4669 1242 4703 1276
rect 4669 1174 4703 1208
rect 4669 1105 4703 1139
rect 4757 1378 4791 1412
rect 4757 1310 4791 1344
rect 4757 1242 4791 1276
rect 4757 1174 4791 1208
rect 4845 1378 4879 1412
rect 4845 1310 4879 1344
rect 4845 1242 4879 1276
rect 4845 1174 4879 1208
rect 4845 1105 4879 1139
rect 4933 1378 4967 1412
rect 4933 1310 4967 1344
rect 4933 1242 4967 1276
rect 4933 1174 4967 1208
rect 5223 1378 5257 1412
rect 5223 1310 5257 1344
rect 5223 1242 5257 1276
rect 5223 1174 5257 1208
rect 5223 1105 5257 1139
rect 5311 1378 5345 1412
rect 5311 1310 5345 1344
rect 5311 1242 5345 1276
rect 5311 1174 5345 1208
rect 5311 1105 5345 1139
rect 5399 1378 5433 1412
rect 5399 1310 5433 1344
rect 5399 1242 5433 1276
rect 5399 1174 5433 1208
rect 5399 1105 5433 1139
rect 5691 1378 5725 1412
rect 5691 1310 5725 1344
rect 5691 1242 5725 1276
rect 5691 1174 5725 1208
rect 5691 1105 5725 1139
rect 5779 1378 5813 1412
rect 5779 1310 5813 1344
rect 5779 1242 5813 1276
rect 5779 1174 5813 1208
rect 5779 1105 5813 1139
rect 5867 1378 5901 1412
rect 5867 1310 5901 1344
rect 5867 1242 5901 1276
rect 5867 1174 5901 1208
rect 5955 1378 5989 1412
rect 5955 1310 5989 1344
rect 5955 1242 5989 1276
rect 5955 1174 5989 1208
rect 5955 1105 5989 1139
rect 6043 1378 6077 1412
rect 6043 1310 6077 1344
rect 6043 1242 6077 1276
rect 6043 1174 6077 1208
rect 6333 1378 6367 1412
rect 6333 1310 6367 1344
rect 6333 1242 6367 1276
rect 6333 1174 6367 1208
rect 6333 1105 6367 1139
rect 6421 1378 6455 1412
rect 6421 1310 6455 1344
rect 6421 1242 6455 1276
rect 6421 1174 6455 1208
rect 6421 1105 6455 1139
rect 6509 1378 6543 1412
rect 6509 1310 6543 1344
rect 6509 1242 6543 1276
rect 6509 1174 6543 1208
rect 6509 1105 6543 1139
rect 6801 1377 6835 1411
rect 6801 1309 6835 1343
rect 6801 1241 6835 1275
rect 6801 1173 6835 1207
rect 6801 1105 6835 1139
rect 6889 1377 6923 1411
rect 6889 1309 6923 1343
rect 6889 1241 6923 1275
rect 6889 1173 6923 1207
rect 6977 1377 7011 1411
rect 6977 1309 7011 1343
rect 6977 1241 7011 1275
rect 6977 1173 7011 1207
rect 6977 1105 7011 1139
rect 7065 1309 7099 1343
rect 7065 1241 7099 1275
rect 7065 1173 7099 1207
rect 7065 1105 7099 1139
rect 7153 1377 7187 1411
rect 7153 1309 7187 1343
rect 7153 1241 7187 1275
rect 7153 1173 7187 1207
rect 7443 1378 7477 1412
rect 7443 1310 7477 1344
rect 7443 1242 7477 1276
rect 7443 1174 7477 1208
rect 7443 1105 7477 1139
rect 7531 1378 7565 1412
rect 7531 1310 7565 1344
rect 7531 1242 7565 1276
rect 7531 1174 7565 1208
rect 7531 1105 7565 1139
rect 7619 1378 7653 1412
rect 7619 1310 7653 1344
rect 7619 1242 7653 1276
rect 7619 1174 7653 1208
rect 7619 1105 7653 1139
<< psubdiff >>
rect -31 546 7801 572
rect -31 512 -17 546
rect 17 512 427 546
rect 461 512 1093 546
rect 1127 512 1759 546
rect 1793 512 2203 546
rect 2237 512 2647 546
rect 2681 512 3313 546
rect 3347 512 3979 546
rect 4013 512 4423 546
rect 4457 512 5089 546
rect 5123 512 5533 546
rect 5567 512 6199 546
rect 6233 512 6643 546
rect 6677 512 7309 546
rect 7343 512 7753 546
rect 7787 512 7801 546
rect -31 510 7801 512
rect -31 474 31 510
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect 413 474 475 510
rect -31 368 -17 402
rect 17 368 31 402
rect 413 440 427 474
rect 461 440 475 474
rect 413 402 475 440
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect 413 368 427 402
rect 461 368 475 402
rect 1079 474 1141 510
rect 1079 440 1093 474
rect 1127 440 1141 474
rect 1079 402 1141 440
rect 413 330 475 368
rect 413 296 427 330
rect 461 296 475 330
rect 413 258 475 296
rect 413 224 427 258
rect 461 224 475 258
rect 413 186 475 224
rect 413 152 427 186
rect 461 152 475 186
rect 413 114 475 152
rect -31 47 31 80
rect 413 80 427 114
rect 461 80 475 114
rect 1079 368 1093 402
rect 1127 368 1141 402
rect 1745 474 1807 510
rect 1745 440 1759 474
rect 1793 440 1807 474
rect 1745 402 1807 440
rect 1079 330 1141 368
rect 1079 296 1093 330
rect 1127 296 1141 330
rect 1079 258 1141 296
rect 1079 224 1093 258
rect 1127 224 1141 258
rect 1079 186 1141 224
rect 1079 152 1093 186
rect 1127 152 1141 186
rect 1079 114 1141 152
rect 413 47 475 80
rect 1079 80 1093 114
rect 1127 80 1141 114
rect 1745 368 1759 402
rect 1793 368 1807 402
rect 2189 474 2251 510
rect 2189 440 2203 474
rect 2237 440 2251 474
rect 2189 402 2251 440
rect 2633 474 2695 510
rect 1745 330 1807 368
rect 1745 296 1759 330
rect 1793 296 1807 330
rect 1745 258 1807 296
rect 1745 224 1759 258
rect 1793 224 1807 258
rect 1745 186 1807 224
rect 1745 152 1759 186
rect 1793 152 1807 186
rect 1745 114 1807 152
rect 1079 47 1141 80
rect 1745 80 1759 114
rect 1793 80 1807 114
rect 2189 368 2203 402
rect 2237 368 2251 402
rect 2633 440 2647 474
rect 2681 440 2695 474
rect 2633 402 2695 440
rect 2189 330 2251 368
rect 2189 296 2203 330
rect 2237 296 2251 330
rect 2189 258 2251 296
rect 2189 224 2203 258
rect 2237 224 2251 258
rect 2189 186 2251 224
rect 2189 152 2203 186
rect 2237 152 2251 186
rect 2189 114 2251 152
rect 1745 47 1807 80
rect 2189 80 2203 114
rect 2237 80 2251 114
rect 2633 368 2647 402
rect 2681 368 2695 402
rect 3299 474 3361 510
rect 3299 440 3313 474
rect 3347 440 3361 474
rect 3299 402 3361 440
rect 2633 330 2695 368
rect 2633 296 2647 330
rect 2681 296 2695 330
rect 2633 258 2695 296
rect 2633 224 2647 258
rect 2681 224 2695 258
rect 2633 186 2695 224
rect 2633 152 2647 186
rect 2681 152 2695 186
rect 2633 114 2695 152
rect 2189 47 2251 80
rect 2633 80 2647 114
rect 2681 80 2695 114
rect 3299 368 3313 402
rect 3347 368 3361 402
rect 3965 474 4027 510
rect 3965 440 3979 474
rect 4013 440 4027 474
rect 3965 402 4027 440
rect 3299 330 3361 368
rect 3299 296 3313 330
rect 3347 296 3361 330
rect 3299 258 3361 296
rect 3299 224 3313 258
rect 3347 224 3361 258
rect 3299 186 3361 224
rect 3299 152 3313 186
rect 3347 152 3361 186
rect 3299 114 3361 152
rect 2633 47 2695 80
rect 3299 80 3313 114
rect 3347 80 3361 114
rect 3965 368 3979 402
rect 4013 368 4027 402
rect 4409 474 4471 510
rect 4409 440 4423 474
rect 4457 440 4471 474
rect 4409 402 4471 440
rect 3965 330 4027 368
rect 3965 296 3979 330
rect 4013 296 4027 330
rect 3965 258 4027 296
rect 3965 224 3979 258
rect 4013 224 4027 258
rect 3965 186 4027 224
rect 3965 152 3979 186
rect 4013 152 4027 186
rect 3965 114 4027 152
rect 3299 47 3361 80
rect 3965 80 3979 114
rect 4013 80 4027 114
rect 4409 368 4423 402
rect 4457 368 4471 402
rect 5075 474 5137 510
rect 5075 440 5089 474
rect 5123 440 5137 474
rect 5075 402 5137 440
rect 5519 474 5581 510
rect 4409 330 4471 368
rect 4409 296 4423 330
rect 4457 296 4471 330
rect 4409 258 4471 296
rect 4409 224 4423 258
rect 4457 224 4471 258
rect 4409 186 4471 224
rect 4409 152 4423 186
rect 4457 152 4471 186
rect 4409 114 4471 152
rect 3965 47 4027 80
rect 4409 80 4423 114
rect 4457 80 4471 114
rect 5075 368 5089 402
rect 5123 368 5137 402
rect 5519 440 5533 474
rect 5567 440 5581 474
rect 5519 402 5581 440
rect 5075 330 5137 368
rect 5075 296 5089 330
rect 5123 296 5137 330
rect 5075 258 5137 296
rect 5075 224 5089 258
rect 5123 224 5137 258
rect 5075 186 5137 224
rect 5075 152 5089 186
rect 5123 152 5137 186
rect 5075 114 5137 152
rect 4409 47 4471 80
rect 5075 80 5089 114
rect 5123 80 5137 114
rect 5519 368 5533 402
rect 5567 368 5581 402
rect 6185 474 6247 510
rect 6185 440 6199 474
rect 6233 440 6247 474
rect 6185 402 6247 440
rect 6629 474 6691 510
rect 5519 330 5581 368
rect 5519 296 5533 330
rect 5567 296 5581 330
rect 5519 258 5581 296
rect 5519 224 5533 258
rect 5567 224 5581 258
rect 5519 186 5581 224
rect 5519 152 5533 186
rect 5567 152 5581 186
rect 5519 114 5581 152
rect 5075 47 5137 80
rect 5519 80 5533 114
rect 5567 80 5581 114
rect 6185 368 6199 402
rect 6233 368 6247 402
rect 6629 440 6643 474
rect 6677 440 6691 474
rect 6629 402 6691 440
rect 6185 330 6247 368
rect 6185 296 6199 330
rect 6233 296 6247 330
rect 6185 258 6247 296
rect 6185 224 6199 258
rect 6233 224 6247 258
rect 6185 186 6247 224
rect 6185 152 6199 186
rect 6233 152 6247 186
rect 6185 114 6247 152
rect 5519 47 5581 80
rect 6185 80 6199 114
rect 6233 80 6247 114
rect 6629 368 6643 402
rect 6677 368 6691 402
rect 7295 474 7357 510
rect 7295 440 7309 474
rect 7343 440 7357 474
rect 7295 402 7357 440
rect 7739 474 7801 510
rect 6629 330 6691 368
rect 6629 296 6643 330
rect 6677 296 6691 330
rect 6629 258 6691 296
rect 6629 224 6643 258
rect 6677 224 6691 258
rect 6629 186 6691 224
rect 6629 152 6643 186
rect 6677 152 6691 186
rect 6629 114 6691 152
rect 6185 47 6247 80
rect 6629 80 6643 114
rect 6677 80 6691 114
rect 7295 368 7309 402
rect 7343 368 7357 402
rect 7739 440 7753 474
rect 7787 440 7801 474
rect 7739 402 7801 440
rect 7295 330 7357 368
rect 7295 296 7309 330
rect 7343 296 7357 330
rect 7295 258 7357 296
rect 7295 224 7309 258
rect 7343 224 7357 258
rect 7295 186 7357 224
rect 7295 152 7309 186
rect 7343 152 7357 186
rect 7295 114 7357 152
rect 6629 47 6691 80
rect 7295 80 7309 114
rect 7343 80 7357 114
rect 7739 368 7753 402
rect 7787 368 7801 402
rect 7739 330 7801 368
rect 7739 296 7753 330
rect 7787 296 7801 330
rect 7739 258 7801 296
rect 7739 224 7753 258
rect 7787 224 7801 258
rect 7739 186 7801 224
rect 7739 152 7753 186
rect 7787 152 7801 186
rect 7739 114 7801 152
rect 7295 47 7357 80
rect 7739 80 7753 114
rect 7787 80 7801 114
rect 7739 47 7801 80
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 205 47
rect 239 13 283 47
rect 317 13 355 47
rect 389 13 499 47
rect 533 13 571 47
rect 605 13 643 47
rect 677 13 715 47
rect 749 13 805 47
rect 839 13 877 47
rect 911 13 949 47
rect 983 13 1021 47
rect 1055 13 1165 47
rect 1199 13 1237 47
rect 1271 13 1309 47
rect 1343 13 1381 47
rect 1415 13 1471 47
rect 1505 13 1543 47
rect 1577 13 1615 47
rect 1649 13 1687 47
rect 1721 13 1831 47
rect 1865 13 1903 47
rect 1937 13 1981 47
rect 2015 13 2059 47
rect 2093 13 2131 47
rect 2165 13 2275 47
rect 2309 13 2347 47
rect 2381 13 2425 47
rect 2459 13 2503 47
rect 2537 13 2575 47
rect 2609 13 2719 47
rect 2753 13 2791 47
rect 2825 13 2863 47
rect 2897 13 2935 47
rect 2969 13 3025 47
rect 3059 13 3097 47
rect 3131 13 3169 47
rect 3203 13 3241 47
rect 3275 13 3385 47
rect 3419 13 3457 47
rect 3491 13 3529 47
rect 3563 13 3601 47
rect 3635 13 3691 47
rect 3725 13 3763 47
rect 3797 13 3835 47
rect 3869 13 3907 47
rect 3941 13 4051 47
rect 4085 13 4123 47
rect 4157 13 4201 47
rect 4235 13 4279 47
rect 4313 13 4351 47
rect 4385 13 4495 47
rect 4529 13 4567 47
rect 4601 13 4639 47
rect 4673 13 4711 47
rect 4745 13 4801 47
rect 4835 13 4873 47
rect 4907 13 4945 47
rect 4979 13 5017 47
rect 5051 13 5161 47
rect 5195 13 5233 47
rect 5267 13 5311 47
rect 5345 13 5389 47
rect 5423 13 5461 47
rect 5495 13 5605 47
rect 5639 13 5677 47
rect 5711 13 5749 47
rect 5783 13 5821 47
rect 5855 13 5911 47
rect 5945 13 5983 47
rect 6017 13 6055 47
rect 6089 13 6127 47
rect 6161 13 6271 47
rect 6305 13 6343 47
rect 6377 13 6421 47
rect 6455 13 6499 47
rect 6533 13 6571 47
rect 6605 13 6715 47
rect 6749 13 6787 47
rect 6821 13 6859 47
rect 6893 13 6931 47
rect 6965 13 7021 47
rect 7055 13 7093 47
rect 7127 13 7165 47
rect 7199 13 7237 47
rect 7271 13 7381 47
rect 7415 13 7453 47
rect 7487 13 7531 47
rect 7565 13 7609 47
rect 7643 13 7681 47
rect 7715 13 7801 47
rect -31 11 31 13
rect 413 11 475 13
rect 1079 11 1141 13
rect 1745 11 1807 13
rect 2189 11 2251 13
rect 2633 11 2695 13
rect 3299 11 3361 13
rect 3965 11 4027 13
rect 4409 11 4471 13
rect 5075 11 5137 13
rect 5519 11 5581 13
rect 6185 11 6247 13
rect 6629 11 6691 13
rect 7295 11 7357 13
rect 7739 11 7801 13
<< nsubdiff >>
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 205 1539
rect 239 1505 283 1539
rect 317 1505 355 1539
rect 389 1505 499 1539
rect 533 1505 571 1539
rect 605 1505 643 1539
rect 677 1505 715 1539
rect 749 1505 805 1539
rect 839 1505 877 1539
rect 911 1505 949 1539
rect 983 1505 1021 1539
rect 1055 1505 1165 1539
rect 1199 1505 1237 1539
rect 1271 1505 1309 1539
rect 1343 1505 1381 1539
rect 1415 1505 1471 1539
rect 1505 1505 1543 1539
rect 1577 1505 1615 1539
rect 1649 1505 1687 1539
rect 1721 1505 1831 1539
rect 1865 1505 1903 1539
rect 1937 1505 1981 1539
rect 2015 1505 2059 1539
rect 2093 1505 2131 1539
rect 2165 1505 2275 1539
rect 2309 1505 2347 1539
rect 2381 1505 2425 1539
rect 2459 1505 2503 1539
rect 2537 1505 2575 1539
rect 2609 1505 2719 1539
rect 2753 1505 2791 1539
rect 2825 1505 2863 1539
rect 2897 1505 2935 1539
rect 2969 1505 3025 1539
rect 3059 1505 3097 1539
rect 3131 1505 3169 1539
rect 3203 1505 3241 1539
rect 3275 1505 3385 1539
rect 3419 1505 3457 1539
rect 3491 1505 3529 1539
rect 3563 1505 3601 1539
rect 3635 1505 3691 1539
rect 3725 1505 3763 1539
rect 3797 1505 3835 1539
rect 3869 1505 3907 1539
rect 3941 1505 4051 1539
rect 4085 1505 4123 1539
rect 4157 1505 4201 1539
rect 4235 1505 4279 1539
rect 4313 1505 4351 1539
rect 4385 1505 4495 1539
rect 4529 1505 4567 1539
rect 4601 1505 4639 1539
rect 4673 1505 4711 1539
rect 4745 1505 4801 1539
rect 4835 1505 4873 1539
rect 4907 1505 4945 1539
rect 4979 1505 5017 1539
rect 5051 1505 5161 1539
rect 5195 1505 5233 1539
rect 5267 1505 5311 1539
rect 5345 1505 5389 1539
rect 5423 1505 5461 1539
rect 5495 1505 5605 1539
rect 5639 1505 5677 1539
rect 5711 1505 5749 1539
rect 5783 1505 5821 1539
rect 5855 1505 5911 1539
rect 5945 1505 5983 1539
rect 6017 1505 6055 1539
rect 6089 1505 6127 1539
rect 6161 1505 6271 1539
rect 6305 1505 6343 1539
rect 6377 1505 6421 1539
rect 6455 1505 6499 1539
rect 6533 1505 6571 1539
rect 6605 1505 6715 1539
rect 6749 1505 6787 1539
rect 6821 1505 6859 1539
rect 6893 1505 6931 1539
rect 6965 1505 7021 1539
rect 7055 1505 7093 1539
rect 7127 1505 7165 1539
rect 7199 1505 7237 1539
rect 7271 1505 7381 1539
rect 7415 1505 7453 1539
rect 7487 1505 7531 1539
rect 7565 1505 7609 1539
rect 7643 1505 7681 1539
rect 7715 1505 7801 1539
rect -31 1470 31 1505
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect 413 1470 475 1505
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect -31 1038 31 1076
rect 413 1436 427 1470
rect 461 1436 475 1470
rect 1079 1470 1141 1505
rect 413 1398 475 1436
rect 413 1364 427 1398
rect 461 1364 475 1398
rect 413 1326 475 1364
rect 413 1292 427 1326
rect 461 1292 475 1326
rect 413 1254 475 1292
rect 413 1220 427 1254
rect 461 1220 475 1254
rect 413 1182 475 1220
rect 413 1148 427 1182
rect 461 1148 475 1182
rect 413 1110 475 1148
rect 413 1076 427 1110
rect 461 1076 475 1110
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect 413 1038 475 1076
rect 1079 1436 1093 1470
rect 1127 1436 1141 1470
rect 1745 1470 1807 1505
rect 1079 1398 1141 1436
rect 1079 1364 1093 1398
rect 1127 1364 1141 1398
rect 1079 1326 1141 1364
rect 1079 1292 1093 1326
rect 1127 1292 1141 1326
rect 1079 1254 1141 1292
rect 1079 1220 1093 1254
rect 1127 1220 1141 1254
rect 1079 1182 1141 1220
rect 1079 1148 1093 1182
rect 1127 1148 1141 1182
rect 1079 1110 1141 1148
rect 1079 1076 1093 1110
rect 1127 1076 1141 1110
rect 413 1004 427 1038
rect 461 1004 475 1038
rect 413 966 475 1004
rect -31 930 31 932
rect 413 932 427 966
rect 461 932 475 966
rect 1079 1038 1141 1076
rect 1745 1436 1759 1470
rect 1793 1436 1807 1470
rect 2189 1470 2251 1505
rect 1745 1398 1807 1436
rect 1745 1364 1759 1398
rect 1793 1364 1807 1398
rect 1745 1326 1807 1364
rect 1745 1292 1759 1326
rect 1793 1292 1807 1326
rect 1745 1254 1807 1292
rect 1745 1220 1759 1254
rect 1793 1220 1807 1254
rect 1745 1182 1807 1220
rect 1745 1148 1759 1182
rect 1793 1148 1807 1182
rect 1745 1110 1807 1148
rect 1745 1076 1759 1110
rect 1793 1076 1807 1110
rect 1079 1004 1093 1038
rect 1127 1004 1141 1038
rect 1079 966 1141 1004
rect 413 930 475 932
rect 1079 932 1093 966
rect 1127 932 1141 966
rect 1745 1038 1807 1076
rect 2189 1436 2203 1470
rect 2237 1436 2251 1470
rect 2633 1470 2695 1505
rect 2189 1398 2251 1436
rect 2189 1364 2203 1398
rect 2237 1364 2251 1398
rect 2189 1326 2251 1364
rect 2189 1292 2203 1326
rect 2237 1292 2251 1326
rect 2189 1254 2251 1292
rect 2189 1220 2203 1254
rect 2237 1220 2251 1254
rect 2189 1182 2251 1220
rect 2189 1148 2203 1182
rect 2237 1148 2251 1182
rect 2189 1110 2251 1148
rect 2189 1076 2203 1110
rect 2237 1076 2251 1110
rect 1745 1004 1759 1038
rect 1793 1004 1807 1038
rect 1745 966 1807 1004
rect 2189 1038 2251 1076
rect 2633 1436 2647 1470
rect 2681 1436 2695 1470
rect 3299 1470 3361 1505
rect 2633 1398 2695 1436
rect 2633 1364 2647 1398
rect 2681 1364 2695 1398
rect 2633 1326 2695 1364
rect 2633 1292 2647 1326
rect 2681 1292 2695 1326
rect 2633 1254 2695 1292
rect 2633 1220 2647 1254
rect 2681 1220 2695 1254
rect 2633 1182 2695 1220
rect 2633 1148 2647 1182
rect 2681 1148 2695 1182
rect 2633 1110 2695 1148
rect 2633 1076 2647 1110
rect 2681 1076 2695 1110
rect 1079 930 1141 932
rect 1745 932 1759 966
rect 1793 932 1807 966
rect 2189 1004 2203 1038
rect 2237 1004 2251 1038
rect 2189 966 2251 1004
rect 1745 930 1807 932
rect 2189 932 2203 966
rect 2237 932 2251 966
rect 2633 1038 2695 1076
rect 3299 1436 3313 1470
rect 3347 1436 3361 1470
rect 3965 1470 4027 1505
rect 3299 1398 3361 1436
rect 3299 1364 3313 1398
rect 3347 1364 3361 1398
rect 3299 1326 3361 1364
rect 3299 1292 3313 1326
rect 3347 1292 3361 1326
rect 3299 1254 3361 1292
rect 3299 1220 3313 1254
rect 3347 1220 3361 1254
rect 3299 1182 3361 1220
rect 3299 1148 3313 1182
rect 3347 1148 3361 1182
rect 3299 1110 3361 1148
rect 3299 1076 3313 1110
rect 3347 1076 3361 1110
rect 2633 1004 2647 1038
rect 2681 1004 2695 1038
rect 2633 966 2695 1004
rect 2189 930 2251 932
rect 2633 932 2647 966
rect 2681 932 2695 966
rect 3299 1038 3361 1076
rect 3965 1436 3979 1470
rect 4013 1436 4027 1470
rect 4409 1470 4471 1505
rect 3965 1398 4027 1436
rect 3965 1364 3979 1398
rect 4013 1364 4027 1398
rect 3965 1326 4027 1364
rect 3965 1292 3979 1326
rect 4013 1292 4027 1326
rect 3965 1254 4027 1292
rect 3965 1220 3979 1254
rect 4013 1220 4027 1254
rect 3965 1182 4027 1220
rect 3965 1148 3979 1182
rect 4013 1148 4027 1182
rect 3965 1110 4027 1148
rect 3965 1076 3979 1110
rect 4013 1076 4027 1110
rect 3299 1004 3313 1038
rect 3347 1004 3361 1038
rect 3299 966 3361 1004
rect 2633 930 2695 932
rect 3299 932 3313 966
rect 3347 932 3361 966
rect 3965 1038 4027 1076
rect 4409 1436 4423 1470
rect 4457 1436 4471 1470
rect 5075 1470 5137 1505
rect 4409 1398 4471 1436
rect 4409 1364 4423 1398
rect 4457 1364 4471 1398
rect 4409 1326 4471 1364
rect 4409 1292 4423 1326
rect 4457 1292 4471 1326
rect 4409 1254 4471 1292
rect 4409 1220 4423 1254
rect 4457 1220 4471 1254
rect 4409 1182 4471 1220
rect 4409 1148 4423 1182
rect 4457 1148 4471 1182
rect 4409 1110 4471 1148
rect 4409 1076 4423 1110
rect 4457 1076 4471 1110
rect 3965 1004 3979 1038
rect 4013 1004 4027 1038
rect 3965 966 4027 1004
rect 4409 1038 4471 1076
rect 5075 1436 5089 1470
rect 5123 1436 5137 1470
rect 5519 1470 5581 1505
rect 5075 1398 5137 1436
rect 5075 1364 5089 1398
rect 5123 1364 5137 1398
rect 5075 1326 5137 1364
rect 5075 1292 5089 1326
rect 5123 1292 5137 1326
rect 5075 1254 5137 1292
rect 5075 1220 5089 1254
rect 5123 1220 5137 1254
rect 5075 1182 5137 1220
rect 5075 1148 5089 1182
rect 5123 1148 5137 1182
rect 5075 1110 5137 1148
rect 5075 1076 5089 1110
rect 5123 1076 5137 1110
rect 3299 930 3361 932
rect 3965 932 3979 966
rect 4013 932 4027 966
rect 4409 1004 4423 1038
rect 4457 1004 4471 1038
rect 4409 966 4471 1004
rect 3965 930 4027 932
rect 4409 932 4423 966
rect 4457 932 4471 966
rect 5075 1038 5137 1076
rect 5519 1436 5533 1470
rect 5567 1436 5581 1470
rect 6185 1470 6247 1505
rect 5519 1398 5581 1436
rect 5519 1364 5533 1398
rect 5567 1364 5581 1398
rect 5519 1326 5581 1364
rect 5519 1292 5533 1326
rect 5567 1292 5581 1326
rect 5519 1254 5581 1292
rect 5519 1220 5533 1254
rect 5567 1220 5581 1254
rect 5519 1182 5581 1220
rect 5519 1148 5533 1182
rect 5567 1148 5581 1182
rect 5519 1110 5581 1148
rect 5519 1076 5533 1110
rect 5567 1076 5581 1110
rect 5075 1004 5089 1038
rect 5123 1004 5137 1038
rect 5075 966 5137 1004
rect 4409 930 4471 932
rect 5075 932 5089 966
rect 5123 932 5137 966
rect 5519 1038 5581 1076
rect 6185 1436 6199 1470
rect 6233 1436 6247 1470
rect 6629 1470 6691 1505
rect 6185 1398 6247 1436
rect 6185 1364 6199 1398
rect 6233 1364 6247 1398
rect 6185 1326 6247 1364
rect 6185 1292 6199 1326
rect 6233 1292 6247 1326
rect 6185 1254 6247 1292
rect 6185 1220 6199 1254
rect 6233 1220 6247 1254
rect 6185 1182 6247 1220
rect 6185 1148 6199 1182
rect 6233 1148 6247 1182
rect 6185 1110 6247 1148
rect 6185 1076 6199 1110
rect 6233 1076 6247 1110
rect 5519 1004 5533 1038
rect 5567 1004 5581 1038
rect 5519 966 5581 1004
rect 5075 930 5137 932
rect 5519 932 5533 966
rect 5567 932 5581 966
rect 6185 1038 6247 1076
rect 6629 1436 6643 1470
rect 6677 1436 6691 1470
rect 7295 1470 7357 1505
rect 6629 1398 6691 1436
rect 6629 1364 6643 1398
rect 6677 1364 6691 1398
rect 6629 1326 6691 1364
rect 6629 1292 6643 1326
rect 6677 1292 6691 1326
rect 6629 1254 6691 1292
rect 6629 1220 6643 1254
rect 6677 1220 6691 1254
rect 6629 1182 6691 1220
rect 6629 1148 6643 1182
rect 6677 1148 6691 1182
rect 6629 1110 6691 1148
rect 6629 1076 6643 1110
rect 6677 1076 6691 1110
rect 6185 1004 6199 1038
rect 6233 1004 6247 1038
rect 6185 966 6247 1004
rect 5519 930 5581 932
rect 6185 932 6199 966
rect 6233 932 6247 966
rect 6629 1038 6691 1076
rect 7295 1436 7309 1470
rect 7343 1436 7357 1470
rect 7739 1470 7801 1505
rect 7295 1398 7357 1436
rect 7295 1364 7309 1398
rect 7343 1364 7357 1398
rect 7295 1326 7357 1364
rect 7295 1292 7309 1326
rect 7343 1292 7357 1326
rect 7295 1254 7357 1292
rect 7295 1220 7309 1254
rect 7343 1220 7357 1254
rect 7295 1182 7357 1220
rect 7295 1148 7309 1182
rect 7343 1148 7357 1182
rect 7295 1110 7357 1148
rect 7295 1076 7309 1110
rect 7343 1076 7357 1110
rect 6629 1004 6643 1038
rect 6677 1004 6691 1038
rect 6629 966 6691 1004
rect 6185 930 6247 932
rect 6629 932 6643 966
rect 6677 932 6691 966
rect 7295 1038 7357 1076
rect 7739 1436 7753 1470
rect 7787 1436 7801 1470
rect 7739 1398 7801 1436
rect 7739 1364 7753 1398
rect 7787 1364 7801 1398
rect 7739 1326 7801 1364
rect 7739 1292 7753 1326
rect 7787 1292 7801 1326
rect 7739 1254 7801 1292
rect 7739 1220 7753 1254
rect 7787 1220 7801 1254
rect 7739 1182 7801 1220
rect 7739 1148 7753 1182
rect 7787 1148 7801 1182
rect 7739 1110 7801 1148
rect 7739 1076 7753 1110
rect 7787 1076 7801 1110
rect 7295 1004 7309 1038
rect 7343 1004 7357 1038
rect 7295 966 7357 1004
rect 6629 930 6691 932
rect 7295 932 7309 966
rect 7343 932 7357 966
rect 7739 1038 7801 1076
rect 7739 1004 7753 1038
rect 7787 1004 7801 1038
rect 7739 966 7801 1004
rect 7295 930 7357 932
rect 7739 932 7753 966
rect 7787 932 7801 966
rect 7739 930 7801 932
rect -31 868 7801 930
<< psubdiffcont >>
rect -17 512 17 546
rect 427 512 461 546
rect 1093 512 1127 546
rect 1759 512 1793 546
rect 2203 512 2237 546
rect 2647 512 2681 546
rect 3313 512 3347 546
rect 3979 512 4013 546
rect 4423 512 4457 546
rect 5089 512 5123 546
rect 5533 512 5567 546
rect 6199 512 6233 546
rect 6643 512 6677 546
rect 7309 512 7343 546
rect 7753 512 7787 546
rect -17 440 17 474
rect -17 368 17 402
rect 427 440 461 474
rect -17 296 17 330
rect -17 224 17 258
rect -17 152 17 186
rect -17 80 17 114
rect 427 368 461 402
rect 1093 440 1127 474
rect 427 296 461 330
rect 427 224 461 258
rect 427 152 461 186
rect 427 80 461 114
rect 1093 368 1127 402
rect 1759 440 1793 474
rect 1093 296 1127 330
rect 1093 224 1127 258
rect 1093 152 1127 186
rect 1093 80 1127 114
rect 1759 368 1793 402
rect 2203 440 2237 474
rect 1759 296 1793 330
rect 1759 224 1793 258
rect 1759 152 1793 186
rect 1759 80 1793 114
rect 2203 368 2237 402
rect 2647 440 2681 474
rect 2203 296 2237 330
rect 2203 224 2237 258
rect 2203 152 2237 186
rect 2203 80 2237 114
rect 2647 368 2681 402
rect 3313 440 3347 474
rect 2647 296 2681 330
rect 2647 224 2681 258
rect 2647 152 2681 186
rect 2647 80 2681 114
rect 3313 368 3347 402
rect 3979 440 4013 474
rect 3313 296 3347 330
rect 3313 224 3347 258
rect 3313 152 3347 186
rect 3313 80 3347 114
rect 3979 368 4013 402
rect 4423 440 4457 474
rect 3979 296 4013 330
rect 3979 224 4013 258
rect 3979 152 4013 186
rect 3979 80 4013 114
rect 4423 368 4457 402
rect 5089 440 5123 474
rect 4423 296 4457 330
rect 4423 224 4457 258
rect 4423 152 4457 186
rect 4423 80 4457 114
rect 5089 368 5123 402
rect 5533 440 5567 474
rect 5089 296 5123 330
rect 5089 224 5123 258
rect 5089 152 5123 186
rect 5089 80 5123 114
rect 5533 368 5567 402
rect 6199 440 6233 474
rect 5533 296 5567 330
rect 5533 224 5567 258
rect 5533 152 5567 186
rect 5533 80 5567 114
rect 6199 368 6233 402
rect 6643 440 6677 474
rect 6199 296 6233 330
rect 6199 224 6233 258
rect 6199 152 6233 186
rect 6199 80 6233 114
rect 6643 368 6677 402
rect 7309 440 7343 474
rect 6643 296 6677 330
rect 6643 224 6677 258
rect 6643 152 6677 186
rect 6643 80 6677 114
rect 7309 368 7343 402
rect 7753 440 7787 474
rect 7309 296 7343 330
rect 7309 224 7343 258
rect 7309 152 7343 186
rect 7309 80 7343 114
rect 7753 368 7787 402
rect 7753 296 7787 330
rect 7753 224 7787 258
rect 7753 152 7787 186
rect 7753 80 7787 114
rect 55 13 89 47
rect 127 13 161 47
rect 205 13 239 47
rect 283 13 317 47
rect 355 13 389 47
rect 499 13 533 47
rect 571 13 605 47
rect 643 13 677 47
rect 715 13 749 47
rect 805 13 839 47
rect 877 13 911 47
rect 949 13 983 47
rect 1021 13 1055 47
rect 1165 13 1199 47
rect 1237 13 1271 47
rect 1309 13 1343 47
rect 1381 13 1415 47
rect 1471 13 1505 47
rect 1543 13 1577 47
rect 1615 13 1649 47
rect 1687 13 1721 47
rect 1831 13 1865 47
rect 1903 13 1937 47
rect 1981 13 2015 47
rect 2059 13 2093 47
rect 2131 13 2165 47
rect 2275 13 2309 47
rect 2347 13 2381 47
rect 2425 13 2459 47
rect 2503 13 2537 47
rect 2575 13 2609 47
rect 2719 13 2753 47
rect 2791 13 2825 47
rect 2863 13 2897 47
rect 2935 13 2969 47
rect 3025 13 3059 47
rect 3097 13 3131 47
rect 3169 13 3203 47
rect 3241 13 3275 47
rect 3385 13 3419 47
rect 3457 13 3491 47
rect 3529 13 3563 47
rect 3601 13 3635 47
rect 3691 13 3725 47
rect 3763 13 3797 47
rect 3835 13 3869 47
rect 3907 13 3941 47
rect 4051 13 4085 47
rect 4123 13 4157 47
rect 4201 13 4235 47
rect 4279 13 4313 47
rect 4351 13 4385 47
rect 4495 13 4529 47
rect 4567 13 4601 47
rect 4639 13 4673 47
rect 4711 13 4745 47
rect 4801 13 4835 47
rect 4873 13 4907 47
rect 4945 13 4979 47
rect 5017 13 5051 47
rect 5161 13 5195 47
rect 5233 13 5267 47
rect 5311 13 5345 47
rect 5389 13 5423 47
rect 5461 13 5495 47
rect 5605 13 5639 47
rect 5677 13 5711 47
rect 5749 13 5783 47
rect 5821 13 5855 47
rect 5911 13 5945 47
rect 5983 13 6017 47
rect 6055 13 6089 47
rect 6127 13 6161 47
rect 6271 13 6305 47
rect 6343 13 6377 47
rect 6421 13 6455 47
rect 6499 13 6533 47
rect 6571 13 6605 47
rect 6715 13 6749 47
rect 6787 13 6821 47
rect 6859 13 6893 47
rect 6931 13 6965 47
rect 7021 13 7055 47
rect 7093 13 7127 47
rect 7165 13 7199 47
rect 7237 13 7271 47
rect 7381 13 7415 47
rect 7453 13 7487 47
rect 7531 13 7565 47
rect 7609 13 7643 47
rect 7681 13 7715 47
<< nsubdiffcont >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 205 1505 239 1539
rect 283 1505 317 1539
rect 355 1505 389 1539
rect 499 1505 533 1539
rect 571 1505 605 1539
rect 643 1505 677 1539
rect 715 1505 749 1539
rect 805 1505 839 1539
rect 877 1505 911 1539
rect 949 1505 983 1539
rect 1021 1505 1055 1539
rect 1165 1505 1199 1539
rect 1237 1505 1271 1539
rect 1309 1505 1343 1539
rect 1381 1505 1415 1539
rect 1471 1505 1505 1539
rect 1543 1505 1577 1539
rect 1615 1505 1649 1539
rect 1687 1505 1721 1539
rect 1831 1505 1865 1539
rect 1903 1505 1937 1539
rect 1981 1505 2015 1539
rect 2059 1505 2093 1539
rect 2131 1505 2165 1539
rect 2275 1505 2309 1539
rect 2347 1505 2381 1539
rect 2425 1505 2459 1539
rect 2503 1505 2537 1539
rect 2575 1505 2609 1539
rect 2719 1505 2753 1539
rect 2791 1505 2825 1539
rect 2863 1505 2897 1539
rect 2935 1505 2969 1539
rect 3025 1505 3059 1539
rect 3097 1505 3131 1539
rect 3169 1505 3203 1539
rect 3241 1505 3275 1539
rect 3385 1505 3419 1539
rect 3457 1505 3491 1539
rect 3529 1505 3563 1539
rect 3601 1505 3635 1539
rect 3691 1505 3725 1539
rect 3763 1505 3797 1539
rect 3835 1505 3869 1539
rect 3907 1505 3941 1539
rect 4051 1505 4085 1539
rect 4123 1505 4157 1539
rect 4201 1505 4235 1539
rect 4279 1505 4313 1539
rect 4351 1505 4385 1539
rect 4495 1505 4529 1539
rect 4567 1505 4601 1539
rect 4639 1505 4673 1539
rect 4711 1505 4745 1539
rect 4801 1505 4835 1539
rect 4873 1505 4907 1539
rect 4945 1505 4979 1539
rect 5017 1505 5051 1539
rect 5161 1505 5195 1539
rect 5233 1505 5267 1539
rect 5311 1505 5345 1539
rect 5389 1505 5423 1539
rect 5461 1505 5495 1539
rect 5605 1505 5639 1539
rect 5677 1505 5711 1539
rect 5749 1505 5783 1539
rect 5821 1505 5855 1539
rect 5911 1505 5945 1539
rect 5983 1505 6017 1539
rect 6055 1505 6089 1539
rect 6127 1505 6161 1539
rect 6271 1505 6305 1539
rect 6343 1505 6377 1539
rect 6421 1505 6455 1539
rect 6499 1505 6533 1539
rect 6571 1505 6605 1539
rect 6715 1505 6749 1539
rect 6787 1505 6821 1539
rect 6859 1505 6893 1539
rect 6931 1505 6965 1539
rect 7021 1505 7055 1539
rect 7093 1505 7127 1539
rect 7165 1505 7199 1539
rect 7237 1505 7271 1539
rect 7381 1505 7415 1539
rect 7453 1505 7487 1539
rect 7531 1505 7565 1539
rect 7609 1505 7643 1539
rect 7681 1505 7715 1539
rect -17 1436 17 1470
rect -17 1364 17 1398
rect -17 1292 17 1326
rect -17 1220 17 1254
rect -17 1148 17 1182
rect -17 1076 17 1110
rect 427 1436 461 1470
rect 427 1364 461 1398
rect 427 1292 461 1326
rect 427 1220 461 1254
rect 427 1148 461 1182
rect 427 1076 461 1110
rect -17 1004 17 1038
rect -17 932 17 966
rect 1093 1436 1127 1470
rect 1093 1364 1127 1398
rect 1093 1292 1127 1326
rect 1093 1220 1127 1254
rect 1093 1148 1127 1182
rect 1093 1076 1127 1110
rect 427 1004 461 1038
rect 427 932 461 966
rect 1759 1436 1793 1470
rect 1759 1364 1793 1398
rect 1759 1292 1793 1326
rect 1759 1220 1793 1254
rect 1759 1148 1793 1182
rect 1759 1076 1793 1110
rect 1093 1004 1127 1038
rect 1093 932 1127 966
rect 2203 1436 2237 1470
rect 2203 1364 2237 1398
rect 2203 1292 2237 1326
rect 2203 1220 2237 1254
rect 2203 1148 2237 1182
rect 2203 1076 2237 1110
rect 1759 1004 1793 1038
rect 2647 1436 2681 1470
rect 2647 1364 2681 1398
rect 2647 1292 2681 1326
rect 2647 1220 2681 1254
rect 2647 1148 2681 1182
rect 2647 1076 2681 1110
rect 1759 932 1793 966
rect 2203 1004 2237 1038
rect 2203 932 2237 966
rect 3313 1436 3347 1470
rect 3313 1364 3347 1398
rect 3313 1292 3347 1326
rect 3313 1220 3347 1254
rect 3313 1148 3347 1182
rect 3313 1076 3347 1110
rect 2647 1004 2681 1038
rect 2647 932 2681 966
rect 3979 1436 4013 1470
rect 3979 1364 4013 1398
rect 3979 1292 4013 1326
rect 3979 1220 4013 1254
rect 3979 1148 4013 1182
rect 3979 1076 4013 1110
rect 3313 1004 3347 1038
rect 3313 932 3347 966
rect 4423 1436 4457 1470
rect 4423 1364 4457 1398
rect 4423 1292 4457 1326
rect 4423 1220 4457 1254
rect 4423 1148 4457 1182
rect 4423 1076 4457 1110
rect 3979 1004 4013 1038
rect 5089 1436 5123 1470
rect 5089 1364 5123 1398
rect 5089 1292 5123 1326
rect 5089 1220 5123 1254
rect 5089 1148 5123 1182
rect 5089 1076 5123 1110
rect 3979 932 4013 966
rect 4423 1004 4457 1038
rect 4423 932 4457 966
rect 5533 1436 5567 1470
rect 5533 1364 5567 1398
rect 5533 1292 5567 1326
rect 5533 1220 5567 1254
rect 5533 1148 5567 1182
rect 5533 1076 5567 1110
rect 5089 1004 5123 1038
rect 5089 932 5123 966
rect 6199 1436 6233 1470
rect 6199 1364 6233 1398
rect 6199 1292 6233 1326
rect 6199 1220 6233 1254
rect 6199 1148 6233 1182
rect 6199 1076 6233 1110
rect 5533 1004 5567 1038
rect 5533 932 5567 966
rect 6643 1436 6677 1470
rect 6643 1364 6677 1398
rect 6643 1292 6677 1326
rect 6643 1220 6677 1254
rect 6643 1148 6677 1182
rect 6643 1076 6677 1110
rect 6199 1004 6233 1038
rect 6199 932 6233 966
rect 7309 1436 7343 1470
rect 7309 1364 7343 1398
rect 7309 1292 7343 1326
rect 7309 1220 7343 1254
rect 7309 1148 7343 1182
rect 7309 1076 7343 1110
rect 6643 1004 6677 1038
rect 6643 932 6677 966
rect 7753 1436 7787 1470
rect 7753 1364 7787 1398
rect 7753 1292 7787 1326
rect 7753 1220 7787 1254
rect 7753 1148 7787 1182
rect 7753 1076 7787 1110
rect 7309 1004 7343 1038
rect 7309 932 7343 966
rect 7753 1004 7787 1038
rect 7753 932 7787 966
<< poly >>
rect 163 1450 193 1476
rect 251 1450 281 1476
rect 631 1451 661 1477
rect 719 1451 749 1477
rect 807 1451 837 1477
rect 895 1451 925 1477
rect 163 1019 193 1050
rect 251 1019 281 1050
rect 121 1003 281 1019
rect 121 969 131 1003
rect 165 989 281 1003
rect 1297 1451 1327 1477
rect 1385 1451 1415 1477
rect 1473 1451 1503 1477
rect 1561 1451 1591 1477
rect 165 969 175 989
rect 121 953 175 969
rect 631 1020 661 1051
rect 719 1020 749 1051
rect 631 1004 749 1020
rect 631 990 649 1004
rect 639 970 649 990
rect 683 990 749 1004
rect 807 1020 837 1051
rect 895 1020 925 1051
rect 807 1004 925 1020
rect 807 990 871 1004
rect 683 970 693 990
rect 639 954 693 970
rect 861 970 871 990
rect 905 990 925 1004
rect 1939 1450 1969 1476
rect 2027 1450 2057 1476
rect 905 970 915 990
rect 861 954 915 970
rect 1297 1020 1327 1051
rect 1385 1020 1415 1051
rect 1297 1004 1415 1020
rect 1297 990 1315 1004
rect 1305 970 1315 990
rect 1349 990 1415 1004
rect 1473 1020 1503 1051
rect 1561 1020 1591 1051
rect 1473 1004 1591 1020
rect 1473 990 1537 1004
rect 1349 970 1359 990
rect 1305 954 1359 970
rect 1527 970 1537 990
rect 1571 990 1591 1004
rect 2383 1450 2413 1476
rect 2471 1450 2501 1476
rect 1571 970 1581 990
rect 1527 954 1581 970
rect 1939 1019 1969 1050
rect 2027 1019 2057 1050
rect 2851 1451 2881 1477
rect 2939 1451 2969 1477
rect 3027 1451 3057 1477
rect 3115 1451 3145 1477
rect 1939 1003 2099 1019
rect 1939 989 2055 1003
rect 2045 969 2055 989
rect 2089 969 2099 1003
rect 2045 953 2099 969
rect 2383 1019 2413 1050
rect 2471 1019 2501 1050
rect 2341 1003 2501 1019
rect 2341 969 2351 1003
rect 2385 989 2501 1003
rect 3517 1451 3547 1477
rect 3605 1451 3635 1477
rect 3693 1451 3723 1477
rect 3781 1451 3811 1477
rect 2385 969 2395 989
rect 2341 953 2395 969
rect 2851 1020 2881 1051
rect 2939 1020 2969 1051
rect 2851 1004 2969 1020
rect 2851 990 2869 1004
rect 2859 970 2869 990
rect 2903 990 2969 1004
rect 3027 1020 3057 1051
rect 3115 1020 3145 1051
rect 3027 1004 3145 1020
rect 3027 990 3091 1004
rect 2903 970 2913 990
rect 2859 954 2913 970
rect 3081 970 3091 990
rect 3125 990 3145 1004
rect 4159 1450 4189 1476
rect 4247 1450 4277 1476
rect 3125 970 3135 990
rect 3081 954 3135 970
rect 3517 1020 3547 1051
rect 3605 1020 3635 1051
rect 3517 1004 3635 1020
rect 3517 990 3535 1004
rect 3525 970 3535 990
rect 3569 990 3635 1004
rect 3693 1020 3723 1051
rect 3781 1020 3811 1051
rect 3693 1004 3811 1020
rect 3693 990 3757 1004
rect 3569 970 3579 990
rect 3525 954 3579 970
rect 3747 970 3757 990
rect 3791 990 3811 1004
rect 4627 1450 4657 1476
rect 4715 1450 4745 1476
rect 4803 1450 4833 1476
rect 4891 1450 4921 1476
rect 3791 970 3801 990
rect 3747 954 3801 970
rect 4159 1019 4189 1050
rect 4247 1019 4277 1050
rect 5269 1450 5299 1476
rect 5357 1450 5387 1476
rect 4159 1003 4319 1019
rect 4159 989 4275 1003
rect 4265 969 4275 989
rect 4309 969 4319 1003
rect 4265 953 4319 969
rect 4627 1019 4657 1050
rect 4715 1019 4745 1050
rect 4803 1019 4833 1050
rect 4891 1019 4921 1050
rect 4627 1003 4745 1019
rect 4627 989 4645 1003
rect 4635 969 4645 989
rect 4679 989 4745 1003
rect 4789 1003 4921 1019
rect 4679 969 4689 989
rect 4635 953 4689 969
rect 4789 969 4799 1003
rect 4833 989 4921 1003
rect 5737 1450 5767 1476
rect 5825 1450 5855 1476
rect 5913 1450 5943 1476
rect 6001 1450 6031 1476
rect 5269 1019 5299 1050
rect 5357 1019 5387 1050
rect 4833 969 4843 989
rect 4789 953 4843 969
rect 5227 1003 5387 1019
rect 5227 969 5237 1003
rect 5271 989 5387 1003
rect 6379 1450 6409 1476
rect 6467 1450 6497 1476
rect 5271 969 5281 989
rect 5227 953 5281 969
rect 5737 1019 5767 1050
rect 5825 1019 5855 1050
rect 5913 1019 5943 1050
rect 6001 1019 6031 1050
rect 5737 1003 5855 1019
rect 5737 989 5755 1003
rect 5745 969 5755 989
rect 5789 989 5855 1003
rect 5899 1003 6031 1019
rect 5789 969 5799 989
rect 5745 953 5799 969
rect 5899 969 5909 1003
rect 5943 989 6031 1003
rect 6847 1451 6877 1477
rect 6935 1451 6965 1477
rect 7023 1451 7053 1477
rect 7111 1451 7141 1477
rect 6379 1019 6409 1050
rect 6467 1019 6497 1050
rect 5943 969 5953 989
rect 5899 953 5953 969
rect 6337 1003 6497 1019
rect 6337 969 6347 1003
rect 6381 989 6497 1003
rect 7489 1450 7519 1476
rect 7577 1450 7607 1476
rect 6847 1020 6877 1051
rect 6935 1020 6965 1051
rect 7023 1020 7053 1051
rect 7111 1020 7141 1051
rect 6381 969 6391 989
rect 6337 953 6391 969
rect 6824 1004 6965 1020
rect 6824 970 6834 1004
rect 6868 990 6965 1004
rect 7010 1004 7141 1020
rect 6868 970 6878 990
rect 6824 954 6878 970
rect 7010 970 7020 1004
rect 7054 990 7141 1004
rect 7489 1019 7519 1050
rect 7577 1019 7607 1050
rect 7054 970 7064 990
rect 7010 954 7064 970
rect 7447 1003 7607 1019
rect 7447 969 7457 1003
rect 7491 989 7607 1003
rect 7491 969 7501 989
rect 7447 953 7501 969
rect 121 461 175 477
rect 121 427 131 461
rect 165 441 175 461
rect 165 427 185 441
rect 121 411 185 427
rect 155 377 185 411
rect 639 461 693 477
rect 639 441 649 461
rect 612 427 649 441
rect 683 427 693 461
rect 861 461 915 477
rect 861 441 871 461
rect 612 411 693 427
rect 806 427 871 441
rect 905 427 915 461
rect 806 411 915 427
rect 1305 461 1359 477
rect 1305 441 1315 461
rect 612 377 642 411
rect 806 377 836 411
rect 1278 427 1315 441
rect 1349 427 1359 461
rect 1527 461 1581 477
rect 1527 441 1537 461
rect 1278 411 1359 427
rect 1472 427 1537 441
rect 1571 427 1581 461
rect 1472 411 1581 427
rect 2045 461 2099 477
rect 2045 441 2055 461
rect 1278 377 1308 411
rect 1472 377 1502 411
rect 2035 427 2055 441
rect 2089 427 2099 461
rect 2035 411 2099 427
rect 2035 377 2065 411
rect 2341 461 2395 477
rect 2341 427 2351 461
rect 2385 441 2395 461
rect 2385 427 2405 441
rect 2341 411 2405 427
rect 2375 377 2405 411
rect 2859 461 2913 477
rect 2859 441 2869 461
rect 2832 427 2869 441
rect 2903 427 2913 461
rect 3081 461 3135 477
rect 3081 441 3091 461
rect 2832 411 2913 427
rect 3026 427 3091 441
rect 3125 427 3135 461
rect 3026 411 3135 427
rect 3525 461 3579 477
rect 3525 441 3535 461
rect 2832 377 2862 411
rect 3026 377 3056 411
rect 3498 427 3535 441
rect 3569 427 3579 461
rect 3747 461 3801 477
rect 3747 441 3757 461
rect 3498 411 3579 427
rect 3692 427 3757 441
rect 3791 427 3801 461
rect 3692 411 3801 427
rect 4265 461 4319 477
rect 4265 441 4275 461
rect 3498 377 3528 411
rect 3692 377 3722 411
rect 4255 427 4275 441
rect 4309 427 4319 461
rect 4255 411 4319 427
rect 4635 461 4689 477
rect 4635 441 4645 461
rect 4255 377 4285 411
rect 4608 427 4645 441
rect 4679 427 4689 461
rect 4608 411 4689 427
rect 4783 461 4837 477
rect 4783 427 4793 461
rect 4827 427 4837 461
rect 4783 411 4837 427
rect 4608 377 4638 411
rect 4802 377 4832 411
rect 5227 461 5281 477
rect 5227 427 5237 461
rect 5271 441 5281 461
rect 5271 427 5291 441
rect 5227 411 5291 427
rect 5261 377 5291 411
rect 5745 461 5799 477
rect 5745 441 5755 461
rect 5718 427 5755 441
rect 5789 427 5799 461
rect 5718 411 5799 427
rect 5893 461 5947 477
rect 5893 427 5903 461
rect 5937 427 5947 461
rect 5893 411 5947 427
rect 5718 377 5748 411
rect 5912 377 5942 411
rect 6337 461 6391 477
rect 6337 427 6347 461
rect 6381 441 6391 461
rect 6381 427 6401 441
rect 6337 411 6401 427
rect 6371 377 6401 411
rect 6855 461 6909 477
rect 6855 441 6865 461
rect 6828 427 6865 441
rect 6899 427 6909 461
rect 6828 411 6909 427
rect 7003 461 7057 477
rect 7003 427 7013 461
rect 7047 427 7057 461
rect 7003 411 7057 427
rect 6828 377 6858 411
rect 7022 377 7052 411
rect 7447 461 7501 477
rect 7447 427 7457 461
rect 7491 441 7501 461
rect 7491 427 7511 441
rect 7447 411 7511 427
rect 7481 377 7511 411
<< polycont >>
rect 131 969 165 1003
rect 649 970 683 1004
rect 871 970 905 1004
rect 1315 970 1349 1004
rect 1537 970 1571 1004
rect 2055 969 2089 1003
rect 2351 969 2385 1003
rect 2869 970 2903 1004
rect 3091 970 3125 1004
rect 3535 970 3569 1004
rect 3757 970 3791 1004
rect 4275 969 4309 1003
rect 4645 969 4679 1003
rect 4799 969 4833 1003
rect 5237 969 5271 1003
rect 5755 969 5789 1003
rect 5909 969 5943 1003
rect 6347 969 6381 1003
rect 6834 970 6868 1004
rect 7020 970 7054 1004
rect 7457 969 7491 1003
rect 131 427 165 461
rect 649 427 683 461
rect 871 427 905 461
rect 1315 427 1349 461
rect 1537 427 1571 461
rect 2055 427 2089 461
rect 2351 427 2385 461
rect 2869 427 2903 461
rect 3091 427 3125 461
rect 3535 427 3569 461
rect 3757 427 3791 461
rect 4275 427 4309 461
rect 4645 427 4679 461
rect 4793 427 4827 461
rect 5237 427 5271 461
rect 5755 427 5789 461
rect 5903 427 5937 461
rect 6347 427 6381 461
rect 6865 427 6899 461
rect 7013 427 7047 461
rect 7457 427 7491 461
<< locali >>
rect -31 1539 7801 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 205 1539
rect 239 1505 283 1539
rect 317 1505 355 1539
rect 389 1505 499 1539
rect 533 1505 571 1539
rect 605 1505 643 1539
rect 677 1505 715 1539
rect 749 1505 805 1539
rect 839 1505 877 1539
rect 911 1505 949 1539
rect 983 1505 1021 1539
rect 1055 1505 1165 1539
rect 1199 1505 1237 1539
rect 1271 1505 1309 1539
rect 1343 1505 1381 1539
rect 1415 1505 1471 1539
rect 1505 1505 1543 1539
rect 1577 1505 1615 1539
rect 1649 1505 1687 1539
rect 1721 1505 1831 1539
rect 1865 1505 1903 1539
rect 1937 1505 1981 1539
rect 2015 1505 2059 1539
rect 2093 1505 2131 1539
rect 2165 1505 2275 1539
rect 2309 1505 2347 1539
rect 2381 1505 2425 1539
rect 2459 1505 2503 1539
rect 2537 1505 2575 1539
rect 2609 1505 2719 1539
rect 2753 1505 2791 1539
rect 2825 1505 2863 1539
rect 2897 1505 2935 1539
rect 2969 1505 3025 1539
rect 3059 1505 3097 1539
rect 3131 1505 3169 1539
rect 3203 1505 3241 1539
rect 3275 1505 3385 1539
rect 3419 1505 3457 1539
rect 3491 1505 3529 1539
rect 3563 1505 3601 1539
rect 3635 1505 3691 1539
rect 3725 1505 3763 1539
rect 3797 1505 3835 1539
rect 3869 1505 3907 1539
rect 3941 1505 4051 1539
rect 4085 1505 4123 1539
rect 4157 1505 4201 1539
rect 4235 1505 4279 1539
rect 4313 1505 4351 1539
rect 4385 1505 4495 1539
rect 4529 1505 4567 1539
rect 4601 1505 4639 1539
rect 4673 1505 4711 1539
rect 4745 1505 4801 1539
rect 4835 1505 4873 1539
rect 4907 1505 4945 1539
rect 4979 1505 5017 1539
rect 5051 1505 5161 1539
rect 5195 1505 5233 1539
rect 5267 1505 5311 1539
rect 5345 1505 5389 1539
rect 5423 1505 5461 1539
rect 5495 1505 5605 1539
rect 5639 1505 5677 1539
rect 5711 1505 5749 1539
rect 5783 1505 5821 1539
rect 5855 1505 5911 1539
rect 5945 1505 5983 1539
rect 6017 1505 6055 1539
rect 6089 1505 6127 1539
rect 6161 1505 6271 1539
rect 6305 1505 6343 1539
rect 6377 1505 6421 1539
rect 6455 1505 6499 1539
rect 6533 1505 6571 1539
rect 6605 1505 6715 1539
rect 6749 1505 6787 1539
rect 6821 1505 6859 1539
rect 6893 1505 6931 1539
rect 6965 1505 7021 1539
rect 7055 1505 7093 1539
rect 7127 1505 7165 1539
rect 7199 1505 7237 1539
rect 7271 1505 7381 1539
rect 7415 1505 7453 1539
rect 7487 1505 7531 1539
rect 7565 1505 7609 1539
rect 7643 1505 7681 1539
rect 7715 1505 7801 1539
rect -31 1492 7801 1505
rect -31 1470 31 1492
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect 117 1412 151 1492
rect 117 1344 151 1378
rect 117 1276 151 1310
rect 117 1208 151 1242
rect 117 1139 151 1174
rect 117 1083 151 1105
rect 205 1412 239 1450
rect 205 1344 239 1378
rect 205 1276 239 1310
rect 205 1208 239 1242
rect 205 1139 239 1174
rect -31 1038 31 1076
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect -31 868 31 932
rect 131 1003 165 1019
rect 131 905 165 969
rect 205 979 239 1105
rect 293 1412 327 1492
rect 293 1344 327 1378
rect 293 1276 327 1310
rect 293 1208 327 1242
rect 293 1139 327 1174
rect 293 1083 327 1105
rect 413 1470 475 1492
rect 413 1436 427 1470
rect 461 1436 475 1470
rect 413 1398 475 1436
rect 413 1364 427 1398
rect 461 1364 475 1398
rect 413 1326 475 1364
rect 413 1292 427 1326
rect 461 1292 475 1326
rect 413 1254 475 1292
rect 413 1220 427 1254
rect 461 1220 475 1254
rect 413 1182 475 1220
rect 413 1148 427 1182
rect 461 1148 475 1182
rect 413 1110 475 1148
rect 413 1076 427 1110
rect 461 1076 475 1110
rect 413 1038 475 1076
rect 585 1411 619 1427
rect 585 1343 619 1377
rect 585 1275 619 1309
rect 585 1207 619 1241
rect 585 1139 619 1173
rect 673 1343 707 1492
rect 1079 1470 1141 1492
rect 673 1275 707 1309
rect 673 1207 707 1241
rect 673 1157 707 1173
rect 761 1411 971 1445
rect 761 1343 795 1377
rect 761 1275 795 1309
rect 761 1207 795 1241
rect 761 1139 795 1173
rect 585 1071 795 1105
rect 849 1343 883 1359
rect 849 1275 883 1309
rect 849 1207 883 1241
rect 849 1139 883 1173
rect 937 1343 971 1377
rect 937 1275 971 1309
rect 937 1207 971 1241
rect 937 1157 971 1173
rect 1079 1436 1093 1470
rect 1127 1436 1141 1470
rect 1079 1398 1141 1436
rect 1079 1364 1093 1398
rect 1127 1364 1141 1398
rect 1079 1326 1141 1364
rect 1079 1292 1093 1326
rect 1127 1292 1141 1326
rect 1079 1254 1141 1292
rect 1079 1220 1093 1254
rect 1127 1220 1141 1254
rect 1079 1182 1141 1220
rect 1079 1148 1093 1182
rect 1127 1148 1141 1182
rect 1079 1110 1141 1148
rect 849 1071 979 1105
rect 413 1004 427 1038
rect 461 1004 475 1038
rect 205 945 313 979
rect -31 546 31 572
rect -31 512 -17 546
rect 17 512 31 546
rect -31 474 31 512
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect 131 461 165 871
rect 279 683 313 945
rect 413 966 475 1004
rect 413 932 427 966
rect 461 932 475 966
rect 413 868 475 932
rect 649 1004 683 1020
rect 649 905 683 970
rect 279 461 313 649
rect 131 411 165 427
rect 205 427 313 461
rect 413 546 475 572
rect 413 512 427 546
rect 461 512 475 546
rect 413 474 475 512
rect 413 440 427 474
rect 461 440 475 474
rect 649 461 683 871
rect 871 1004 905 1020
rect 871 831 905 970
rect 871 781 905 797
rect 945 757 979 1071
rect 1079 1076 1093 1110
rect 1127 1076 1141 1110
rect 1079 1038 1141 1076
rect 1251 1411 1285 1427
rect 1251 1343 1285 1377
rect 1251 1275 1285 1309
rect 1251 1207 1285 1241
rect 1251 1139 1285 1173
rect 1339 1343 1373 1492
rect 1745 1470 1807 1492
rect 1339 1275 1373 1309
rect 1339 1207 1373 1241
rect 1339 1157 1373 1173
rect 1427 1411 1637 1445
rect 1427 1343 1461 1377
rect 1427 1275 1461 1309
rect 1427 1207 1461 1241
rect 1427 1139 1461 1173
rect 1251 1071 1461 1105
rect 1515 1343 1549 1359
rect 1515 1275 1549 1309
rect 1515 1207 1549 1241
rect 1515 1139 1549 1173
rect 1603 1343 1637 1377
rect 1603 1275 1637 1309
rect 1603 1207 1637 1241
rect 1603 1157 1637 1173
rect 1745 1436 1759 1470
rect 1793 1436 1807 1470
rect 1745 1398 1807 1436
rect 1745 1364 1759 1398
rect 1793 1364 1807 1398
rect 1745 1326 1807 1364
rect 1745 1292 1759 1326
rect 1793 1292 1807 1326
rect 1745 1254 1807 1292
rect 1745 1220 1759 1254
rect 1793 1220 1807 1254
rect 1745 1182 1807 1220
rect 1745 1148 1759 1182
rect 1793 1148 1807 1182
rect 1745 1110 1807 1148
rect 1515 1071 1645 1105
rect 1079 1004 1093 1038
rect 1127 1004 1141 1038
rect 1079 966 1141 1004
rect 1079 932 1093 966
rect 1127 932 1141 966
rect 1079 868 1141 932
rect 1315 1004 1349 1020
rect 1315 905 1349 970
rect 1315 855 1349 871
rect 1537 1004 1571 1020
rect 871 535 905 551
rect 871 461 905 501
rect -31 368 -17 402
rect 17 368 31 402
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect -31 62 31 80
rect 109 361 143 377
rect 109 289 143 327
rect 109 221 143 255
rect 205 245 239 427
rect 413 402 475 440
rect 633 427 649 461
rect 683 427 699 461
rect 649 411 683 427
rect 871 411 905 427
rect 205 195 239 211
rect 303 361 337 377
rect 303 289 337 327
rect 303 221 337 255
rect 109 151 143 187
rect 303 151 337 187
rect 143 117 205 151
rect 239 117 303 151
rect 109 62 143 117
rect 206 62 240 117
rect 303 62 337 117
rect 413 368 427 402
rect 461 368 475 402
rect 413 330 475 368
rect 413 296 427 330
rect 461 296 475 330
rect 413 258 475 296
rect 413 224 427 258
rect 461 224 475 258
rect 413 186 475 224
rect 413 152 427 186
rect 461 152 475 186
rect 413 114 475 152
rect 413 80 427 114
rect 461 80 475 114
rect 566 361 600 377
rect 760 361 794 377
rect 945 375 979 723
rect 1537 683 1571 970
rect 1315 609 1349 625
rect 600 327 663 361
rect 697 327 760 361
rect 566 289 600 327
rect 566 221 600 255
rect 760 289 794 327
rect 566 151 600 187
rect 566 101 600 117
rect 663 236 697 252
rect 413 62 475 80
rect 663 62 697 202
rect 760 221 794 255
rect 857 341 979 375
rect 1079 546 1141 572
rect 1079 512 1093 546
rect 1127 512 1141 546
rect 1079 474 1141 512
rect 1079 440 1093 474
rect 1127 440 1141 474
rect 1079 402 1141 440
rect 1315 461 1349 575
rect 1315 411 1349 427
rect 1537 461 1571 649
rect 1537 411 1571 427
rect 1611 757 1645 1071
rect 1745 1076 1759 1110
rect 1793 1076 1807 1110
rect 1893 1412 1927 1492
rect 1893 1344 1927 1378
rect 1893 1276 1927 1310
rect 1893 1208 1927 1242
rect 1893 1139 1927 1174
rect 1893 1083 1927 1105
rect 1981 1412 2015 1450
rect 1981 1344 2015 1378
rect 1981 1276 2015 1310
rect 1981 1208 2015 1242
rect 1981 1139 2015 1174
rect 1745 1038 1807 1076
rect 1745 1004 1759 1038
rect 1793 1004 1807 1038
rect 1745 966 1807 1004
rect 1981 979 2015 1105
rect 2069 1412 2103 1492
rect 2069 1344 2103 1378
rect 2069 1276 2103 1310
rect 2069 1208 2103 1242
rect 2069 1139 2103 1174
rect 2069 1083 2103 1105
rect 2189 1470 2251 1492
rect 2189 1436 2203 1470
rect 2237 1436 2251 1470
rect 2189 1398 2251 1436
rect 2189 1364 2203 1398
rect 2237 1364 2251 1398
rect 2189 1326 2251 1364
rect 2189 1292 2203 1326
rect 2237 1292 2251 1326
rect 2189 1254 2251 1292
rect 2189 1220 2203 1254
rect 2237 1220 2251 1254
rect 2189 1182 2251 1220
rect 2189 1148 2203 1182
rect 2237 1148 2251 1182
rect 2189 1110 2251 1148
rect 2189 1076 2203 1110
rect 2237 1076 2251 1110
rect 2337 1412 2371 1492
rect 2337 1344 2371 1378
rect 2337 1276 2371 1310
rect 2337 1208 2371 1242
rect 2337 1139 2371 1174
rect 2337 1083 2371 1105
rect 2425 1412 2459 1450
rect 2425 1344 2459 1378
rect 2425 1276 2459 1310
rect 2425 1208 2459 1242
rect 2425 1139 2459 1174
rect 2189 1038 2251 1076
rect 1745 932 1759 966
rect 1793 932 1807 966
rect 1745 868 1807 932
rect 1907 945 2015 979
rect 2055 1003 2089 1019
rect 1079 368 1093 402
rect 1127 368 1141 402
rect 857 245 891 341
rect 1079 330 1141 368
rect 857 195 891 211
rect 954 289 988 305
rect 954 221 988 255
rect 760 151 794 187
rect 954 151 988 187
rect 794 117 857 151
rect 891 117 954 151
rect 760 101 794 117
rect 954 101 988 117
rect 1079 296 1093 330
rect 1127 296 1141 330
rect 1079 258 1141 296
rect 1079 224 1093 258
rect 1127 224 1141 258
rect 1079 186 1141 224
rect 1079 152 1093 186
rect 1127 152 1141 186
rect 1079 114 1141 152
rect 1079 80 1093 114
rect 1127 80 1141 114
rect 1232 361 1266 377
rect 1426 361 1460 377
rect 1611 375 1645 723
rect 1907 831 1941 945
rect 1907 609 1941 797
rect 1266 327 1329 361
rect 1363 327 1426 361
rect 1232 289 1266 327
rect 1232 221 1266 255
rect 1426 289 1460 327
rect 1232 151 1266 187
rect 1232 101 1266 117
rect 1329 236 1363 252
rect 1079 62 1141 80
rect 1329 62 1363 202
rect 1426 221 1460 255
rect 1523 341 1645 375
rect 1745 546 1807 572
rect 1745 512 1759 546
rect 1793 512 1807 546
rect 1745 474 1807 512
rect 1745 440 1759 474
rect 1793 440 1807 474
rect 1745 402 1807 440
rect 1907 461 1941 575
rect 2055 905 2089 945
rect 2055 535 2089 871
rect 2189 1004 2203 1038
rect 2237 1004 2251 1038
rect 2189 966 2251 1004
rect 2189 932 2203 966
rect 2237 932 2251 966
rect 2189 868 2251 932
rect 2351 1003 2385 1019
rect 2351 905 2385 969
rect 2425 979 2459 1105
rect 2513 1412 2547 1492
rect 2513 1344 2547 1378
rect 2513 1276 2547 1310
rect 2513 1208 2547 1242
rect 2513 1139 2547 1174
rect 2513 1083 2547 1105
rect 2633 1470 2695 1492
rect 2633 1436 2647 1470
rect 2681 1436 2695 1470
rect 2633 1398 2695 1436
rect 2633 1364 2647 1398
rect 2681 1364 2695 1398
rect 2633 1326 2695 1364
rect 2633 1292 2647 1326
rect 2681 1292 2695 1326
rect 2633 1254 2695 1292
rect 2633 1220 2647 1254
rect 2681 1220 2695 1254
rect 2633 1182 2695 1220
rect 2633 1148 2647 1182
rect 2681 1148 2695 1182
rect 2633 1110 2695 1148
rect 2633 1076 2647 1110
rect 2681 1076 2695 1110
rect 2633 1038 2695 1076
rect 2805 1411 2839 1427
rect 2805 1343 2839 1377
rect 2805 1275 2839 1309
rect 2805 1207 2839 1241
rect 2805 1139 2839 1173
rect 2893 1343 2927 1492
rect 3299 1470 3361 1492
rect 2893 1275 2927 1309
rect 2893 1207 2927 1241
rect 2893 1157 2927 1173
rect 2981 1411 3191 1445
rect 2981 1343 3015 1377
rect 2981 1275 3015 1309
rect 2981 1207 3015 1241
rect 2981 1139 3015 1173
rect 2805 1071 3015 1105
rect 3069 1343 3103 1359
rect 3069 1275 3103 1309
rect 3069 1207 3103 1241
rect 3069 1139 3103 1173
rect 3157 1343 3191 1377
rect 3157 1275 3191 1309
rect 3157 1207 3191 1241
rect 3157 1157 3191 1173
rect 3299 1436 3313 1470
rect 3347 1436 3361 1470
rect 3299 1398 3361 1436
rect 3299 1364 3313 1398
rect 3347 1364 3361 1398
rect 3299 1326 3361 1364
rect 3299 1292 3313 1326
rect 3347 1292 3361 1326
rect 3299 1254 3361 1292
rect 3299 1220 3313 1254
rect 3347 1220 3361 1254
rect 3299 1182 3361 1220
rect 3299 1148 3313 1182
rect 3347 1148 3361 1182
rect 3299 1110 3361 1148
rect 3069 1071 3199 1105
rect 2633 1004 2647 1038
rect 2681 1004 2695 1038
rect 2425 945 2533 979
rect 2351 757 2385 871
rect 2055 461 2089 501
rect 1907 427 2015 461
rect 1745 368 1759 402
rect 1793 368 1807 402
rect 1523 245 1557 341
rect 1745 330 1807 368
rect 1523 195 1557 211
rect 1620 289 1654 305
rect 1620 221 1654 255
rect 1426 151 1460 187
rect 1620 151 1654 187
rect 1460 117 1523 151
rect 1557 117 1620 151
rect 1426 101 1460 117
rect 1620 101 1654 117
rect 1745 296 1759 330
rect 1793 296 1807 330
rect 1745 258 1807 296
rect 1745 224 1759 258
rect 1793 224 1807 258
rect 1745 186 1807 224
rect 1745 152 1759 186
rect 1793 152 1807 186
rect 1745 114 1807 152
rect 1745 80 1759 114
rect 1793 80 1807 114
rect 1745 62 1807 80
rect 1883 361 1917 377
rect 1883 289 1917 327
rect 1883 221 1917 255
rect 1981 245 2015 427
rect 2055 411 2089 427
rect 2189 546 2251 572
rect 2189 512 2203 546
rect 2237 512 2251 546
rect 2189 474 2251 512
rect 2189 440 2203 474
rect 2237 440 2251 474
rect 2189 402 2251 440
rect 2351 461 2385 723
rect 2499 683 2533 945
rect 2633 966 2695 1004
rect 2633 932 2647 966
rect 2681 932 2695 966
rect 2633 868 2695 932
rect 2869 1004 2903 1020
rect 2869 905 2903 970
rect 2499 461 2533 649
rect 2351 411 2385 427
rect 2425 427 2533 461
rect 2633 546 2695 572
rect 2633 512 2647 546
rect 2681 512 2695 546
rect 2633 474 2695 512
rect 2633 440 2647 474
rect 2681 440 2695 474
rect 1981 195 2015 211
rect 2077 361 2111 377
rect 2077 289 2111 327
rect 2077 221 2111 255
rect 1883 151 1917 187
rect 2077 151 2111 187
rect 1917 117 1981 151
rect 2015 117 2077 151
rect 1883 62 1917 117
rect 1980 62 2014 117
rect 2077 62 2111 117
rect 2189 368 2203 402
rect 2237 368 2251 402
rect 2189 330 2251 368
rect 2189 296 2203 330
rect 2237 296 2251 330
rect 2189 258 2251 296
rect 2189 224 2203 258
rect 2237 224 2251 258
rect 2189 186 2251 224
rect 2189 152 2203 186
rect 2237 152 2251 186
rect 2189 114 2251 152
rect 2189 80 2203 114
rect 2237 80 2251 114
rect 2189 62 2251 80
rect 2329 361 2363 377
rect 2329 289 2363 327
rect 2329 221 2363 255
rect 2425 245 2459 427
rect 2633 402 2695 440
rect 2869 461 2903 871
rect 3091 1004 3125 1020
rect 3091 831 3125 970
rect 3091 781 3125 797
rect 3165 757 3199 1071
rect 3299 1076 3313 1110
rect 3347 1076 3361 1110
rect 3299 1038 3361 1076
rect 3471 1411 3505 1427
rect 3471 1343 3505 1377
rect 3471 1275 3505 1309
rect 3471 1207 3505 1241
rect 3471 1139 3505 1173
rect 3559 1343 3593 1492
rect 3965 1470 4027 1492
rect 3559 1275 3593 1309
rect 3559 1207 3593 1241
rect 3559 1157 3593 1173
rect 3647 1411 3857 1445
rect 3647 1343 3681 1377
rect 3647 1275 3681 1309
rect 3647 1207 3681 1241
rect 3647 1139 3681 1173
rect 3471 1071 3681 1105
rect 3735 1343 3769 1359
rect 3735 1275 3769 1309
rect 3735 1207 3769 1241
rect 3735 1139 3769 1173
rect 3823 1343 3857 1377
rect 3823 1275 3857 1309
rect 3823 1207 3857 1241
rect 3823 1157 3857 1173
rect 3965 1436 3979 1470
rect 4013 1436 4027 1470
rect 3965 1398 4027 1436
rect 3965 1364 3979 1398
rect 4013 1364 4027 1398
rect 3965 1326 4027 1364
rect 3965 1292 3979 1326
rect 4013 1292 4027 1326
rect 3965 1254 4027 1292
rect 3965 1220 3979 1254
rect 4013 1220 4027 1254
rect 3965 1182 4027 1220
rect 3965 1148 3979 1182
rect 4013 1148 4027 1182
rect 3965 1110 4027 1148
rect 3735 1071 3865 1105
rect 3299 1004 3313 1038
rect 3347 1004 3361 1038
rect 3299 966 3361 1004
rect 3299 932 3313 966
rect 3347 932 3361 966
rect 3299 868 3361 932
rect 3535 1004 3569 1020
rect 3535 905 3569 970
rect 3535 855 3569 871
rect 3757 1004 3791 1020
rect 2869 411 2903 427
rect 3091 535 3125 551
rect 3091 461 3125 501
rect 3091 411 3125 427
rect 2425 195 2459 211
rect 2523 361 2557 377
rect 2523 289 2557 327
rect 2523 221 2557 255
rect 2329 151 2363 187
rect 2523 151 2557 187
rect 2363 117 2425 151
rect 2459 117 2523 151
rect 2329 62 2363 117
rect 2426 62 2460 117
rect 2523 62 2557 117
rect 2633 368 2647 402
rect 2681 368 2695 402
rect 2633 330 2695 368
rect 2633 296 2647 330
rect 2681 296 2695 330
rect 2633 258 2695 296
rect 2633 224 2647 258
rect 2681 224 2695 258
rect 2633 186 2695 224
rect 2633 152 2647 186
rect 2681 152 2695 186
rect 2633 114 2695 152
rect 2633 80 2647 114
rect 2681 80 2695 114
rect 2786 361 2820 377
rect 2980 361 3014 377
rect 3165 375 3199 723
rect 3757 683 3791 970
rect 3535 609 3569 625
rect 2820 327 2883 361
rect 2917 327 2980 361
rect 2786 289 2820 327
rect 2786 221 2820 255
rect 2980 289 3014 327
rect 2786 151 2820 187
rect 2786 101 2820 117
rect 2883 236 2917 252
rect 2633 62 2695 80
rect 2883 62 2917 202
rect 2980 221 3014 255
rect 3077 341 3199 375
rect 3299 546 3361 572
rect 3299 512 3313 546
rect 3347 512 3361 546
rect 3299 474 3361 512
rect 3299 440 3313 474
rect 3347 440 3361 474
rect 3299 402 3361 440
rect 3535 461 3569 575
rect 3535 411 3569 427
rect 3757 461 3791 649
rect 3757 411 3791 427
rect 3831 757 3865 1071
rect 3965 1076 3979 1110
rect 4013 1076 4027 1110
rect 4113 1412 4147 1492
rect 4113 1344 4147 1378
rect 4113 1276 4147 1310
rect 4113 1208 4147 1242
rect 4113 1139 4147 1174
rect 4113 1083 4147 1105
rect 4201 1412 4235 1450
rect 4201 1344 4235 1378
rect 4201 1276 4235 1310
rect 4201 1208 4235 1242
rect 4201 1139 4235 1174
rect 3965 1038 4027 1076
rect 3965 1004 3979 1038
rect 4013 1004 4027 1038
rect 3965 966 4027 1004
rect 4201 979 4235 1105
rect 4289 1412 4323 1492
rect 4289 1344 4323 1378
rect 4289 1276 4323 1310
rect 4289 1208 4323 1242
rect 4289 1139 4323 1174
rect 4289 1083 4323 1105
rect 4409 1470 4471 1492
rect 4409 1436 4423 1470
rect 4457 1436 4471 1470
rect 4409 1398 4471 1436
rect 4409 1364 4423 1398
rect 4457 1364 4471 1398
rect 4409 1326 4471 1364
rect 4409 1292 4423 1326
rect 4457 1292 4471 1326
rect 4409 1254 4471 1292
rect 4409 1220 4423 1254
rect 4457 1220 4471 1254
rect 4409 1182 4471 1220
rect 4409 1148 4423 1182
rect 4457 1148 4471 1182
rect 4409 1110 4471 1148
rect 4409 1076 4423 1110
rect 4457 1076 4471 1110
rect 4409 1038 4471 1076
rect 4581 1412 4615 1492
rect 4581 1344 4615 1378
rect 4581 1276 4615 1310
rect 4581 1208 4615 1242
rect 4581 1139 4615 1174
rect 4581 1073 4615 1105
rect 4669 1412 4703 1450
rect 4669 1344 4703 1378
rect 4669 1276 4703 1310
rect 4669 1208 4703 1242
rect 4669 1139 4703 1174
rect 4757 1412 4791 1492
rect 4757 1344 4791 1378
rect 4757 1276 4791 1310
rect 4757 1208 4791 1242
rect 4757 1157 4791 1174
rect 4845 1412 4879 1450
rect 4845 1344 4879 1378
rect 4845 1276 4879 1310
rect 4845 1208 4879 1242
rect 4669 1103 4703 1105
rect 4845 1139 4879 1174
rect 4933 1412 4967 1492
rect 4933 1344 4967 1378
rect 4933 1276 4967 1310
rect 4933 1208 4967 1242
rect 4933 1157 4967 1174
rect 5075 1470 5137 1492
rect 5075 1436 5089 1470
rect 5123 1436 5137 1470
rect 5075 1398 5137 1436
rect 5075 1364 5089 1398
rect 5123 1364 5137 1398
rect 5075 1326 5137 1364
rect 5075 1292 5089 1326
rect 5123 1292 5137 1326
rect 5075 1254 5137 1292
rect 5075 1220 5089 1254
rect 5123 1220 5137 1254
rect 5075 1182 5137 1220
rect 4845 1103 4879 1105
rect 5075 1148 5089 1182
rect 5123 1148 5137 1182
rect 5075 1110 5137 1148
rect 4669 1069 4975 1103
rect 3965 932 3979 966
rect 4013 932 4027 966
rect 3965 868 4027 932
rect 4127 945 4235 979
rect 4275 1003 4309 1019
rect 3299 368 3313 402
rect 3347 368 3361 402
rect 3077 245 3111 341
rect 3299 330 3361 368
rect 3077 195 3111 211
rect 3174 289 3208 305
rect 3174 221 3208 255
rect 2980 151 3014 187
rect 3174 151 3208 187
rect 3014 117 3077 151
rect 3111 117 3174 151
rect 2980 101 3014 117
rect 3174 101 3208 117
rect 3299 296 3313 330
rect 3347 296 3361 330
rect 3299 258 3361 296
rect 3299 224 3313 258
rect 3347 224 3361 258
rect 3299 186 3361 224
rect 3299 152 3313 186
rect 3347 152 3361 186
rect 3299 114 3361 152
rect 3299 80 3313 114
rect 3347 80 3361 114
rect 3452 361 3486 377
rect 3646 361 3680 377
rect 3831 375 3865 723
rect 4127 831 4161 945
rect 4127 609 4161 797
rect 3486 327 3549 361
rect 3583 327 3646 361
rect 3452 289 3486 327
rect 3452 221 3486 255
rect 3646 289 3680 327
rect 3452 151 3486 187
rect 3452 101 3486 117
rect 3549 236 3583 252
rect 3299 62 3361 80
rect 3549 62 3583 202
rect 3646 221 3680 255
rect 3743 341 3865 375
rect 3965 546 4027 572
rect 3965 512 3979 546
rect 4013 512 4027 546
rect 3965 474 4027 512
rect 3965 440 3979 474
rect 4013 440 4027 474
rect 3965 402 4027 440
rect 4127 461 4161 575
rect 4275 905 4309 969
rect 4275 535 4309 871
rect 4409 1004 4423 1038
rect 4457 1004 4471 1038
rect 4409 966 4471 1004
rect 4409 932 4423 966
rect 4457 932 4471 966
rect 4409 868 4471 932
rect 4645 1003 4679 1019
rect 4799 1003 4833 1019
rect 4645 905 4679 969
rect 4275 461 4309 501
rect 4127 427 4235 461
rect 3965 368 3979 402
rect 4013 368 4027 402
rect 3743 245 3777 341
rect 3965 330 4027 368
rect 3743 195 3777 211
rect 3840 289 3874 305
rect 3840 221 3874 255
rect 3646 151 3680 187
rect 3840 151 3874 187
rect 3680 117 3743 151
rect 3777 117 3840 151
rect 3646 101 3680 117
rect 3840 101 3874 117
rect 3965 296 3979 330
rect 4013 296 4027 330
rect 3965 258 4027 296
rect 3965 224 3979 258
rect 4013 224 4027 258
rect 3965 186 4027 224
rect 3965 152 3979 186
rect 4013 152 4027 186
rect 3965 114 4027 152
rect 3965 80 3979 114
rect 4013 80 4027 114
rect 3965 62 4027 80
rect 4103 361 4137 377
rect 4103 289 4137 327
rect 4103 221 4137 255
rect 4201 245 4235 427
rect 4275 411 4309 427
rect 4409 546 4471 572
rect 4409 512 4423 546
rect 4457 512 4471 546
rect 4409 474 4471 512
rect 4409 440 4423 474
rect 4457 440 4471 474
rect 4409 402 4471 440
rect 4645 461 4679 871
rect 4645 411 4679 427
rect 4793 969 4799 988
rect 4793 953 4833 969
rect 4793 461 4827 953
rect 4793 411 4827 427
rect 4941 683 4975 1069
rect 5075 1076 5089 1110
rect 5123 1076 5137 1110
rect 5223 1412 5257 1492
rect 5223 1344 5257 1378
rect 5223 1276 5257 1310
rect 5223 1208 5257 1242
rect 5223 1139 5257 1174
rect 5223 1083 5257 1105
rect 5311 1412 5345 1450
rect 5311 1344 5345 1378
rect 5311 1276 5345 1310
rect 5311 1208 5345 1242
rect 5311 1139 5345 1174
rect 5075 1038 5137 1076
rect 5075 1004 5089 1038
rect 5123 1004 5137 1038
rect 5075 966 5137 1004
rect 5075 932 5089 966
rect 5123 932 5137 966
rect 5075 868 5137 932
rect 5237 1003 5271 1019
rect 4201 195 4235 211
rect 4297 361 4331 377
rect 4297 289 4331 327
rect 4297 221 4331 255
rect 4103 151 4137 187
rect 4297 151 4331 187
rect 4137 117 4201 151
rect 4235 117 4297 151
rect 4103 62 4137 117
rect 4200 62 4234 117
rect 4297 62 4331 117
rect 4409 368 4423 402
rect 4457 368 4471 402
rect 4409 330 4471 368
rect 4409 296 4423 330
rect 4457 296 4471 330
rect 4409 258 4471 296
rect 4409 224 4423 258
rect 4457 224 4471 258
rect 4409 186 4471 224
rect 4409 152 4423 186
rect 4457 152 4471 186
rect 4409 114 4471 152
rect 4409 80 4423 114
rect 4457 80 4471 114
rect 4562 361 4596 377
rect 4756 361 4790 377
rect 4941 376 4975 649
rect 5237 683 5271 969
rect 5311 979 5345 1105
rect 5399 1412 5433 1492
rect 5399 1344 5433 1378
rect 5399 1276 5433 1310
rect 5399 1208 5433 1242
rect 5399 1139 5433 1174
rect 5399 1083 5433 1105
rect 5519 1470 5581 1492
rect 5519 1436 5533 1470
rect 5567 1436 5581 1470
rect 5519 1398 5581 1436
rect 5519 1364 5533 1398
rect 5567 1364 5581 1398
rect 5519 1326 5581 1364
rect 5519 1292 5533 1326
rect 5567 1292 5581 1326
rect 5519 1254 5581 1292
rect 5519 1220 5533 1254
rect 5567 1220 5581 1254
rect 5519 1182 5581 1220
rect 5519 1148 5533 1182
rect 5567 1148 5581 1182
rect 5519 1110 5581 1148
rect 5519 1076 5533 1110
rect 5567 1076 5581 1110
rect 5519 1038 5581 1076
rect 5691 1412 5725 1492
rect 5691 1344 5725 1378
rect 5691 1276 5725 1310
rect 5691 1208 5725 1242
rect 5691 1139 5725 1174
rect 5691 1073 5725 1105
rect 5779 1412 5813 1450
rect 5779 1344 5813 1378
rect 5779 1276 5813 1310
rect 5779 1208 5813 1242
rect 5779 1139 5813 1174
rect 5867 1412 5901 1492
rect 5867 1344 5901 1378
rect 5867 1276 5901 1310
rect 5867 1208 5901 1242
rect 5867 1157 5901 1174
rect 5955 1412 5989 1450
rect 5955 1344 5989 1378
rect 5955 1276 5989 1310
rect 5955 1208 5989 1242
rect 5779 1103 5813 1105
rect 5955 1139 5989 1174
rect 6043 1412 6077 1492
rect 6043 1344 6077 1378
rect 6043 1276 6077 1310
rect 6043 1208 6077 1242
rect 6043 1157 6077 1174
rect 6185 1470 6247 1492
rect 6185 1436 6199 1470
rect 6233 1436 6247 1470
rect 6185 1398 6247 1436
rect 6185 1364 6199 1398
rect 6233 1364 6247 1398
rect 6185 1326 6247 1364
rect 6185 1292 6199 1326
rect 6233 1292 6247 1326
rect 6185 1254 6247 1292
rect 6185 1220 6199 1254
rect 6233 1220 6247 1254
rect 6185 1182 6247 1220
rect 5955 1103 5989 1105
rect 6185 1148 6199 1182
rect 6233 1148 6247 1182
rect 6185 1110 6247 1148
rect 5779 1069 6085 1103
rect 5519 1004 5533 1038
rect 5567 1004 5581 1038
rect 5311 945 5419 979
rect 4596 327 4659 361
rect 4693 327 4756 361
rect 4562 289 4596 327
rect 4562 221 4596 255
rect 4756 289 4790 327
rect 4562 151 4596 187
rect 4562 101 4596 117
rect 4659 236 4693 252
rect 4409 62 4471 80
rect 4659 62 4693 202
rect 4756 221 4790 255
rect 4853 342 4975 376
rect 5075 546 5137 572
rect 5075 512 5089 546
rect 5123 512 5137 546
rect 5075 474 5137 512
rect 5075 440 5089 474
rect 5123 440 5137 474
rect 5075 402 5137 440
rect 5237 461 5271 649
rect 5385 609 5419 945
rect 5519 966 5581 1004
rect 5519 932 5533 966
rect 5567 932 5581 966
rect 5519 868 5581 932
rect 5755 1003 5789 1019
rect 5909 1003 5943 1019
rect 5385 461 5419 575
rect 5237 411 5271 427
rect 5311 427 5419 461
rect 5519 546 5581 572
rect 5519 512 5533 546
rect 5567 512 5581 546
rect 5519 474 5581 512
rect 5519 440 5533 474
rect 5567 440 5581 474
rect 5075 368 5089 402
rect 5123 368 5137 402
rect 4853 245 4887 342
rect 5075 330 5137 368
rect 4853 195 4887 211
rect 4950 289 4984 305
rect 4950 221 4984 255
rect 4756 151 4790 187
rect 4950 151 4984 187
rect 4790 117 4853 151
rect 4887 117 4950 151
rect 4756 101 4790 117
rect 4950 101 4984 117
rect 5075 296 5089 330
rect 5123 296 5137 330
rect 5075 258 5137 296
rect 5075 224 5089 258
rect 5123 224 5137 258
rect 5075 186 5137 224
rect 5075 152 5089 186
rect 5123 152 5137 186
rect 5075 114 5137 152
rect 5075 80 5089 114
rect 5123 80 5137 114
rect 5075 62 5137 80
rect 5215 361 5249 377
rect 5215 289 5249 327
rect 5215 221 5249 255
rect 5311 245 5345 427
rect 5519 402 5581 440
rect 5755 461 5789 945
rect 5903 969 5909 988
rect 5903 953 5943 969
rect 5903 461 5937 953
rect 6051 683 6085 1069
rect 6185 1076 6199 1110
rect 6233 1076 6247 1110
rect 6333 1412 6367 1492
rect 6333 1344 6367 1378
rect 6333 1276 6367 1310
rect 6333 1208 6367 1242
rect 6333 1139 6367 1174
rect 6333 1083 6367 1105
rect 6421 1412 6455 1450
rect 6421 1344 6455 1378
rect 6421 1276 6455 1310
rect 6421 1208 6455 1242
rect 6421 1139 6455 1174
rect 6185 1038 6247 1076
rect 6185 1004 6199 1038
rect 6233 1004 6247 1038
rect 6185 966 6247 1004
rect 6185 932 6199 966
rect 6233 932 6247 966
rect 6185 868 6247 932
rect 6347 1003 6381 1019
rect 5887 427 5903 461
rect 5937 427 5953 461
rect 5755 411 5789 427
rect 5903 411 5937 427
rect 5311 195 5345 211
rect 5409 361 5443 377
rect 5409 289 5443 327
rect 5409 221 5443 255
rect 5215 151 5249 187
rect 5409 151 5443 187
rect 5249 117 5311 151
rect 5345 117 5409 151
rect 5215 62 5249 117
rect 5312 62 5346 117
rect 5409 62 5443 117
rect 5519 368 5533 402
rect 5567 368 5581 402
rect 5519 330 5581 368
rect 5519 296 5533 330
rect 5567 296 5581 330
rect 5519 258 5581 296
rect 5519 224 5533 258
rect 5567 224 5581 258
rect 5519 186 5581 224
rect 5519 152 5533 186
rect 5567 152 5581 186
rect 5519 114 5581 152
rect 5519 80 5533 114
rect 5567 80 5581 114
rect 5672 361 5706 377
rect 5866 361 5900 377
rect 6051 376 6085 649
rect 6347 683 6381 969
rect 6421 979 6455 1105
rect 6509 1412 6543 1492
rect 6509 1344 6543 1378
rect 6509 1276 6543 1310
rect 6509 1208 6543 1242
rect 6509 1139 6543 1174
rect 6509 1083 6543 1105
rect 6629 1470 6691 1492
rect 6629 1436 6643 1470
rect 6677 1436 6691 1470
rect 6629 1398 6691 1436
rect 6629 1364 6643 1398
rect 6677 1364 6691 1398
rect 6629 1326 6691 1364
rect 6629 1292 6643 1326
rect 6677 1292 6691 1326
rect 6629 1254 6691 1292
rect 6629 1220 6643 1254
rect 6677 1220 6691 1254
rect 6629 1182 6691 1220
rect 6629 1148 6643 1182
rect 6677 1148 6691 1182
rect 6629 1110 6691 1148
rect 6629 1076 6643 1110
rect 6677 1076 6691 1110
rect 6629 1038 6691 1076
rect 6801 1411 6835 1451
rect 6801 1343 6835 1377
rect 6801 1275 6835 1309
rect 6801 1207 6835 1241
rect 6801 1139 6835 1173
rect 6889 1411 6923 1492
rect 7295 1470 7357 1492
rect 6889 1343 6923 1377
rect 6889 1275 6923 1309
rect 6889 1207 6923 1241
rect 6889 1157 6923 1173
rect 6977 1411 7187 1445
rect 6977 1343 7011 1377
rect 6977 1275 7011 1309
rect 6977 1207 7011 1241
rect 6977 1139 7011 1173
rect 6801 1071 7011 1105
rect 7065 1343 7099 1359
rect 7065 1275 7099 1309
rect 7065 1207 7099 1241
rect 7065 1139 7099 1173
rect 7153 1343 7187 1377
rect 7153 1275 7187 1309
rect 7153 1207 7187 1241
rect 7153 1157 7187 1173
rect 7295 1436 7309 1470
rect 7343 1436 7357 1470
rect 7295 1398 7357 1436
rect 7295 1364 7309 1398
rect 7343 1364 7357 1398
rect 7295 1326 7357 1364
rect 7295 1292 7309 1326
rect 7343 1292 7357 1326
rect 7295 1254 7357 1292
rect 7295 1220 7309 1254
rect 7343 1220 7357 1254
rect 7295 1182 7357 1220
rect 7295 1148 7309 1182
rect 7343 1148 7357 1182
rect 7295 1110 7357 1148
rect 7065 1071 7195 1105
rect 6629 1004 6643 1038
rect 6677 1004 6691 1038
rect 6421 945 6529 979
rect 5706 327 5769 361
rect 5803 327 5866 361
rect 5672 289 5706 327
rect 5672 221 5706 255
rect 5866 289 5900 327
rect 5672 151 5706 187
rect 5672 101 5706 117
rect 5769 236 5803 252
rect 5519 62 5581 80
rect 5769 62 5803 202
rect 5866 221 5900 255
rect 5963 342 6085 376
rect 6185 546 6247 572
rect 6185 512 6199 546
rect 6233 512 6247 546
rect 6185 474 6247 512
rect 6185 440 6199 474
rect 6233 440 6247 474
rect 6185 402 6247 440
rect 6347 461 6381 649
rect 6495 683 6529 945
rect 6629 966 6691 1004
rect 6629 932 6643 966
rect 6677 932 6691 966
rect 6834 1004 6868 1020
rect 7020 1004 7054 1020
rect 6868 970 6899 988
rect 6834 954 6899 970
rect 6629 868 6691 932
rect 6495 461 6529 649
rect 6865 609 6899 954
rect 6347 411 6381 427
rect 6421 427 6529 461
rect 6629 546 6691 572
rect 6629 512 6643 546
rect 6677 512 6691 546
rect 6629 474 6691 512
rect 6629 440 6643 474
rect 6677 440 6691 474
rect 6185 368 6199 402
rect 6233 368 6247 402
rect 5963 245 5997 342
rect 6185 330 6247 368
rect 5963 195 5997 211
rect 6060 289 6094 305
rect 6060 221 6094 255
rect 5866 151 5900 187
rect 6060 151 6094 187
rect 5900 117 5963 151
rect 5997 117 6060 151
rect 5866 101 5900 117
rect 6060 101 6094 117
rect 6185 296 6199 330
rect 6233 296 6247 330
rect 6185 258 6247 296
rect 6185 224 6199 258
rect 6233 224 6247 258
rect 6185 186 6247 224
rect 6185 152 6199 186
rect 6233 152 6247 186
rect 6185 114 6247 152
rect 6185 80 6199 114
rect 6233 80 6247 114
rect 6185 62 6247 80
rect 6325 361 6359 377
rect 6325 289 6359 327
rect 6325 221 6359 255
rect 6421 245 6455 427
rect 6629 402 6691 440
rect 6865 461 6899 575
rect 6865 411 6899 427
rect 7013 970 7020 988
rect 7013 954 7054 970
rect 7013 683 7047 954
rect 7013 461 7047 649
rect 7013 411 7047 427
rect 7161 683 7195 1071
rect 7295 1076 7309 1110
rect 7343 1076 7357 1110
rect 7443 1412 7477 1492
rect 7443 1344 7477 1378
rect 7443 1276 7477 1310
rect 7443 1208 7477 1242
rect 7443 1139 7477 1174
rect 7443 1083 7477 1105
rect 7531 1412 7565 1450
rect 7531 1344 7565 1378
rect 7531 1276 7565 1310
rect 7531 1208 7565 1242
rect 7531 1139 7565 1174
rect 7295 1038 7357 1076
rect 7295 1004 7309 1038
rect 7343 1004 7357 1038
rect 7295 966 7357 1004
rect 7295 932 7309 966
rect 7343 932 7357 966
rect 7295 868 7357 932
rect 7457 1003 7491 1019
rect 6421 195 6455 211
rect 6519 361 6553 377
rect 6519 289 6553 327
rect 6519 221 6553 255
rect 6325 151 6359 187
rect 6519 151 6553 187
rect 6359 117 6421 151
rect 6455 117 6519 151
rect 6325 62 6359 117
rect 6422 62 6456 117
rect 6519 62 6553 117
rect 6629 368 6643 402
rect 6677 368 6691 402
rect 6629 330 6691 368
rect 6629 296 6643 330
rect 6677 296 6691 330
rect 6629 258 6691 296
rect 6629 224 6643 258
rect 6677 224 6691 258
rect 6629 186 6691 224
rect 6629 152 6643 186
rect 6677 152 6691 186
rect 6629 114 6691 152
rect 6629 80 6643 114
rect 6677 80 6691 114
rect 6629 62 6691 80
rect 6782 361 6816 377
rect 7161 376 7195 649
rect 7457 683 7491 969
rect 7531 979 7565 1105
rect 7619 1412 7653 1492
rect 7619 1344 7653 1378
rect 7619 1276 7653 1310
rect 7619 1208 7653 1242
rect 7619 1139 7653 1174
rect 7619 1083 7653 1105
rect 7739 1470 7801 1492
rect 7739 1436 7753 1470
rect 7787 1436 7801 1470
rect 7739 1398 7801 1436
rect 7739 1364 7753 1398
rect 7787 1364 7801 1398
rect 7739 1326 7801 1364
rect 7739 1292 7753 1326
rect 7787 1292 7801 1326
rect 7739 1254 7801 1292
rect 7739 1220 7753 1254
rect 7787 1220 7801 1254
rect 7739 1182 7801 1220
rect 7739 1148 7753 1182
rect 7787 1148 7801 1182
rect 7739 1110 7801 1148
rect 7739 1076 7753 1110
rect 7787 1076 7801 1110
rect 7739 1038 7801 1076
rect 7739 1004 7753 1038
rect 7787 1004 7801 1038
rect 7531 945 7639 979
rect 6782 289 6816 327
rect 6782 221 6816 255
rect 6879 342 7195 376
rect 7295 546 7357 572
rect 7295 512 7309 546
rect 7343 512 7357 546
rect 7295 474 7357 512
rect 7295 440 7309 474
rect 7343 440 7357 474
rect 7295 402 7357 440
rect 7457 461 7491 649
rect 7605 683 7639 945
rect 7739 966 7801 1004
rect 7739 932 7753 966
rect 7787 932 7801 966
rect 7739 868 7801 932
rect 7605 461 7639 649
rect 7457 411 7491 427
rect 7531 427 7639 461
rect 7739 546 7801 572
rect 7739 512 7753 546
rect 7787 512 7801 546
rect 7739 474 7801 512
rect 7739 440 7753 474
rect 7787 440 7801 474
rect 7295 368 7309 402
rect 7343 368 7357 402
rect 6879 245 6913 342
rect 6879 195 6913 211
rect 6976 289 7010 306
rect 6976 221 7010 255
rect 6782 151 6816 187
rect 7073 245 7107 342
rect 7295 330 7357 368
rect 7073 195 7107 211
rect 7170 289 7204 306
rect 7170 221 7204 255
rect 6976 151 7010 187
rect 7170 151 7204 187
rect 6816 117 6879 151
rect 6913 117 6976 151
rect 7010 117 7073 151
rect 7107 117 7170 151
rect 6782 62 6816 117
rect 6879 62 6913 117
rect 6976 62 7010 117
rect 7073 62 7107 117
rect 7170 62 7204 117
rect 7295 296 7309 330
rect 7343 296 7357 330
rect 7295 258 7357 296
rect 7295 224 7309 258
rect 7343 224 7357 258
rect 7295 186 7357 224
rect 7295 152 7309 186
rect 7343 152 7357 186
rect 7295 114 7357 152
rect 7295 80 7309 114
rect 7343 80 7357 114
rect 7295 62 7357 80
rect 7435 361 7469 377
rect 7435 289 7469 327
rect 7435 221 7469 255
rect 7531 245 7565 427
rect 7739 402 7801 440
rect 7531 195 7565 211
rect 7629 361 7663 377
rect 7629 289 7663 327
rect 7629 221 7663 255
rect 7435 151 7469 187
rect 7629 151 7663 187
rect 7469 117 7531 151
rect 7565 117 7629 151
rect 7435 62 7469 117
rect 7532 62 7566 117
rect 7629 62 7663 117
rect 7739 368 7753 402
rect 7787 368 7801 402
rect 7739 330 7801 368
rect 7739 296 7753 330
rect 7787 296 7801 330
rect 7739 258 7801 296
rect 7739 224 7753 258
rect 7787 224 7801 258
rect 7739 186 7801 224
rect 7739 152 7753 186
rect 7787 152 7801 186
rect 7739 114 7801 152
rect 7739 80 7753 114
rect 7787 80 7801 114
rect 7739 62 7801 80
rect -31 47 7801 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 205 47
rect 239 13 283 47
rect 317 13 355 47
rect 389 13 499 47
rect 533 13 571 47
rect 605 13 643 47
rect 677 13 715 47
rect 749 13 805 47
rect 839 13 877 47
rect 911 13 949 47
rect 983 13 1021 47
rect 1055 13 1165 47
rect 1199 13 1237 47
rect 1271 13 1309 47
rect 1343 13 1381 47
rect 1415 13 1471 47
rect 1505 13 1543 47
rect 1577 13 1615 47
rect 1649 13 1687 47
rect 1721 13 1831 47
rect 1865 13 1903 47
rect 1937 13 1981 47
rect 2015 13 2059 47
rect 2093 13 2131 47
rect 2165 13 2275 47
rect 2309 13 2347 47
rect 2381 13 2425 47
rect 2459 13 2503 47
rect 2537 13 2575 47
rect 2609 13 2719 47
rect 2753 13 2791 47
rect 2825 13 2863 47
rect 2897 13 2935 47
rect 2969 13 3025 47
rect 3059 13 3097 47
rect 3131 13 3169 47
rect 3203 13 3241 47
rect 3275 13 3385 47
rect 3419 13 3457 47
rect 3491 13 3529 47
rect 3563 13 3601 47
rect 3635 13 3691 47
rect 3725 13 3763 47
rect 3797 13 3835 47
rect 3869 13 3907 47
rect 3941 13 4051 47
rect 4085 13 4123 47
rect 4157 13 4201 47
rect 4235 13 4279 47
rect 4313 13 4351 47
rect 4385 13 4495 47
rect 4529 13 4567 47
rect 4601 13 4639 47
rect 4673 13 4711 47
rect 4745 13 4801 47
rect 4835 13 4873 47
rect 4907 13 4945 47
rect 4979 13 5017 47
rect 5051 13 5161 47
rect 5195 13 5233 47
rect 5267 13 5311 47
rect 5345 13 5389 47
rect 5423 13 5461 47
rect 5495 13 5605 47
rect 5639 13 5677 47
rect 5711 13 5749 47
rect 5783 13 5821 47
rect 5855 13 5911 47
rect 5945 13 5983 47
rect 6017 13 6055 47
rect 6089 13 6127 47
rect 6161 13 6271 47
rect 6305 13 6343 47
rect 6377 13 6421 47
rect 6455 13 6499 47
rect 6533 13 6571 47
rect 6605 13 6715 47
rect 6749 13 6787 47
rect 6821 13 6859 47
rect 6893 13 6931 47
rect 6965 13 7021 47
rect 7055 13 7093 47
rect 7127 13 7165 47
rect 7199 13 7237 47
rect 7271 13 7381 47
rect 7415 13 7453 47
rect 7487 13 7531 47
rect 7565 13 7609 47
rect 7643 13 7681 47
rect 7715 13 7801 47
rect -31 0 7801 13
<< viali >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 205 1505 239 1539
rect 283 1505 317 1539
rect 355 1505 389 1539
rect 499 1505 533 1539
rect 571 1505 605 1539
rect 643 1505 677 1539
rect 715 1505 749 1539
rect 805 1505 839 1539
rect 877 1505 911 1539
rect 949 1505 983 1539
rect 1021 1505 1055 1539
rect 1165 1505 1199 1539
rect 1237 1505 1271 1539
rect 1309 1505 1343 1539
rect 1381 1505 1415 1539
rect 1471 1505 1505 1539
rect 1543 1505 1577 1539
rect 1615 1505 1649 1539
rect 1687 1505 1721 1539
rect 1831 1505 1865 1539
rect 1903 1505 1937 1539
rect 1981 1505 2015 1539
rect 2059 1505 2093 1539
rect 2131 1505 2165 1539
rect 2275 1505 2309 1539
rect 2347 1505 2381 1539
rect 2425 1505 2459 1539
rect 2503 1505 2537 1539
rect 2575 1505 2609 1539
rect 2719 1505 2753 1539
rect 2791 1505 2825 1539
rect 2863 1505 2897 1539
rect 2935 1505 2969 1539
rect 3025 1505 3059 1539
rect 3097 1505 3131 1539
rect 3169 1505 3203 1539
rect 3241 1505 3275 1539
rect 3385 1505 3419 1539
rect 3457 1505 3491 1539
rect 3529 1505 3563 1539
rect 3601 1505 3635 1539
rect 3691 1505 3725 1539
rect 3763 1505 3797 1539
rect 3835 1505 3869 1539
rect 3907 1505 3941 1539
rect 4051 1505 4085 1539
rect 4123 1505 4157 1539
rect 4201 1505 4235 1539
rect 4279 1505 4313 1539
rect 4351 1505 4385 1539
rect 4495 1505 4529 1539
rect 4567 1505 4601 1539
rect 4639 1505 4673 1539
rect 4711 1505 4745 1539
rect 4801 1505 4835 1539
rect 4873 1505 4907 1539
rect 4945 1505 4979 1539
rect 5017 1505 5051 1539
rect 5161 1505 5195 1539
rect 5233 1505 5267 1539
rect 5311 1505 5345 1539
rect 5389 1505 5423 1539
rect 5461 1505 5495 1539
rect 5605 1505 5639 1539
rect 5677 1505 5711 1539
rect 5749 1505 5783 1539
rect 5821 1505 5855 1539
rect 5911 1505 5945 1539
rect 5983 1505 6017 1539
rect 6055 1505 6089 1539
rect 6127 1505 6161 1539
rect 6271 1505 6305 1539
rect 6343 1505 6377 1539
rect 6421 1505 6455 1539
rect 6499 1505 6533 1539
rect 6571 1505 6605 1539
rect 6715 1505 6749 1539
rect 6787 1505 6821 1539
rect 6859 1505 6893 1539
rect 6931 1505 6965 1539
rect 7021 1505 7055 1539
rect 7093 1505 7127 1539
rect 7165 1505 7199 1539
rect 7237 1505 7271 1539
rect 7381 1505 7415 1539
rect 7453 1505 7487 1539
rect 7531 1505 7565 1539
rect 7609 1505 7643 1539
rect 7681 1505 7715 1539
rect 131 871 165 905
rect 649 871 683 905
rect 279 649 313 683
rect 871 797 905 831
rect 1315 871 1349 905
rect 945 723 979 757
rect 871 501 905 535
rect 649 427 683 461
rect 1537 649 1571 683
rect 1315 575 1349 609
rect 2055 969 2089 979
rect 2055 945 2089 969
rect 1611 723 1645 757
rect 1907 797 1941 831
rect 1907 575 1941 609
rect 2055 871 2089 905
rect 2351 871 2385 905
rect 2351 723 2385 757
rect 2055 501 2089 535
rect 2869 871 2903 905
rect 2499 649 2533 683
rect 2351 427 2385 461
rect 3091 797 3125 831
rect 3535 871 3569 905
rect 3165 723 3199 757
rect 3091 501 3125 535
rect 3757 649 3791 683
rect 3535 575 3569 609
rect 3831 723 3865 757
rect 4127 797 4161 831
rect 4127 575 4161 609
rect 4275 871 4309 905
rect 4645 871 4679 905
rect 4275 501 4309 535
rect 4793 427 4827 461
rect 4941 649 4975 683
rect 5237 649 5271 683
rect 5755 969 5789 979
rect 5755 945 5789 969
rect 5385 575 5419 609
rect 6051 649 6085 683
rect 5903 427 5937 461
rect 6347 649 6381 683
rect 6495 649 6529 683
rect 6865 575 6899 609
rect 7013 649 7047 683
rect 7161 649 7195 683
rect 7457 649 7491 683
rect 7605 649 7639 683
rect 55 13 89 47
rect 127 13 161 47
rect 205 13 239 47
rect 283 13 317 47
rect 355 13 389 47
rect 499 13 533 47
rect 571 13 605 47
rect 643 13 677 47
rect 715 13 749 47
rect 805 13 839 47
rect 877 13 911 47
rect 949 13 983 47
rect 1021 13 1055 47
rect 1165 13 1199 47
rect 1237 13 1271 47
rect 1309 13 1343 47
rect 1381 13 1415 47
rect 1471 13 1505 47
rect 1543 13 1577 47
rect 1615 13 1649 47
rect 1687 13 1721 47
rect 1831 13 1865 47
rect 1903 13 1937 47
rect 1981 13 2015 47
rect 2059 13 2093 47
rect 2131 13 2165 47
rect 2275 13 2309 47
rect 2347 13 2381 47
rect 2425 13 2459 47
rect 2503 13 2537 47
rect 2575 13 2609 47
rect 2719 13 2753 47
rect 2791 13 2825 47
rect 2863 13 2897 47
rect 2935 13 2969 47
rect 3025 13 3059 47
rect 3097 13 3131 47
rect 3169 13 3203 47
rect 3241 13 3275 47
rect 3385 13 3419 47
rect 3457 13 3491 47
rect 3529 13 3563 47
rect 3601 13 3635 47
rect 3691 13 3725 47
rect 3763 13 3797 47
rect 3835 13 3869 47
rect 3907 13 3941 47
rect 4051 13 4085 47
rect 4123 13 4157 47
rect 4201 13 4235 47
rect 4279 13 4313 47
rect 4351 13 4385 47
rect 4495 13 4529 47
rect 4567 13 4601 47
rect 4639 13 4673 47
rect 4711 13 4745 47
rect 4801 13 4835 47
rect 4873 13 4907 47
rect 4945 13 4979 47
rect 5017 13 5051 47
rect 5161 13 5195 47
rect 5233 13 5267 47
rect 5311 13 5345 47
rect 5389 13 5423 47
rect 5461 13 5495 47
rect 5605 13 5639 47
rect 5677 13 5711 47
rect 5749 13 5783 47
rect 5821 13 5855 47
rect 5911 13 5945 47
rect 5983 13 6017 47
rect 6055 13 6089 47
rect 6127 13 6161 47
rect 6271 13 6305 47
rect 6343 13 6377 47
rect 6421 13 6455 47
rect 6499 13 6533 47
rect 6571 13 6605 47
rect 6715 13 6749 47
rect 6787 13 6821 47
rect 6859 13 6893 47
rect 6931 13 6965 47
rect 7021 13 7055 47
rect 7093 13 7127 47
rect 7165 13 7199 47
rect 7237 13 7271 47
rect 7381 13 7415 47
rect 7453 13 7487 47
rect 7531 13 7565 47
rect 7609 13 7643 47
rect 7681 13 7715 47
<< metal1 >>
rect -31 1539 7801 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 205 1539
rect 239 1505 283 1539
rect 317 1505 355 1539
rect 389 1505 499 1539
rect 533 1505 571 1539
rect 605 1505 643 1539
rect 677 1505 715 1539
rect 749 1505 805 1539
rect 839 1505 877 1539
rect 911 1505 949 1539
rect 983 1505 1021 1539
rect 1055 1505 1165 1539
rect 1199 1505 1237 1539
rect 1271 1505 1309 1539
rect 1343 1505 1381 1539
rect 1415 1505 1471 1539
rect 1505 1505 1543 1539
rect 1577 1505 1615 1539
rect 1649 1505 1687 1539
rect 1721 1505 1831 1539
rect 1865 1505 1903 1539
rect 1937 1505 1981 1539
rect 2015 1505 2059 1539
rect 2093 1505 2131 1539
rect 2165 1505 2275 1539
rect 2309 1505 2347 1539
rect 2381 1505 2425 1539
rect 2459 1505 2503 1539
rect 2537 1505 2575 1539
rect 2609 1505 2719 1539
rect 2753 1505 2791 1539
rect 2825 1505 2863 1539
rect 2897 1505 2935 1539
rect 2969 1505 3025 1539
rect 3059 1505 3097 1539
rect 3131 1505 3169 1539
rect 3203 1505 3241 1539
rect 3275 1505 3385 1539
rect 3419 1505 3457 1539
rect 3491 1505 3529 1539
rect 3563 1505 3601 1539
rect 3635 1505 3691 1539
rect 3725 1505 3763 1539
rect 3797 1505 3835 1539
rect 3869 1505 3907 1539
rect 3941 1505 4051 1539
rect 4085 1505 4123 1539
rect 4157 1505 4201 1539
rect 4235 1505 4279 1539
rect 4313 1505 4351 1539
rect 4385 1505 4495 1539
rect 4529 1505 4567 1539
rect 4601 1505 4639 1539
rect 4673 1505 4711 1539
rect 4745 1505 4801 1539
rect 4835 1505 4873 1539
rect 4907 1505 4945 1539
rect 4979 1505 5017 1539
rect 5051 1505 5161 1539
rect 5195 1505 5233 1539
rect 5267 1505 5311 1539
rect 5345 1505 5389 1539
rect 5423 1505 5461 1539
rect 5495 1505 5605 1539
rect 5639 1505 5677 1539
rect 5711 1505 5749 1539
rect 5783 1505 5821 1539
rect 5855 1505 5911 1539
rect 5945 1505 5983 1539
rect 6017 1505 6055 1539
rect 6089 1505 6127 1539
rect 6161 1505 6271 1539
rect 6305 1505 6343 1539
rect 6377 1505 6421 1539
rect 6455 1505 6499 1539
rect 6533 1505 6571 1539
rect 6605 1505 6715 1539
rect 6749 1505 6787 1539
rect 6821 1505 6859 1539
rect 6893 1505 6931 1539
rect 6965 1505 7021 1539
rect 7055 1505 7093 1539
rect 7127 1505 7165 1539
rect 7199 1505 7237 1539
rect 7271 1505 7381 1539
rect 7415 1505 7453 1539
rect 7487 1505 7531 1539
rect 7565 1505 7609 1539
rect 7643 1505 7681 1539
rect 7715 1505 7801 1539
rect -31 1492 7801 1505
rect 2049 979 2095 985
rect 5749 979 5795 985
rect 2043 945 2055 979
rect 2089 945 5755 979
rect 5789 945 5801 979
rect 2049 939 2095 945
rect 5749 939 5795 945
rect 125 905 171 911
rect 643 905 689 911
rect 1309 905 1355 911
rect 2049 905 2095 911
rect 2345 905 2391 911
rect 2863 905 2909 911
rect 3529 905 3575 911
rect 4269 905 4315 911
rect 4639 905 4685 911
rect 119 871 131 905
rect 165 871 649 905
rect 683 871 695 905
rect 1303 871 1315 905
rect 1349 871 2055 905
rect 2089 871 2101 905
rect 2339 871 2351 905
rect 2385 871 2869 905
rect 2903 871 2915 905
rect 3523 871 3535 905
rect 3569 871 4275 905
rect 4309 871 4645 905
rect 4679 871 4691 905
rect 125 865 171 871
rect 643 865 689 871
rect 1309 865 1355 871
rect 2049 865 2095 871
rect 2345 865 2391 871
rect 2863 865 2909 871
rect 3529 865 3575 871
rect 4269 865 4315 871
rect 4639 865 4685 871
rect 865 831 911 837
rect 1901 831 1947 837
rect 3085 831 3131 837
rect 4121 831 4167 837
rect 859 797 871 831
rect 905 797 1907 831
rect 1941 797 1953 831
rect 3079 797 3091 831
rect 3125 797 4127 831
rect 4161 797 4173 831
rect 865 791 911 797
rect 1901 791 1947 797
rect 3085 791 3131 797
rect 4121 791 4167 797
rect 939 757 985 763
rect 1605 757 1651 763
rect 2345 757 2391 763
rect 3159 757 3205 763
rect 3825 757 3871 763
rect 933 723 945 757
rect 979 723 1611 757
rect 1645 723 2351 757
rect 2385 723 2397 757
rect 3153 723 3165 757
rect 3199 723 3831 757
rect 3865 723 3877 757
rect 939 717 985 723
rect 1605 717 1651 723
rect 2345 717 2391 723
rect 3159 717 3205 723
rect 3825 717 3871 723
rect 273 683 319 689
rect 1531 683 1577 689
rect 2493 683 2539 689
rect 3751 683 3797 689
rect 4935 683 4981 689
rect 5231 683 5277 689
rect 6045 683 6091 689
rect 6341 683 6387 689
rect 6489 683 6535 689
rect 7007 683 7053 689
rect 7155 683 7201 689
rect 7451 683 7497 689
rect 7599 683 7645 689
rect 267 649 279 683
rect 313 649 1537 683
rect 1571 649 1583 683
rect 2487 649 2499 683
rect 2533 649 3757 683
rect 3791 649 3803 683
rect 4929 649 4941 683
rect 4975 649 5237 683
rect 5271 649 5283 683
rect 6039 649 6051 683
rect 6085 649 6347 683
rect 6381 649 6393 683
rect 6483 649 6495 683
rect 6529 649 7013 683
rect 7047 649 7059 683
rect 7149 649 7161 683
rect 7195 649 7457 683
rect 7491 649 7503 683
rect 7593 649 7605 683
rect 7639 649 7675 683
rect 273 643 319 649
rect 1531 643 1577 649
rect 2493 643 2539 649
rect 3751 643 3797 649
rect 4935 643 4981 649
rect 5231 643 5277 649
rect 6045 643 6091 649
rect 6341 643 6387 649
rect 6489 643 6535 649
rect 7007 643 7053 649
rect 7155 643 7201 649
rect 7451 643 7497 649
rect 7599 643 7645 649
rect 1309 609 1355 615
rect 1901 609 1947 615
rect 3529 609 3575 615
rect 4121 609 4167 615
rect 5379 609 5425 615
rect 6859 609 6905 615
rect 1303 575 1315 609
rect 1349 575 1907 609
rect 1941 575 1953 609
rect 3523 575 3535 609
rect 3569 575 4127 609
rect 4161 575 4173 609
rect 5373 575 5385 609
rect 5419 575 6865 609
rect 6899 575 6911 609
rect 1309 569 1355 575
rect 1901 569 1947 575
rect 3529 569 3575 575
rect 4121 569 4167 575
rect 5379 569 5425 575
rect 6859 569 6905 575
rect 865 535 911 541
rect 2049 535 2095 541
rect 3085 535 3131 541
rect 4269 535 4315 541
rect 859 501 871 535
rect 905 501 2055 535
rect 2089 501 2101 535
rect 3079 501 3091 535
rect 3125 501 4275 535
rect 4309 501 4321 535
rect 865 495 911 501
rect 2049 495 2095 501
rect 3085 495 3131 501
rect 4269 495 4315 501
rect 649 467 683 473
rect 5903 467 5937 473
rect 643 461 689 467
rect 2345 461 2391 467
rect 4787 461 4833 467
rect 5897 461 5943 467
rect 643 427 649 461
rect 683 427 689 461
rect 2339 427 2351 461
rect 2385 427 4793 461
rect 4827 427 4839 461
rect 5897 427 5903 461
rect 5937 427 5943 461
rect 643 421 689 427
rect 2345 421 2391 427
rect 4787 421 4833 427
rect 5897 421 5943 427
rect 649 387 683 421
rect 5903 387 5937 421
rect 649 353 5937 387
rect -31 47 7801 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 205 47
rect 239 13 283 47
rect 317 13 355 47
rect 389 13 499 47
rect 533 13 571 47
rect 605 13 643 47
rect 677 13 715 47
rect 749 13 805 47
rect 839 13 877 47
rect 911 13 949 47
rect 983 13 1021 47
rect 1055 13 1165 47
rect 1199 13 1237 47
rect 1271 13 1309 47
rect 1343 13 1381 47
rect 1415 13 1471 47
rect 1505 13 1543 47
rect 1577 13 1615 47
rect 1649 13 1687 47
rect 1721 13 1831 47
rect 1865 13 1903 47
rect 1937 13 1981 47
rect 2015 13 2059 47
rect 2093 13 2131 47
rect 2165 13 2275 47
rect 2309 13 2347 47
rect 2381 13 2425 47
rect 2459 13 2503 47
rect 2537 13 2575 47
rect 2609 13 2719 47
rect 2753 13 2791 47
rect 2825 13 2863 47
rect 2897 13 2935 47
rect 2969 13 3025 47
rect 3059 13 3097 47
rect 3131 13 3169 47
rect 3203 13 3241 47
rect 3275 13 3385 47
rect 3419 13 3457 47
rect 3491 13 3529 47
rect 3563 13 3601 47
rect 3635 13 3691 47
rect 3725 13 3763 47
rect 3797 13 3835 47
rect 3869 13 3907 47
rect 3941 13 4051 47
rect 4085 13 4123 47
rect 4157 13 4201 47
rect 4235 13 4279 47
rect 4313 13 4351 47
rect 4385 13 4495 47
rect 4529 13 4567 47
rect 4601 13 4639 47
rect 4673 13 4711 47
rect 4745 13 4801 47
rect 4835 13 4873 47
rect 4907 13 4945 47
rect 4979 13 5017 47
rect 5051 13 5161 47
rect 5195 13 5233 47
rect 5267 13 5311 47
rect 5345 13 5389 47
rect 5423 13 5461 47
rect 5495 13 5605 47
rect 5639 13 5677 47
rect 5711 13 5749 47
rect 5783 13 5821 47
rect 5855 13 5911 47
rect 5945 13 5983 47
rect 6017 13 6055 47
rect 6089 13 6127 47
rect 6161 13 6271 47
rect 6305 13 6343 47
rect 6377 13 6421 47
rect 6455 13 6499 47
rect 6533 13 6571 47
rect 6605 13 6715 47
rect 6749 13 6787 47
rect 6821 13 6859 47
rect 6893 13 6931 47
rect 6965 13 7021 47
rect 7055 13 7093 47
rect 7127 13 7165 47
rect 7199 13 7237 47
rect 7271 13 7381 47
rect 7415 13 7453 47
rect 7487 13 7531 47
rect 7565 13 7609 47
rect 7643 13 7681 47
rect 7715 13 7801 47
rect -31 0 7801 13
<< labels >>
rlabel metal1 3831 723 3865 757 1 SUM
port 1 n
rlabel metal1 7605 649 7639 683 1 COUT
port 2 n
rlabel metal1 131 871 165 905 1 A
port 3 n
rlabel metal1 1315 871 1349 905 1 B
port 4 n
rlabel metal1 4645 871 4679 905 1 CIN
port 5 n
rlabel metal1 -31 1492 7801 1554 1 VDD
port 6 n
rlabel metal1 -31 0 7801 62 1 GND
port 7 n
<< end >>
