* SPICE3 file created from INVX1.ext - technology: sky130A

.subckt INVX1 VDD A VSS Y
M1000 Y A VDD VDD pshort w=3u l=0.15u
+  ad=0.87p pd=6.58u as=1.65p ps=13.1u
M1001 Y A VSS VSS nshort w=3u l=0.15u
+  ad=0.1588p pd=1.5u as=1.16175p ps=8.02u
M1002 VDD A Y VDD pshort w=3u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
.ends
