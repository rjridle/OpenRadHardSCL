* NGSPICE file created from OR2X1.ext - technology: sky130A

.subckt nmos_top a_85_108# a_55_92# a_n1_0# VSUBS
X0 a_85_108# a_55_92# a_n1_0# VSUBS sky130_fd_pr__nfet_01v8 ad=1.772p pd=1.56u as=1.15725p ps=8.12u w=3u l=0.15u
.ends

.subckt pmos2 a_144_n460# a_262_n399# a_88_n399# w_52_n435# a_174_n399#
X0 a_174_n399# a_144_n460# a_88_n399# w_52_n435# sky130_fd_pr__pfet_01v8 ad=5.8p pd=4.58u as=5.6p ps=4.56u w=2u l=0.15u
X1 a_262_n399# a_144_n460# a_174_n399# w_52_n435# sky130_fd_pr__pfet_01v8 ad=5.4p pd=4.54u as=0p ps=0u w=2u l=0.15u
.ends

.subckt invx1_pcell VSS VDD a_154_410# a_205_1105#
Xnmos_top_0 a_205_1105# a_154_410# VSS VSS nmos_top
Xpmos2_0 a_154_410# VDD VDD VDD a_205_1105# pmos2
.ends

.subckt pmos2_1 a_144_n460# a_262_n399# a_88_n399# w_52_n435# a_174_n399#
X0 a_174_n399# a_144_n460# a_88_n399# w_52_n435# sky130_fd_pr__pfet_01v8 ad=5.8p pd=4.58u as=5.6p ps=4.56u w=2u l=0.15u
X1 a_262_n399# a_144_n460# a_174_n399# w_52_n435# sky130_fd_pr__pfet_01v8 ad=5.4p pd=4.54u as=0p ps=0u w=2u l=0.15u
.ends

.subckt nmos_top_trim1 a_56_92# a_86_108# a_0_0# VSUBS
X0 a_86_108# a_56_92# a_0_0# VSUBS sky130_fd_pr__nfet_01v8 ad=1.772p pd=1.56u as=1.15725p ps=8.12u w=3u l=0.15u
.ends

.subckt nmos_top_trim2 a_56_92# a_86_108# a_0_0# VSUBS
X0 a_86_108# a_56_92# a_0_0# VSUBS sky130_fd_pr__nfet_01v8 ad=1.772p pd=1.56u as=1.15725p ps=8.12u w=3u l=0.15u
.ends

.subckt nor2x1_pcell VDD VSS a_168_403# a_362_410# a_405_1105#
Xpmos2_1_0 a_168_403# a_317_1377# a_317_1377# VDD VDD pmos2_1
Xpmos2_1_1 a_362_410# a_317_1377# a_317_1377# VDD a_405_1105# pmos2_1
Xnmos_top_trim1_1 a_168_403# a_405_1105# VSS VSS nmos_top_trim1
Xnmos_top_trim2_0 a_362_410# a_405_1105# VSS VSS nmos_top_trim2
.ends

.subckt or2x1_pcell VSS VDD invx1_pcell_0/a_205_1105# nor2x1_pcell_0/a_168_403# nor2x1_pcell_0/a_362_410#
Xinvx1_pcell_0 VSS VDD m1_547_649# invx1_pcell_0/a_205_1105# invx1_pcell
Xnor2x1_pcell_0 VDD VSS nor2x1_pcell_0/a_168_403# nor2x1_pcell_0/a_362_410# m1_547_649#
+ nor2x1_pcell
.ends

.subckt OR2X1 Y A B VDD VSS
Xor2x1_pcell_0 VSS VDD Y A B or2x1_pcell
.ends

