* NGSPICE file created from NAND3X1.ext - technology: sky130A

.subckt NAND3X1 VDD VSS B A C Y
X0 VSS A nmos_bottom_0/a_0_0# VSS sky130_fd_pr__nfet_01v8 ad=1.772e+11p pd=1.56e+06u as=0p ps=0u w=3e+06u l=150000u
X1 Y C li_393_210# VSS sky130_fd_pr__nfet_01v8 ad=1.772e+11p pd=1.56e+06u as=0p ps=0u w=3e+06u l=150000u
X2 li_393_210# B nmos_bottom_0/a_0_0# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X3 Y A VDD VDD sky130_fd_pr__pfet_01v8 ad=-1.3025e+10p pd=1.3745e+07u as=4.00705e+12p ps=1.8265e+07u w=2e+06u l=150000u M=2
X4 Y B VDD VDD sky130_fd_pr__pfet_01v8 ad=-0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X5 Y C VDD VDD sky130_fd_pr__pfet_01v8 ad=-0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
.ends
