* SPICE3 file created from INVX1_diff_ring.ext - technology: sky130A

.subckt INVX1_diff_ring VDD Y A VSS
M1000 VDD A Y VDD pshort w=2u l=0.15u
+  ad=1.1p pd=9.1u as=0.58p ps=4.58u
M1001 Y A VSS VSS nshort w=3u l=0.15u
+  ad=0.1588p pd=1.5u as=1.16175p ps=8.02u
M1002 Y A VDD VDD pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
.ends
