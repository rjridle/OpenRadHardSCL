* SPICE3 file created from TIELO.ext - technology: sky130A

.subckt TIELO YN VDD GND
X0 YN a_121_411.t4 GND.t0 GND sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=0p ps=0u w=0u l=0u
X1 a_121_411.t3 a_121_411.t2 VDD.t3  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X2 VDD.t1 a_121_411.t0 a_121_411.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
R0 a_121_411.n0 a_121_411.t0 512.525
R1 a_121_411.n1 a_121_411.t4 396.923
R2 a_121_411.n0 a_121_411.t2 371.139
R3 a_121_411.n2 a_121_411.n1 157.398
R4 a_121_411.n1 a_121_411.n0 126.877
R5 a_121_411.n2 a_121_411.t1 14.282
R6 a_121_411.t3 a_121_411.n2 14.282
R7 VDD.n55 VDD.t3 135.162
R8 VDD.n24 VDD.t1 135.162
R9 VDD.n38 VDD.n37 92.5
R10 VDD.n36 VDD.n35 92.5
R11 VDD.n34 VDD.n33 92.5
R12 VDD.n32 VDD.n31 92.5
R13 VDD.n40 VDD.n39 92.5
R14 VDD.n14 VDD.n1 92.5
R15 VDD.n5 VDD.n4 92.5
R16 VDD.n7 VDD.n6 92.5
R17 VDD.n9 VDD.n8 92.5
R18 VDD.n11 VDD.n10 92.5
R19 VDD.n13 VDD.n12 92.5
R20 VDD.n21 VDD.n20 92.059
R21 VDD.n49 VDD.n48 92.059
R22 VDD.n20 VDD.n16 67.194
R23 VDD.n20 VDD.n17 67.194
R24 VDD.n20 VDD.n18 67.194
R25 VDD.n20 VDD.n19 67.194
R26 VDD.n5 VDD.n3 44.141
R27 VDD.n3 VDD.n2 44.107
R28 VDD.n25 VDD.t0 43.472
R29 VDD.n53 ���߫U 43.472
R30 VDD.n20 VDD.n15 41.052
R31 VDD.n47 VDD.n45 39.742
R32 VDD.n47 VDD.n46 39.742
R33 VDD.n44 VDD.n43 39.742
R34 VDD.n1 VDD.n0 30.923
R35 VDD.n48 VDD.n47 26.38
R36 VDD.n48 VDD.n44 26.38
R37 VDD.n48 VDD.n42 26.38
R38 VDD.n48 VDD.n41 26.38
R39 VDD.n51 VDD.n40 22.915
R40 VDD.n23 VDD.n14 22.915
R41 VDD.n40 VDD.n38 14.864
R42 VDD.n38 VDD.n36 14.864
R43 VDD.n36 VDD.n34 14.864
R44 VDD.n34 VDD.n32 14.864
R45 VDD.n32 VDD.n30 14.864
R46 VDD.n30 VDD.n29 14.864
R47 VDD.n14 VDD.n13 14.864
R48 VDD.n13 VDD.n11 14.864
R49 VDD.n11 VDD.n9 14.864
R50 VDD.n9 VDD.n7 14.864
R51 VDD.n7 VDD.n5 14.864
R52 VDD.n23 VDD.n22 8.855
R53 VDD.n22 VDD.n21 8.855
R54 VDD.n27 VDD.n26 8.855
R55 VDD.n26 VDD.n25 8.855
R56 VDD.n60 VDD.n59 8.855
R57 VDD.n59 VDD.n58 8.855
R58 VDD.n56 VDD.n54 8.855
R59 VDD.n54 VDD.n53 8.855
R60 VDD.n51 VDD.n50 8.855
R61 VDD.n50 VDD.n49 8.855
R62 VDD.n28 VDD.n23 4.795
R63 VDD.n28 VDD.n27 4.65
R64 VDD.n61 VDD.n60 4.65
R65 VDD.n57 VDD.n56 4.65
R66 VDD.n52 VDD.n51 4.65
R67 VDD.n27 VDD.n24 2.064
R68 VDD.n56 VDD.n55 2.064
R69 VDD.n52 VDD 0.207
R70 VDD.n61 VDD.n28 0.157
R71 VDD.n61 VDD.n57 0.157
R72 VDD.n57 VDD.n52 0.145
R73 GND.n5 GND.n4 120.01
R74 GND.n3 GND.n2 92.5
R75 GND.n24 GND.n23 92.5
R76 GND.n17 GND.t0 45.413
R77 GND.n17 GND.n16 39.307
R78 GND.n18 GND.n17 23.77
R79 GND.n26 GND.n24 20.705
R80 GND.n6 GND.n5 20.705
R81 GND.n19 GND.n18 20.705
R82 GND.n5 GND.n3 19.952
R83 GND.n20 GND.n13 9.154
R84 GND.n26 GND.n25 9.154
R85 GND.n8 GND.n7 9.154
R86 GND.n9 GND.n1 4.795
R87 GND.n12 GND.n11 4.65
R88 GND.n9 GND.n8 4.65
R89 GND.n27 GND.n26 4.65
R90 GND.n21 GND.n20 4.65
R91 GND.n15 GND.n14 4.504
R92 GND.n8 GND.n6 4.129
R93 GND.n20 GND.n19 3.716
R94 GND.t0 GND.n15 2.452
R95 GND.n23 GND.n22 1.935
R96 GND.n1 GND.n0 0.474
R97 GND.n11 GND.n10 0.474
R98 GND.n12 GND 0.207
R99 GND.n27 GND.n9 0.157
R100 GND.n27 GND.n21 0.157
R101 GND.n21 GND.n12 0.145
R102 YN.n1 YN.n0 255.924
R103 YN.n1 YN 0.046
C0 VDD GND 0.96fF
C1 YN.n0 GND 0.35fF
C2 YN.n1 GND 0.37fF
C3 VDD.n1 GND 0.02fF
C4 VDD.n2 GND 0.06fF
C5 VDD.n3 GND 0.02fF
C6 VDD.n4 GND 0.01fF
C7 VDD.n5 GND 0.03fF
C8 VDD.n6 GND 0.01fF
C9 VDD.n7 GND 0.01fF
C10 VDD.n8 GND 0.01fF
C11 VDD.n9 GND 0.01fF
C12 VDD.n10 GND 0.01fF
C13 VDD.n11 GND 0.01fF
C14 VDD.n12 GND 0.01fF
C15 VDD.n13 GND 0.01fF
C16 VDD.n14 GND 0.02fF
C17 VDD.n15 GND 0.01fF
C18 VDD.n20 GND 0.25fF
C19 VDD.n21 GND 0.15fF
C20 VDD.n22 GND 0.01fF
C21 VDD.n23 GND 0.02fF
C22 VDD.n24 GND 0.04fF
C23 VDD.n25 GND 0.11fF
C24 VDD.n26 GND 0.01fF
C25 VDD.n27 GND 0.01fF
C26 VDD.n28 GND 0.04fF
C27 VDD.n29 GND 0.03fF
C28 VDD.n30 GND 0.01fF
C29 VDD.n31 GND 0.01fF
C30 VDD.n32 GND 0.01fF
C31 VDD.n33 GND 0.01fF
C32 VDD.n34 GND 0.01fF
C33 VDD.n35 GND 0.01fF
C34 VDD.n36 GND 0.01fF
C35 VDD.n37 GND 0.01fF
C36 VDD.n38 GND 0.01fF
C37 VDD.n39 GND 0.02fF
C38 VDD.n40 GND 0.02fF
C39 VDD.n43 GND 0.01fF
C40 VDD.n45 GND 0.01fF
C41 VDD.n46 GND 0.06fF
C42 VDD.n48 GND 0.25fF
C43 VDD.n49 GND 0.15fF
C44 VDD.n50 GND 0.01fF
C45 VDD.n51 GND 0.02fF
C46 VDD.n52 GND 0.02fF
C47 VDD.n53 GND 0.11fF
C48 VDD.n54 GND 0.01fF
C49 VDD.n55 GND 0.04fF
C50 VDD.n56 GND 0.01fF
C51 VDD.n57 GND 0.01fF
C52 VDD.n58 GND 0.09fF
C53 VDD.n59 GND 0.01fF
C54 VDD.n60 GND 0.01fF
C55 VDD.n61 GND 0.01fF
C56 a_121_411.n0 GND 0.16fF
C57 a_121_411.n1 GND 0.37fF
C58 a_121_411.n2 GND 0.29fF
.ends
