magic
tech sky130A
magscale 1 2
timestamp 1649530828
<< nwell >>
rect -84 832 16734 1575
<< nmos >>
rect 168 316 198 377
tri 198 316 214 332 sw
rect 362 324 392 377
tri 392 324 408 340 sw
rect 168 286 274 316
tri 274 286 304 316 sw
rect 362 294 468 324
tri 468 294 498 324 sw
rect 168 185 198 286
tri 198 270 214 286 nw
tri 258 270 274 286 ne
tri 198 185 214 201 sw
tri 258 185 274 201 se
rect 274 185 304 286
rect 362 193 392 294
tri 392 278 408 294 nw
tri 452 278 468 294 ne
tri 392 193 408 209 sw
tri 452 193 468 209 se
rect 468 193 498 294
tri 168 155 198 185 ne
rect 198 155 274 185
tri 274 155 304 185 nw
tri 362 163 392 193 ne
rect 392 163 468 193
tri 468 163 498 193 nw
rect 813 318 843 379
tri 843 318 859 334 sw
rect 1113 318 1143 379
rect 813 288 919 318
tri 919 288 949 318 sw
rect 813 187 843 288
tri 843 272 859 288 nw
tri 903 272 919 288 ne
tri 843 187 859 203 sw
tri 903 187 919 203 se
rect 919 187 949 288
tri 1008 288 1038 318 se
rect 1038 288 1143 318
rect 1008 194 1038 288
tri 1038 272 1054 288 nw
tri 1097 272 1113 288 ne
tri 1038 194 1054 210 sw
tri 1097 194 1113 210 se
rect 1113 194 1143 288
tri 813 157 843 187 ne
rect 843 157 919 187
tri 919 157 949 187 nw
tri 1008 164 1038 194 ne
rect 1038 164 1113 194
tri 1113 164 1143 194 nw
rect 1315 326 1345 379
tri 1345 326 1361 342 sw
rect 1315 296 1421 326
tri 1421 296 1451 326 sw
rect 1315 195 1345 296
tri 1345 280 1361 296 nw
tri 1405 280 1421 296 ne
tri 1345 195 1361 211 sw
tri 1405 195 1421 211 se
rect 1421 195 1451 296
tri 1315 165 1345 195 ne
rect 1345 165 1421 195
tri 1421 165 1451 195 nw
rect 1775 318 1805 379
tri 1805 318 1821 334 sw
rect 2075 318 2105 379
rect 1775 288 1881 318
tri 1881 288 1911 318 sw
rect 1775 187 1805 288
tri 1805 272 1821 288 nw
tri 1865 272 1881 288 ne
tri 1805 187 1821 203 sw
tri 1865 187 1881 203 se
rect 1881 187 1911 288
tri 1970 288 2000 318 se
rect 2000 288 2105 318
rect 1970 194 2000 288
tri 2000 272 2016 288 nw
tri 2059 272 2075 288 ne
tri 2000 194 2016 210 sw
tri 2059 194 2075 210 se
rect 2075 194 2105 288
tri 1775 157 1805 187 ne
rect 1805 157 1881 187
tri 1881 157 1911 187 nw
tri 1970 164 2000 194 ne
rect 2000 164 2075 194
tri 2075 164 2105 194 nw
rect 2277 326 2307 379
tri 2307 326 2323 342 sw
rect 2277 296 2383 326
tri 2383 296 2413 326 sw
rect 2277 195 2307 296
tri 2307 280 2323 296 nw
tri 2367 280 2383 296 ne
tri 2307 195 2323 211 sw
tri 2367 195 2383 211 se
rect 2383 195 2413 296
tri 2277 165 2307 195 ne
rect 2307 165 2383 195
tri 2383 165 2413 195 nw
rect 2758 316 2788 377
tri 2788 316 2804 332 sw
rect 2952 324 2982 377
tri 2982 324 2998 340 sw
rect 2758 286 2864 316
tri 2864 286 2894 316 sw
rect 2952 294 3058 324
tri 3058 294 3088 324 sw
rect 2758 185 2788 286
tri 2788 270 2804 286 nw
tri 2848 270 2864 286 ne
tri 2788 185 2804 201 sw
tri 2848 185 2864 201 se
rect 2864 185 2894 286
rect 2952 193 2982 294
tri 2982 278 2998 294 nw
tri 3042 278 3058 294 ne
tri 2982 193 2998 209 sw
tri 3042 193 3058 209 se
rect 3058 193 3088 294
tri 2758 155 2788 185 ne
rect 2788 155 2864 185
tri 2864 155 2894 185 nw
tri 2952 163 2982 193 ne
rect 2982 163 3058 193
tri 3058 163 3088 193 nw
rect 3424 316 3454 377
tri 3454 316 3470 332 sw
rect 3618 324 3648 377
tri 3648 324 3664 340 sw
rect 3424 286 3530 316
tri 3530 286 3560 316 sw
rect 3618 294 3724 324
tri 3724 294 3754 324 sw
rect 3424 185 3454 286
tri 3454 270 3470 286 nw
tri 3514 270 3530 286 ne
tri 3454 185 3470 201 sw
tri 3514 185 3530 201 se
rect 3530 185 3560 286
rect 3618 193 3648 294
tri 3648 278 3664 294 nw
tri 3708 278 3724 294 ne
tri 3648 193 3664 209 sw
tri 3708 193 3724 209 se
rect 3724 193 3754 294
tri 3424 155 3454 185 ne
rect 3454 155 3530 185
tri 3530 155 3560 185 nw
tri 3618 163 3648 193 ne
rect 3648 163 3724 193
tri 3724 163 3754 193 nw
rect 4069 318 4099 379
tri 4099 318 4115 334 sw
rect 4369 318 4399 379
rect 4069 288 4175 318
tri 4175 288 4205 318 sw
rect 4069 187 4099 288
tri 4099 272 4115 288 nw
tri 4159 272 4175 288 ne
tri 4099 187 4115 203 sw
tri 4159 187 4175 203 se
rect 4175 187 4205 288
tri 4264 288 4294 318 se
rect 4294 288 4399 318
rect 4264 194 4294 288
tri 4294 272 4310 288 nw
tri 4353 272 4369 288 ne
tri 4294 194 4310 210 sw
tri 4353 194 4369 210 se
rect 4369 194 4399 288
tri 4069 157 4099 187 ne
rect 4099 157 4175 187
tri 4175 157 4205 187 nw
tri 4264 164 4294 194 ne
rect 4294 164 4369 194
tri 4369 164 4399 194 nw
rect 4571 326 4601 379
tri 4601 326 4617 342 sw
rect 4571 296 4677 326
tri 4677 296 4707 326 sw
rect 4571 195 4601 296
tri 4601 280 4617 296 nw
tri 4661 280 4677 296 ne
tri 4601 195 4617 211 sw
tri 4661 195 4677 211 se
rect 4677 195 4707 296
tri 4571 165 4601 195 ne
rect 4601 165 4677 195
tri 4677 165 4707 195 nw
rect 5052 316 5082 377
tri 5082 316 5098 332 sw
rect 5246 324 5276 377
tri 5276 324 5292 340 sw
rect 5052 286 5158 316
tri 5158 286 5188 316 sw
rect 5246 294 5352 324
tri 5352 294 5382 324 sw
rect 5052 185 5082 286
tri 5082 270 5098 286 nw
tri 5142 270 5158 286 ne
tri 5082 185 5098 201 sw
tri 5142 185 5158 201 se
rect 5158 185 5188 286
rect 5246 193 5276 294
tri 5276 278 5292 294 nw
tri 5336 278 5352 294 ne
tri 5276 193 5292 209 sw
tri 5336 193 5352 209 se
rect 5352 193 5382 294
tri 5052 155 5082 185 ne
rect 5082 155 5158 185
tri 5158 155 5188 185 nw
tri 5246 163 5276 193 ne
rect 5276 163 5352 193
tri 5352 163 5382 193 nw
rect 5697 318 5727 379
tri 5727 318 5743 334 sw
rect 5997 318 6027 379
rect 5697 288 5803 318
tri 5803 288 5833 318 sw
rect 5697 187 5727 288
tri 5727 272 5743 288 nw
tri 5787 272 5803 288 ne
tri 5727 187 5743 203 sw
tri 5787 187 5803 203 se
rect 5803 187 5833 288
tri 5892 288 5922 318 se
rect 5922 288 6027 318
rect 5892 194 5922 288
tri 5922 272 5938 288 nw
tri 5981 272 5997 288 ne
tri 5922 194 5938 210 sw
tri 5981 194 5997 210 se
rect 5997 194 6027 288
tri 5697 157 5727 187 ne
rect 5727 157 5803 187
tri 5803 157 5833 187 nw
tri 5892 164 5922 194 ne
rect 5922 164 5997 194
tri 5997 164 6027 194 nw
rect 6199 326 6229 379
tri 6229 326 6245 342 sw
rect 6199 296 6305 326
tri 6305 296 6335 326 sw
rect 6199 195 6229 296
tri 6229 280 6245 296 nw
tri 6289 280 6305 296 ne
tri 6229 195 6245 211 sw
tri 6289 195 6305 211 se
rect 6305 195 6335 296
tri 6199 165 6229 195 ne
rect 6229 165 6305 195
tri 6305 165 6335 195 nw
rect 6659 318 6689 379
tri 6689 318 6705 334 sw
rect 6959 318 6989 379
rect 6659 288 6765 318
tri 6765 288 6795 318 sw
rect 6659 187 6689 288
tri 6689 272 6705 288 nw
tri 6749 272 6765 288 ne
tri 6689 187 6705 203 sw
tri 6749 187 6765 203 se
rect 6765 187 6795 288
tri 6854 288 6884 318 se
rect 6884 288 6989 318
rect 6854 194 6884 288
tri 6884 272 6900 288 nw
tri 6943 272 6959 288 ne
tri 6884 194 6900 210 sw
tri 6943 194 6959 210 se
rect 6959 194 6989 288
tri 6659 157 6689 187 ne
rect 6689 157 6765 187
tri 6765 157 6795 187 nw
tri 6854 164 6884 194 ne
rect 6884 164 6959 194
tri 6959 164 6989 194 nw
rect 7161 326 7191 379
tri 7191 326 7207 342 sw
rect 7161 296 7267 326
tri 7267 296 7297 326 sw
rect 7161 195 7191 296
tri 7191 280 7207 296 nw
tri 7251 280 7267 296 ne
tri 7191 195 7207 211 sw
tri 7251 195 7267 211 se
rect 7267 195 7297 296
tri 7161 165 7191 195 ne
rect 7191 165 7267 195
tri 7267 165 7297 195 nw
rect 7642 316 7672 377
tri 7672 316 7688 332 sw
rect 7836 324 7866 377
tri 7866 324 7882 340 sw
rect 7642 286 7748 316
tri 7748 286 7778 316 sw
rect 7836 294 7942 324
tri 7942 294 7972 324 sw
rect 7642 185 7672 286
tri 7672 270 7688 286 nw
tri 7732 270 7748 286 ne
tri 7672 185 7688 201 sw
tri 7732 185 7748 201 se
rect 7748 185 7778 286
rect 7836 193 7866 294
tri 7866 278 7882 294 nw
tri 7926 278 7942 294 ne
tri 7866 193 7882 209 sw
tri 7926 193 7942 209 se
rect 7942 193 7972 294
tri 7642 155 7672 185 ne
rect 7672 155 7748 185
tri 7748 155 7778 185 nw
tri 7836 163 7866 193 ne
rect 7866 163 7942 193
tri 7942 163 7972 193 nw
rect 8308 316 8338 377
tri 8338 316 8354 332 sw
rect 8502 324 8532 377
tri 8532 324 8548 340 sw
rect 8308 286 8414 316
tri 8414 286 8444 316 sw
rect 8502 294 8608 324
tri 8608 294 8638 324 sw
rect 8308 185 8338 286
tri 8338 270 8354 286 nw
tri 8398 270 8414 286 ne
tri 8338 185 8354 201 sw
tri 8398 185 8414 201 se
rect 8414 185 8444 286
rect 8502 193 8532 294
tri 8532 278 8548 294 nw
tri 8592 278 8608 294 ne
tri 8532 193 8548 209 sw
tri 8592 193 8608 209 se
rect 8608 193 8638 294
tri 8308 155 8338 185 ne
rect 8338 155 8414 185
tri 8414 155 8444 185 nw
tri 8502 163 8532 193 ne
rect 8532 163 8608 193
tri 8608 163 8638 193 nw
rect 8953 318 8983 379
tri 8983 318 8999 334 sw
rect 9253 318 9283 379
rect 8953 288 9059 318
tri 9059 288 9089 318 sw
rect 8953 187 8983 288
tri 8983 272 8999 288 nw
tri 9043 272 9059 288 ne
tri 8983 187 8999 203 sw
tri 9043 187 9059 203 se
rect 9059 187 9089 288
tri 9148 288 9178 318 se
rect 9178 288 9283 318
rect 9148 194 9178 288
tri 9178 272 9194 288 nw
tri 9237 272 9253 288 ne
tri 9178 194 9194 210 sw
tri 9237 194 9253 210 se
rect 9253 194 9283 288
tri 8953 157 8983 187 ne
rect 8983 157 9059 187
tri 9059 157 9089 187 nw
tri 9148 164 9178 194 ne
rect 9178 164 9253 194
tri 9253 164 9283 194 nw
rect 9455 326 9485 379
tri 9485 326 9501 342 sw
rect 9455 296 9561 326
tri 9561 296 9591 326 sw
rect 9455 195 9485 296
tri 9485 280 9501 296 nw
tri 9545 280 9561 296 ne
tri 9485 195 9501 211 sw
tri 9545 195 9561 211 se
rect 9561 195 9591 296
tri 9455 165 9485 195 ne
rect 9485 165 9561 195
tri 9561 165 9591 195 nw
rect 9936 316 9966 377
tri 9966 316 9982 332 sw
rect 10130 324 10160 377
tri 10160 324 10176 340 sw
rect 9936 286 10042 316
tri 10042 286 10072 316 sw
rect 10130 294 10236 324
tri 10236 294 10266 324 sw
rect 9936 185 9966 286
tri 9966 270 9982 286 nw
tri 10026 270 10042 286 ne
tri 9966 185 9982 201 sw
tri 10026 185 10042 201 se
rect 10042 185 10072 286
rect 10130 193 10160 294
tri 10160 278 10176 294 nw
tri 10220 278 10236 294 ne
tri 10160 193 10176 209 sw
tri 10220 193 10236 209 se
rect 10236 193 10266 294
tri 9936 155 9966 185 ne
rect 9966 155 10042 185
tri 10042 155 10072 185 nw
tri 10130 163 10160 193 ne
rect 10160 163 10236 193
tri 10236 163 10266 193 nw
rect 10581 318 10611 379
tri 10611 318 10627 334 sw
rect 10881 318 10911 379
rect 10581 288 10687 318
tri 10687 288 10717 318 sw
rect 10581 187 10611 288
tri 10611 272 10627 288 nw
tri 10671 272 10687 288 ne
tri 10611 187 10627 203 sw
tri 10671 187 10687 203 se
rect 10687 187 10717 288
tri 10776 288 10806 318 se
rect 10806 288 10911 318
rect 10776 194 10806 288
tri 10806 272 10822 288 nw
tri 10865 272 10881 288 ne
tri 10806 194 10822 210 sw
tri 10865 194 10881 210 se
rect 10881 194 10911 288
tri 10581 157 10611 187 ne
rect 10611 157 10687 187
tri 10687 157 10717 187 nw
tri 10776 164 10806 194 ne
rect 10806 164 10881 194
tri 10881 164 10911 194 nw
rect 11083 326 11113 379
tri 11113 326 11129 342 sw
rect 11083 296 11189 326
tri 11189 296 11219 326 sw
rect 11083 195 11113 296
tri 11113 280 11129 296 nw
tri 11173 280 11189 296 ne
tri 11113 195 11129 211 sw
tri 11173 195 11189 211 se
rect 11189 195 11219 296
tri 11083 165 11113 195 ne
rect 11113 165 11189 195
tri 11189 165 11219 195 nw
rect 11543 318 11573 379
tri 11573 318 11589 334 sw
rect 11843 318 11873 379
rect 11543 288 11649 318
tri 11649 288 11679 318 sw
rect 11543 187 11573 288
tri 11573 272 11589 288 nw
tri 11633 272 11649 288 ne
tri 11573 187 11589 203 sw
tri 11633 187 11649 203 se
rect 11649 187 11679 288
tri 11738 288 11768 318 se
rect 11768 288 11873 318
rect 11738 194 11768 288
tri 11768 272 11784 288 nw
tri 11827 272 11843 288 ne
tri 11768 194 11784 210 sw
tri 11827 194 11843 210 se
rect 11843 194 11873 288
tri 11543 157 11573 187 ne
rect 11573 157 11649 187
tri 11649 157 11679 187 nw
tri 11738 164 11768 194 ne
rect 11768 164 11843 194
tri 11843 164 11873 194 nw
rect 12045 326 12075 379
tri 12075 326 12091 342 sw
rect 12045 296 12151 326
tri 12151 296 12181 326 sw
rect 12045 195 12075 296
tri 12075 280 12091 296 nw
tri 12135 280 12151 296 ne
tri 12075 195 12091 211 sw
tri 12135 195 12151 211 se
rect 12151 195 12181 296
tri 12045 165 12075 195 ne
rect 12075 165 12151 195
tri 12151 165 12181 195 nw
rect 12526 316 12556 377
tri 12556 316 12572 332 sw
rect 12720 324 12750 377
tri 12750 324 12766 340 sw
rect 12526 286 12632 316
tri 12632 286 12662 316 sw
rect 12720 294 12826 324
tri 12826 294 12856 324 sw
rect 12526 185 12556 286
tri 12556 270 12572 286 nw
tri 12616 270 12632 286 ne
tri 12556 185 12572 201 sw
tri 12616 185 12632 201 se
rect 12632 185 12662 286
rect 12720 193 12750 294
tri 12750 278 12766 294 nw
tri 12810 278 12826 294 ne
tri 12750 193 12766 209 sw
tri 12810 193 12826 209 se
rect 12826 193 12856 294
tri 12526 155 12556 185 ne
rect 12556 155 12632 185
tri 12632 155 12662 185 nw
tri 12720 163 12750 193 ne
rect 12750 163 12826 193
tri 12826 163 12856 193 nw
rect 13192 316 13222 377
tri 13222 316 13238 332 sw
rect 13386 324 13416 377
tri 13416 324 13432 340 sw
rect 13192 286 13298 316
tri 13298 286 13328 316 sw
rect 13386 294 13492 324
tri 13492 294 13522 324 sw
rect 13192 185 13222 286
tri 13222 270 13238 286 nw
tri 13282 270 13298 286 ne
tri 13222 185 13238 201 sw
tri 13282 185 13298 201 se
rect 13298 185 13328 286
rect 13386 193 13416 294
tri 13416 278 13432 294 nw
tri 13476 278 13492 294 ne
tri 13416 193 13432 209 sw
tri 13476 193 13492 209 se
rect 13492 193 13522 294
tri 13192 155 13222 185 ne
rect 13222 155 13298 185
tri 13298 155 13328 185 nw
tri 13386 163 13416 193 ne
rect 13416 163 13492 193
tri 13492 163 13522 193 nw
rect 13837 318 13867 379
tri 13867 318 13883 334 sw
rect 14137 318 14167 379
rect 13837 288 13943 318
tri 13943 288 13973 318 sw
rect 13837 187 13867 288
tri 13867 272 13883 288 nw
tri 13927 272 13943 288 ne
tri 13867 187 13883 203 sw
tri 13927 187 13943 203 se
rect 13943 187 13973 288
tri 14032 288 14062 318 se
rect 14062 288 14167 318
rect 14032 194 14062 288
tri 14062 272 14078 288 nw
tri 14121 272 14137 288 ne
tri 14062 194 14078 210 sw
tri 14121 194 14137 210 se
rect 14137 194 14167 288
tri 13837 157 13867 187 ne
rect 13867 157 13943 187
tri 13943 157 13973 187 nw
tri 14032 164 14062 194 ne
rect 14062 164 14137 194
tri 14137 164 14167 194 nw
rect 14339 326 14369 379
tri 14369 326 14385 342 sw
rect 14339 296 14445 326
tri 14445 296 14475 326 sw
rect 14339 195 14369 296
tri 14369 280 14385 296 nw
tri 14429 280 14445 296 ne
tri 14369 195 14385 211 sw
tri 14429 195 14445 211 se
rect 14445 195 14475 296
tri 14339 165 14369 195 ne
rect 14369 165 14445 195
tri 14445 165 14475 195 nw
rect 14820 316 14850 377
tri 14850 316 14866 332 sw
rect 15014 324 15044 377
tri 15044 324 15060 340 sw
rect 14820 286 14926 316
tri 14926 286 14956 316 sw
rect 15014 294 15120 324
tri 15120 294 15150 324 sw
rect 14820 185 14850 286
tri 14850 270 14866 286 nw
tri 14910 270 14926 286 ne
tri 14850 185 14866 201 sw
tri 14910 185 14926 201 se
rect 14926 185 14956 286
rect 15014 193 15044 294
tri 15044 278 15060 294 nw
tri 15104 278 15120 294 ne
tri 15044 193 15060 209 sw
tri 15104 193 15120 209 se
rect 15120 193 15150 294
tri 14820 155 14850 185 ne
rect 14850 155 14926 185
tri 14926 155 14956 185 nw
tri 15014 163 15044 193 ne
rect 15044 163 15120 193
tri 15120 163 15150 193 nw
rect 15486 316 15516 377
tri 15516 316 15532 332 sw
tri 15770 324 15786 340 se
rect 15786 324 15816 377
rect 15486 286 15592 316
tri 15592 286 15622 316 sw
tri 15680 294 15710 324 se
rect 15710 294 15816 324
rect 15486 185 15516 286
tri 15516 270 15532 286 nw
tri 15576 270 15592 286 ne
tri 15516 185 15532 201 sw
tri 15576 185 15592 201 se
rect 15592 185 15622 286
rect 15680 193 15710 294
tri 15710 278 15726 294 nw
tri 15770 278 15786 294 ne
tri 15710 193 15726 209 sw
tri 15770 193 15786 209 se
rect 15786 193 15816 294
tri 15486 155 15516 185 ne
rect 15516 155 15592 185
tri 15592 155 15622 185 nw
tri 15680 163 15710 193 ne
rect 15710 163 15786 193
tri 15786 163 15816 193 nw
rect 16152 316 16182 377
tri 16182 316 16198 332 sw
rect 16346 324 16376 377
tri 16376 324 16392 340 sw
rect 16152 286 16258 316
tri 16258 286 16288 316 sw
rect 16346 294 16452 324
tri 16452 294 16482 324 sw
rect 16152 185 16182 286
tri 16182 270 16198 286 nw
tri 16242 270 16258 286 ne
tri 16182 185 16198 201 sw
tri 16242 185 16258 201 se
rect 16258 185 16288 286
rect 16346 279 16377 294
tri 16377 279 16392 294 nw
tri 16436 279 16451 294 ne
rect 16451 279 16482 294
rect 16346 193 16376 279
tri 16376 193 16392 209 sw
tri 16436 193 16452 209 se
rect 16452 193 16482 279
tri 16152 155 16182 185 ne
rect 16182 155 16258 185
tri 16258 155 16288 185 nw
tri 16346 163 16376 193 ne
rect 16376 163 16452 193
tri 16452 163 16482 193 nw
<< pmos >>
rect 187 1050 217 1450
rect 275 1050 305 1450
rect 363 1050 393 1450
rect 451 1050 481 1450
rect 913 1050 943 1450
rect 1001 1050 1031 1450
rect 1089 1050 1119 1450
rect 1177 1050 1207 1450
rect 1265 1050 1295 1450
rect 1353 1050 1383 1450
rect 1875 1050 1905 1450
rect 1963 1050 1993 1450
rect 2051 1050 2081 1450
rect 2139 1050 2169 1450
rect 2227 1050 2257 1450
rect 2315 1050 2345 1450
rect 2777 1050 2807 1450
rect 2865 1050 2895 1450
rect 2953 1050 2983 1450
rect 3041 1050 3071 1450
rect 3443 1050 3473 1450
rect 3531 1050 3561 1450
rect 3619 1050 3649 1450
rect 3707 1050 3737 1450
rect 4169 1050 4199 1450
rect 4257 1050 4287 1450
rect 4345 1050 4375 1450
rect 4433 1050 4463 1450
rect 4521 1050 4551 1450
rect 4609 1050 4639 1450
rect 5071 1050 5101 1450
rect 5159 1050 5189 1450
rect 5247 1050 5277 1450
rect 5335 1050 5365 1450
rect 5797 1050 5827 1450
rect 5885 1050 5915 1450
rect 5973 1050 6003 1450
rect 6061 1050 6091 1450
rect 6149 1050 6179 1450
rect 6237 1050 6267 1450
rect 6759 1050 6789 1450
rect 6847 1050 6877 1450
rect 6935 1050 6965 1450
rect 7023 1050 7053 1450
rect 7111 1050 7141 1450
rect 7199 1050 7229 1450
rect 7661 1050 7691 1450
rect 7749 1050 7779 1450
rect 7837 1050 7867 1450
rect 7925 1050 7955 1450
rect 8327 1050 8357 1450
rect 8415 1050 8445 1450
rect 8503 1050 8533 1450
rect 8591 1050 8621 1450
rect 9053 1050 9083 1450
rect 9141 1050 9171 1450
rect 9229 1050 9259 1450
rect 9317 1050 9347 1450
rect 9405 1050 9435 1450
rect 9493 1050 9523 1450
rect 9955 1050 9985 1450
rect 10043 1050 10073 1450
rect 10131 1050 10161 1450
rect 10219 1050 10249 1450
rect 10681 1050 10711 1450
rect 10769 1050 10799 1450
rect 10857 1050 10887 1450
rect 10945 1050 10975 1450
rect 11033 1050 11063 1450
rect 11121 1050 11151 1450
rect 11643 1050 11673 1450
rect 11731 1050 11761 1450
rect 11819 1050 11849 1450
rect 11907 1050 11937 1450
rect 11995 1050 12025 1450
rect 12083 1050 12113 1450
rect 12545 1050 12575 1450
rect 12633 1050 12663 1450
rect 12721 1050 12751 1450
rect 12809 1050 12839 1450
rect 13211 1050 13241 1450
rect 13299 1050 13329 1450
rect 13387 1050 13417 1450
rect 13475 1050 13505 1450
rect 13937 1050 13967 1450
rect 14025 1050 14055 1450
rect 14113 1050 14143 1450
rect 14201 1050 14231 1450
rect 14289 1050 14319 1450
rect 14377 1050 14407 1450
rect 14839 1051 14869 1451
rect 14927 1051 14957 1451
rect 15015 1051 15045 1451
rect 15103 1051 15133 1451
rect 15503 1051 15533 1451
rect 15591 1051 15621 1451
rect 15679 1051 15709 1451
rect 15767 1051 15797 1451
rect 16171 1051 16201 1451
rect 16259 1051 16289 1451
rect 16347 1051 16377 1451
rect 16435 1051 16465 1451
<< ndiff >>
rect 112 361 168 377
rect 112 327 122 361
rect 156 327 168 361
rect 112 289 168 327
rect 198 361 362 377
rect 198 332 219 361
tri 198 316 214 332 ne
rect 214 327 219 332
rect 253 327 316 361
rect 350 327 362 361
rect 214 316 362 327
rect 392 340 554 377
tri 392 324 408 340 ne
rect 408 324 554 340
rect 112 255 122 289
rect 156 255 168 289
tri 274 286 304 316 ne
rect 304 289 362 316
tri 468 294 498 324 ne
rect 112 221 168 255
rect 112 187 122 221
rect 156 187 168 221
rect 112 155 168 187
tri 198 270 214 286 se
rect 214 270 258 286
tri 258 270 274 286 sw
rect 198 236 274 270
rect 198 202 219 236
rect 253 202 274 236
rect 198 201 274 202
tri 198 185 214 201 ne
rect 214 185 258 201
tri 258 185 274 201 nw
rect 304 255 316 289
rect 350 255 362 289
rect 304 221 362 255
rect 304 187 316 221
rect 350 187 362 221
tri 392 278 408 294 se
rect 408 278 452 294
tri 452 278 468 294 sw
rect 392 245 468 278
rect 392 211 413 245
rect 447 211 468 245
rect 392 209 468 211
tri 392 193 408 209 ne
rect 408 193 452 209
tri 452 193 468 209 nw
rect 498 289 554 324
rect 498 255 510 289
rect 544 255 554 289
rect 498 221 554 255
tri 168 155 198 185 sw
tri 274 155 304 185 se
rect 304 163 362 187
tri 362 163 392 193 sw
tri 468 163 498 193 se
rect 498 187 510 221
rect 544 187 554 221
rect 498 163 554 187
rect 304 155 554 163
rect 112 151 554 155
rect 112 117 122 151
rect 156 117 316 151
rect 350 117 413 151
rect 447 117 510 151
rect 544 117 554 151
rect 112 101 554 117
rect 757 363 813 379
rect 757 329 767 363
rect 801 329 813 363
rect 757 291 813 329
rect 843 363 1113 379
rect 843 334 864 363
tri 843 318 859 334 ne
rect 859 329 864 334
rect 898 329 961 363
rect 995 329 1058 363
rect 1092 329 1113 363
rect 859 318 1113 329
rect 1143 363 1199 379
rect 1143 329 1155 363
rect 1189 329 1199 363
rect 757 257 767 291
rect 801 257 813 291
tri 919 288 949 318 ne
rect 949 291 1008 318
rect 757 223 813 257
rect 757 189 767 223
rect 801 189 813 223
rect 757 157 813 189
tri 843 272 859 288 se
rect 859 272 903 288
tri 903 272 919 288 sw
rect 843 238 919 272
rect 843 204 864 238
rect 898 204 919 238
rect 843 203 919 204
tri 843 187 859 203 ne
rect 859 187 903 203
tri 903 187 919 203 nw
rect 949 257 961 291
rect 995 257 1008 291
tri 1008 288 1038 318 nw
rect 949 223 1008 257
rect 949 189 961 223
rect 995 189 1008 223
tri 1038 272 1054 288 se
rect 1054 272 1097 288
tri 1097 272 1113 288 sw
rect 1038 244 1113 272
rect 1038 210 1059 244
rect 1093 210 1113 244
tri 1038 194 1054 210 ne
rect 1054 194 1097 210
tri 1097 194 1113 210 nw
tri 813 157 843 187 sw
tri 919 157 949 187 se
rect 949 164 1008 189
tri 1008 164 1038 194 sw
tri 1113 164 1143 194 se
rect 1143 164 1199 329
rect 949 157 1199 164
rect 757 153 1199 157
rect 757 119 767 153
rect 801 119 961 153
rect 995 119 1058 153
rect 1092 119 1155 153
rect 1189 119 1199 153
rect 757 103 1199 119
rect 1259 363 1315 379
rect 1259 329 1269 363
rect 1303 329 1315 363
rect 1259 291 1315 329
rect 1345 342 1507 379
tri 1345 326 1361 342 ne
rect 1361 326 1507 342
tri 1421 296 1451 326 ne
rect 1259 257 1269 291
rect 1303 257 1315 291
rect 1259 223 1315 257
rect 1259 189 1269 223
rect 1303 189 1315 223
tri 1345 280 1361 296 se
rect 1361 280 1405 296
tri 1405 280 1421 296 sw
rect 1345 247 1421 280
rect 1345 213 1366 247
rect 1400 213 1421 247
rect 1345 211 1421 213
tri 1345 195 1361 211 ne
rect 1361 195 1405 211
tri 1405 195 1421 211 nw
rect 1451 291 1507 326
rect 1451 257 1463 291
rect 1497 257 1507 291
rect 1451 223 1507 257
rect 1259 165 1315 189
tri 1315 165 1345 195 sw
tri 1421 165 1451 195 se
rect 1451 189 1463 223
rect 1497 189 1507 223
rect 1451 165 1507 189
rect 1259 153 1507 165
rect 1259 119 1269 153
rect 1303 119 1366 153
rect 1400 119 1463 153
rect 1497 119 1507 153
rect 1259 103 1507 119
rect 1719 363 1775 379
rect 1719 329 1729 363
rect 1763 329 1775 363
rect 1719 291 1775 329
rect 1805 363 2075 379
rect 1805 334 1826 363
tri 1805 318 1821 334 ne
rect 1821 329 1826 334
rect 1860 329 1923 363
rect 1957 329 2020 363
rect 2054 329 2075 363
rect 1821 318 2075 329
rect 2105 363 2161 379
rect 2105 329 2117 363
rect 2151 329 2161 363
rect 1719 257 1729 291
rect 1763 257 1775 291
tri 1881 288 1911 318 ne
rect 1911 291 1970 318
rect 1719 223 1775 257
rect 1719 189 1729 223
rect 1763 189 1775 223
rect 1719 157 1775 189
tri 1805 272 1821 288 se
rect 1821 272 1865 288
tri 1865 272 1881 288 sw
rect 1805 238 1881 272
rect 1805 204 1826 238
rect 1860 204 1881 238
rect 1805 203 1881 204
tri 1805 187 1821 203 ne
rect 1821 187 1865 203
tri 1865 187 1881 203 nw
rect 1911 257 1923 291
rect 1957 257 1970 291
tri 1970 288 2000 318 nw
rect 1911 223 1970 257
rect 1911 189 1923 223
rect 1957 189 1970 223
tri 2000 272 2016 288 se
rect 2016 272 2059 288
tri 2059 272 2075 288 sw
rect 2000 244 2075 272
rect 2000 210 2021 244
rect 2055 210 2075 244
tri 2000 194 2016 210 ne
rect 2016 194 2059 210
tri 2059 194 2075 210 nw
tri 1775 157 1805 187 sw
tri 1881 157 1911 187 se
rect 1911 164 1970 189
tri 1970 164 2000 194 sw
tri 2075 164 2105 194 se
rect 2105 164 2161 329
rect 1911 157 2161 164
rect 1719 153 2161 157
rect 1719 119 1729 153
rect 1763 119 1923 153
rect 1957 119 2020 153
rect 2054 119 2117 153
rect 2151 119 2161 153
rect 1719 103 2161 119
rect 2221 363 2277 379
rect 2221 329 2231 363
rect 2265 329 2277 363
rect 2221 291 2277 329
rect 2307 342 2469 379
tri 2307 326 2323 342 ne
rect 2323 326 2469 342
tri 2383 296 2413 326 ne
rect 2221 257 2231 291
rect 2265 257 2277 291
rect 2221 223 2277 257
rect 2221 189 2231 223
rect 2265 189 2277 223
tri 2307 280 2323 296 se
rect 2323 280 2367 296
tri 2367 280 2383 296 sw
rect 2307 247 2383 280
rect 2307 213 2328 247
rect 2362 213 2383 247
rect 2307 211 2383 213
tri 2307 195 2323 211 ne
rect 2323 195 2367 211
tri 2367 195 2383 211 nw
rect 2413 291 2469 326
rect 2413 257 2425 291
rect 2459 257 2469 291
rect 2413 223 2469 257
rect 2221 165 2277 189
tri 2277 165 2307 195 sw
tri 2383 165 2413 195 se
rect 2413 189 2425 223
rect 2459 189 2469 223
rect 2413 165 2469 189
rect 2221 153 2469 165
rect 2221 119 2231 153
rect 2265 119 2328 153
rect 2362 119 2425 153
rect 2459 119 2469 153
rect 2221 103 2469 119
rect 2702 361 2758 377
rect 2702 327 2712 361
rect 2746 327 2758 361
rect 2702 289 2758 327
rect 2788 361 2952 377
rect 2788 332 2809 361
tri 2788 316 2804 332 ne
rect 2804 327 2809 332
rect 2843 327 2906 361
rect 2940 327 2952 361
rect 2804 316 2952 327
rect 2982 340 3144 377
tri 2982 324 2998 340 ne
rect 2998 324 3144 340
rect 2702 255 2712 289
rect 2746 255 2758 289
tri 2864 286 2894 316 ne
rect 2894 289 2952 316
tri 3058 294 3088 324 ne
rect 2702 221 2758 255
rect 2702 187 2712 221
rect 2746 187 2758 221
rect 2702 155 2758 187
tri 2788 270 2804 286 se
rect 2804 270 2848 286
tri 2848 270 2864 286 sw
rect 2788 236 2864 270
rect 2788 202 2809 236
rect 2843 202 2864 236
rect 2788 201 2864 202
tri 2788 185 2804 201 ne
rect 2804 185 2848 201
tri 2848 185 2864 201 nw
rect 2894 255 2906 289
rect 2940 255 2952 289
rect 2894 221 2952 255
rect 2894 187 2906 221
rect 2940 187 2952 221
tri 2982 278 2998 294 se
rect 2998 278 3042 294
tri 3042 278 3058 294 sw
rect 2982 245 3058 278
rect 2982 211 3003 245
rect 3037 211 3058 245
rect 2982 209 3058 211
tri 2982 193 2998 209 ne
rect 2998 193 3042 209
tri 3042 193 3058 209 nw
rect 3088 289 3144 324
rect 3088 255 3100 289
rect 3134 255 3144 289
rect 3088 221 3144 255
tri 2758 155 2788 185 sw
tri 2864 155 2894 185 se
rect 2894 163 2952 187
tri 2952 163 2982 193 sw
tri 3058 163 3088 193 se
rect 3088 187 3100 221
rect 3134 187 3144 221
rect 3088 163 3144 187
rect 2894 155 3144 163
rect 2702 151 3144 155
rect 2702 117 2712 151
rect 2746 117 2906 151
rect 2940 117 3003 151
rect 3037 117 3100 151
rect 3134 117 3144 151
rect 2702 101 3144 117
rect 3368 361 3424 377
rect 3368 327 3378 361
rect 3412 327 3424 361
rect 3368 289 3424 327
rect 3454 361 3618 377
rect 3454 332 3475 361
tri 3454 316 3470 332 ne
rect 3470 327 3475 332
rect 3509 327 3572 361
rect 3606 327 3618 361
rect 3470 316 3618 327
rect 3648 340 3810 377
tri 3648 324 3664 340 ne
rect 3664 324 3810 340
rect 3368 255 3378 289
rect 3412 255 3424 289
tri 3530 286 3560 316 ne
rect 3560 289 3618 316
tri 3724 294 3754 324 ne
rect 3368 221 3424 255
rect 3368 187 3378 221
rect 3412 187 3424 221
rect 3368 155 3424 187
tri 3454 270 3470 286 se
rect 3470 270 3514 286
tri 3514 270 3530 286 sw
rect 3454 236 3530 270
rect 3454 202 3475 236
rect 3509 202 3530 236
rect 3454 201 3530 202
tri 3454 185 3470 201 ne
rect 3470 185 3514 201
tri 3514 185 3530 201 nw
rect 3560 255 3572 289
rect 3606 255 3618 289
rect 3560 221 3618 255
rect 3560 187 3572 221
rect 3606 187 3618 221
tri 3648 278 3664 294 se
rect 3664 278 3708 294
tri 3708 278 3724 294 sw
rect 3648 245 3724 278
rect 3648 211 3669 245
rect 3703 211 3724 245
rect 3648 209 3724 211
tri 3648 193 3664 209 ne
rect 3664 193 3708 209
tri 3708 193 3724 209 nw
rect 3754 289 3810 324
rect 3754 255 3766 289
rect 3800 255 3810 289
rect 3754 221 3810 255
tri 3424 155 3454 185 sw
tri 3530 155 3560 185 se
rect 3560 163 3618 187
tri 3618 163 3648 193 sw
tri 3724 163 3754 193 se
rect 3754 187 3766 221
rect 3800 187 3810 221
rect 3754 163 3810 187
rect 3560 155 3810 163
rect 3368 151 3810 155
rect 3368 117 3378 151
rect 3412 117 3572 151
rect 3606 117 3669 151
rect 3703 117 3766 151
rect 3800 117 3810 151
rect 3368 101 3810 117
rect 4013 363 4069 379
rect 4013 329 4023 363
rect 4057 329 4069 363
rect 4013 291 4069 329
rect 4099 363 4369 379
rect 4099 334 4120 363
tri 4099 318 4115 334 ne
rect 4115 329 4120 334
rect 4154 329 4217 363
rect 4251 329 4314 363
rect 4348 329 4369 363
rect 4115 318 4369 329
rect 4399 363 4455 379
rect 4399 329 4411 363
rect 4445 329 4455 363
rect 4013 257 4023 291
rect 4057 257 4069 291
tri 4175 288 4205 318 ne
rect 4205 291 4264 318
rect 4013 223 4069 257
rect 4013 189 4023 223
rect 4057 189 4069 223
rect 4013 157 4069 189
tri 4099 272 4115 288 se
rect 4115 272 4159 288
tri 4159 272 4175 288 sw
rect 4099 238 4175 272
rect 4099 204 4120 238
rect 4154 204 4175 238
rect 4099 203 4175 204
tri 4099 187 4115 203 ne
rect 4115 187 4159 203
tri 4159 187 4175 203 nw
rect 4205 257 4217 291
rect 4251 257 4264 291
tri 4264 288 4294 318 nw
rect 4205 223 4264 257
rect 4205 189 4217 223
rect 4251 189 4264 223
tri 4294 272 4310 288 se
rect 4310 272 4353 288
tri 4353 272 4369 288 sw
rect 4294 244 4369 272
rect 4294 210 4315 244
rect 4349 210 4369 244
tri 4294 194 4310 210 ne
rect 4310 194 4353 210
tri 4353 194 4369 210 nw
tri 4069 157 4099 187 sw
tri 4175 157 4205 187 se
rect 4205 164 4264 189
tri 4264 164 4294 194 sw
tri 4369 164 4399 194 se
rect 4399 164 4455 329
rect 4205 157 4455 164
rect 4013 153 4455 157
rect 4013 119 4023 153
rect 4057 119 4217 153
rect 4251 119 4314 153
rect 4348 119 4411 153
rect 4445 119 4455 153
rect 4013 103 4455 119
rect 4515 363 4571 379
rect 4515 329 4525 363
rect 4559 329 4571 363
rect 4515 291 4571 329
rect 4601 342 4763 379
tri 4601 326 4617 342 ne
rect 4617 326 4763 342
tri 4677 296 4707 326 ne
rect 4515 257 4525 291
rect 4559 257 4571 291
rect 4515 223 4571 257
rect 4515 189 4525 223
rect 4559 189 4571 223
tri 4601 280 4617 296 se
rect 4617 280 4661 296
tri 4661 280 4677 296 sw
rect 4601 247 4677 280
rect 4601 213 4622 247
rect 4656 213 4677 247
rect 4601 211 4677 213
tri 4601 195 4617 211 ne
rect 4617 195 4661 211
tri 4661 195 4677 211 nw
rect 4707 291 4763 326
rect 4707 257 4719 291
rect 4753 257 4763 291
rect 4707 223 4763 257
rect 4515 165 4571 189
tri 4571 165 4601 195 sw
tri 4677 165 4707 195 se
rect 4707 189 4719 223
rect 4753 189 4763 223
rect 4707 165 4763 189
rect 4515 153 4763 165
rect 4515 119 4525 153
rect 4559 119 4622 153
rect 4656 119 4719 153
rect 4753 119 4763 153
rect 4515 103 4763 119
rect 4996 361 5052 377
rect 4996 327 5006 361
rect 5040 327 5052 361
rect 4996 289 5052 327
rect 5082 361 5246 377
rect 5082 332 5103 361
tri 5082 316 5098 332 ne
rect 5098 327 5103 332
rect 5137 327 5200 361
rect 5234 327 5246 361
rect 5098 316 5246 327
rect 5276 340 5438 377
tri 5276 324 5292 340 ne
rect 5292 324 5438 340
rect 4996 255 5006 289
rect 5040 255 5052 289
tri 5158 286 5188 316 ne
rect 5188 289 5246 316
tri 5352 294 5382 324 ne
rect 4996 221 5052 255
rect 4996 187 5006 221
rect 5040 187 5052 221
rect 4996 155 5052 187
tri 5082 270 5098 286 se
rect 5098 270 5142 286
tri 5142 270 5158 286 sw
rect 5082 236 5158 270
rect 5082 202 5103 236
rect 5137 202 5158 236
rect 5082 201 5158 202
tri 5082 185 5098 201 ne
rect 5098 185 5142 201
tri 5142 185 5158 201 nw
rect 5188 255 5200 289
rect 5234 255 5246 289
rect 5188 221 5246 255
rect 5188 187 5200 221
rect 5234 187 5246 221
tri 5276 278 5292 294 se
rect 5292 278 5336 294
tri 5336 278 5352 294 sw
rect 5276 245 5352 278
rect 5276 211 5297 245
rect 5331 211 5352 245
rect 5276 209 5352 211
tri 5276 193 5292 209 ne
rect 5292 193 5336 209
tri 5336 193 5352 209 nw
rect 5382 289 5438 324
rect 5382 255 5394 289
rect 5428 255 5438 289
rect 5382 221 5438 255
tri 5052 155 5082 185 sw
tri 5158 155 5188 185 se
rect 5188 163 5246 187
tri 5246 163 5276 193 sw
tri 5352 163 5382 193 se
rect 5382 187 5394 221
rect 5428 187 5438 221
rect 5382 163 5438 187
rect 5188 155 5438 163
rect 4996 151 5438 155
rect 4996 117 5006 151
rect 5040 117 5200 151
rect 5234 117 5297 151
rect 5331 117 5394 151
rect 5428 117 5438 151
rect 4996 101 5438 117
rect 5641 363 5697 379
rect 5641 329 5651 363
rect 5685 329 5697 363
rect 5641 291 5697 329
rect 5727 363 5997 379
rect 5727 334 5748 363
tri 5727 318 5743 334 ne
rect 5743 329 5748 334
rect 5782 329 5845 363
rect 5879 329 5942 363
rect 5976 329 5997 363
rect 5743 318 5997 329
rect 6027 363 6083 379
rect 6027 329 6039 363
rect 6073 329 6083 363
rect 5641 257 5651 291
rect 5685 257 5697 291
tri 5803 288 5833 318 ne
rect 5833 291 5892 318
rect 5641 223 5697 257
rect 5641 189 5651 223
rect 5685 189 5697 223
rect 5641 157 5697 189
tri 5727 272 5743 288 se
rect 5743 272 5787 288
tri 5787 272 5803 288 sw
rect 5727 238 5803 272
rect 5727 204 5748 238
rect 5782 204 5803 238
rect 5727 203 5803 204
tri 5727 187 5743 203 ne
rect 5743 187 5787 203
tri 5787 187 5803 203 nw
rect 5833 257 5845 291
rect 5879 257 5892 291
tri 5892 288 5922 318 nw
rect 5833 223 5892 257
rect 5833 189 5845 223
rect 5879 189 5892 223
tri 5922 272 5938 288 se
rect 5938 272 5981 288
tri 5981 272 5997 288 sw
rect 5922 244 5997 272
rect 5922 210 5943 244
rect 5977 210 5997 244
tri 5922 194 5938 210 ne
rect 5938 194 5981 210
tri 5981 194 5997 210 nw
tri 5697 157 5727 187 sw
tri 5803 157 5833 187 se
rect 5833 164 5892 189
tri 5892 164 5922 194 sw
tri 5997 164 6027 194 se
rect 6027 164 6083 329
rect 5833 157 6083 164
rect 5641 153 6083 157
rect 5641 119 5651 153
rect 5685 119 5845 153
rect 5879 119 5942 153
rect 5976 119 6039 153
rect 6073 119 6083 153
rect 5641 103 6083 119
rect 6143 363 6199 379
rect 6143 329 6153 363
rect 6187 329 6199 363
rect 6143 291 6199 329
rect 6229 342 6391 379
tri 6229 326 6245 342 ne
rect 6245 326 6391 342
tri 6305 296 6335 326 ne
rect 6143 257 6153 291
rect 6187 257 6199 291
rect 6143 223 6199 257
rect 6143 189 6153 223
rect 6187 189 6199 223
tri 6229 280 6245 296 se
rect 6245 280 6289 296
tri 6289 280 6305 296 sw
rect 6229 247 6305 280
rect 6229 213 6250 247
rect 6284 213 6305 247
rect 6229 211 6305 213
tri 6229 195 6245 211 ne
rect 6245 195 6289 211
tri 6289 195 6305 211 nw
rect 6335 291 6391 326
rect 6335 257 6347 291
rect 6381 257 6391 291
rect 6335 223 6391 257
rect 6143 165 6199 189
tri 6199 165 6229 195 sw
tri 6305 165 6335 195 se
rect 6335 189 6347 223
rect 6381 189 6391 223
rect 6335 165 6391 189
rect 6143 153 6391 165
rect 6143 119 6153 153
rect 6187 119 6250 153
rect 6284 119 6347 153
rect 6381 119 6391 153
rect 6143 103 6391 119
rect 6603 363 6659 379
rect 6603 329 6613 363
rect 6647 329 6659 363
rect 6603 291 6659 329
rect 6689 363 6959 379
rect 6689 334 6710 363
tri 6689 318 6705 334 ne
rect 6705 329 6710 334
rect 6744 329 6807 363
rect 6841 329 6904 363
rect 6938 329 6959 363
rect 6705 318 6959 329
rect 6989 363 7045 379
rect 6989 329 7001 363
rect 7035 329 7045 363
rect 6603 257 6613 291
rect 6647 257 6659 291
tri 6765 288 6795 318 ne
rect 6795 291 6854 318
rect 6603 223 6659 257
rect 6603 189 6613 223
rect 6647 189 6659 223
rect 6603 157 6659 189
tri 6689 272 6705 288 se
rect 6705 272 6749 288
tri 6749 272 6765 288 sw
rect 6689 238 6765 272
rect 6689 204 6710 238
rect 6744 204 6765 238
rect 6689 203 6765 204
tri 6689 187 6705 203 ne
rect 6705 187 6749 203
tri 6749 187 6765 203 nw
rect 6795 257 6807 291
rect 6841 257 6854 291
tri 6854 288 6884 318 nw
rect 6795 223 6854 257
rect 6795 189 6807 223
rect 6841 189 6854 223
tri 6884 272 6900 288 se
rect 6900 272 6943 288
tri 6943 272 6959 288 sw
rect 6884 244 6959 272
rect 6884 210 6905 244
rect 6939 210 6959 244
tri 6884 194 6900 210 ne
rect 6900 194 6943 210
tri 6943 194 6959 210 nw
tri 6659 157 6689 187 sw
tri 6765 157 6795 187 se
rect 6795 164 6854 189
tri 6854 164 6884 194 sw
tri 6959 164 6989 194 se
rect 6989 164 7045 329
rect 6795 157 7045 164
rect 6603 153 7045 157
rect 6603 119 6613 153
rect 6647 119 6807 153
rect 6841 119 6904 153
rect 6938 119 7001 153
rect 7035 119 7045 153
rect 6603 103 7045 119
rect 7105 363 7161 379
rect 7105 329 7115 363
rect 7149 329 7161 363
rect 7105 291 7161 329
rect 7191 342 7353 379
tri 7191 326 7207 342 ne
rect 7207 326 7353 342
tri 7267 296 7297 326 ne
rect 7105 257 7115 291
rect 7149 257 7161 291
rect 7105 223 7161 257
rect 7105 189 7115 223
rect 7149 189 7161 223
tri 7191 280 7207 296 se
rect 7207 280 7251 296
tri 7251 280 7267 296 sw
rect 7191 247 7267 280
rect 7191 213 7212 247
rect 7246 213 7267 247
rect 7191 211 7267 213
tri 7191 195 7207 211 ne
rect 7207 195 7251 211
tri 7251 195 7267 211 nw
rect 7297 291 7353 326
rect 7297 257 7309 291
rect 7343 257 7353 291
rect 7297 223 7353 257
rect 7105 165 7161 189
tri 7161 165 7191 195 sw
tri 7267 165 7297 195 se
rect 7297 189 7309 223
rect 7343 189 7353 223
rect 7297 165 7353 189
rect 7105 153 7353 165
rect 7105 119 7115 153
rect 7149 119 7212 153
rect 7246 119 7309 153
rect 7343 119 7353 153
rect 7105 103 7353 119
rect 7586 361 7642 377
rect 7586 327 7596 361
rect 7630 327 7642 361
rect 7586 289 7642 327
rect 7672 361 7836 377
rect 7672 332 7693 361
tri 7672 316 7688 332 ne
rect 7688 327 7693 332
rect 7727 327 7790 361
rect 7824 327 7836 361
rect 7688 316 7836 327
rect 7866 340 8028 377
tri 7866 324 7882 340 ne
rect 7882 324 8028 340
rect 7586 255 7596 289
rect 7630 255 7642 289
tri 7748 286 7778 316 ne
rect 7778 289 7836 316
tri 7942 294 7972 324 ne
rect 7586 221 7642 255
rect 7586 187 7596 221
rect 7630 187 7642 221
rect 7586 155 7642 187
tri 7672 270 7688 286 se
rect 7688 270 7732 286
tri 7732 270 7748 286 sw
rect 7672 236 7748 270
rect 7672 202 7693 236
rect 7727 202 7748 236
rect 7672 201 7748 202
tri 7672 185 7688 201 ne
rect 7688 185 7732 201
tri 7732 185 7748 201 nw
rect 7778 255 7790 289
rect 7824 255 7836 289
rect 7778 221 7836 255
rect 7778 187 7790 221
rect 7824 187 7836 221
tri 7866 278 7882 294 se
rect 7882 278 7926 294
tri 7926 278 7942 294 sw
rect 7866 245 7942 278
rect 7866 211 7887 245
rect 7921 211 7942 245
rect 7866 209 7942 211
tri 7866 193 7882 209 ne
rect 7882 193 7926 209
tri 7926 193 7942 209 nw
rect 7972 289 8028 324
rect 7972 255 7984 289
rect 8018 255 8028 289
rect 7972 221 8028 255
tri 7642 155 7672 185 sw
tri 7748 155 7778 185 se
rect 7778 163 7836 187
tri 7836 163 7866 193 sw
tri 7942 163 7972 193 se
rect 7972 187 7984 221
rect 8018 187 8028 221
rect 7972 163 8028 187
rect 7778 155 8028 163
rect 7586 151 8028 155
rect 7586 117 7596 151
rect 7630 117 7790 151
rect 7824 117 7887 151
rect 7921 117 7984 151
rect 8018 117 8028 151
rect 7586 101 8028 117
rect 8252 361 8308 377
rect 8252 327 8262 361
rect 8296 327 8308 361
rect 8252 289 8308 327
rect 8338 361 8502 377
rect 8338 332 8359 361
tri 8338 316 8354 332 ne
rect 8354 327 8359 332
rect 8393 327 8456 361
rect 8490 327 8502 361
rect 8354 316 8502 327
rect 8532 340 8694 377
tri 8532 324 8548 340 ne
rect 8548 324 8694 340
rect 8252 255 8262 289
rect 8296 255 8308 289
tri 8414 286 8444 316 ne
rect 8444 289 8502 316
tri 8608 294 8638 324 ne
rect 8252 221 8308 255
rect 8252 187 8262 221
rect 8296 187 8308 221
rect 8252 155 8308 187
tri 8338 270 8354 286 se
rect 8354 270 8398 286
tri 8398 270 8414 286 sw
rect 8338 236 8414 270
rect 8338 202 8359 236
rect 8393 202 8414 236
rect 8338 201 8414 202
tri 8338 185 8354 201 ne
rect 8354 185 8398 201
tri 8398 185 8414 201 nw
rect 8444 255 8456 289
rect 8490 255 8502 289
rect 8444 221 8502 255
rect 8444 187 8456 221
rect 8490 187 8502 221
tri 8532 278 8548 294 se
rect 8548 278 8592 294
tri 8592 278 8608 294 sw
rect 8532 245 8608 278
rect 8532 211 8553 245
rect 8587 211 8608 245
rect 8532 209 8608 211
tri 8532 193 8548 209 ne
rect 8548 193 8592 209
tri 8592 193 8608 209 nw
rect 8638 289 8694 324
rect 8638 255 8650 289
rect 8684 255 8694 289
rect 8638 221 8694 255
tri 8308 155 8338 185 sw
tri 8414 155 8444 185 se
rect 8444 163 8502 187
tri 8502 163 8532 193 sw
tri 8608 163 8638 193 se
rect 8638 187 8650 221
rect 8684 187 8694 221
rect 8638 163 8694 187
rect 8444 155 8694 163
rect 8252 151 8694 155
rect 8252 117 8262 151
rect 8296 117 8456 151
rect 8490 117 8553 151
rect 8587 117 8650 151
rect 8684 117 8694 151
rect 8252 101 8694 117
rect 8897 363 8953 379
rect 8897 329 8907 363
rect 8941 329 8953 363
rect 8897 291 8953 329
rect 8983 363 9253 379
rect 8983 334 9004 363
tri 8983 318 8999 334 ne
rect 8999 329 9004 334
rect 9038 329 9101 363
rect 9135 329 9198 363
rect 9232 329 9253 363
rect 8999 318 9253 329
rect 9283 363 9339 379
rect 9283 329 9295 363
rect 9329 329 9339 363
rect 8897 257 8907 291
rect 8941 257 8953 291
tri 9059 288 9089 318 ne
rect 9089 291 9148 318
rect 8897 223 8953 257
rect 8897 189 8907 223
rect 8941 189 8953 223
rect 8897 157 8953 189
tri 8983 272 8999 288 se
rect 8999 272 9043 288
tri 9043 272 9059 288 sw
rect 8983 238 9059 272
rect 8983 204 9004 238
rect 9038 204 9059 238
rect 8983 203 9059 204
tri 8983 187 8999 203 ne
rect 8999 187 9043 203
tri 9043 187 9059 203 nw
rect 9089 257 9101 291
rect 9135 257 9148 291
tri 9148 288 9178 318 nw
rect 9089 223 9148 257
rect 9089 189 9101 223
rect 9135 189 9148 223
tri 9178 272 9194 288 se
rect 9194 272 9237 288
tri 9237 272 9253 288 sw
rect 9178 244 9253 272
rect 9178 210 9199 244
rect 9233 210 9253 244
tri 9178 194 9194 210 ne
rect 9194 194 9237 210
tri 9237 194 9253 210 nw
tri 8953 157 8983 187 sw
tri 9059 157 9089 187 se
rect 9089 164 9148 189
tri 9148 164 9178 194 sw
tri 9253 164 9283 194 se
rect 9283 164 9339 329
rect 9089 157 9339 164
rect 8897 153 9339 157
rect 8897 119 8907 153
rect 8941 119 9101 153
rect 9135 119 9198 153
rect 9232 119 9295 153
rect 9329 119 9339 153
rect 8897 103 9339 119
rect 9399 363 9455 379
rect 9399 329 9409 363
rect 9443 329 9455 363
rect 9399 291 9455 329
rect 9485 342 9647 379
tri 9485 326 9501 342 ne
rect 9501 326 9647 342
tri 9561 296 9591 326 ne
rect 9399 257 9409 291
rect 9443 257 9455 291
rect 9399 223 9455 257
rect 9399 189 9409 223
rect 9443 189 9455 223
tri 9485 280 9501 296 se
rect 9501 280 9545 296
tri 9545 280 9561 296 sw
rect 9485 247 9561 280
rect 9485 213 9506 247
rect 9540 213 9561 247
rect 9485 211 9561 213
tri 9485 195 9501 211 ne
rect 9501 195 9545 211
tri 9545 195 9561 211 nw
rect 9591 291 9647 326
rect 9591 257 9603 291
rect 9637 257 9647 291
rect 9591 223 9647 257
rect 9399 165 9455 189
tri 9455 165 9485 195 sw
tri 9561 165 9591 195 se
rect 9591 189 9603 223
rect 9637 189 9647 223
rect 9591 165 9647 189
rect 9399 153 9647 165
rect 9399 119 9409 153
rect 9443 119 9506 153
rect 9540 119 9603 153
rect 9637 119 9647 153
rect 9399 103 9647 119
rect 9880 361 9936 377
rect 9880 327 9890 361
rect 9924 327 9936 361
rect 9880 289 9936 327
rect 9966 361 10130 377
rect 9966 332 9987 361
tri 9966 316 9982 332 ne
rect 9982 327 9987 332
rect 10021 327 10084 361
rect 10118 327 10130 361
rect 9982 316 10130 327
rect 10160 340 10322 377
tri 10160 324 10176 340 ne
rect 10176 324 10322 340
rect 9880 255 9890 289
rect 9924 255 9936 289
tri 10042 286 10072 316 ne
rect 10072 289 10130 316
tri 10236 294 10266 324 ne
rect 9880 221 9936 255
rect 9880 187 9890 221
rect 9924 187 9936 221
rect 9880 155 9936 187
tri 9966 270 9982 286 se
rect 9982 270 10026 286
tri 10026 270 10042 286 sw
rect 9966 236 10042 270
rect 9966 202 9987 236
rect 10021 202 10042 236
rect 9966 201 10042 202
tri 9966 185 9982 201 ne
rect 9982 185 10026 201
tri 10026 185 10042 201 nw
rect 10072 255 10084 289
rect 10118 255 10130 289
rect 10072 221 10130 255
rect 10072 187 10084 221
rect 10118 187 10130 221
tri 10160 278 10176 294 se
rect 10176 278 10220 294
tri 10220 278 10236 294 sw
rect 10160 245 10236 278
rect 10160 211 10181 245
rect 10215 211 10236 245
rect 10160 209 10236 211
tri 10160 193 10176 209 ne
rect 10176 193 10220 209
tri 10220 193 10236 209 nw
rect 10266 289 10322 324
rect 10266 255 10278 289
rect 10312 255 10322 289
rect 10266 221 10322 255
tri 9936 155 9966 185 sw
tri 10042 155 10072 185 se
rect 10072 163 10130 187
tri 10130 163 10160 193 sw
tri 10236 163 10266 193 se
rect 10266 187 10278 221
rect 10312 187 10322 221
rect 10266 163 10322 187
rect 10072 155 10322 163
rect 9880 151 10322 155
rect 9880 117 9890 151
rect 9924 117 10084 151
rect 10118 117 10181 151
rect 10215 117 10278 151
rect 10312 117 10322 151
rect 9880 101 10322 117
rect 10525 363 10581 379
rect 10525 329 10535 363
rect 10569 329 10581 363
rect 10525 291 10581 329
rect 10611 363 10881 379
rect 10611 334 10632 363
tri 10611 318 10627 334 ne
rect 10627 329 10632 334
rect 10666 329 10729 363
rect 10763 329 10826 363
rect 10860 329 10881 363
rect 10627 318 10881 329
rect 10911 363 10967 379
rect 10911 329 10923 363
rect 10957 329 10967 363
rect 10525 257 10535 291
rect 10569 257 10581 291
tri 10687 288 10717 318 ne
rect 10717 291 10776 318
rect 10525 223 10581 257
rect 10525 189 10535 223
rect 10569 189 10581 223
rect 10525 157 10581 189
tri 10611 272 10627 288 se
rect 10627 272 10671 288
tri 10671 272 10687 288 sw
rect 10611 238 10687 272
rect 10611 204 10632 238
rect 10666 204 10687 238
rect 10611 203 10687 204
tri 10611 187 10627 203 ne
rect 10627 187 10671 203
tri 10671 187 10687 203 nw
rect 10717 257 10729 291
rect 10763 257 10776 291
tri 10776 288 10806 318 nw
rect 10717 223 10776 257
rect 10717 189 10729 223
rect 10763 189 10776 223
tri 10806 272 10822 288 se
rect 10822 272 10865 288
tri 10865 272 10881 288 sw
rect 10806 244 10881 272
rect 10806 210 10827 244
rect 10861 210 10881 244
tri 10806 194 10822 210 ne
rect 10822 194 10865 210
tri 10865 194 10881 210 nw
tri 10581 157 10611 187 sw
tri 10687 157 10717 187 se
rect 10717 164 10776 189
tri 10776 164 10806 194 sw
tri 10881 164 10911 194 se
rect 10911 164 10967 329
rect 10717 157 10967 164
rect 10525 153 10967 157
rect 10525 119 10535 153
rect 10569 119 10729 153
rect 10763 119 10826 153
rect 10860 119 10923 153
rect 10957 119 10967 153
rect 10525 103 10967 119
rect 11027 363 11083 379
rect 11027 329 11037 363
rect 11071 329 11083 363
rect 11027 291 11083 329
rect 11113 342 11275 379
tri 11113 326 11129 342 ne
rect 11129 326 11275 342
tri 11189 296 11219 326 ne
rect 11027 257 11037 291
rect 11071 257 11083 291
rect 11027 223 11083 257
rect 11027 189 11037 223
rect 11071 189 11083 223
tri 11113 280 11129 296 se
rect 11129 280 11173 296
tri 11173 280 11189 296 sw
rect 11113 247 11189 280
rect 11113 213 11134 247
rect 11168 213 11189 247
rect 11113 211 11189 213
tri 11113 195 11129 211 ne
rect 11129 195 11173 211
tri 11173 195 11189 211 nw
rect 11219 291 11275 326
rect 11219 257 11231 291
rect 11265 257 11275 291
rect 11219 223 11275 257
rect 11027 165 11083 189
tri 11083 165 11113 195 sw
tri 11189 165 11219 195 se
rect 11219 189 11231 223
rect 11265 189 11275 223
rect 11219 165 11275 189
rect 11027 153 11275 165
rect 11027 119 11037 153
rect 11071 119 11134 153
rect 11168 119 11231 153
rect 11265 119 11275 153
rect 11027 103 11275 119
rect 11487 363 11543 379
rect 11487 329 11497 363
rect 11531 329 11543 363
rect 11487 291 11543 329
rect 11573 363 11843 379
rect 11573 334 11594 363
tri 11573 318 11589 334 ne
rect 11589 329 11594 334
rect 11628 329 11691 363
rect 11725 329 11788 363
rect 11822 329 11843 363
rect 11589 318 11843 329
rect 11873 363 11929 379
rect 11873 329 11885 363
rect 11919 329 11929 363
rect 11487 257 11497 291
rect 11531 257 11543 291
tri 11649 288 11679 318 ne
rect 11679 291 11738 318
rect 11487 223 11543 257
rect 11487 189 11497 223
rect 11531 189 11543 223
rect 11487 157 11543 189
tri 11573 272 11589 288 se
rect 11589 272 11633 288
tri 11633 272 11649 288 sw
rect 11573 238 11649 272
rect 11573 204 11594 238
rect 11628 204 11649 238
rect 11573 203 11649 204
tri 11573 187 11589 203 ne
rect 11589 187 11633 203
tri 11633 187 11649 203 nw
rect 11679 257 11691 291
rect 11725 257 11738 291
tri 11738 288 11768 318 nw
rect 11679 223 11738 257
rect 11679 189 11691 223
rect 11725 189 11738 223
tri 11768 272 11784 288 se
rect 11784 272 11827 288
tri 11827 272 11843 288 sw
rect 11768 244 11843 272
rect 11768 210 11789 244
rect 11823 210 11843 244
tri 11768 194 11784 210 ne
rect 11784 194 11827 210
tri 11827 194 11843 210 nw
tri 11543 157 11573 187 sw
tri 11649 157 11679 187 se
rect 11679 164 11738 189
tri 11738 164 11768 194 sw
tri 11843 164 11873 194 se
rect 11873 164 11929 329
rect 11679 157 11929 164
rect 11487 153 11929 157
rect 11487 119 11497 153
rect 11531 119 11691 153
rect 11725 119 11788 153
rect 11822 119 11885 153
rect 11919 119 11929 153
rect 11487 103 11929 119
rect 11989 363 12045 379
rect 11989 329 11999 363
rect 12033 329 12045 363
rect 11989 291 12045 329
rect 12075 342 12237 379
tri 12075 326 12091 342 ne
rect 12091 326 12237 342
tri 12151 296 12181 326 ne
rect 11989 257 11999 291
rect 12033 257 12045 291
rect 11989 223 12045 257
rect 11989 189 11999 223
rect 12033 189 12045 223
tri 12075 280 12091 296 se
rect 12091 280 12135 296
tri 12135 280 12151 296 sw
rect 12075 247 12151 280
rect 12075 213 12096 247
rect 12130 213 12151 247
rect 12075 211 12151 213
tri 12075 195 12091 211 ne
rect 12091 195 12135 211
tri 12135 195 12151 211 nw
rect 12181 291 12237 326
rect 12181 257 12193 291
rect 12227 257 12237 291
rect 12181 223 12237 257
rect 11989 165 12045 189
tri 12045 165 12075 195 sw
tri 12151 165 12181 195 se
rect 12181 189 12193 223
rect 12227 189 12237 223
rect 12181 165 12237 189
rect 11989 153 12237 165
rect 11989 119 11999 153
rect 12033 119 12096 153
rect 12130 119 12193 153
rect 12227 119 12237 153
rect 11989 103 12237 119
rect 12470 361 12526 377
rect 12470 327 12480 361
rect 12514 327 12526 361
rect 12470 289 12526 327
rect 12556 361 12720 377
rect 12556 332 12577 361
tri 12556 316 12572 332 ne
rect 12572 327 12577 332
rect 12611 327 12674 361
rect 12708 327 12720 361
rect 12572 316 12720 327
rect 12750 340 12912 377
tri 12750 324 12766 340 ne
rect 12766 324 12912 340
rect 12470 255 12480 289
rect 12514 255 12526 289
tri 12632 286 12662 316 ne
rect 12662 289 12720 316
tri 12826 294 12856 324 ne
rect 12470 221 12526 255
rect 12470 187 12480 221
rect 12514 187 12526 221
rect 12470 155 12526 187
tri 12556 270 12572 286 se
rect 12572 270 12616 286
tri 12616 270 12632 286 sw
rect 12556 236 12632 270
rect 12556 202 12577 236
rect 12611 202 12632 236
rect 12556 201 12632 202
tri 12556 185 12572 201 ne
rect 12572 185 12616 201
tri 12616 185 12632 201 nw
rect 12662 255 12674 289
rect 12708 255 12720 289
rect 12662 221 12720 255
rect 12662 187 12674 221
rect 12708 187 12720 221
tri 12750 278 12766 294 se
rect 12766 278 12810 294
tri 12810 278 12826 294 sw
rect 12750 245 12826 278
rect 12750 211 12771 245
rect 12805 211 12826 245
rect 12750 209 12826 211
tri 12750 193 12766 209 ne
rect 12766 193 12810 209
tri 12810 193 12826 209 nw
rect 12856 289 12912 324
rect 12856 255 12868 289
rect 12902 255 12912 289
rect 12856 221 12912 255
tri 12526 155 12556 185 sw
tri 12632 155 12662 185 se
rect 12662 163 12720 187
tri 12720 163 12750 193 sw
tri 12826 163 12856 193 se
rect 12856 187 12868 221
rect 12902 187 12912 221
rect 12856 163 12912 187
rect 12662 155 12912 163
rect 12470 151 12912 155
rect 12470 117 12480 151
rect 12514 117 12674 151
rect 12708 117 12771 151
rect 12805 117 12868 151
rect 12902 117 12912 151
rect 12470 101 12912 117
rect 13136 361 13192 377
rect 13136 327 13146 361
rect 13180 327 13192 361
rect 13136 289 13192 327
rect 13222 361 13386 377
rect 13222 332 13243 361
tri 13222 316 13238 332 ne
rect 13238 327 13243 332
rect 13277 327 13340 361
rect 13374 327 13386 361
rect 13238 316 13386 327
rect 13416 340 13578 377
tri 13416 324 13432 340 ne
rect 13432 324 13578 340
rect 13136 255 13146 289
rect 13180 255 13192 289
tri 13298 286 13328 316 ne
rect 13328 289 13386 316
tri 13492 294 13522 324 ne
rect 13136 221 13192 255
rect 13136 187 13146 221
rect 13180 187 13192 221
rect 13136 155 13192 187
tri 13222 270 13238 286 se
rect 13238 270 13282 286
tri 13282 270 13298 286 sw
rect 13222 236 13298 270
rect 13222 202 13243 236
rect 13277 202 13298 236
rect 13222 201 13298 202
tri 13222 185 13238 201 ne
rect 13238 185 13282 201
tri 13282 185 13298 201 nw
rect 13328 255 13340 289
rect 13374 255 13386 289
rect 13328 221 13386 255
rect 13328 187 13340 221
rect 13374 187 13386 221
tri 13416 278 13432 294 se
rect 13432 278 13476 294
tri 13476 278 13492 294 sw
rect 13416 245 13492 278
rect 13416 211 13437 245
rect 13471 211 13492 245
rect 13416 209 13492 211
tri 13416 193 13432 209 ne
rect 13432 193 13476 209
tri 13476 193 13492 209 nw
rect 13522 289 13578 324
rect 13522 255 13534 289
rect 13568 255 13578 289
rect 13522 221 13578 255
tri 13192 155 13222 185 sw
tri 13298 155 13328 185 se
rect 13328 163 13386 187
tri 13386 163 13416 193 sw
tri 13492 163 13522 193 se
rect 13522 187 13534 221
rect 13568 187 13578 221
rect 13522 163 13578 187
rect 13328 155 13578 163
rect 13136 151 13578 155
rect 13136 117 13146 151
rect 13180 117 13340 151
rect 13374 117 13437 151
rect 13471 117 13534 151
rect 13568 117 13578 151
rect 13136 101 13578 117
rect 13781 363 13837 379
rect 13781 329 13791 363
rect 13825 329 13837 363
rect 13781 291 13837 329
rect 13867 363 14137 379
rect 13867 334 13888 363
tri 13867 318 13883 334 ne
rect 13883 329 13888 334
rect 13922 329 13985 363
rect 14019 329 14082 363
rect 14116 329 14137 363
rect 13883 318 14137 329
rect 14167 363 14223 379
rect 14167 329 14179 363
rect 14213 329 14223 363
rect 13781 257 13791 291
rect 13825 257 13837 291
tri 13943 288 13973 318 ne
rect 13973 291 14032 318
rect 13781 223 13837 257
rect 13781 189 13791 223
rect 13825 189 13837 223
rect 13781 157 13837 189
tri 13867 272 13883 288 se
rect 13883 272 13927 288
tri 13927 272 13943 288 sw
rect 13867 238 13943 272
rect 13867 204 13888 238
rect 13922 204 13943 238
rect 13867 203 13943 204
tri 13867 187 13883 203 ne
rect 13883 187 13927 203
tri 13927 187 13943 203 nw
rect 13973 257 13985 291
rect 14019 257 14032 291
tri 14032 288 14062 318 nw
rect 13973 223 14032 257
rect 13973 189 13985 223
rect 14019 189 14032 223
tri 14062 272 14078 288 se
rect 14078 272 14121 288
tri 14121 272 14137 288 sw
rect 14062 244 14137 272
rect 14062 210 14083 244
rect 14117 210 14137 244
tri 14062 194 14078 210 ne
rect 14078 194 14121 210
tri 14121 194 14137 210 nw
tri 13837 157 13867 187 sw
tri 13943 157 13973 187 se
rect 13973 164 14032 189
tri 14032 164 14062 194 sw
tri 14137 164 14167 194 se
rect 14167 164 14223 329
rect 13973 157 14223 164
rect 13781 153 14223 157
rect 13781 119 13791 153
rect 13825 119 13985 153
rect 14019 119 14082 153
rect 14116 119 14179 153
rect 14213 119 14223 153
rect 13781 103 14223 119
rect 14283 363 14339 379
rect 14283 329 14293 363
rect 14327 329 14339 363
rect 14283 291 14339 329
rect 14369 342 14531 379
tri 14369 326 14385 342 ne
rect 14385 326 14531 342
tri 14445 296 14475 326 ne
rect 14283 257 14293 291
rect 14327 257 14339 291
rect 14283 223 14339 257
rect 14283 189 14293 223
rect 14327 189 14339 223
tri 14369 280 14385 296 se
rect 14385 280 14429 296
tri 14429 280 14445 296 sw
rect 14369 247 14445 280
rect 14369 213 14390 247
rect 14424 213 14445 247
rect 14369 211 14445 213
tri 14369 195 14385 211 ne
rect 14385 195 14429 211
tri 14429 195 14445 211 nw
rect 14475 291 14531 326
rect 14475 257 14487 291
rect 14521 257 14531 291
rect 14475 223 14531 257
rect 14283 165 14339 189
tri 14339 165 14369 195 sw
tri 14445 165 14475 195 se
rect 14475 189 14487 223
rect 14521 189 14531 223
rect 14475 165 14531 189
rect 14283 153 14531 165
rect 14283 119 14293 153
rect 14327 119 14390 153
rect 14424 119 14487 153
rect 14521 119 14531 153
rect 14283 103 14531 119
rect 14764 361 14820 377
rect 14764 327 14774 361
rect 14808 327 14820 361
rect 14764 289 14820 327
rect 14850 361 15014 377
rect 14850 332 14871 361
tri 14850 316 14866 332 ne
rect 14866 327 14871 332
rect 14905 327 14968 361
rect 15002 327 15014 361
rect 14866 316 15014 327
rect 15044 361 15204 377
rect 15044 340 15162 361
tri 15044 324 15060 340 ne
rect 15060 327 15162 340
rect 15196 327 15204 361
rect 15060 324 15204 327
rect 14764 255 14774 289
rect 14808 255 14820 289
tri 14926 286 14956 316 ne
rect 14956 289 15014 316
tri 15120 294 15150 324 ne
rect 14764 221 14820 255
rect 14764 187 14774 221
rect 14808 187 14820 221
rect 14764 155 14820 187
tri 14850 270 14866 286 se
rect 14866 270 14910 286
tri 14910 270 14926 286 sw
rect 14850 236 14926 270
rect 14850 202 14871 236
rect 14905 202 14926 236
rect 14850 201 14926 202
tri 14850 185 14866 201 ne
rect 14866 185 14910 201
tri 14910 185 14926 201 nw
rect 14956 255 14968 289
rect 15002 255 15014 289
rect 14956 221 15014 255
rect 14956 187 14968 221
rect 15002 187 15014 221
tri 15044 278 15060 294 se
rect 15060 278 15104 294
tri 15104 278 15120 294 sw
rect 15044 245 15120 278
rect 15044 211 15064 245
rect 15098 211 15120 245
rect 15044 209 15120 211
tri 15044 193 15060 209 ne
rect 15060 193 15104 209
tri 15104 193 15120 209 nw
rect 15150 289 15204 324
rect 15150 255 15162 289
rect 15196 255 15204 289
rect 15150 221 15204 255
tri 14820 155 14850 185 sw
tri 14926 155 14956 185 se
rect 14956 163 15014 187
tri 15014 163 15044 193 sw
tri 15120 163 15150 193 se
rect 15150 187 15162 221
rect 15196 187 15204 221
rect 15150 163 15204 187
rect 14956 155 15204 163
rect 14764 151 15204 155
rect 14764 117 14774 151
rect 14808 117 14968 151
rect 15002 117 15064 151
rect 15098 117 15162 151
rect 15196 117 15204 151
rect 14764 101 15204 117
rect 15430 361 15486 377
rect 15430 327 15440 361
rect 15474 327 15486 361
rect 15430 289 15486 327
rect 15516 361 15786 377
rect 15516 332 15537 361
tri 15516 316 15532 332 ne
rect 15532 327 15537 332
rect 15571 327 15634 361
rect 15668 340 15786 361
rect 15668 327 15770 340
rect 15532 324 15770 327
tri 15770 324 15786 340 nw
rect 15816 361 15872 377
rect 15816 327 15828 361
rect 15862 327 15872 361
rect 15532 316 15680 324
rect 15430 255 15440 289
rect 15474 255 15486 289
tri 15592 286 15622 316 ne
rect 15622 289 15680 316
tri 15680 294 15710 324 nw
rect 15430 221 15486 255
rect 15430 187 15440 221
rect 15474 187 15486 221
rect 15430 155 15486 187
tri 15516 270 15532 286 se
rect 15532 270 15576 286
tri 15576 270 15592 286 sw
rect 15516 236 15592 270
rect 15516 202 15537 236
rect 15571 202 15592 236
rect 15516 201 15592 202
tri 15516 185 15532 201 ne
rect 15532 185 15576 201
tri 15576 185 15592 201 nw
rect 15622 255 15634 289
rect 15668 255 15680 289
rect 15622 221 15680 255
rect 15622 187 15634 221
rect 15668 187 15680 221
tri 15710 278 15726 294 se
rect 15726 278 15770 294
tri 15770 278 15786 294 sw
rect 15710 245 15786 278
rect 15710 211 15731 245
rect 15765 211 15786 245
rect 15710 209 15786 211
tri 15710 193 15726 209 ne
rect 15726 193 15770 209
tri 15770 193 15786 209 nw
rect 15816 289 15872 327
rect 15816 255 15828 289
rect 15862 255 15872 289
rect 15816 221 15872 255
tri 15486 155 15516 185 sw
tri 15592 155 15622 185 se
rect 15622 163 15680 187
tri 15680 163 15710 193 sw
tri 15786 163 15816 193 se
rect 15816 187 15828 221
rect 15862 187 15872 221
rect 15816 163 15872 187
rect 15622 155 15872 163
rect 15430 151 15872 155
rect 15430 117 15440 151
rect 15474 117 15634 151
rect 15668 117 15731 151
rect 15765 117 15828 151
rect 15862 117 15872 151
rect 15430 101 15872 117
rect 16096 361 16152 377
rect 16096 327 16106 361
rect 16140 327 16152 361
rect 16096 289 16152 327
rect 16182 361 16346 377
rect 16182 332 16203 361
tri 16182 316 16198 332 ne
rect 16198 327 16203 332
rect 16237 327 16300 361
rect 16334 327 16346 361
rect 16198 316 16346 327
rect 16376 340 16538 377
tri 16376 324 16392 340 ne
rect 16392 324 16538 340
rect 16096 255 16106 289
rect 16140 255 16152 289
tri 16258 286 16288 316 ne
rect 16288 289 16346 316
tri 16452 294 16482 324 ne
rect 16096 221 16152 255
rect 16096 187 16106 221
rect 16140 187 16152 221
rect 16096 155 16152 187
tri 16182 270 16198 286 se
rect 16198 270 16242 286
tri 16242 270 16258 286 sw
rect 16182 236 16258 270
rect 16182 202 16203 236
rect 16237 202 16258 236
rect 16182 201 16258 202
tri 16182 185 16198 201 ne
rect 16198 185 16242 201
tri 16242 185 16258 201 nw
rect 16288 255 16300 289
rect 16334 255 16346 289
tri 16377 279 16392 294 se
rect 16392 279 16436 294
tri 16436 279 16451 294 sw
rect 16482 289 16538 324
rect 16288 221 16346 255
rect 16288 187 16300 221
rect 16334 187 16346 221
rect 16376 245 16452 279
rect 16376 211 16397 245
rect 16431 211 16452 245
rect 16376 209 16452 211
tri 16376 193 16392 209 ne
rect 16392 193 16436 209
tri 16436 193 16452 209 nw
rect 16482 255 16494 289
rect 16528 255 16538 289
rect 16482 221 16538 255
tri 16152 155 16182 185 sw
tri 16258 155 16288 185 se
rect 16288 163 16346 187
tri 16346 163 16376 193 sw
tri 16452 163 16482 193 se
rect 16482 187 16494 221
rect 16528 187 16538 221
rect 16482 163 16538 187
rect 16288 155 16538 163
rect 16096 151 16538 155
rect 16096 117 16106 151
rect 16140 117 16300 151
rect 16334 117 16397 151
rect 16431 117 16494 151
rect 16528 117 16538 151
rect 16096 101 16538 117
<< pdiff >>
rect 131 1412 187 1450
rect 131 1378 141 1412
rect 175 1378 187 1412
rect 131 1344 187 1378
rect 131 1310 141 1344
rect 175 1310 187 1344
rect 131 1276 187 1310
rect 131 1242 141 1276
rect 175 1242 187 1276
rect 131 1208 187 1242
rect 131 1174 141 1208
rect 175 1174 187 1208
rect 131 1139 187 1174
rect 131 1105 141 1139
rect 175 1105 187 1139
rect 131 1050 187 1105
rect 217 1412 275 1450
rect 217 1378 229 1412
rect 263 1378 275 1412
rect 217 1344 275 1378
rect 217 1310 229 1344
rect 263 1310 275 1344
rect 217 1276 275 1310
rect 217 1242 229 1276
rect 263 1242 275 1276
rect 217 1208 275 1242
rect 217 1174 229 1208
rect 263 1174 275 1208
rect 217 1139 275 1174
rect 217 1105 229 1139
rect 263 1105 275 1139
rect 217 1050 275 1105
rect 305 1412 363 1450
rect 305 1378 317 1412
rect 351 1378 363 1412
rect 305 1344 363 1378
rect 305 1310 317 1344
rect 351 1310 363 1344
rect 305 1276 363 1310
rect 305 1242 317 1276
rect 351 1242 363 1276
rect 305 1208 363 1242
rect 305 1174 317 1208
rect 351 1174 363 1208
rect 305 1050 363 1174
rect 393 1412 451 1450
rect 393 1378 405 1412
rect 439 1378 451 1412
rect 393 1344 451 1378
rect 393 1310 405 1344
rect 439 1310 451 1344
rect 393 1276 451 1310
rect 393 1242 405 1276
rect 439 1242 451 1276
rect 393 1208 451 1242
rect 393 1174 405 1208
rect 439 1174 451 1208
rect 393 1139 451 1174
rect 393 1105 405 1139
rect 439 1105 451 1139
rect 393 1050 451 1105
rect 481 1412 535 1450
rect 481 1378 493 1412
rect 527 1378 535 1412
rect 481 1344 535 1378
rect 481 1310 493 1344
rect 527 1310 535 1344
rect 481 1276 535 1310
rect 481 1242 493 1276
rect 527 1242 535 1276
rect 481 1208 535 1242
rect 481 1174 493 1208
rect 527 1174 535 1208
rect 481 1050 535 1174
rect 857 1412 913 1450
rect 857 1378 867 1412
rect 901 1378 913 1412
rect 857 1344 913 1378
rect 857 1310 867 1344
rect 901 1310 913 1344
rect 857 1276 913 1310
rect 857 1242 867 1276
rect 901 1242 913 1276
rect 857 1208 913 1242
rect 857 1174 867 1208
rect 901 1174 913 1208
rect 857 1139 913 1174
rect 857 1105 867 1139
rect 901 1105 913 1139
rect 857 1050 913 1105
rect 943 1412 1001 1450
rect 943 1378 955 1412
rect 989 1378 1001 1412
rect 943 1344 1001 1378
rect 943 1310 955 1344
rect 989 1310 1001 1344
rect 943 1276 1001 1310
rect 943 1242 955 1276
rect 989 1242 1001 1276
rect 943 1208 1001 1242
rect 943 1174 955 1208
rect 989 1174 1001 1208
rect 943 1139 1001 1174
rect 943 1105 955 1139
rect 989 1105 1001 1139
rect 943 1050 1001 1105
rect 1031 1412 1089 1450
rect 1031 1378 1043 1412
rect 1077 1378 1089 1412
rect 1031 1344 1089 1378
rect 1031 1310 1043 1344
rect 1077 1310 1089 1344
rect 1031 1276 1089 1310
rect 1031 1242 1043 1276
rect 1077 1242 1089 1276
rect 1031 1208 1089 1242
rect 1031 1174 1043 1208
rect 1077 1174 1089 1208
rect 1031 1050 1089 1174
rect 1119 1412 1177 1450
rect 1119 1378 1131 1412
rect 1165 1378 1177 1412
rect 1119 1344 1177 1378
rect 1119 1310 1131 1344
rect 1165 1310 1177 1344
rect 1119 1276 1177 1310
rect 1119 1242 1131 1276
rect 1165 1242 1177 1276
rect 1119 1208 1177 1242
rect 1119 1174 1131 1208
rect 1165 1174 1177 1208
rect 1119 1139 1177 1174
rect 1119 1105 1131 1139
rect 1165 1105 1177 1139
rect 1119 1050 1177 1105
rect 1207 1412 1265 1450
rect 1207 1378 1219 1412
rect 1253 1378 1265 1412
rect 1207 1344 1265 1378
rect 1207 1310 1219 1344
rect 1253 1310 1265 1344
rect 1207 1276 1265 1310
rect 1207 1242 1219 1276
rect 1253 1242 1265 1276
rect 1207 1208 1265 1242
rect 1207 1174 1219 1208
rect 1253 1174 1265 1208
rect 1207 1050 1265 1174
rect 1295 1412 1353 1450
rect 1295 1378 1307 1412
rect 1341 1378 1353 1412
rect 1295 1344 1353 1378
rect 1295 1310 1307 1344
rect 1341 1310 1353 1344
rect 1295 1276 1353 1310
rect 1295 1242 1307 1276
rect 1341 1242 1353 1276
rect 1295 1208 1353 1242
rect 1295 1174 1307 1208
rect 1341 1174 1353 1208
rect 1295 1139 1353 1174
rect 1295 1105 1307 1139
rect 1341 1105 1353 1139
rect 1295 1050 1353 1105
rect 1383 1412 1437 1450
rect 1383 1378 1395 1412
rect 1429 1378 1437 1412
rect 1383 1344 1437 1378
rect 1383 1310 1395 1344
rect 1429 1310 1437 1344
rect 1383 1276 1437 1310
rect 1383 1242 1395 1276
rect 1429 1242 1437 1276
rect 1383 1208 1437 1242
rect 1383 1174 1395 1208
rect 1429 1174 1437 1208
rect 1383 1050 1437 1174
rect 1819 1412 1875 1450
rect 1819 1378 1829 1412
rect 1863 1378 1875 1412
rect 1819 1344 1875 1378
rect 1819 1310 1829 1344
rect 1863 1310 1875 1344
rect 1819 1276 1875 1310
rect 1819 1242 1829 1276
rect 1863 1242 1875 1276
rect 1819 1208 1875 1242
rect 1819 1174 1829 1208
rect 1863 1174 1875 1208
rect 1819 1139 1875 1174
rect 1819 1105 1829 1139
rect 1863 1105 1875 1139
rect 1819 1050 1875 1105
rect 1905 1412 1963 1450
rect 1905 1378 1917 1412
rect 1951 1378 1963 1412
rect 1905 1344 1963 1378
rect 1905 1310 1917 1344
rect 1951 1310 1963 1344
rect 1905 1276 1963 1310
rect 1905 1242 1917 1276
rect 1951 1242 1963 1276
rect 1905 1208 1963 1242
rect 1905 1174 1917 1208
rect 1951 1174 1963 1208
rect 1905 1139 1963 1174
rect 1905 1105 1917 1139
rect 1951 1105 1963 1139
rect 1905 1050 1963 1105
rect 1993 1412 2051 1450
rect 1993 1378 2005 1412
rect 2039 1378 2051 1412
rect 1993 1344 2051 1378
rect 1993 1310 2005 1344
rect 2039 1310 2051 1344
rect 1993 1276 2051 1310
rect 1993 1242 2005 1276
rect 2039 1242 2051 1276
rect 1993 1208 2051 1242
rect 1993 1174 2005 1208
rect 2039 1174 2051 1208
rect 1993 1050 2051 1174
rect 2081 1412 2139 1450
rect 2081 1378 2093 1412
rect 2127 1378 2139 1412
rect 2081 1344 2139 1378
rect 2081 1310 2093 1344
rect 2127 1310 2139 1344
rect 2081 1276 2139 1310
rect 2081 1242 2093 1276
rect 2127 1242 2139 1276
rect 2081 1208 2139 1242
rect 2081 1174 2093 1208
rect 2127 1174 2139 1208
rect 2081 1139 2139 1174
rect 2081 1105 2093 1139
rect 2127 1105 2139 1139
rect 2081 1050 2139 1105
rect 2169 1412 2227 1450
rect 2169 1378 2181 1412
rect 2215 1378 2227 1412
rect 2169 1344 2227 1378
rect 2169 1310 2181 1344
rect 2215 1310 2227 1344
rect 2169 1276 2227 1310
rect 2169 1242 2181 1276
rect 2215 1242 2227 1276
rect 2169 1208 2227 1242
rect 2169 1174 2181 1208
rect 2215 1174 2227 1208
rect 2169 1050 2227 1174
rect 2257 1412 2315 1450
rect 2257 1378 2269 1412
rect 2303 1378 2315 1412
rect 2257 1344 2315 1378
rect 2257 1310 2269 1344
rect 2303 1310 2315 1344
rect 2257 1276 2315 1310
rect 2257 1242 2269 1276
rect 2303 1242 2315 1276
rect 2257 1208 2315 1242
rect 2257 1174 2269 1208
rect 2303 1174 2315 1208
rect 2257 1139 2315 1174
rect 2257 1105 2269 1139
rect 2303 1105 2315 1139
rect 2257 1050 2315 1105
rect 2345 1412 2399 1450
rect 2345 1378 2357 1412
rect 2391 1378 2399 1412
rect 2345 1344 2399 1378
rect 2345 1310 2357 1344
rect 2391 1310 2399 1344
rect 2345 1276 2399 1310
rect 2345 1242 2357 1276
rect 2391 1242 2399 1276
rect 2345 1208 2399 1242
rect 2345 1174 2357 1208
rect 2391 1174 2399 1208
rect 2345 1050 2399 1174
rect 2721 1412 2777 1450
rect 2721 1378 2731 1412
rect 2765 1378 2777 1412
rect 2721 1344 2777 1378
rect 2721 1310 2731 1344
rect 2765 1310 2777 1344
rect 2721 1276 2777 1310
rect 2721 1242 2731 1276
rect 2765 1242 2777 1276
rect 2721 1208 2777 1242
rect 2721 1174 2731 1208
rect 2765 1174 2777 1208
rect 2721 1139 2777 1174
rect 2721 1105 2731 1139
rect 2765 1105 2777 1139
rect 2721 1050 2777 1105
rect 2807 1412 2865 1450
rect 2807 1378 2819 1412
rect 2853 1378 2865 1412
rect 2807 1344 2865 1378
rect 2807 1310 2819 1344
rect 2853 1310 2865 1344
rect 2807 1276 2865 1310
rect 2807 1242 2819 1276
rect 2853 1242 2865 1276
rect 2807 1208 2865 1242
rect 2807 1174 2819 1208
rect 2853 1174 2865 1208
rect 2807 1139 2865 1174
rect 2807 1105 2819 1139
rect 2853 1105 2865 1139
rect 2807 1050 2865 1105
rect 2895 1412 2953 1450
rect 2895 1378 2907 1412
rect 2941 1378 2953 1412
rect 2895 1344 2953 1378
rect 2895 1310 2907 1344
rect 2941 1310 2953 1344
rect 2895 1276 2953 1310
rect 2895 1242 2907 1276
rect 2941 1242 2953 1276
rect 2895 1208 2953 1242
rect 2895 1174 2907 1208
rect 2941 1174 2953 1208
rect 2895 1050 2953 1174
rect 2983 1412 3041 1450
rect 2983 1378 2995 1412
rect 3029 1378 3041 1412
rect 2983 1344 3041 1378
rect 2983 1310 2995 1344
rect 3029 1310 3041 1344
rect 2983 1276 3041 1310
rect 2983 1242 2995 1276
rect 3029 1242 3041 1276
rect 2983 1208 3041 1242
rect 2983 1174 2995 1208
rect 3029 1174 3041 1208
rect 2983 1139 3041 1174
rect 2983 1105 2995 1139
rect 3029 1105 3041 1139
rect 2983 1050 3041 1105
rect 3071 1412 3125 1450
rect 3071 1378 3083 1412
rect 3117 1378 3125 1412
rect 3071 1344 3125 1378
rect 3071 1310 3083 1344
rect 3117 1310 3125 1344
rect 3071 1276 3125 1310
rect 3071 1242 3083 1276
rect 3117 1242 3125 1276
rect 3071 1208 3125 1242
rect 3071 1174 3083 1208
rect 3117 1174 3125 1208
rect 3071 1050 3125 1174
rect 3387 1412 3443 1450
rect 3387 1378 3397 1412
rect 3431 1378 3443 1412
rect 3387 1344 3443 1378
rect 3387 1310 3397 1344
rect 3431 1310 3443 1344
rect 3387 1276 3443 1310
rect 3387 1242 3397 1276
rect 3431 1242 3443 1276
rect 3387 1208 3443 1242
rect 3387 1174 3397 1208
rect 3431 1174 3443 1208
rect 3387 1139 3443 1174
rect 3387 1105 3397 1139
rect 3431 1105 3443 1139
rect 3387 1050 3443 1105
rect 3473 1412 3531 1450
rect 3473 1378 3485 1412
rect 3519 1378 3531 1412
rect 3473 1344 3531 1378
rect 3473 1310 3485 1344
rect 3519 1310 3531 1344
rect 3473 1276 3531 1310
rect 3473 1242 3485 1276
rect 3519 1242 3531 1276
rect 3473 1208 3531 1242
rect 3473 1174 3485 1208
rect 3519 1174 3531 1208
rect 3473 1139 3531 1174
rect 3473 1105 3485 1139
rect 3519 1105 3531 1139
rect 3473 1050 3531 1105
rect 3561 1412 3619 1450
rect 3561 1378 3573 1412
rect 3607 1378 3619 1412
rect 3561 1344 3619 1378
rect 3561 1310 3573 1344
rect 3607 1310 3619 1344
rect 3561 1276 3619 1310
rect 3561 1242 3573 1276
rect 3607 1242 3619 1276
rect 3561 1208 3619 1242
rect 3561 1174 3573 1208
rect 3607 1174 3619 1208
rect 3561 1050 3619 1174
rect 3649 1412 3707 1450
rect 3649 1378 3661 1412
rect 3695 1378 3707 1412
rect 3649 1344 3707 1378
rect 3649 1310 3661 1344
rect 3695 1310 3707 1344
rect 3649 1276 3707 1310
rect 3649 1242 3661 1276
rect 3695 1242 3707 1276
rect 3649 1208 3707 1242
rect 3649 1174 3661 1208
rect 3695 1174 3707 1208
rect 3649 1139 3707 1174
rect 3649 1105 3661 1139
rect 3695 1105 3707 1139
rect 3649 1050 3707 1105
rect 3737 1412 3791 1450
rect 3737 1378 3749 1412
rect 3783 1378 3791 1412
rect 3737 1344 3791 1378
rect 3737 1310 3749 1344
rect 3783 1310 3791 1344
rect 3737 1276 3791 1310
rect 3737 1242 3749 1276
rect 3783 1242 3791 1276
rect 3737 1208 3791 1242
rect 3737 1174 3749 1208
rect 3783 1174 3791 1208
rect 3737 1050 3791 1174
rect 4113 1412 4169 1450
rect 4113 1378 4123 1412
rect 4157 1378 4169 1412
rect 4113 1344 4169 1378
rect 4113 1310 4123 1344
rect 4157 1310 4169 1344
rect 4113 1276 4169 1310
rect 4113 1242 4123 1276
rect 4157 1242 4169 1276
rect 4113 1208 4169 1242
rect 4113 1174 4123 1208
rect 4157 1174 4169 1208
rect 4113 1139 4169 1174
rect 4113 1105 4123 1139
rect 4157 1105 4169 1139
rect 4113 1050 4169 1105
rect 4199 1412 4257 1450
rect 4199 1378 4211 1412
rect 4245 1378 4257 1412
rect 4199 1344 4257 1378
rect 4199 1310 4211 1344
rect 4245 1310 4257 1344
rect 4199 1276 4257 1310
rect 4199 1242 4211 1276
rect 4245 1242 4257 1276
rect 4199 1208 4257 1242
rect 4199 1174 4211 1208
rect 4245 1174 4257 1208
rect 4199 1139 4257 1174
rect 4199 1105 4211 1139
rect 4245 1105 4257 1139
rect 4199 1050 4257 1105
rect 4287 1412 4345 1450
rect 4287 1378 4299 1412
rect 4333 1378 4345 1412
rect 4287 1344 4345 1378
rect 4287 1310 4299 1344
rect 4333 1310 4345 1344
rect 4287 1276 4345 1310
rect 4287 1242 4299 1276
rect 4333 1242 4345 1276
rect 4287 1208 4345 1242
rect 4287 1174 4299 1208
rect 4333 1174 4345 1208
rect 4287 1050 4345 1174
rect 4375 1412 4433 1450
rect 4375 1378 4387 1412
rect 4421 1378 4433 1412
rect 4375 1344 4433 1378
rect 4375 1310 4387 1344
rect 4421 1310 4433 1344
rect 4375 1276 4433 1310
rect 4375 1242 4387 1276
rect 4421 1242 4433 1276
rect 4375 1208 4433 1242
rect 4375 1174 4387 1208
rect 4421 1174 4433 1208
rect 4375 1139 4433 1174
rect 4375 1105 4387 1139
rect 4421 1105 4433 1139
rect 4375 1050 4433 1105
rect 4463 1412 4521 1450
rect 4463 1378 4475 1412
rect 4509 1378 4521 1412
rect 4463 1344 4521 1378
rect 4463 1310 4475 1344
rect 4509 1310 4521 1344
rect 4463 1276 4521 1310
rect 4463 1242 4475 1276
rect 4509 1242 4521 1276
rect 4463 1208 4521 1242
rect 4463 1174 4475 1208
rect 4509 1174 4521 1208
rect 4463 1050 4521 1174
rect 4551 1412 4609 1450
rect 4551 1378 4563 1412
rect 4597 1378 4609 1412
rect 4551 1344 4609 1378
rect 4551 1310 4563 1344
rect 4597 1310 4609 1344
rect 4551 1276 4609 1310
rect 4551 1242 4563 1276
rect 4597 1242 4609 1276
rect 4551 1208 4609 1242
rect 4551 1174 4563 1208
rect 4597 1174 4609 1208
rect 4551 1139 4609 1174
rect 4551 1105 4563 1139
rect 4597 1105 4609 1139
rect 4551 1050 4609 1105
rect 4639 1412 4693 1450
rect 4639 1378 4651 1412
rect 4685 1378 4693 1412
rect 4639 1344 4693 1378
rect 4639 1310 4651 1344
rect 4685 1310 4693 1344
rect 4639 1276 4693 1310
rect 4639 1242 4651 1276
rect 4685 1242 4693 1276
rect 4639 1208 4693 1242
rect 4639 1174 4651 1208
rect 4685 1174 4693 1208
rect 4639 1050 4693 1174
rect 5015 1412 5071 1450
rect 5015 1378 5025 1412
rect 5059 1378 5071 1412
rect 5015 1344 5071 1378
rect 5015 1310 5025 1344
rect 5059 1310 5071 1344
rect 5015 1276 5071 1310
rect 5015 1242 5025 1276
rect 5059 1242 5071 1276
rect 5015 1208 5071 1242
rect 5015 1174 5025 1208
rect 5059 1174 5071 1208
rect 5015 1139 5071 1174
rect 5015 1105 5025 1139
rect 5059 1105 5071 1139
rect 5015 1050 5071 1105
rect 5101 1412 5159 1450
rect 5101 1378 5113 1412
rect 5147 1378 5159 1412
rect 5101 1344 5159 1378
rect 5101 1310 5113 1344
rect 5147 1310 5159 1344
rect 5101 1276 5159 1310
rect 5101 1242 5113 1276
rect 5147 1242 5159 1276
rect 5101 1208 5159 1242
rect 5101 1174 5113 1208
rect 5147 1174 5159 1208
rect 5101 1139 5159 1174
rect 5101 1105 5113 1139
rect 5147 1105 5159 1139
rect 5101 1050 5159 1105
rect 5189 1412 5247 1450
rect 5189 1378 5201 1412
rect 5235 1378 5247 1412
rect 5189 1344 5247 1378
rect 5189 1310 5201 1344
rect 5235 1310 5247 1344
rect 5189 1276 5247 1310
rect 5189 1242 5201 1276
rect 5235 1242 5247 1276
rect 5189 1208 5247 1242
rect 5189 1174 5201 1208
rect 5235 1174 5247 1208
rect 5189 1050 5247 1174
rect 5277 1412 5335 1450
rect 5277 1378 5289 1412
rect 5323 1378 5335 1412
rect 5277 1344 5335 1378
rect 5277 1310 5289 1344
rect 5323 1310 5335 1344
rect 5277 1276 5335 1310
rect 5277 1242 5289 1276
rect 5323 1242 5335 1276
rect 5277 1208 5335 1242
rect 5277 1174 5289 1208
rect 5323 1174 5335 1208
rect 5277 1139 5335 1174
rect 5277 1105 5289 1139
rect 5323 1105 5335 1139
rect 5277 1050 5335 1105
rect 5365 1412 5419 1450
rect 5365 1378 5377 1412
rect 5411 1378 5419 1412
rect 5365 1344 5419 1378
rect 5365 1310 5377 1344
rect 5411 1310 5419 1344
rect 5365 1276 5419 1310
rect 5365 1242 5377 1276
rect 5411 1242 5419 1276
rect 5365 1208 5419 1242
rect 5365 1174 5377 1208
rect 5411 1174 5419 1208
rect 5365 1050 5419 1174
rect 5741 1412 5797 1450
rect 5741 1378 5751 1412
rect 5785 1378 5797 1412
rect 5741 1344 5797 1378
rect 5741 1310 5751 1344
rect 5785 1310 5797 1344
rect 5741 1276 5797 1310
rect 5741 1242 5751 1276
rect 5785 1242 5797 1276
rect 5741 1208 5797 1242
rect 5741 1174 5751 1208
rect 5785 1174 5797 1208
rect 5741 1139 5797 1174
rect 5741 1105 5751 1139
rect 5785 1105 5797 1139
rect 5741 1050 5797 1105
rect 5827 1412 5885 1450
rect 5827 1378 5839 1412
rect 5873 1378 5885 1412
rect 5827 1344 5885 1378
rect 5827 1310 5839 1344
rect 5873 1310 5885 1344
rect 5827 1276 5885 1310
rect 5827 1242 5839 1276
rect 5873 1242 5885 1276
rect 5827 1208 5885 1242
rect 5827 1174 5839 1208
rect 5873 1174 5885 1208
rect 5827 1139 5885 1174
rect 5827 1105 5839 1139
rect 5873 1105 5885 1139
rect 5827 1050 5885 1105
rect 5915 1412 5973 1450
rect 5915 1378 5927 1412
rect 5961 1378 5973 1412
rect 5915 1344 5973 1378
rect 5915 1310 5927 1344
rect 5961 1310 5973 1344
rect 5915 1276 5973 1310
rect 5915 1242 5927 1276
rect 5961 1242 5973 1276
rect 5915 1208 5973 1242
rect 5915 1174 5927 1208
rect 5961 1174 5973 1208
rect 5915 1050 5973 1174
rect 6003 1412 6061 1450
rect 6003 1378 6015 1412
rect 6049 1378 6061 1412
rect 6003 1344 6061 1378
rect 6003 1310 6015 1344
rect 6049 1310 6061 1344
rect 6003 1276 6061 1310
rect 6003 1242 6015 1276
rect 6049 1242 6061 1276
rect 6003 1208 6061 1242
rect 6003 1174 6015 1208
rect 6049 1174 6061 1208
rect 6003 1139 6061 1174
rect 6003 1105 6015 1139
rect 6049 1105 6061 1139
rect 6003 1050 6061 1105
rect 6091 1412 6149 1450
rect 6091 1378 6103 1412
rect 6137 1378 6149 1412
rect 6091 1344 6149 1378
rect 6091 1310 6103 1344
rect 6137 1310 6149 1344
rect 6091 1276 6149 1310
rect 6091 1242 6103 1276
rect 6137 1242 6149 1276
rect 6091 1208 6149 1242
rect 6091 1174 6103 1208
rect 6137 1174 6149 1208
rect 6091 1050 6149 1174
rect 6179 1412 6237 1450
rect 6179 1378 6191 1412
rect 6225 1378 6237 1412
rect 6179 1344 6237 1378
rect 6179 1310 6191 1344
rect 6225 1310 6237 1344
rect 6179 1276 6237 1310
rect 6179 1242 6191 1276
rect 6225 1242 6237 1276
rect 6179 1208 6237 1242
rect 6179 1174 6191 1208
rect 6225 1174 6237 1208
rect 6179 1139 6237 1174
rect 6179 1105 6191 1139
rect 6225 1105 6237 1139
rect 6179 1050 6237 1105
rect 6267 1412 6321 1450
rect 6267 1378 6279 1412
rect 6313 1378 6321 1412
rect 6267 1344 6321 1378
rect 6267 1310 6279 1344
rect 6313 1310 6321 1344
rect 6267 1276 6321 1310
rect 6267 1242 6279 1276
rect 6313 1242 6321 1276
rect 6267 1208 6321 1242
rect 6267 1174 6279 1208
rect 6313 1174 6321 1208
rect 6267 1050 6321 1174
rect 6703 1412 6759 1450
rect 6703 1378 6713 1412
rect 6747 1378 6759 1412
rect 6703 1344 6759 1378
rect 6703 1310 6713 1344
rect 6747 1310 6759 1344
rect 6703 1276 6759 1310
rect 6703 1242 6713 1276
rect 6747 1242 6759 1276
rect 6703 1208 6759 1242
rect 6703 1174 6713 1208
rect 6747 1174 6759 1208
rect 6703 1139 6759 1174
rect 6703 1105 6713 1139
rect 6747 1105 6759 1139
rect 6703 1050 6759 1105
rect 6789 1412 6847 1450
rect 6789 1378 6801 1412
rect 6835 1378 6847 1412
rect 6789 1344 6847 1378
rect 6789 1310 6801 1344
rect 6835 1310 6847 1344
rect 6789 1276 6847 1310
rect 6789 1242 6801 1276
rect 6835 1242 6847 1276
rect 6789 1208 6847 1242
rect 6789 1174 6801 1208
rect 6835 1174 6847 1208
rect 6789 1139 6847 1174
rect 6789 1105 6801 1139
rect 6835 1105 6847 1139
rect 6789 1050 6847 1105
rect 6877 1412 6935 1450
rect 6877 1378 6889 1412
rect 6923 1378 6935 1412
rect 6877 1344 6935 1378
rect 6877 1310 6889 1344
rect 6923 1310 6935 1344
rect 6877 1276 6935 1310
rect 6877 1242 6889 1276
rect 6923 1242 6935 1276
rect 6877 1208 6935 1242
rect 6877 1174 6889 1208
rect 6923 1174 6935 1208
rect 6877 1050 6935 1174
rect 6965 1412 7023 1450
rect 6965 1378 6977 1412
rect 7011 1378 7023 1412
rect 6965 1344 7023 1378
rect 6965 1310 6977 1344
rect 7011 1310 7023 1344
rect 6965 1276 7023 1310
rect 6965 1242 6977 1276
rect 7011 1242 7023 1276
rect 6965 1208 7023 1242
rect 6965 1174 6977 1208
rect 7011 1174 7023 1208
rect 6965 1139 7023 1174
rect 6965 1105 6977 1139
rect 7011 1105 7023 1139
rect 6965 1050 7023 1105
rect 7053 1412 7111 1450
rect 7053 1378 7065 1412
rect 7099 1378 7111 1412
rect 7053 1344 7111 1378
rect 7053 1310 7065 1344
rect 7099 1310 7111 1344
rect 7053 1276 7111 1310
rect 7053 1242 7065 1276
rect 7099 1242 7111 1276
rect 7053 1208 7111 1242
rect 7053 1174 7065 1208
rect 7099 1174 7111 1208
rect 7053 1050 7111 1174
rect 7141 1412 7199 1450
rect 7141 1378 7153 1412
rect 7187 1378 7199 1412
rect 7141 1344 7199 1378
rect 7141 1310 7153 1344
rect 7187 1310 7199 1344
rect 7141 1276 7199 1310
rect 7141 1242 7153 1276
rect 7187 1242 7199 1276
rect 7141 1208 7199 1242
rect 7141 1174 7153 1208
rect 7187 1174 7199 1208
rect 7141 1139 7199 1174
rect 7141 1105 7153 1139
rect 7187 1105 7199 1139
rect 7141 1050 7199 1105
rect 7229 1412 7283 1450
rect 7229 1378 7241 1412
rect 7275 1378 7283 1412
rect 7229 1344 7283 1378
rect 7229 1310 7241 1344
rect 7275 1310 7283 1344
rect 7229 1276 7283 1310
rect 7229 1242 7241 1276
rect 7275 1242 7283 1276
rect 7229 1208 7283 1242
rect 7229 1174 7241 1208
rect 7275 1174 7283 1208
rect 7229 1050 7283 1174
rect 7605 1412 7661 1450
rect 7605 1378 7615 1412
rect 7649 1378 7661 1412
rect 7605 1344 7661 1378
rect 7605 1310 7615 1344
rect 7649 1310 7661 1344
rect 7605 1276 7661 1310
rect 7605 1242 7615 1276
rect 7649 1242 7661 1276
rect 7605 1208 7661 1242
rect 7605 1174 7615 1208
rect 7649 1174 7661 1208
rect 7605 1139 7661 1174
rect 7605 1105 7615 1139
rect 7649 1105 7661 1139
rect 7605 1050 7661 1105
rect 7691 1412 7749 1450
rect 7691 1378 7703 1412
rect 7737 1378 7749 1412
rect 7691 1344 7749 1378
rect 7691 1310 7703 1344
rect 7737 1310 7749 1344
rect 7691 1276 7749 1310
rect 7691 1242 7703 1276
rect 7737 1242 7749 1276
rect 7691 1208 7749 1242
rect 7691 1174 7703 1208
rect 7737 1174 7749 1208
rect 7691 1139 7749 1174
rect 7691 1105 7703 1139
rect 7737 1105 7749 1139
rect 7691 1050 7749 1105
rect 7779 1412 7837 1450
rect 7779 1378 7791 1412
rect 7825 1378 7837 1412
rect 7779 1344 7837 1378
rect 7779 1310 7791 1344
rect 7825 1310 7837 1344
rect 7779 1276 7837 1310
rect 7779 1242 7791 1276
rect 7825 1242 7837 1276
rect 7779 1208 7837 1242
rect 7779 1174 7791 1208
rect 7825 1174 7837 1208
rect 7779 1050 7837 1174
rect 7867 1412 7925 1450
rect 7867 1378 7879 1412
rect 7913 1378 7925 1412
rect 7867 1344 7925 1378
rect 7867 1310 7879 1344
rect 7913 1310 7925 1344
rect 7867 1276 7925 1310
rect 7867 1242 7879 1276
rect 7913 1242 7925 1276
rect 7867 1208 7925 1242
rect 7867 1174 7879 1208
rect 7913 1174 7925 1208
rect 7867 1139 7925 1174
rect 7867 1105 7879 1139
rect 7913 1105 7925 1139
rect 7867 1050 7925 1105
rect 7955 1412 8009 1450
rect 7955 1378 7967 1412
rect 8001 1378 8009 1412
rect 7955 1344 8009 1378
rect 7955 1310 7967 1344
rect 8001 1310 8009 1344
rect 7955 1276 8009 1310
rect 7955 1242 7967 1276
rect 8001 1242 8009 1276
rect 7955 1208 8009 1242
rect 7955 1174 7967 1208
rect 8001 1174 8009 1208
rect 7955 1050 8009 1174
rect 8271 1412 8327 1450
rect 8271 1378 8281 1412
rect 8315 1378 8327 1412
rect 8271 1344 8327 1378
rect 8271 1310 8281 1344
rect 8315 1310 8327 1344
rect 8271 1276 8327 1310
rect 8271 1242 8281 1276
rect 8315 1242 8327 1276
rect 8271 1208 8327 1242
rect 8271 1174 8281 1208
rect 8315 1174 8327 1208
rect 8271 1139 8327 1174
rect 8271 1105 8281 1139
rect 8315 1105 8327 1139
rect 8271 1050 8327 1105
rect 8357 1412 8415 1450
rect 8357 1378 8369 1412
rect 8403 1378 8415 1412
rect 8357 1344 8415 1378
rect 8357 1310 8369 1344
rect 8403 1310 8415 1344
rect 8357 1276 8415 1310
rect 8357 1242 8369 1276
rect 8403 1242 8415 1276
rect 8357 1208 8415 1242
rect 8357 1174 8369 1208
rect 8403 1174 8415 1208
rect 8357 1139 8415 1174
rect 8357 1105 8369 1139
rect 8403 1105 8415 1139
rect 8357 1050 8415 1105
rect 8445 1412 8503 1450
rect 8445 1378 8457 1412
rect 8491 1378 8503 1412
rect 8445 1344 8503 1378
rect 8445 1310 8457 1344
rect 8491 1310 8503 1344
rect 8445 1276 8503 1310
rect 8445 1242 8457 1276
rect 8491 1242 8503 1276
rect 8445 1208 8503 1242
rect 8445 1174 8457 1208
rect 8491 1174 8503 1208
rect 8445 1050 8503 1174
rect 8533 1412 8591 1450
rect 8533 1378 8545 1412
rect 8579 1378 8591 1412
rect 8533 1344 8591 1378
rect 8533 1310 8545 1344
rect 8579 1310 8591 1344
rect 8533 1276 8591 1310
rect 8533 1242 8545 1276
rect 8579 1242 8591 1276
rect 8533 1208 8591 1242
rect 8533 1174 8545 1208
rect 8579 1174 8591 1208
rect 8533 1139 8591 1174
rect 8533 1105 8545 1139
rect 8579 1105 8591 1139
rect 8533 1050 8591 1105
rect 8621 1412 8675 1450
rect 8621 1378 8633 1412
rect 8667 1378 8675 1412
rect 8621 1344 8675 1378
rect 8621 1310 8633 1344
rect 8667 1310 8675 1344
rect 8621 1276 8675 1310
rect 8621 1242 8633 1276
rect 8667 1242 8675 1276
rect 8621 1208 8675 1242
rect 8621 1174 8633 1208
rect 8667 1174 8675 1208
rect 8621 1050 8675 1174
rect 8997 1412 9053 1450
rect 8997 1378 9007 1412
rect 9041 1378 9053 1412
rect 8997 1344 9053 1378
rect 8997 1310 9007 1344
rect 9041 1310 9053 1344
rect 8997 1276 9053 1310
rect 8997 1242 9007 1276
rect 9041 1242 9053 1276
rect 8997 1208 9053 1242
rect 8997 1174 9007 1208
rect 9041 1174 9053 1208
rect 8997 1139 9053 1174
rect 8997 1105 9007 1139
rect 9041 1105 9053 1139
rect 8997 1050 9053 1105
rect 9083 1412 9141 1450
rect 9083 1378 9095 1412
rect 9129 1378 9141 1412
rect 9083 1344 9141 1378
rect 9083 1310 9095 1344
rect 9129 1310 9141 1344
rect 9083 1276 9141 1310
rect 9083 1242 9095 1276
rect 9129 1242 9141 1276
rect 9083 1208 9141 1242
rect 9083 1174 9095 1208
rect 9129 1174 9141 1208
rect 9083 1139 9141 1174
rect 9083 1105 9095 1139
rect 9129 1105 9141 1139
rect 9083 1050 9141 1105
rect 9171 1412 9229 1450
rect 9171 1378 9183 1412
rect 9217 1378 9229 1412
rect 9171 1344 9229 1378
rect 9171 1310 9183 1344
rect 9217 1310 9229 1344
rect 9171 1276 9229 1310
rect 9171 1242 9183 1276
rect 9217 1242 9229 1276
rect 9171 1208 9229 1242
rect 9171 1174 9183 1208
rect 9217 1174 9229 1208
rect 9171 1050 9229 1174
rect 9259 1412 9317 1450
rect 9259 1378 9271 1412
rect 9305 1378 9317 1412
rect 9259 1344 9317 1378
rect 9259 1310 9271 1344
rect 9305 1310 9317 1344
rect 9259 1276 9317 1310
rect 9259 1242 9271 1276
rect 9305 1242 9317 1276
rect 9259 1208 9317 1242
rect 9259 1174 9271 1208
rect 9305 1174 9317 1208
rect 9259 1139 9317 1174
rect 9259 1105 9271 1139
rect 9305 1105 9317 1139
rect 9259 1050 9317 1105
rect 9347 1412 9405 1450
rect 9347 1378 9359 1412
rect 9393 1378 9405 1412
rect 9347 1344 9405 1378
rect 9347 1310 9359 1344
rect 9393 1310 9405 1344
rect 9347 1276 9405 1310
rect 9347 1242 9359 1276
rect 9393 1242 9405 1276
rect 9347 1208 9405 1242
rect 9347 1174 9359 1208
rect 9393 1174 9405 1208
rect 9347 1050 9405 1174
rect 9435 1412 9493 1450
rect 9435 1378 9447 1412
rect 9481 1378 9493 1412
rect 9435 1344 9493 1378
rect 9435 1310 9447 1344
rect 9481 1310 9493 1344
rect 9435 1276 9493 1310
rect 9435 1242 9447 1276
rect 9481 1242 9493 1276
rect 9435 1208 9493 1242
rect 9435 1174 9447 1208
rect 9481 1174 9493 1208
rect 9435 1139 9493 1174
rect 9435 1105 9447 1139
rect 9481 1105 9493 1139
rect 9435 1050 9493 1105
rect 9523 1412 9577 1450
rect 9523 1378 9535 1412
rect 9569 1378 9577 1412
rect 9523 1344 9577 1378
rect 9523 1310 9535 1344
rect 9569 1310 9577 1344
rect 9523 1276 9577 1310
rect 9523 1242 9535 1276
rect 9569 1242 9577 1276
rect 9523 1208 9577 1242
rect 9523 1174 9535 1208
rect 9569 1174 9577 1208
rect 9523 1050 9577 1174
rect 9899 1412 9955 1450
rect 9899 1378 9909 1412
rect 9943 1378 9955 1412
rect 9899 1344 9955 1378
rect 9899 1310 9909 1344
rect 9943 1310 9955 1344
rect 9899 1276 9955 1310
rect 9899 1242 9909 1276
rect 9943 1242 9955 1276
rect 9899 1208 9955 1242
rect 9899 1174 9909 1208
rect 9943 1174 9955 1208
rect 9899 1139 9955 1174
rect 9899 1105 9909 1139
rect 9943 1105 9955 1139
rect 9899 1050 9955 1105
rect 9985 1412 10043 1450
rect 9985 1378 9997 1412
rect 10031 1378 10043 1412
rect 9985 1344 10043 1378
rect 9985 1310 9997 1344
rect 10031 1310 10043 1344
rect 9985 1276 10043 1310
rect 9985 1242 9997 1276
rect 10031 1242 10043 1276
rect 9985 1208 10043 1242
rect 9985 1174 9997 1208
rect 10031 1174 10043 1208
rect 9985 1139 10043 1174
rect 9985 1105 9997 1139
rect 10031 1105 10043 1139
rect 9985 1050 10043 1105
rect 10073 1412 10131 1450
rect 10073 1378 10085 1412
rect 10119 1378 10131 1412
rect 10073 1344 10131 1378
rect 10073 1310 10085 1344
rect 10119 1310 10131 1344
rect 10073 1276 10131 1310
rect 10073 1242 10085 1276
rect 10119 1242 10131 1276
rect 10073 1208 10131 1242
rect 10073 1174 10085 1208
rect 10119 1174 10131 1208
rect 10073 1050 10131 1174
rect 10161 1412 10219 1450
rect 10161 1378 10173 1412
rect 10207 1378 10219 1412
rect 10161 1344 10219 1378
rect 10161 1310 10173 1344
rect 10207 1310 10219 1344
rect 10161 1276 10219 1310
rect 10161 1242 10173 1276
rect 10207 1242 10219 1276
rect 10161 1208 10219 1242
rect 10161 1174 10173 1208
rect 10207 1174 10219 1208
rect 10161 1139 10219 1174
rect 10161 1105 10173 1139
rect 10207 1105 10219 1139
rect 10161 1050 10219 1105
rect 10249 1412 10303 1450
rect 10249 1378 10261 1412
rect 10295 1378 10303 1412
rect 10249 1344 10303 1378
rect 10249 1310 10261 1344
rect 10295 1310 10303 1344
rect 10249 1276 10303 1310
rect 10249 1242 10261 1276
rect 10295 1242 10303 1276
rect 10249 1208 10303 1242
rect 10249 1174 10261 1208
rect 10295 1174 10303 1208
rect 10249 1050 10303 1174
rect 10625 1412 10681 1450
rect 10625 1378 10635 1412
rect 10669 1378 10681 1412
rect 10625 1344 10681 1378
rect 10625 1310 10635 1344
rect 10669 1310 10681 1344
rect 10625 1276 10681 1310
rect 10625 1242 10635 1276
rect 10669 1242 10681 1276
rect 10625 1208 10681 1242
rect 10625 1174 10635 1208
rect 10669 1174 10681 1208
rect 10625 1139 10681 1174
rect 10625 1105 10635 1139
rect 10669 1105 10681 1139
rect 10625 1050 10681 1105
rect 10711 1412 10769 1450
rect 10711 1378 10723 1412
rect 10757 1378 10769 1412
rect 10711 1344 10769 1378
rect 10711 1310 10723 1344
rect 10757 1310 10769 1344
rect 10711 1276 10769 1310
rect 10711 1242 10723 1276
rect 10757 1242 10769 1276
rect 10711 1208 10769 1242
rect 10711 1174 10723 1208
rect 10757 1174 10769 1208
rect 10711 1139 10769 1174
rect 10711 1105 10723 1139
rect 10757 1105 10769 1139
rect 10711 1050 10769 1105
rect 10799 1412 10857 1450
rect 10799 1378 10811 1412
rect 10845 1378 10857 1412
rect 10799 1344 10857 1378
rect 10799 1310 10811 1344
rect 10845 1310 10857 1344
rect 10799 1276 10857 1310
rect 10799 1242 10811 1276
rect 10845 1242 10857 1276
rect 10799 1208 10857 1242
rect 10799 1174 10811 1208
rect 10845 1174 10857 1208
rect 10799 1050 10857 1174
rect 10887 1412 10945 1450
rect 10887 1378 10899 1412
rect 10933 1378 10945 1412
rect 10887 1344 10945 1378
rect 10887 1310 10899 1344
rect 10933 1310 10945 1344
rect 10887 1276 10945 1310
rect 10887 1242 10899 1276
rect 10933 1242 10945 1276
rect 10887 1208 10945 1242
rect 10887 1174 10899 1208
rect 10933 1174 10945 1208
rect 10887 1139 10945 1174
rect 10887 1105 10899 1139
rect 10933 1105 10945 1139
rect 10887 1050 10945 1105
rect 10975 1412 11033 1450
rect 10975 1378 10987 1412
rect 11021 1378 11033 1412
rect 10975 1344 11033 1378
rect 10975 1310 10987 1344
rect 11021 1310 11033 1344
rect 10975 1276 11033 1310
rect 10975 1242 10987 1276
rect 11021 1242 11033 1276
rect 10975 1208 11033 1242
rect 10975 1174 10987 1208
rect 11021 1174 11033 1208
rect 10975 1050 11033 1174
rect 11063 1412 11121 1450
rect 11063 1378 11075 1412
rect 11109 1378 11121 1412
rect 11063 1344 11121 1378
rect 11063 1310 11075 1344
rect 11109 1310 11121 1344
rect 11063 1276 11121 1310
rect 11063 1242 11075 1276
rect 11109 1242 11121 1276
rect 11063 1208 11121 1242
rect 11063 1174 11075 1208
rect 11109 1174 11121 1208
rect 11063 1139 11121 1174
rect 11063 1105 11075 1139
rect 11109 1105 11121 1139
rect 11063 1050 11121 1105
rect 11151 1412 11205 1450
rect 11151 1378 11163 1412
rect 11197 1378 11205 1412
rect 11151 1344 11205 1378
rect 11151 1310 11163 1344
rect 11197 1310 11205 1344
rect 11151 1276 11205 1310
rect 11151 1242 11163 1276
rect 11197 1242 11205 1276
rect 11151 1208 11205 1242
rect 11151 1174 11163 1208
rect 11197 1174 11205 1208
rect 11151 1050 11205 1174
rect 11587 1412 11643 1450
rect 11587 1378 11597 1412
rect 11631 1378 11643 1412
rect 11587 1344 11643 1378
rect 11587 1310 11597 1344
rect 11631 1310 11643 1344
rect 11587 1276 11643 1310
rect 11587 1242 11597 1276
rect 11631 1242 11643 1276
rect 11587 1208 11643 1242
rect 11587 1174 11597 1208
rect 11631 1174 11643 1208
rect 11587 1139 11643 1174
rect 11587 1105 11597 1139
rect 11631 1105 11643 1139
rect 11587 1050 11643 1105
rect 11673 1412 11731 1450
rect 11673 1378 11685 1412
rect 11719 1378 11731 1412
rect 11673 1344 11731 1378
rect 11673 1310 11685 1344
rect 11719 1310 11731 1344
rect 11673 1276 11731 1310
rect 11673 1242 11685 1276
rect 11719 1242 11731 1276
rect 11673 1208 11731 1242
rect 11673 1174 11685 1208
rect 11719 1174 11731 1208
rect 11673 1139 11731 1174
rect 11673 1105 11685 1139
rect 11719 1105 11731 1139
rect 11673 1050 11731 1105
rect 11761 1412 11819 1450
rect 11761 1378 11773 1412
rect 11807 1378 11819 1412
rect 11761 1344 11819 1378
rect 11761 1310 11773 1344
rect 11807 1310 11819 1344
rect 11761 1276 11819 1310
rect 11761 1242 11773 1276
rect 11807 1242 11819 1276
rect 11761 1208 11819 1242
rect 11761 1174 11773 1208
rect 11807 1174 11819 1208
rect 11761 1050 11819 1174
rect 11849 1412 11907 1450
rect 11849 1378 11861 1412
rect 11895 1378 11907 1412
rect 11849 1344 11907 1378
rect 11849 1310 11861 1344
rect 11895 1310 11907 1344
rect 11849 1276 11907 1310
rect 11849 1242 11861 1276
rect 11895 1242 11907 1276
rect 11849 1208 11907 1242
rect 11849 1174 11861 1208
rect 11895 1174 11907 1208
rect 11849 1139 11907 1174
rect 11849 1105 11861 1139
rect 11895 1105 11907 1139
rect 11849 1050 11907 1105
rect 11937 1412 11995 1450
rect 11937 1378 11949 1412
rect 11983 1378 11995 1412
rect 11937 1344 11995 1378
rect 11937 1310 11949 1344
rect 11983 1310 11995 1344
rect 11937 1276 11995 1310
rect 11937 1242 11949 1276
rect 11983 1242 11995 1276
rect 11937 1208 11995 1242
rect 11937 1174 11949 1208
rect 11983 1174 11995 1208
rect 11937 1050 11995 1174
rect 12025 1412 12083 1450
rect 12025 1378 12037 1412
rect 12071 1378 12083 1412
rect 12025 1344 12083 1378
rect 12025 1310 12037 1344
rect 12071 1310 12083 1344
rect 12025 1276 12083 1310
rect 12025 1242 12037 1276
rect 12071 1242 12083 1276
rect 12025 1208 12083 1242
rect 12025 1174 12037 1208
rect 12071 1174 12083 1208
rect 12025 1139 12083 1174
rect 12025 1105 12037 1139
rect 12071 1105 12083 1139
rect 12025 1050 12083 1105
rect 12113 1412 12167 1450
rect 12113 1378 12125 1412
rect 12159 1378 12167 1412
rect 12113 1344 12167 1378
rect 12113 1310 12125 1344
rect 12159 1310 12167 1344
rect 12113 1276 12167 1310
rect 12113 1242 12125 1276
rect 12159 1242 12167 1276
rect 12113 1208 12167 1242
rect 12113 1174 12125 1208
rect 12159 1174 12167 1208
rect 12113 1050 12167 1174
rect 12489 1412 12545 1450
rect 12489 1378 12499 1412
rect 12533 1378 12545 1412
rect 12489 1344 12545 1378
rect 12489 1310 12499 1344
rect 12533 1310 12545 1344
rect 12489 1276 12545 1310
rect 12489 1242 12499 1276
rect 12533 1242 12545 1276
rect 12489 1208 12545 1242
rect 12489 1174 12499 1208
rect 12533 1174 12545 1208
rect 12489 1139 12545 1174
rect 12489 1105 12499 1139
rect 12533 1105 12545 1139
rect 12489 1050 12545 1105
rect 12575 1412 12633 1450
rect 12575 1378 12587 1412
rect 12621 1378 12633 1412
rect 12575 1344 12633 1378
rect 12575 1310 12587 1344
rect 12621 1310 12633 1344
rect 12575 1276 12633 1310
rect 12575 1242 12587 1276
rect 12621 1242 12633 1276
rect 12575 1208 12633 1242
rect 12575 1174 12587 1208
rect 12621 1174 12633 1208
rect 12575 1139 12633 1174
rect 12575 1105 12587 1139
rect 12621 1105 12633 1139
rect 12575 1050 12633 1105
rect 12663 1412 12721 1450
rect 12663 1378 12675 1412
rect 12709 1378 12721 1412
rect 12663 1344 12721 1378
rect 12663 1310 12675 1344
rect 12709 1310 12721 1344
rect 12663 1276 12721 1310
rect 12663 1242 12675 1276
rect 12709 1242 12721 1276
rect 12663 1208 12721 1242
rect 12663 1174 12675 1208
rect 12709 1174 12721 1208
rect 12663 1050 12721 1174
rect 12751 1412 12809 1450
rect 12751 1378 12763 1412
rect 12797 1378 12809 1412
rect 12751 1344 12809 1378
rect 12751 1310 12763 1344
rect 12797 1310 12809 1344
rect 12751 1276 12809 1310
rect 12751 1242 12763 1276
rect 12797 1242 12809 1276
rect 12751 1208 12809 1242
rect 12751 1174 12763 1208
rect 12797 1174 12809 1208
rect 12751 1139 12809 1174
rect 12751 1105 12763 1139
rect 12797 1105 12809 1139
rect 12751 1050 12809 1105
rect 12839 1412 12893 1450
rect 12839 1378 12851 1412
rect 12885 1378 12893 1412
rect 12839 1344 12893 1378
rect 12839 1310 12851 1344
rect 12885 1310 12893 1344
rect 12839 1276 12893 1310
rect 12839 1242 12851 1276
rect 12885 1242 12893 1276
rect 12839 1208 12893 1242
rect 12839 1174 12851 1208
rect 12885 1174 12893 1208
rect 12839 1050 12893 1174
rect 13155 1412 13211 1450
rect 13155 1378 13165 1412
rect 13199 1378 13211 1412
rect 13155 1344 13211 1378
rect 13155 1310 13165 1344
rect 13199 1310 13211 1344
rect 13155 1276 13211 1310
rect 13155 1242 13165 1276
rect 13199 1242 13211 1276
rect 13155 1208 13211 1242
rect 13155 1174 13165 1208
rect 13199 1174 13211 1208
rect 13155 1139 13211 1174
rect 13155 1105 13165 1139
rect 13199 1105 13211 1139
rect 13155 1050 13211 1105
rect 13241 1412 13299 1450
rect 13241 1378 13253 1412
rect 13287 1378 13299 1412
rect 13241 1344 13299 1378
rect 13241 1310 13253 1344
rect 13287 1310 13299 1344
rect 13241 1276 13299 1310
rect 13241 1242 13253 1276
rect 13287 1242 13299 1276
rect 13241 1208 13299 1242
rect 13241 1174 13253 1208
rect 13287 1174 13299 1208
rect 13241 1139 13299 1174
rect 13241 1105 13253 1139
rect 13287 1105 13299 1139
rect 13241 1050 13299 1105
rect 13329 1412 13387 1450
rect 13329 1378 13341 1412
rect 13375 1378 13387 1412
rect 13329 1344 13387 1378
rect 13329 1310 13341 1344
rect 13375 1310 13387 1344
rect 13329 1276 13387 1310
rect 13329 1242 13341 1276
rect 13375 1242 13387 1276
rect 13329 1208 13387 1242
rect 13329 1174 13341 1208
rect 13375 1174 13387 1208
rect 13329 1050 13387 1174
rect 13417 1412 13475 1450
rect 13417 1378 13429 1412
rect 13463 1378 13475 1412
rect 13417 1344 13475 1378
rect 13417 1310 13429 1344
rect 13463 1310 13475 1344
rect 13417 1276 13475 1310
rect 13417 1242 13429 1276
rect 13463 1242 13475 1276
rect 13417 1208 13475 1242
rect 13417 1174 13429 1208
rect 13463 1174 13475 1208
rect 13417 1139 13475 1174
rect 13417 1105 13429 1139
rect 13463 1105 13475 1139
rect 13417 1050 13475 1105
rect 13505 1412 13559 1450
rect 13505 1378 13517 1412
rect 13551 1378 13559 1412
rect 13505 1344 13559 1378
rect 13505 1310 13517 1344
rect 13551 1310 13559 1344
rect 13505 1276 13559 1310
rect 13505 1242 13517 1276
rect 13551 1242 13559 1276
rect 13505 1208 13559 1242
rect 13505 1174 13517 1208
rect 13551 1174 13559 1208
rect 13505 1050 13559 1174
rect 13881 1412 13937 1450
rect 13881 1378 13891 1412
rect 13925 1378 13937 1412
rect 13881 1344 13937 1378
rect 13881 1310 13891 1344
rect 13925 1310 13937 1344
rect 13881 1276 13937 1310
rect 13881 1242 13891 1276
rect 13925 1242 13937 1276
rect 13881 1208 13937 1242
rect 13881 1174 13891 1208
rect 13925 1174 13937 1208
rect 13881 1139 13937 1174
rect 13881 1105 13891 1139
rect 13925 1105 13937 1139
rect 13881 1050 13937 1105
rect 13967 1412 14025 1450
rect 13967 1378 13979 1412
rect 14013 1378 14025 1412
rect 13967 1344 14025 1378
rect 13967 1310 13979 1344
rect 14013 1310 14025 1344
rect 13967 1276 14025 1310
rect 13967 1242 13979 1276
rect 14013 1242 14025 1276
rect 13967 1208 14025 1242
rect 13967 1174 13979 1208
rect 14013 1174 14025 1208
rect 13967 1139 14025 1174
rect 13967 1105 13979 1139
rect 14013 1105 14025 1139
rect 13967 1050 14025 1105
rect 14055 1412 14113 1450
rect 14055 1378 14067 1412
rect 14101 1378 14113 1412
rect 14055 1344 14113 1378
rect 14055 1310 14067 1344
rect 14101 1310 14113 1344
rect 14055 1276 14113 1310
rect 14055 1242 14067 1276
rect 14101 1242 14113 1276
rect 14055 1208 14113 1242
rect 14055 1174 14067 1208
rect 14101 1174 14113 1208
rect 14055 1050 14113 1174
rect 14143 1412 14201 1450
rect 14143 1378 14155 1412
rect 14189 1378 14201 1412
rect 14143 1344 14201 1378
rect 14143 1310 14155 1344
rect 14189 1310 14201 1344
rect 14143 1276 14201 1310
rect 14143 1242 14155 1276
rect 14189 1242 14201 1276
rect 14143 1208 14201 1242
rect 14143 1174 14155 1208
rect 14189 1174 14201 1208
rect 14143 1139 14201 1174
rect 14143 1105 14155 1139
rect 14189 1105 14201 1139
rect 14143 1050 14201 1105
rect 14231 1412 14289 1450
rect 14231 1378 14243 1412
rect 14277 1378 14289 1412
rect 14231 1344 14289 1378
rect 14231 1310 14243 1344
rect 14277 1310 14289 1344
rect 14231 1276 14289 1310
rect 14231 1242 14243 1276
rect 14277 1242 14289 1276
rect 14231 1208 14289 1242
rect 14231 1174 14243 1208
rect 14277 1174 14289 1208
rect 14231 1050 14289 1174
rect 14319 1412 14377 1450
rect 14319 1378 14331 1412
rect 14365 1378 14377 1412
rect 14319 1344 14377 1378
rect 14319 1310 14331 1344
rect 14365 1310 14377 1344
rect 14319 1276 14377 1310
rect 14319 1242 14331 1276
rect 14365 1242 14377 1276
rect 14319 1208 14377 1242
rect 14319 1174 14331 1208
rect 14365 1174 14377 1208
rect 14319 1139 14377 1174
rect 14319 1105 14331 1139
rect 14365 1105 14377 1139
rect 14319 1050 14377 1105
rect 14407 1412 14461 1450
rect 14407 1378 14419 1412
rect 14453 1378 14461 1412
rect 14407 1344 14461 1378
rect 14407 1310 14419 1344
rect 14453 1310 14461 1344
rect 14407 1276 14461 1310
rect 14407 1242 14419 1276
rect 14453 1242 14461 1276
rect 14407 1208 14461 1242
rect 14407 1174 14419 1208
rect 14453 1174 14461 1208
rect 14407 1050 14461 1174
rect 14783 1411 14839 1451
rect 14783 1377 14793 1411
rect 14827 1377 14839 1411
rect 14783 1343 14839 1377
rect 14783 1309 14793 1343
rect 14827 1309 14839 1343
rect 14783 1275 14839 1309
rect 14783 1241 14793 1275
rect 14827 1241 14839 1275
rect 14783 1207 14839 1241
rect 14783 1173 14793 1207
rect 14827 1173 14839 1207
rect 14783 1139 14839 1173
rect 14783 1105 14793 1139
rect 14827 1105 14839 1139
rect 14783 1051 14839 1105
rect 14869 1411 14927 1451
rect 14869 1377 14881 1411
rect 14915 1377 14927 1411
rect 14869 1343 14927 1377
rect 14869 1309 14881 1343
rect 14915 1309 14927 1343
rect 14869 1275 14927 1309
rect 14869 1241 14881 1275
rect 14915 1241 14927 1275
rect 14869 1207 14927 1241
rect 14869 1173 14881 1207
rect 14915 1173 14927 1207
rect 14869 1139 14927 1173
rect 14869 1105 14881 1139
rect 14915 1105 14927 1139
rect 14869 1051 14927 1105
rect 14957 1411 15015 1451
rect 14957 1377 14969 1411
rect 15003 1377 15015 1411
rect 14957 1343 15015 1377
rect 14957 1309 14969 1343
rect 15003 1309 15015 1343
rect 14957 1275 15015 1309
rect 14957 1241 14969 1275
rect 15003 1241 15015 1275
rect 14957 1207 15015 1241
rect 14957 1173 14969 1207
rect 15003 1173 15015 1207
rect 14957 1051 15015 1173
rect 15045 1411 15103 1451
rect 15045 1377 15057 1411
rect 15091 1377 15103 1411
rect 15045 1343 15103 1377
rect 15045 1309 15057 1343
rect 15091 1309 15103 1343
rect 15045 1275 15103 1309
rect 15045 1241 15057 1275
rect 15091 1241 15103 1275
rect 15045 1207 15103 1241
rect 15045 1173 15057 1207
rect 15091 1173 15103 1207
rect 15045 1051 15103 1173
rect 15133 1411 15187 1451
rect 15133 1377 15145 1411
rect 15179 1377 15187 1411
rect 15133 1343 15187 1377
rect 15133 1309 15145 1343
rect 15179 1309 15187 1343
rect 15133 1275 15187 1309
rect 15133 1241 15145 1275
rect 15179 1241 15187 1275
rect 15133 1207 15187 1241
rect 15133 1173 15145 1207
rect 15179 1173 15187 1207
rect 15133 1139 15187 1173
rect 15133 1105 15145 1139
rect 15179 1105 15187 1139
rect 15133 1051 15187 1105
rect 15449 1411 15503 1451
rect 15449 1377 15457 1411
rect 15491 1377 15503 1411
rect 15449 1343 15503 1377
rect 15449 1309 15457 1343
rect 15491 1309 15503 1343
rect 15449 1275 15503 1309
rect 15449 1241 15457 1275
rect 15491 1241 15503 1275
rect 15449 1207 15503 1241
rect 15449 1173 15457 1207
rect 15491 1173 15503 1207
rect 15449 1051 15503 1173
rect 15533 1343 15591 1451
rect 15533 1309 15545 1343
rect 15579 1309 15591 1343
rect 15533 1275 15591 1309
rect 15533 1241 15545 1275
rect 15579 1241 15591 1275
rect 15533 1207 15591 1241
rect 15533 1173 15545 1207
rect 15579 1173 15591 1207
rect 15533 1139 15591 1173
rect 15533 1105 15545 1139
rect 15579 1105 15591 1139
rect 15533 1051 15591 1105
rect 15621 1411 15679 1451
rect 15621 1377 15633 1411
rect 15667 1377 15679 1411
rect 15621 1343 15679 1377
rect 15621 1309 15633 1343
rect 15667 1309 15679 1343
rect 15621 1275 15679 1309
rect 15621 1241 15633 1275
rect 15667 1241 15679 1275
rect 15621 1207 15679 1241
rect 15621 1173 15633 1207
rect 15667 1173 15679 1207
rect 15621 1051 15679 1173
rect 15709 1343 15767 1451
rect 15709 1309 15721 1343
rect 15755 1309 15767 1343
rect 15709 1275 15767 1309
rect 15709 1241 15721 1275
rect 15755 1241 15767 1275
rect 15709 1207 15767 1241
rect 15709 1173 15721 1207
rect 15755 1173 15767 1207
rect 15709 1051 15767 1173
rect 15797 1411 15853 1451
rect 15797 1377 15809 1411
rect 15843 1377 15853 1411
rect 15797 1343 15853 1377
rect 15797 1309 15809 1343
rect 15843 1309 15853 1343
rect 15797 1275 15853 1309
rect 15797 1241 15809 1275
rect 15843 1241 15853 1275
rect 15797 1207 15853 1241
rect 15797 1173 15809 1207
rect 15843 1173 15853 1207
rect 15797 1051 15853 1173
rect 16115 1411 16171 1451
rect 16115 1377 16125 1411
rect 16159 1377 16171 1411
rect 16115 1343 16171 1377
rect 16115 1309 16125 1343
rect 16159 1309 16171 1343
rect 16115 1275 16171 1309
rect 16115 1241 16125 1275
rect 16159 1241 16171 1275
rect 16115 1207 16171 1241
rect 16115 1173 16125 1207
rect 16159 1173 16171 1207
rect 16115 1051 16171 1173
rect 16201 1343 16259 1451
rect 16201 1309 16213 1343
rect 16247 1309 16259 1343
rect 16201 1275 16259 1309
rect 16201 1241 16213 1275
rect 16247 1241 16259 1275
rect 16201 1207 16259 1241
rect 16201 1173 16213 1207
rect 16247 1173 16259 1207
rect 16201 1139 16259 1173
rect 16201 1105 16213 1139
rect 16247 1105 16259 1139
rect 16201 1051 16259 1105
rect 16289 1411 16347 1451
rect 16289 1377 16301 1411
rect 16335 1377 16347 1411
rect 16289 1343 16347 1377
rect 16289 1309 16301 1343
rect 16335 1309 16347 1343
rect 16289 1275 16347 1309
rect 16289 1241 16301 1275
rect 16335 1241 16347 1275
rect 16289 1207 16347 1241
rect 16289 1173 16301 1207
rect 16335 1173 16347 1207
rect 16289 1051 16347 1173
rect 16377 1343 16435 1451
rect 16377 1309 16389 1343
rect 16423 1309 16435 1343
rect 16377 1275 16435 1309
rect 16377 1241 16389 1275
rect 16423 1241 16435 1275
rect 16377 1207 16435 1241
rect 16377 1173 16389 1207
rect 16423 1173 16435 1207
rect 16377 1139 16435 1173
rect 16377 1105 16389 1139
rect 16423 1105 16435 1139
rect 16377 1051 16435 1105
rect 16465 1411 16519 1451
rect 16465 1377 16477 1411
rect 16511 1377 16519 1411
rect 16465 1343 16519 1377
rect 16465 1309 16477 1343
rect 16511 1309 16519 1343
rect 16465 1275 16519 1309
rect 16465 1241 16477 1275
rect 16511 1241 16519 1275
rect 16465 1207 16519 1241
rect 16465 1173 16477 1207
rect 16511 1173 16519 1207
rect 16465 1051 16519 1173
<< ndiffc >>
rect 122 327 156 361
rect 219 327 253 361
rect 316 327 350 361
rect 122 255 156 289
rect 122 187 156 221
rect 219 202 253 236
rect 316 255 350 289
rect 316 187 350 221
rect 413 211 447 245
rect 510 255 544 289
rect 510 187 544 221
rect 122 117 156 151
rect 316 117 350 151
rect 413 117 447 151
rect 510 117 544 151
rect 767 329 801 363
rect 864 329 898 363
rect 961 329 995 363
rect 1058 329 1092 363
rect 1155 329 1189 363
rect 767 257 801 291
rect 767 189 801 223
rect 864 204 898 238
rect 961 257 995 291
rect 961 189 995 223
rect 1059 210 1093 244
rect 767 119 801 153
rect 961 119 995 153
rect 1058 119 1092 153
rect 1155 119 1189 153
rect 1269 329 1303 363
rect 1269 257 1303 291
rect 1269 189 1303 223
rect 1366 213 1400 247
rect 1463 257 1497 291
rect 1463 189 1497 223
rect 1269 119 1303 153
rect 1366 119 1400 153
rect 1463 119 1497 153
rect 1729 329 1763 363
rect 1826 329 1860 363
rect 1923 329 1957 363
rect 2020 329 2054 363
rect 2117 329 2151 363
rect 1729 257 1763 291
rect 1729 189 1763 223
rect 1826 204 1860 238
rect 1923 257 1957 291
rect 1923 189 1957 223
rect 2021 210 2055 244
rect 1729 119 1763 153
rect 1923 119 1957 153
rect 2020 119 2054 153
rect 2117 119 2151 153
rect 2231 329 2265 363
rect 2231 257 2265 291
rect 2231 189 2265 223
rect 2328 213 2362 247
rect 2425 257 2459 291
rect 2425 189 2459 223
rect 2231 119 2265 153
rect 2328 119 2362 153
rect 2425 119 2459 153
rect 2712 327 2746 361
rect 2809 327 2843 361
rect 2906 327 2940 361
rect 2712 255 2746 289
rect 2712 187 2746 221
rect 2809 202 2843 236
rect 2906 255 2940 289
rect 2906 187 2940 221
rect 3003 211 3037 245
rect 3100 255 3134 289
rect 3100 187 3134 221
rect 2712 117 2746 151
rect 2906 117 2940 151
rect 3003 117 3037 151
rect 3100 117 3134 151
rect 3378 327 3412 361
rect 3475 327 3509 361
rect 3572 327 3606 361
rect 3378 255 3412 289
rect 3378 187 3412 221
rect 3475 202 3509 236
rect 3572 255 3606 289
rect 3572 187 3606 221
rect 3669 211 3703 245
rect 3766 255 3800 289
rect 3766 187 3800 221
rect 3378 117 3412 151
rect 3572 117 3606 151
rect 3669 117 3703 151
rect 3766 117 3800 151
rect 4023 329 4057 363
rect 4120 329 4154 363
rect 4217 329 4251 363
rect 4314 329 4348 363
rect 4411 329 4445 363
rect 4023 257 4057 291
rect 4023 189 4057 223
rect 4120 204 4154 238
rect 4217 257 4251 291
rect 4217 189 4251 223
rect 4315 210 4349 244
rect 4023 119 4057 153
rect 4217 119 4251 153
rect 4314 119 4348 153
rect 4411 119 4445 153
rect 4525 329 4559 363
rect 4525 257 4559 291
rect 4525 189 4559 223
rect 4622 213 4656 247
rect 4719 257 4753 291
rect 4719 189 4753 223
rect 4525 119 4559 153
rect 4622 119 4656 153
rect 4719 119 4753 153
rect 5006 327 5040 361
rect 5103 327 5137 361
rect 5200 327 5234 361
rect 5006 255 5040 289
rect 5006 187 5040 221
rect 5103 202 5137 236
rect 5200 255 5234 289
rect 5200 187 5234 221
rect 5297 211 5331 245
rect 5394 255 5428 289
rect 5394 187 5428 221
rect 5006 117 5040 151
rect 5200 117 5234 151
rect 5297 117 5331 151
rect 5394 117 5428 151
rect 5651 329 5685 363
rect 5748 329 5782 363
rect 5845 329 5879 363
rect 5942 329 5976 363
rect 6039 329 6073 363
rect 5651 257 5685 291
rect 5651 189 5685 223
rect 5748 204 5782 238
rect 5845 257 5879 291
rect 5845 189 5879 223
rect 5943 210 5977 244
rect 5651 119 5685 153
rect 5845 119 5879 153
rect 5942 119 5976 153
rect 6039 119 6073 153
rect 6153 329 6187 363
rect 6153 257 6187 291
rect 6153 189 6187 223
rect 6250 213 6284 247
rect 6347 257 6381 291
rect 6347 189 6381 223
rect 6153 119 6187 153
rect 6250 119 6284 153
rect 6347 119 6381 153
rect 6613 329 6647 363
rect 6710 329 6744 363
rect 6807 329 6841 363
rect 6904 329 6938 363
rect 7001 329 7035 363
rect 6613 257 6647 291
rect 6613 189 6647 223
rect 6710 204 6744 238
rect 6807 257 6841 291
rect 6807 189 6841 223
rect 6905 210 6939 244
rect 6613 119 6647 153
rect 6807 119 6841 153
rect 6904 119 6938 153
rect 7001 119 7035 153
rect 7115 329 7149 363
rect 7115 257 7149 291
rect 7115 189 7149 223
rect 7212 213 7246 247
rect 7309 257 7343 291
rect 7309 189 7343 223
rect 7115 119 7149 153
rect 7212 119 7246 153
rect 7309 119 7343 153
rect 7596 327 7630 361
rect 7693 327 7727 361
rect 7790 327 7824 361
rect 7596 255 7630 289
rect 7596 187 7630 221
rect 7693 202 7727 236
rect 7790 255 7824 289
rect 7790 187 7824 221
rect 7887 211 7921 245
rect 7984 255 8018 289
rect 7984 187 8018 221
rect 7596 117 7630 151
rect 7790 117 7824 151
rect 7887 117 7921 151
rect 7984 117 8018 151
rect 8262 327 8296 361
rect 8359 327 8393 361
rect 8456 327 8490 361
rect 8262 255 8296 289
rect 8262 187 8296 221
rect 8359 202 8393 236
rect 8456 255 8490 289
rect 8456 187 8490 221
rect 8553 211 8587 245
rect 8650 255 8684 289
rect 8650 187 8684 221
rect 8262 117 8296 151
rect 8456 117 8490 151
rect 8553 117 8587 151
rect 8650 117 8684 151
rect 8907 329 8941 363
rect 9004 329 9038 363
rect 9101 329 9135 363
rect 9198 329 9232 363
rect 9295 329 9329 363
rect 8907 257 8941 291
rect 8907 189 8941 223
rect 9004 204 9038 238
rect 9101 257 9135 291
rect 9101 189 9135 223
rect 9199 210 9233 244
rect 8907 119 8941 153
rect 9101 119 9135 153
rect 9198 119 9232 153
rect 9295 119 9329 153
rect 9409 329 9443 363
rect 9409 257 9443 291
rect 9409 189 9443 223
rect 9506 213 9540 247
rect 9603 257 9637 291
rect 9603 189 9637 223
rect 9409 119 9443 153
rect 9506 119 9540 153
rect 9603 119 9637 153
rect 9890 327 9924 361
rect 9987 327 10021 361
rect 10084 327 10118 361
rect 9890 255 9924 289
rect 9890 187 9924 221
rect 9987 202 10021 236
rect 10084 255 10118 289
rect 10084 187 10118 221
rect 10181 211 10215 245
rect 10278 255 10312 289
rect 10278 187 10312 221
rect 9890 117 9924 151
rect 10084 117 10118 151
rect 10181 117 10215 151
rect 10278 117 10312 151
rect 10535 329 10569 363
rect 10632 329 10666 363
rect 10729 329 10763 363
rect 10826 329 10860 363
rect 10923 329 10957 363
rect 10535 257 10569 291
rect 10535 189 10569 223
rect 10632 204 10666 238
rect 10729 257 10763 291
rect 10729 189 10763 223
rect 10827 210 10861 244
rect 10535 119 10569 153
rect 10729 119 10763 153
rect 10826 119 10860 153
rect 10923 119 10957 153
rect 11037 329 11071 363
rect 11037 257 11071 291
rect 11037 189 11071 223
rect 11134 213 11168 247
rect 11231 257 11265 291
rect 11231 189 11265 223
rect 11037 119 11071 153
rect 11134 119 11168 153
rect 11231 119 11265 153
rect 11497 329 11531 363
rect 11594 329 11628 363
rect 11691 329 11725 363
rect 11788 329 11822 363
rect 11885 329 11919 363
rect 11497 257 11531 291
rect 11497 189 11531 223
rect 11594 204 11628 238
rect 11691 257 11725 291
rect 11691 189 11725 223
rect 11789 210 11823 244
rect 11497 119 11531 153
rect 11691 119 11725 153
rect 11788 119 11822 153
rect 11885 119 11919 153
rect 11999 329 12033 363
rect 11999 257 12033 291
rect 11999 189 12033 223
rect 12096 213 12130 247
rect 12193 257 12227 291
rect 12193 189 12227 223
rect 11999 119 12033 153
rect 12096 119 12130 153
rect 12193 119 12227 153
rect 12480 327 12514 361
rect 12577 327 12611 361
rect 12674 327 12708 361
rect 12480 255 12514 289
rect 12480 187 12514 221
rect 12577 202 12611 236
rect 12674 255 12708 289
rect 12674 187 12708 221
rect 12771 211 12805 245
rect 12868 255 12902 289
rect 12868 187 12902 221
rect 12480 117 12514 151
rect 12674 117 12708 151
rect 12771 117 12805 151
rect 12868 117 12902 151
rect 13146 327 13180 361
rect 13243 327 13277 361
rect 13340 327 13374 361
rect 13146 255 13180 289
rect 13146 187 13180 221
rect 13243 202 13277 236
rect 13340 255 13374 289
rect 13340 187 13374 221
rect 13437 211 13471 245
rect 13534 255 13568 289
rect 13534 187 13568 221
rect 13146 117 13180 151
rect 13340 117 13374 151
rect 13437 117 13471 151
rect 13534 117 13568 151
rect 13791 329 13825 363
rect 13888 329 13922 363
rect 13985 329 14019 363
rect 14082 329 14116 363
rect 14179 329 14213 363
rect 13791 257 13825 291
rect 13791 189 13825 223
rect 13888 204 13922 238
rect 13985 257 14019 291
rect 13985 189 14019 223
rect 14083 210 14117 244
rect 13791 119 13825 153
rect 13985 119 14019 153
rect 14082 119 14116 153
rect 14179 119 14213 153
rect 14293 329 14327 363
rect 14293 257 14327 291
rect 14293 189 14327 223
rect 14390 213 14424 247
rect 14487 257 14521 291
rect 14487 189 14521 223
rect 14293 119 14327 153
rect 14390 119 14424 153
rect 14487 119 14521 153
rect 14774 327 14808 361
rect 14871 327 14905 361
rect 14968 327 15002 361
rect 15162 327 15196 361
rect 14774 255 14808 289
rect 14774 187 14808 221
rect 14871 202 14905 236
rect 14968 255 15002 289
rect 14968 187 15002 221
rect 15064 211 15098 245
rect 15162 255 15196 289
rect 15162 187 15196 221
rect 14774 117 14808 151
rect 14968 117 15002 151
rect 15064 117 15098 151
rect 15162 117 15196 151
rect 15440 327 15474 361
rect 15537 327 15571 361
rect 15634 327 15668 361
rect 15828 327 15862 361
rect 15440 255 15474 289
rect 15440 187 15474 221
rect 15537 202 15571 236
rect 15634 255 15668 289
rect 15634 187 15668 221
rect 15731 211 15765 245
rect 15828 255 15862 289
rect 15828 187 15862 221
rect 15440 117 15474 151
rect 15634 117 15668 151
rect 15731 117 15765 151
rect 15828 117 15862 151
rect 16106 327 16140 361
rect 16203 327 16237 361
rect 16300 327 16334 361
rect 16106 255 16140 289
rect 16106 187 16140 221
rect 16203 202 16237 236
rect 16300 255 16334 289
rect 16300 187 16334 221
rect 16397 211 16431 245
rect 16494 255 16528 289
rect 16494 187 16528 221
rect 16106 117 16140 151
rect 16300 117 16334 151
rect 16397 117 16431 151
rect 16494 117 16528 151
<< pdiffc >>
rect 141 1378 175 1412
rect 141 1310 175 1344
rect 141 1242 175 1276
rect 141 1174 175 1208
rect 141 1105 175 1139
rect 229 1378 263 1412
rect 229 1310 263 1344
rect 229 1242 263 1276
rect 229 1174 263 1208
rect 229 1105 263 1139
rect 317 1378 351 1412
rect 317 1310 351 1344
rect 317 1242 351 1276
rect 317 1174 351 1208
rect 405 1378 439 1412
rect 405 1310 439 1344
rect 405 1242 439 1276
rect 405 1174 439 1208
rect 405 1105 439 1139
rect 493 1378 527 1412
rect 493 1310 527 1344
rect 493 1242 527 1276
rect 493 1174 527 1208
rect 867 1378 901 1412
rect 867 1310 901 1344
rect 867 1242 901 1276
rect 867 1174 901 1208
rect 867 1105 901 1139
rect 955 1378 989 1412
rect 955 1310 989 1344
rect 955 1242 989 1276
rect 955 1174 989 1208
rect 955 1105 989 1139
rect 1043 1378 1077 1412
rect 1043 1310 1077 1344
rect 1043 1242 1077 1276
rect 1043 1174 1077 1208
rect 1131 1378 1165 1412
rect 1131 1310 1165 1344
rect 1131 1242 1165 1276
rect 1131 1174 1165 1208
rect 1131 1105 1165 1139
rect 1219 1378 1253 1412
rect 1219 1310 1253 1344
rect 1219 1242 1253 1276
rect 1219 1174 1253 1208
rect 1307 1378 1341 1412
rect 1307 1310 1341 1344
rect 1307 1242 1341 1276
rect 1307 1174 1341 1208
rect 1307 1105 1341 1139
rect 1395 1378 1429 1412
rect 1395 1310 1429 1344
rect 1395 1242 1429 1276
rect 1395 1174 1429 1208
rect 1829 1378 1863 1412
rect 1829 1310 1863 1344
rect 1829 1242 1863 1276
rect 1829 1174 1863 1208
rect 1829 1105 1863 1139
rect 1917 1378 1951 1412
rect 1917 1310 1951 1344
rect 1917 1242 1951 1276
rect 1917 1174 1951 1208
rect 1917 1105 1951 1139
rect 2005 1378 2039 1412
rect 2005 1310 2039 1344
rect 2005 1242 2039 1276
rect 2005 1174 2039 1208
rect 2093 1378 2127 1412
rect 2093 1310 2127 1344
rect 2093 1242 2127 1276
rect 2093 1174 2127 1208
rect 2093 1105 2127 1139
rect 2181 1378 2215 1412
rect 2181 1310 2215 1344
rect 2181 1242 2215 1276
rect 2181 1174 2215 1208
rect 2269 1378 2303 1412
rect 2269 1310 2303 1344
rect 2269 1242 2303 1276
rect 2269 1174 2303 1208
rect 2269 1105 2303 1139
rect 2357 1378 2391 1412
rect 2357 1310 2391 1344
rect 2357 1242 2391 1276
rect 2357 1174 2391 1208
rect 2731 1378 2765 1412
rect 2731 1310 2765 1344
rect 2731 1242 2765 1276
rect 2731 1174 2765 1208
rect 2731 1105 2765 1139
rect 2819 1378 2853 1412
rect 2819 1310 2853 1344
rect 2819 1242 2853 1276
rect 2819 1174 2853 1208
rect 2819 1105 2853 1139
rect 2907 1378 2941 1412
rect 2907 1310 2941 1344
rect 2907 1242 2941 1276
rect 2907 1174 2941 1208
rect 2995 1378 3029 1412
rect 2995 1310 3029 1344
rect 2995 1242 3029 1276
rect 2995 1174 3029 1208
rect 2995 1105 3029 1139
rect 3083 1378 3117 1412
rect 3083 1310 3117 1344
rect 3083 1242 3117 1276
rect 3083 1174 3117 1208
rect 3397 1378 3431 1412
rect 3397 1310 3431 1344
rect 3397 1242 3431 1276
rect 3397 1174 3431 1208
rect 3397 1105 3431 1139
rect 3485 1378 3519 1412
rect 3485 1310 3519 1344
rect 3485 1242 3519 1276
rect 3485 1174 3519 1208
rect 3485 1105 3519 1139
rect 3573 1378 3607 1412
rect 3573 1310 3607 1344
rect 3573 1242 3607 1276
rect 3573 1174 3607 1208
rect 3661 1378 3695 1412
rect 3661 1310 3695 1344
rect 3661 1242 3695 1276
rect 3661 1174 3695 1208
rect 3661 1105 3695 1139
rect 3749 1378 3783 1412
rect 3749 1310 3783 1344
rect 3749 1242 3783 1276
rect 3749 1174 3783 1208
rect 4123 1378 4157 1412
rect 4123 1310 4157 1344
rect 4123 1242 4157 1276
rect 4123 1174 4157 1208
rect 4123 1105 4157 1139
rect 4211 1378 4245 1412
rect 4211 1310 4245 1344
rect 4211 1242 4245 1276
rect 4211 1174 4245 1208
rect 4211 1105 4245 1139
rect 4299 1378 4333 1412
rect 4299 1310 4333 1344
rect 4299 1242 4333 1276
rect 4299 1174 4333 1208
rect 4387 1378 4421 1412
rect 4387 1310 4421 1344
rect 4387 1242 4421 1276
rect 4387 1174 4421 1208
rect 4387 1105 4421 1139
rect 4475 1378 4509 1412
rect 4475 1310 4509 1344
rect 4475 1242 4509 1276
rect 4475 1174 4509 1208
rect 4563 1378 4597 1412
rect 4563 1310 4597 1344
rect 4563 1242 4597 1276
rect 4563 1174 4597 1208
rect 4563 1105 4597 1139
rect 4651 1378 4685 1412
rect 4651 1310 4685 1344
rect 4651 1242 4685 1276
rect 4651 1174 4685 1208
rect 5025 1378 5059 1412
rect 5025 1310 5059 1344
rect 5025 1242 5059 1276
rect 5025 1174 5059 1208
rect 5025 1105 5059 1139
rect 5113 1378 5147 1412
rect 5113 1310 5147 1344
rect 5113 1242 5147 1276
rect 5113 1174 5147 1208
rect 5113 1105 5147 1139
rect 5201 1378 5235 1412
rect 5201 1310 5235 1344
rect 5201 1242 5235 1276
rect 5201 1174 5235 1208
rect 5289 1378 5323 1412
rect 5289 1310 5323 1344
rect 5289 1242 5323 1276
rect 5289 1174 5323 1208
rect 5289 1105 5323 1139
rect 5377 1378 5411 1412
rect 5377 1310 5411 1344
rect 5377 1242 5411 1276
rect 5377 1174 5411 1208
rect 5751 1378 5785 1412
rect 5751 1310 5785 1344
rect 5751 1242 5785 1276
rect 5751 1174 5785 1208
rect 5751 1105 5785 1139
rect 5839 1378 5873 1412
rect 5839 1310 5873 1344
rect 5839 1242 5873 1276
rect 5839 1174 5873 1208
rect 5839 1105 5873 1139
rect 5927 1378 5961 1412
rect 5927 1310 5961 1344
rect 5927 1242 5961 1276
rect 5927 1174 5961 1208
rect 6015 1378 6049 1412
rect 6015 1310 6049 1344
rect 6015 1242 6049 1276
rect 6015 1174 6049 1208
rect 6015 1105 6049 1139
rect 6103 1378 6137 1412
rect 6103 1310 6137 1344
rect 6103 1242 6137 1276
rect 6103 1174 6137 1208
rect 6191 1378 6225 1412
rect 6191 1310 6225 1344
rect 6191 1242 6225 1276
rect 6191 1174 6225 1208
rect 6191 1105 6225 1139
rect 6279 1378 6313 1412
rect 6279 1310 6313 1344
rect 6279 1242 6313 1276
rect 6279 1174 6313 1208
rect 6713 1378 6747 1412
rect 6713 1310 6747 1344
rect 6713 1242 6747 1276
rect 6713 1174 6747 1208
rect 6713 1105 6747 1139
rect 6801 1378 6835 1412
rect 6801 1310 6835 1344
rect 6801 1242 6835 1276
rect 6801 1174 6835 1208
rect 6801 1105 6835 1139
rect 6889 1378 6923 1412
rect 6889 1310 6923 1344
rect 6889 1242 6923 1276
rect 6889 1174 6923 1208
rect 6977 1378 7011 1412
rect 6977 1310 7011 1344
rect 6977 1242 7011 1276
rect 6977 1174 7011 1208
rect 6977 1105 7011 1139
rect 7065 1378 7099 1412
rect 7065 1310 7099 1344
rect 7065 1242 7099 1276
rect 7065 1174 7099 1208
rect 7153 1378 7187 1412
rect 7153 1310 7187 1344
rect 7153 1242 7187 1276
rect 7153 1174 7187 1208
rect 7153 1105 7187 1139
rect 7241 1378 7275 1412
rect 7241 1310 7275 1344
rect 7241 1242 7275 1276
rect 7241 1174 7275 1208
rect 7615 1378 7649 1412
rect 7615 1310 7649 1344
rect 7615 1242 7649 1276
rect 7615 1174 7649 1208
rect 7615 1105 7649 1139
rect 7703 1378 7737 1412
rect 7703 1310 7737 1344
rect 7703 1242 7737 1276
rect 7703 1174 7737 1208
rect 7703 1105 7737 1139
rect 7791 1378 7825 1412
rect 7791 1310 7825 1344
rect 7791 1242 7825 1276
rect 7791 1174 7825 1208
rect 7879 1378 7913 1412
rect 7879 1310 7913 1344
rect 7879 1242 7913 1276
rect 7879 1174 7913 1208
rect 7879 1105 7913 1139
rect 7967 1378 8001 1412
rect 7967 1310 8001 1344
rect 7967 1242 8001 1276
rect 7967 1174 8001 1208
rect 8281 1378 8315 1412
rect 8281 1310 8315 1344
rect 8281 1242 8315 1276
rect 8281 1174 8315 1208
rect 8281 1105 8315 1139
rect 8369 1378 8403 1412
rect 8369 1310 8403 1344
rect 8369 1242 8403 1276
rect 8369 1174 8403 1208
rect 8369 1105 8403 1139
rect 8457 1378 8491 1412
rect 8457 1310 8491 1344
rect 8457 1242 8491 1276
rect 8457 1174 8491 1208
rect 8545 1378 8579 1412
rect 8545 1310 8579 1344
rect 8545 1242 8579 1276
rect 8545 1174 8579 1208
rect 8545 1105 8579 1139
rect 8633 1378 8667 1412
rect 8633 1310 8667 1344
rect 8633 1242 8667 1276
rect 8633 1174 8667 1208
rect 9007 1378 9041 1412
rect 9007 1310 9041 1344
rect 9007 1242 9041 1276
rect 9007 1174 9041 1208
rect 9007 1105 9041 1139
rect 9095 1378 9129 1412
rect 9095 1310 9129 1344
rect 9095 1242 9129 1276
rect 9095 1174 9129 1208
rect 9095 1105 9129 1139
rect 9183 1378 9217 1412
rect 9183 1310 9217 1344
rect 9183 1242 9217 1276
rect 9183 1174 9217 1208
rect 9271 1378 9305 1412
rect 9271 1310 9305 1344
rect 9271 1242 9305 1276
rect 9271 1174 9305 1208
rect 9271 1105 9305 1139
rect 9359 1378 9393 1412
rect 9359 1310 9393 1344
rect 9359 1242 9393 1276
rect 9359 1174 9393 1208
rect 9447 1378 9481 1412
rect 9447 1310 9481 1344
rect 9447 1242 9481 1276
rect 9447 1174 9481 1208
rect 9447 1105 9481 1139
rect 9535 1378 9569 1412
rect 9535 1310 9569 1344
rect 9535 1242 9569 1276
rect 9535 1174 9569 1208
rect 9909 1378 9943 1412
rect 9909 1310 9943 1344
rect 9909 1242 9943 1276
rect 9909 1174 9943 1208
rect 9909 1105 9943 1139
rect 9997 1378 10031 1412
rect 9997 1310 10031 1344
rect 9997 1242 10031 1276
rect 9997 1174 10031 1208
rect 9997 1105 10031 1139
rect 10085 1378 10119 1412
rect 10085 1310 10119 1344
rect 10085 1242 10119 1276
rect 10085 1174 10119 1208
rect 10173 1378 10207 1412
rect 10173 1310 10207 1344
rect 10173 1242 10207 1276
rect 10173 1174 10207 1208
rect 10173 1105 10207 1139
rect 10261 1378 10295 1412
rect 10261 1310 10295 1344
rect 10261 1242 10295 1276
rect 10261 1174 10295 1208
rect 10635 1378 10669 1412
rect 10635 1310 10669 1344
rect 10635 1242 10669 1276
rect 10635 1174 10669 1208
rect 10635 1105 10669 1139
rect 10723 1378 10757 1412
rect 10723 1310 10757 1344
rect 10723 1242 10757 1276
rect 10723 1174 10757 1208
rect 10723 1105 10757 1139
rect 10811 1378 10845 1412
rect 10811 1310 10845 1344
rect 10811 1242 10845 1276
rect 10811 1174 10845 1208
rect 10899 1378 10933 1412
rect 10899 1310 10933 1344
rect 10899 1242 10933 1276
rect 10899 1174 10933 1208
rect 10899 1105 10933 1139
rect 10987 1378 11021 1412
rect 10987 1310 11021 1344
rect 10987 1242 11021 1276
rect 10987 1174 11021 1208
rect 11075 1378 11109 1412
rect 11075 1310 11109 1344
rect 11075 1242 11109 1276
rect 11075 1174 11109 1208
rect 11075 1105 11109 1139
rect 11163 1378 11197 1412
rect 11163 1310 11197 1344
rect 11163 1242 11197 1276
rect 11163 1174 11197 1208
rect 11597 1378 11631 1412
rect 11597 1310 11631 1344
rect 11597 1242 11631 1276
rect 11597 1174 11631 1208
rect 11597 1105 11631 1139
rect 11685 1378 11719 1412
rect 11685 1310 11719 1344
rect 11685 1242 11719 1276
rect 11685 1174 11719 1208
rect 11685 1105 11719 1139
rect 11773 1378 11807 1412
rect 11773 1310 11807 1344
rect 11773 1242 11807 1276
rect 11773 1174 11807 1208
rect 11861 1378 11895 1412
rect 11861 1310 11895 1344
rect 11861 1242 11895 1276
rect 11861 1174 11895 1208
rect 11861 1105 11895 1139
rect 11949 1378 11983 1412
rect 11949 1310 11983 1344
rect 11949 1242 11983 1276
rect 11949 1174 11983 1208
rect 12037 1378 12071 1412
rect 12037 1310 12071 1344
rect 12037 1242 12071 1276
rect 12037 1174 12071 1208
rect 12037 1105 12071 1139
rect 12125 1378 12159 1412
rect 12125 1310 12159 1344
rect 12125 1242 12159 1276
rect 12125 1174 12159 1208
rect 12499 1378 12533 1412
rect 12499 1310 12533 1344
rect 12499 1242 12533 1276
rect 12499 1174 12533 1208
rect 12499 1105 12533 1139
rect 12587 1378 12621 1412
rect 12587 1310 12621 1344
rect 12587 1242 12621 1276
rect 12587 1174 12621 1208
rect 12587 1105 12621 1139
rect 12675 1378 12709 1412
rect 12675 1310 12709 1344
rect 12675 1242 12709 1276
rect 12675 1174 12709 1208
rect 12763 1378 12797 1412
rect 12763 1310 12797 1344
rect 12763 1242 12797 1276
rect 12763 1174 12797 1208
rect 12763 1105 12797 1139
rect 12851 1378 12885 1412
rect 12851 1310 12885 1344
rect 12851 1242 12885 1276
rect 12851 1174 12885 1208
rect 13165 1378 13199 1412
rect 13165 1310 13199 1344
rect 13165 1242 13199 1276
rect 13165 1174 13199 1208
rect 13165 1105 13199 1139
rect 13253 1378 13287 1412
rect 13253 1310 13287 1344
rect 13253 1242 13287 1276
rect 13253 1174 13287 1208
rect 13253 1105 13287 1139
rect 13341 1378 13375 1412
rect 13341 1310 13375 1344
rect 13341 1242 13375 1276
rect 13341 1174 13375 1208
rect 13429 1378 13463 1412
rect 13429 1310 13463 1344
rect 13429 1242 13463 1276
rect 13429 1174 13463 1208
rect 13429 1105 13463 1139
rect 13517 1378 13551 1412
rect 13517 1310 13551 1344
rect 13517 1242 13551 1276
rect 13517 1174 13551 1208
rect 13891 1378 13925 1412
rect 13891 1310 13925 1344
rect 13891 1242 13925 1276
rect 13891 1174 13925 1208
rect 13891 1105 13925 1139
rect 13979 1378 14013 1412
rect 13979 1310 14013 1344
rect 13979 1242 14013 1276
rect 13979 1174 14013 1208
rect 13979 1105 14013 1139
rect 14067 1378 14101 1412
rect 14067 1310 14101 1344
rect 14067 1242 14101 1276
rect 14067 1174 14101 1208
rect 14155 1378 14189 1412
rect 14155 1310 14189 1344
rect 14155 1242 14189 1276
rect 14155 1174 14189 1208
rect 14155 1105 14189 1139
rect 14243 1378 14277 1412
rect 14243 1310 14277 1344
rect 14243 1242 14277 1276
rect 14243 1174 14277 1208
rect 14331 1378 14365 1412
rect 14331 1310 14365 1344
rect 14331 1242 14365 1276
rect 14331 1174 14365 1208
rect 14331 1105 14365 1139
rect 14419 1378 14453 1412
rect 14419 1310 14453 1344
rect 14419 1242 14453 1276
rect 14419 1174 14453 1208
rect 14793 1377 14827 1411
rect 14793 1309 14827 1343
rect 14793 1241 14827 1275
rect 14793 1173 14827 1207
rect 14793 1105 14827 1139
rect 14881 1377 14915 1411
rect 14881 1309 14915 1343
rect 14881 1241 14915 1275
rect 14881 1173 14915 1207
rect 14881 1105 14915 1139
rect 14969 1377 15003 1411
rect 14969 1309 15003 1343
rect 14969 1241 15003 1275
rect 14969 1173 15003 1207
rect 15057 1377 15091 1411
rect 15057 1309 15091 1343
rect 15057 1241 15091 1275
rect 15057 1173 15091 1207
rect 15145 1377 15179 1411
rect 15145 1309 15179 1343
rect 15145 1241 15179 1275
rect 15145 1173 15179 1207
rect 15145 1105 15179 1139
rect 15457 1377 15491 1411
rect 15457 1309 15491 1343
rect 15457 1241 15491 1275
rect 15457 1173 15491 1207
rect 15545 1309 15579 1343
rect 15545 1241 15579 1275
rect 15545 1173 15579 1207
rect 15545 1105 15579 1139
rect 15633 1377 15667 1411
rect 15633 1309 15667 1343
rect 15633 1241 15667 1275
rect 15633 1173 15667 1207
rect 15721 1309 15755 1343
rect 15721 1241 15755 1275
rect 15721 1173 15755 1207
rect 15809 1377 15843 1411
rect 15809 1309 15843 1343
rect 15809 1241 15843 1275
rect 15809 1173 15843 1207
rect 16125 1377 16159 1411
rect 16125 1309 16159 1343
rect 16125 1241 16159 1275
rect 16125 1173 16159 1207
rect 16213 1309 16247 1343
rect 16213 1241 16247 1275
rect 16213 1173 16247 1207
rect 16213 1105 16247 1139
rect 16301 1377 16335 1411
rect 16301 1309 16335 1343
rect 16301 1241 16335 1275
rect 16301 1173 16335 1207
rect 16389 1309 16423 1343
rect 16389 1241 16423 1275
rect 16389 1173 16423 1207
rect 16389 1105 16423 1139
rect 16477 1377 16511 1411
rect 16477 1309 16511 1343
rect 16477 1241 16511 1275
rect 16477 1173 16511 1207
<< psubdiff >>
rect -31 546 16681 572
rect -31 512 -17 546
rect 17 512 649 546
rect 683 512 1611 546
rect 1645 512 2573 546
rect 2607 512 3239 546
rect 3273 512 3905 546
rect 3939 512 4867 546
rect 4901 512 5533 546
rect 5567 512 6495 546
rect 6529 512 7457 546
rect 7491 512 8123 546
rect 8157 512 8789 546
rect 8823 512 9751 546
rect 9785 512 10417 546
rect 10451 512 11379 546
rect 11413 512 12341 546
rect 12375 512 13007 546
rect 13041 512 13673 546
rect 13707 512 14635 546
rect 14669 512 15301 546
rect 15335 512 15967 546
rect 16001 512 16633 546
rect 16667 512 16681 546
rect -31 510 16681 512
rect -31 474 31 510
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect -31 368 -17 402
rect 17 368 31 402
rect 635 474 697 510
rect 635 440 649 474
rect 683 440 697 474
rect 635 402 697 440
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect 635 368 649 402
rect 683 368 697 402
rect 1597 474 1659 510
rect 1597 440 1611 474
rect 1645 440 1659 474
rect 1597 402 1659 440
rect 635 330 697 368
rect 635 296 649 330
rect 683 296 697 330
rect 635 258 697 296
rect 635 224 649 258
rect 683 224 697 258
rect 635 186 697 224
rect 635 152 649 186
rect 683 152 697 186
rect 635 114 697 152
rect -31 47 31 80
rect 635 80 649 114
rect 683 80 697 114
rect 1597 368 1611 402
rect 1645 368 1659 402
rect 2559 474 2621 510
rect 2559 440 2573 474
rect 2607 440 2621 474
rect 2559 402 2621 440
rect 1597 330 1659 368
rect 1597 296 1611 330
rect 1645 296 1659 330
rect 1597 258 1659 296
rect 1597 224 1611 258
rect 1645 224 1659 258
rect 1597 186 1659 224
rect 1597 152 1611 186
rect 1645 152 1659 186
rect 1597 114 1659 152
rect 635 47 697 80
rect 1597 80 1611 114
rect 1645 80 1659 114
rect 2559 368 2573 402
rect 2607 368 2621 402
rect 3225 474 3287 510
rect 3225 440 3239 474
rect 3273 440 3287 474
rect 3225 402 3287 440
rect 2559 330 2621 368
rect 2559 296 2573 330
rect 2607 296 2621 330
rect 2559 258 2621 296
rect 2559 224 2573 258
rect 2607 224 2621 258
rect 2559 186 2621 224
rect 2559 152 2573 186
rect 2607 152 2621 186
rect 2559 114 2621 152
rect 1597 47 1659 80
rect 2559 80 2573 114
rect 2607 80 2621 114
rect 3225 368 3239 402
rect 3273 368 3287 402
rect 3891 474 3953 510
rect 3891 440 3905 474
rect 3939 440 3953 474
rect 3891 402 3953 440
rect 3225 330 3287 368
rect 3225 296 3239 330
rect 3273 296 3287 330
rect 3225 258 3287 296
rect 3225 224 3239 258
rect 3273 224 3287 258
rect 3225 186 3287 224
rect 3225 152 3239 186
rect 3273 152 3287 186
rect 3225 114 3287 152
rect 2559 47 2621 80
rect 3225 80 3239 114
rect 3273 80 3287 114
rect 3891 368 3905 402
rect 3939 368 3953 402
rect 4853 474 4915 510
rect 4853 440 4867 474
rect 4901 440 4915 474
rect 4853 402 4915 440
rect 3891 330 3953 368
rect 3891 296 3905 330
rect 3939 296 3953 330
rect 3891 258 3953 296
rect 3891 224 3905 258
rect 3939 224 3953 258
rect 3891 186 3953 224
rect 3891 152 3905 186
rect 3939 152 3953 186
rect 3891 114 3953 152
rect 3225 47 3287 80
rect 3891 80 3905 114
rect 3939 80 3953 114
rect 4853 368 4867 402
rect 4901 368 4915 402
rect 5519 474 5581 510
rect 5519 440 5533 474
rect 5567 440 5581 474
rect 5519 402 5581 440
rect 4853 330 4915 368
rect 4853 296 4867 330
rect 4901 296 4915 330
rect 4853 258 4915 296
rect 4853 224 4867 258
rect 4901 224 4915 258
rect 4853 186 4915 224
rect 4853 152 4867 186
rect 4901 152 4915 186
rect 4853 114 4915 152
rect 3891 47 3953 80
rect 4853 80 4867 114
rect 4901 80 4915 114
rect 5519 368 5533 402
rect 5567 368 5581 402
rect 6481 474 6543 510
rect 6481 440 6495 474
rect 6529 440 6543 474
rect 6481 402 6543 440
rect 5519 330 5581 368
rect 5519 296 5533 330
rect 5567 296 5581 330
rect 5519 258 5581 296
rect 5519 224 5533 258
rect 5567 224 5581 258
rect 5519 186 5581 224
rect 5519 152 5533 186
rect 5567 152 5581 186
rect 5519 114 5581 152
rect 4853 47 4915 80
rect 5519 80 5533 114
rect 5567 80 5581 114
rect 6481 368 6495 402
rect 6529 368 6543 402
rect 7443 474 7505 510
rect 7443 440 7457 474
rect 7491 440 7505 474
rect 7443 402 7505 440
rect 6481 330 6543 368
rect 6481 296 6495 330
rect 6529 296 6543 330
rect 6481 258 6543 296
rect 6481 224 6495 258
rect 6529 224 6543 258
rect 6481 186 6543 224
rect 6481 152 6495 186
rect 6529 152 6543 186
rect 6481 114 6543 152
rect 5519 47 5581 80
rect 6481 80 6495 114
rect 6529 80 6543 114
rect 7443 368 7457 402
rect 7491 368 7505 402
rect 8109 474 8171 510
rect 8109 440 8123 474
rect 8157 440 8171 474
rect 8109 402 8171 440
rect 7443 330 7505 368
rect 7443 296 7457 330
rect 7491 296 7505 330
rect 7443 258 7505 296
rect 7443 224 7457 258
rect 7491 224 7505 258
rect 7443 186 7505 224
rect 7443 152 7457 186
rect 7491 152 7505 186
rect 7443 114 7505 152
rect 6481 47 6543 80
rect 7443 80 7457 114
rect 7491 80 7505 114
rect 8109 368 8123 402
rect 8157 368 8171 402
rect 8775 474 8837 510
rect 8775 440 8789 474
rect 8823 440 8837 474
rect 8775 402 8837 440
rect 8109 330 8171 368
rect 8109 296 8123 330
rect 8157 296 8171 330
rect 8109 258 8171 296
rect 8109 224 8123 258
rect 8157 224 8171 258
rect 8109 186 8171 224
rect 8109 152 8123 186
rect 8157 152 8171 186
rect 8109 114 8171 152
rect 7443 47 7505 80
rect 8109 80 8123 114
rect 8157 80 8171 114
rect 8775 368 8789 402
rect 8823 368 8837 402
rect 9737 474 9799 510
rect 9737 440 9751 474
rect 9785 440 9799 474
rect 9737 402 9799 440
rect 8775 330 8837 368
rect 8775 296 8789 330
rect 8823 296 8837 330
rect 8775 258 8837 296
rect 8775 224 8789 258
rect 8823 224 8837 258
rect 8775 186 8837 224
rect 8775 152 8789 186
rect 8823 152 8837 186
rect 8775 114 8837 152
rect 8109 47 8171 80
rect 8775 80 8789 114
rect 8823 80 8837 114
rect 9737 368 9751 402
rect 9785 368 9799 402
rect 10403 474 10465 510
rect 10403 440 10417 474
rect 10451 440 10465 474
rect 10403 402 10465 440
rect 9737 330 9799 368
rect 9737 296 9751 330
rect 9785 296 9799 330
rect 9737 258 9799 296
rect 9737 224 9751 258
rect 9785 224 9799 258
rect 9737 186 9799 224
rect 9737 152 9751 186
rect 9785 152 9799 186
rect 9737 114 9799 152
rect 8775 47 8837 80
rect 9737 80 9751 114
rect 9785 80 9799 114
rect 10403 368 10417 402
rect 10451 368 10465 402
rect 11365 474 11427 510
rect 11365 440 11379 474
rect 11413 440 11427 474
rect 11365 402 11427 440
rect 10403 330 10465 368
rect 10403 296 10417 330
rect 10451 296 10465 330
rect 10403 258 10465 296
rect 10403 224 10417 258
rect 10451 224 10465 258
rect 10403 186 10465 224
rect 10403 152 10417 186
rect 10451 152 10465 186
rect 10403 114 10465 152
rect 9737 47 9799 80
rect 10403 80 10417 114
rect 10451 80 10465 114
rect 11365 368 11379 402
rect 11413 368 11427 402
rect 12327 474 12389 510
rect 12327 440 12341 474
rect 12375 440 12389 474
rect 12327 402 12389 440
rect 11365 330 11427 368
rect 11365 296 11379 330
rect 11413 296 11427 330
rect 11365 258 11427 296
rect 11365 224 11379 258
rect 11413 224 11427 258
rect 11365 186 11427 224
rect 11365 152 11379 186
rect 11413 152 11427 186
rect 11365 114 11427 152
rect 10403 47 10465 80
rect 11365 80 11379 114
rect 11413 80 11427 114
rect 12327 368 12341 402
rect 12375 368 12389 402
rect 12993 474 13055 510
rect 12993 440 13007 474
rect 13041 440 13055 474
rect 12993 402 13055 440
rect 12327 330 12389 368
rect 12327 296 12341 330
rect 12375 296 12389 330
rect 12327 258 12389 296
rect 12327 224 12341 258
rect 12375 224 12389 258
rect 12327 186 12389 224
rect 12327 152 12341 186
rect 12375 152 12389 186
rect 12327 114 12389 152
rect 11365 47 11427 80
rect 12327 80 12341 114
rect 12375 80 12389 114
rect 12993 368 13007 402
rect 13041 368 13055 402
rect 13659 474 13721 510
rect 13659 440 13673 474
rect 13707 440 13721 474
rect 13659 402 13721 440
rect 12993 330 13055 368
rect 12993 296 13007 330
rect 13041 296 13055 330
rect 12993 258 13055 296
rect 12993 224 13007 258
rect 13041 224 13055 258
rect 12993 186 13055 224
rect 12993 152 13007 186
rect 13041 152 13055 186
rect 12993 114 13055 152
rect 12327 47 12389 80
rect 12993 80 13007 114
rect 13041 80 13055 114
rect 13659 368 13673 402
rect 13707 368 13721 402
rect 14621 474 14683 510
rect 14621 440 14635 474
rect 14669 440 14683 474
rect 14621 402 14683 440
rect 15287 474 15349 510
rect 15287 440 15301 474
rect 15335 440 15349 474
rect 13659 330 13721 368
rect 13659 296 13673 330
rect 13707 296 13721 330
rect 13659 258 13721 296
rect 13659 224 13673 258
rect 13707 224 13721 258
rect 13659 186 13721 224
rect 13659 152 13673 186
rect 13707 152 13721 186
rect 13659 114 13721 152
rect 12993 47 13055 80
rect 13659 80 13673 114
rect 13707 80 13721 114
rect 14621 368 14635 402
rect 14669 368 14683 402
rect 15287 402 15349 440
rect 14621 330 14683 368
rect 14621 296 14635 330
rect 14669 296 14683 330
rect 14621 258 14683 296
rect 14621 224 14635 258
rect 14669 224 14683 258
rect 14621 186 14683 224
rect 14621 152 14635 186
rect 14669 152 14683 186
rect 14621 114 14683 152
rect 13659 47 13721 80
rect 14621 80 14635 114
rect 14669 80 14683 114
rect 15287 368 15301 402
rect 15335 368 15349 402
rect 15953 474 16015 510
rect 15953 440 15967 474
rect 16001 440 16015 474
rect 15953 402 16015 440
rect 16619 474 16681 510
rect 16619 440 16633 474
rect 16667 440 16681 474
rect 15287 330 15349 368
rect 15287 296 15301 330
rect 15335 296 15349 330
rect 15287 258 15349 296
rect 15287 224 15301 258
rect 15335 224 15349 258
rect 15287 186 15349 224
rect 15287 152 15301 186
rect 15335 152 15349 186
rect 15287 114 15349 152
rect 14621 47 14683 80
rect 15287 80 15301 114
rect 15335 80 15349 114
rect 15953 368 15967 402
rect 16001 368 16015 402
rect 16619 402 16681 440
rect 15953 330 16015 368
rect 15953 296 15967 330
rect 16001 296 16015 330
rect 15953 258 16015 296
rect 15953 224 15967 258
rect 16001 224 16015 258
rect 15953 186 16015 224
rect 15953 152 15967 186
rect 16001 152 16015 186
rect 15953 114 16015 152
rect 15287 47 15349 80
rect 15953 80 15967 114
rect 16001 80 16015 114
rect 16619 368 16633 402
rect 16667 368 16681 402
rect 16619 330 16681 368
rect 16619 296 16633 330
rect 16667 296 16681 330
rect 16619 258 16681 296
rect 16619 224 16633 258
rect 16667 224 16681 258
rect 16619 186 16681 224
rect 16619 152 16633 186
rect 16667 152 16681 186
rect 16619 114 16681 152
rect 15953 47 16015 80
rect 16619 80 16633 114
rect 16667 80 16681 114
rect 16619 47 16681 80
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 361 47
rect 395 13 433 47
rect 467 13 505 47
rect 539 13 577 47
rect 611 13 721 47
rect 755 13 793 47
rect 827 13 865 47
rect 899 13 937 47
rect 971 13 1009 47
rect 1043 13 1081 47
rect 1115 13 1179 47
rect 1213 13 1251 47
rect 1285 13 1323 47
rect 1357 13 1395 47
rect 1429 13 1467 47
rect 1501 13 1539 47
rect 1573 13 1683 47
rect 1717 13 1755 47
rect 1789 13 1827 47
rect 1861 13 1899 47
rect 1933 13 1971 47
rect 2005 13 2043 47
rect 2077 13 2141 47
rect 2175 13 2213 47
rect 2247 13 2285 47
rect 2319 13 2357 47
rect 2391 13 2429 47
rect 2463 13 2501 47
rect 2535 13 2645 47
rect 2679 13 2717 47
rect 2751 13 2789 47
rect 2823 13 2861 47
rect 2895 13 2951 47
rect 2985 13 3023 47
rect 3057 13 3095 47
rect 3129 13 3167 47
rect 3201 13 3311 47
rect 3345 13 3383 47
rect 3417 13 3455 47
rect 3489 13 3527 47
rect 3561 13 3617 47
rect 3651 13 3689 47
rect 3723 13 3761 47
rect 3795 13 3833 47
rect 3867 13 3977 47
rect 4011 13 4049 47
rect 4083 13 4121 47
rect 4155 13 4193 47
rect 4227 13 4265 47
rect 4299 13 4337 47
rect 4371 13 4435 47
rect 4469 13 4507 47
rect 4541 13 4579 47
rect 4613 13 4651 47
rect 4685 13 4723 47
rect 4757 13 4795 47
rect 4829 13 4939 47
rect 4973 13 5011 47
rect 5045 13 5083 47
rect 5117 13 5155 47
rect 5189 13 5245 47
rect 5279 13 5317 47
rect 5351 13 5389 47
rect 5423 13 5461 47
rect 5495 13 5605 47
rect 5639 13 5677 47
rect 5711 13 5749 47
rect 5783 13 5821 47
rect 5855 13 5893 47
rect 5927 13 5965 47
rect 5999 13 6063 47
rect 6097 13 6135 47
rect 6169 13 6207 47
rect 6241 13 6279 47
rect 6313 13 6351 47
rect 6385 13 6423 47
rect 6457 13 6567 47
rect 6601 13 6639 47
rect 6673 13 6711 47
rect 6745 13 6783 47
rect 6817 13 6855 47
rect 6889 13 6927 47
rect 6961 13 7025 47
rect 7059 13 7097 47
rect 7131 13 7169 47
rect 7203 13 7241 47
rect 7275 13 7313 47
rect 7347 13 7385 47
rect 7419 13 7529 47
rect 7563 13 7601 47
rect 7635 13 7673 47
rect 7707 13 7745 47
rect 7779 13 7835 47
rect 7869 13 7907 47
rect 7941 13 7979 47
rect 8013 13 8051 47
rect 8085 13 8195 47
rect 8229 13 8267 47
rect 8301 13 8339 47
rect 8373 13 8411 47
rect 8445 13 8501 47
rect 8535 13 8573 47
rect 8607 13 8645 47
rect 8679 13 8717 47
rect 8751 13 8861 47
rect 8895 13 8933 47
rect 8967 13 9005 47
rect 9039 13 9077 47
rect 9111 13 9149 47
rect 9183 13 9221 47
rect 9255 13 9319 47
rect 9353 13 9391 47
rect 9425 13 9463 47
rect 9497 13 9535 47
rect 9569 13 9607 47
rect 9641 13 9679 47
rect 9713 13 9823 47
rect 9857 13 9895 47
rect 9929 13 9967 47
rect 10001 13 10039 47
rect 10073 13 10129 47
rect 10163 13 10201 47
rect 10235 13 10273 47
rect 10307 13 10345 47
rect 10379 13 10489 47
rect 10523 13 10561 47
rect 10595 13 10633 47
rect 10667 13 10705 47
rect 10739 13 10777 47
rect 10811 13 10849 47
rect 10883 13 10947 47
rect 10981 13 11019 47
rect 11053 13 11091 47
rect 11125 13 11163 47
rect 11197 13 11235 47
rect 11269 13 11307 47
rect 11341 13 11451 47
rect 11485 13 11523 47
rect 11557 13 11595 47
rect 11629 13 11667 47
rect 11701 13 11739 47
rect 11773 13 11811 47
rect 11845 13 11909 47
rect 11943 13 11981 47
rect 12015 13 12053 47
rect 12087 13 12125 47
rect 12159 13 12197 47
rect 12231 13 12269 47
rect 12303 13 12413 47
rect 12447 13 12485 47
rect 12519 13 12557 47
rect 12591 13 12629 47
rect 12663 13 12719 47
rect 12753 13 12791 47
rect 12825 13 12863 47
rect 12897 13 12935 47
rect 12969 13 13079 47
rect 13113 13 13151 47
rect 13185 13 13223 47
rect 13257 13 13295 47
rect 13329 13 13385 47
rect 13419 13 13457 47
rect 13491 13 13529 47
rect 13563 13 13601 47
rect 13635 13 13745 47
rect 13779 13 13817 47
rect 13851 13 13889 47
rect 13923 13 13961 47
rect 13995 13 14033 47
rect 14067 13 14105 47
rect 14139 13 14203 47
rect 14237 13 14275 47
rect 14309 13 14347 47
rect 14381 13 14419 47
rect 14453 13 14491 47
rect 14525 13 14563 47
rect 14597 13 14707 47
rect 14741 13 14779 47
rect 14813 13 14851 47
rect 14885 13 14923 47
rect 14957 13 15013 47
rect 15047 13 15085 47
rect 15119 13 15157 47
rect 15191 13 15229 47
rect 15263 13 15373 47
rect 15407 13 15445 47
rect 15479 13 15517 47
rect 15551 13 15589 47
rect 15623 13 15679 47
rect 15713 13 15751 47
rect 15785 13 15823 47
rect 15857 13 15895 47
rect 15929 13 16039 47
rect 16073 13 16111 47
rect 16145 13 16183 47
rect 16217 13 16255 47
rect 16289 13 16345 47
rect 16379 13 16417 47
rect 16451 13 16489 47
rect 16523 13 16561 47
rect 16595 13 16681 47
rect -31 11 31 13
rect 635 11 697 13
rect 1597 11 1659 13
rect 2559 11 2621 13
rect 3225 11 3287 13
rect 3891 11 3953 13
rect 4853 11 4915 13
rect 5519 11 5581 13
rect 6481 11 6543 13
rect 7443 11 7505 13
rect 8109 11 8171 13
rect 8775 11 8837 13
rect 9737 11 9799 13
rect 10403 11 10465 13
rect 11365 11 11427 13
rect 12327 11 12389 13
rect 12993 11 13055 13
rect 13659 11 13721 13
rect 14621 11 14683 13
rect 15287 11 15349 13
rect 15953 11 16015 13
rect 16619 11 16681 13
<< nsubdiff >>
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 361 1539
rect 395 1505 433 1539
rect 467 1505 505 1539
rect 539 1505 577 1539
rect 611 1505 721 1539
rect 755 1505 793 1539
rect 827 1505 865 1539
rect 899 1505 937 1539
rect 971 1505 1009 1539
rect 1043 1505 1081 1539
rect 1115 1505 1179 1539
rect 1213 1505 1251 1539
rect 1285 1505 1323 1539
rect 1357 1505 1395 1539
rect 1429 1505 1467 1539
rect 1501 1505 1539 1539
rect 1573 1505 1683 1539
rect 1717 1505 1755 1539
rect 1789 1505 1827 1539
rect 1861 1505 1899 1539
rect 1933 1505 1971 1539
rect 2005 1505 2043 1539
rect 2077 1505 2141 1539
rect 2175 1505 2213 1539
rect 2247 1505 2285 1539
rect 2319 1505 2357 1539
rect 2391 1505 2429 1539
rect 2463 1505 2501 1539
rect 2535 1505 2645 1539
rect 2679 1505 2717 1539
rect 2751 1505 2789 1539
rect 2823 1505 2861 1539
rect 2895 1505 2951 1539
rect 2985 1505 3023 1539
rect 3057 1505 3095 1539
rect 3129 1505 3167 1539
rect 3201 1505 3311 1539
rect 3345 1505 3383 1539
rect 3417 1505 3455 1539
rect 3489 1505 3527 1539
rect 3561 1505 3617 1539
rect 3651 1505 3689 1539
rect 3723 1505 3761 1539
rect 3795 1505 3833 1539
rect 3867 1505 3977 1539
rect 4011 1505 4049 1539
rect 4083 1505 4121 1539
rect 4155 1505 4193 1539
rect 4227 1505 4265 1539
rect 4299 1505 4337 1539
rect 4371 1505 4435 1539
rect 4469 1505 4507 1539
rect 4541 1505 4579 1539
rect 4613 1505 4651 1539
rect 4685 1505 4723 1539
rect 4757 1505 4795 1539
rect 4829 1505 4939 1539
rect 4973 1505 5011 1539
rect 5045 1505 5083 1539
rect 5117 1505 5155 1539
rect 5189 1505 5245 1539
rect 5279 1505 5317 1539
rect 5351 1505 5389 1539
rect 5423 1505 5461 1539
rect 5495 1505 5605 1539
rect 5639 1505 5677 1539
rect 5711 1505 5749 1539
rect 5783 1505 5821 1539
rect 5855 1505 5893 1539
rect 5927 1505 5965 1539
rect 5999 1505 6063 1539
rect 6097 1505 6135 1539
rect 6169 1505 6207 1539
rect 6241 1505 6279 1539
rect 6313 1505 6351 1539
rect 6385 1505 6423 1539
rect 6457 1505 6567 1539
rect 6601 1505 6639 1539
rect 6673 1505 6711 1539
rect 6745 1505 6783 1539
rect 6817 1505 6855 1539
rect 6889 1505 6927 1539
rect 6961 1505 7025 1539
rect 7059 1505 7097 1539
rect 7131 1505 7169 1539
rect 7203 1505 7241 1539
rect 7275 1505 7313 1539
rect 7347 1505 7385 1539
rect 7419 1505 7529 1539
rect 7563 1505 7601 1539
rect 7635 1505 7673 1539
rect 7707 1505 7745 1539
rect 7779 1505 7835 1539
rect 7869 1505 7907 1539
rect 7941 1505 7979 1539
rect 8013 1505 8051 1539
rect 8085 1505 8195 1539
rect 8229 1505 8267 1539
rect 8301 1505 8339 1539
rect 8373 1505 8411 1539
rect 8445 1505 8501 1539
rect 8535 1505 8573 1539
rect 8607 1505 8645 1539
rect 8679 1505 8717 1539
rect 8751 1505 8861 1539
rect 8895 1505 8933 1539
rect 8967 1505 9005 1539
rect 9039 1505 9077 1539
rect 9111 1505 9149 1539
rect 9183 1505 9221 1539
rect 9255 1505 9319 1539
rect 9353 1505 9391 1539
rect 9425 1505 9463 1539
rect 9497 1505 9535 1539
rect 9569 1505 9607 1539
rect 9641 1505 9679 1539
rect 9713 1505 9823 1539
rect 9857 1505 9895 1539
rect 9929 1505 9967 1539
rect 10001 1505 10039 1539
rect 10073 1505 10129 1539
rect 10163 1505 10201 1539
rect 10235 1505 10273 1539
rect 10307 1505 10345 1539
rect 10379 1505 10489 1539
rect 10523 1505 10561 1539
rect 10595 1505 10633 1539
rect 10667 1505 10705 1539
rect 10739 1505 10777 1539
rect 10811 1505 10849 1539
rect 10883 1505 10947 1539
rect 10981 1505 11019 1539
rect 11053 1505 11091 1539
rect 11125 1505 11163 1539
rect 11197 1505 11235 1539
rect 11269 1505 11307 1539
rect 11341 1505 11451 1539
rect 11485 1505 11523 1539
rect 11557 1505 11595 1539
rect 11629 1505 11667 1539
rect 11701 1505 11739 1539
rect 11773 1505 11811 1539
rect 11845 1505 11909 1539
rect 11943 1505 11981 1539
rect 12015 1505 12053 1539
rect 12087 1505 12125 1539
rect 12159 1505 12197 1539
rect 12231 1505 12269 1539
rect 12303 1505 12413 1539
rect 12447 1505 12485 1539
rect 12519 1505 12557 1539
rect 12591 1505 12629 1539
rect 12663 1505 12719 1539
rect 12753 1505 12791 1539
rect 12825 1505 12863 1539
rect 12897 1505 12935 1539
rect 12969 1505 13079 1539
rect 13113 1505 13151 1539
rect 13185 1505 13223 1539
rect 13257 1505 13295 1539
rect 13329 1505 13385 1539
rect 13419 1505 13457 1539
rect 13491 1505 13529 1539
rect 13563 1505 13601 1539
rect 13635 1505 13745 1539
rect 13779 1505 13817 1539
rect 13851 1505 13889 1539
rect 13923 1505 13961 1539
rect 13995 1505 14033 1539
rect 14067 1505 14105 1539
rect 14139 1505 14203 1539
rect 14237 1505 14275 1539
rect 14309 1505 14347 1539
rect 14381 1505 14419 1539
rect 14453 1505 14491 1539
rect 14525 1505 14563 1539
rect 14597 1505 14707 1539
rect 14741 1505 14779 1539
rect 14813 1505 14851 1539
rect 14885 1505 14923 1539
rect 14957 1505 15013 1539
rect 15047 1505 15085 1539
rect 15119 1505 15157 1539
rect 15191 1505 15229 1539
rect 15263 1505 15373 1539
rect 15407 1505 15445 1539
rect 15479 1505 15517 1539
rect 15551 1505 15589 1539
rect 15623 1505 15679 1539
rect 15713 1505 15751 1539
rect 15785 1505 15823 1539
rect 15857 1505 15895 1539
rect 15929 1505 16039 1539
rect 16073 1505 16111 1539
rect 16145 1505 16183 1539
rect 16217 1505 16255 1539
rect 16289 1505 16345 1539
rect 16379 1505 16417 1539
rect 16451 1505 16489 1539
rect 16523 1505 16561 1539
rect 16595 1505 16681 1539
rect -31 1470 31 1505
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect 635 1470 697 1505
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect -31 1038 31 1076
rect 635 1436 649 1470
rect 683 1436 697 1470
rect 1597 1470 1659 1505
rect 635 1398 697 1436
rect 635 1364 649 1398
rect 683 1364 697 1398
rect 635 1326 697 1364
rect 635 1292 649 1326
rect 683 1292 697 1326
rect 635 1254 697 1292
rect 635 1220 649 1254
rect 683 1220 697 1254
rect 635 1182 697 1220
rect 635 1148 649 1182
rect 683 1148 697 1182
rect 635 1110 697 1148
rect 635 1076 649 1110
rect 683 1076 697 1110
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect 635 1038 697 1076
rect 1597 1436 1611 1470
rect 1645 1436 1659 1470
rect 2559 1470 2621 1505
rect 1597 1398 1659 1436
rect 1597 1364 1611 1398
rect 1645 1364 1659 1398
rect 1597 1326 1659 1364
rect 1597 1292 1611 1326
rect 1645 1292 1659 1326
rect 1597 1254 1659 1292
rect 1597 1220 1611 1254
rect 1645 1220 1659 1254
rect 1597 1182 1659 1220
rect 1597 1148 1611 1182
rect 1645 1148 1659 1182
rect 1597 1110 1659 1148
rect 1597 1076 1611 1110
rect 1645 1076 1659 1110
rect 635 1004 649 1038
rect 683 1004 697 1038
rect 635 966 697 1004
rect -31 930 31 932
rect 635 932 649 966
rect 683 932 697 966
rect 1597 1038 1659 1076
rect 2559 1436 2573 1470
rect 2607 1436 2621 1470
rect 3225 1470 3287 1505
rect 2559 1398 2621 1436
rect 2559 1364 2573 1398
rect 2607 1364 2621 1398
rect 2559 1326 2621 1364
rect 2559 1292 2573 1326
rect 2607 1292 2621 1326
rect 2559 1254 2621 1292
rect 2559 1220 2573 1254
rect 2607 1220 2621 1254
rect 2559 1182 2621 1220
rect 2559 1148 2573 1182
rect 2607 1148 2621 1182
rect 2559 1110 2621 1148
rect 2559 1076 2573 1110
rect 2607 1076 2621 1110
rect 1597 1004 1611 1038
rect 1645 1004 1659 1038
rect 1597 966 1659 1004
rect 635 930 697 932
rect 1597 932 1611 966
rect 1645 932 1659 966
rect 2559 1038 2621 1076
rect 3225 1436 3239 1470
rect 3273 1436 3287 1470
rect 3891 1470 3953 1505
rect 3225 1398 3287 1436
rect 3225 1364 3239 1398
rect 3273 1364 3287 1398
rect 3225 1326 3287 1364
rect 3225 1292 3239 1326
rect 3273 1292 3287 1326
rect 3225 1254 3287 1292
rect 3225 1220 3239 1254
rect 3273 1220 3287 1254
rect 3225 1182 3287 1220
rect 3225 1148 3239 1182
rect 3273 1148 3287 1182
rect 3225 1110 3287 1148
rect 3225 1076 3239 1110
rect 3273 1076 3287 1110
rect 2559 1004 2573 1038
rect 2607 1004 2621 1038
rect 2559 966 2621 1004
rect 1597 930 1659 932
rect 2559 932 2573 966
rect 2607 932 2621 966
rect 3225 1038 3287 1076
rect 3891 1436 3905 1470
rect 3939 1436 3953 1470
rect 4853 1470 4915 1505
rect 3891 1398 3953 1436
rect 3891 1364 3905 1398
rect 3939 1364 3953 1398
rect 3891 1326 3953 1364
rect 3891 1292 3905 1326
rect 3939 1292 3953 1326
rect 3891 1254 3953 1292
rect 3891 1220 3905 1254
rect 3939 1220 3953 1254
rect 3891 1182 3953 1220
rect 3891 1148 3905 1182
rect 3939 1148 3953 1182
rect 3891 1110 3953 1148
rect 3891 1076 3905 1110
rect 3939 1076 3953 1110
rect 3225 1004 3239 1038
rect 3273 1004 3287 1038
rect 3225 966 3287 1004
rect 2559 930 2621 932
rect 3225 932 3239 966
rect 3273 932 3287 966
rect 3891 1038 3953 1076
rect 4853 1436 4867 1470
rect 4901 1436 4915 1470
rect 5519 1470 5581 1505
rect 4853 1398 4915 1436
rect 4853 1364 4867 1398
rect 4901 1364 4915 1398
rect 4853 1326 4915 1364
rect 4853 1292 4867 1326
rect 4901 1292 4915 1326
rect 4853 1254 4915 1292
rect 4853 1220 4867 1254
rect 4901 1220 4915 1254
rect 4853 1182 4915 1220
rect 4853 1148 4867 1182
rect 4901 1148 4915 1182
rect 4853 1110 4915 1148
rect 4853 1076 4867 1110
rect 4901 1076 4915 1110
rect 3891 1004 3905 1038
rect 3939 1004 3953 1038
rect 3891 966 3953 1004
rect 3225 930 3287 932
rect 3891 932 3905 966
rect 3939 932 3953 966
rect 4853 1038 4915 1076
rect 5519 1436 5533 1470
rect 5567 1436 5581 1470
rect 6481 1470 6543 1505
rect 5519 1398 5581 1436
rect 5519 1364 5533 1398
rect 5567 1364 5581 1398
rect 5519 1326 5581 1364
rect 5519 1292 5533 1326
rect 5567 1292 5581 1326
rect 5519 1254 5581 1292
rect 5519 1220 5533 1254
rect 5567 1220 5581 1254
rect 5519 1182 5581 1220
rect 5519 1148 5533 1182
rect 5567 1148 5581 1182
rect 5519 1110 5581 1148
rect 5519 1076 5533 1110
rect 5567 1076 5581 1110
rect 4853 1004 4867 1038
rect 4901 1004 4915 1038
rect 4853 966 4915 1004
rect 3891 930 3953 932
rect 4853 932 4867 966
rect 4901 932 4915 966
rect 5519 1038 5581 1076
rect 6481 1436 6495 1470
rect 6529 1436 6543 1470
rect 7443 1470 7505 1505
rect 6481 1398 6543 1436
rect 6481 1364 6495 1398
rect 6529 1364 6543 1398
rect 6481 1326 6543 1364
rect 6481 1292 6495 1326
rect 6529 1292 6543 1326
rect 6481 1254 6543 1292
rect 6481 1220 6495 1254
rect 6529 1220 6543 1254
rect 6481 1182 6543 1220
rect 6481 1148 6495 1182
rect 6529 1148 6543 1182
rect 6481 1110 6543 1148
rect 6481 1076 6495 1110
rect 6529 1076 6543 1110
rect 5519 1004 5533 1038
rect 5567 1004 5581 1038
rect 5519 966 5581 1004
rect 4853 930 4915 932
rect 5519 932 5533 966
rect 5567 932 5581 966
rect 6481 1038 6543 1076
rect 7443 1436 7457 1470
rect 7491 1436 7505 1470
rect 8109 1470 8171 1505
rect 7443 1398 7505 1436
rect 7443 1364 7457 1398
rect 7491 1364 7505 1398
rect 7443 1326 7505 1364
rect 7443 1292 7457 1326
rect 7491 1292 7505 1326
rect 7443 1254 7505 1292
rect 7443 1220 7457 1254
rect 7491 1220 7505 1254
rect 7443 1182 7505 1220
rect 7443 1148 7457 1182
rect 7491 1148 7505 1182
rect 7443 1110 7505 1148
rect 7443 1076 7457 1110
rect 7491 1076 7505 1110
rect 6481 1004 6495 1038
rect 6529 1004 6543 1038
rect 6481 966 6543 1004
rect 5519 930 5581 932
rect 6481 932 6495 966
rect 6529 932 6543 966
rect 7443 1038 7505 1076
rect 8109 1436 8123 1470
rect 8157 1436 8171 1470
rect 8775 1470 8837 1505
rect 8109 1398 8171 1436
rect 8109 1364 8123 1398
rect 8157 1364 8171 1398
rect 8109 1326 8171 1364
rect 8109 1292 8123 1326
rect 8157 1292 8171 1326
rect 8109 1254 8171 1292
rect 8109 1220 8123 1254
rect 8157 1220 8171 1254
rect 8109 1182 8171 1220
rect 8109 1148 8123 1182
rect 8157 1148 8171 1182
rect 8109 1110 8171 1148
rect 8109 1076 8123 1110
rect 8157 1076 8171 1110
rect 7443 1004 7457 1038
rect 7491 1004 7505 1038
rect 7443 966 7505 1004
rect 6481 930 6543 932
rect 7443 932 7457 966
rect 7491 932 7505 966
rect 8109 1038 8171 1076
rect 8775 1436 8789 1470
rect 8823 1436 8837 1470
rect 9737 1470 9799 1505
rect 8775 1398 8837 1436
rect 8775 1364 8789 1398
rect 8823 1364 8837 1398
rect 8775 1326 8837 1364
rect 8775 1292 8789 1326
rect 8823 1292 8837 1326
rect 8775 1254 8837 1292
rect 8775 1220 8789 1254
rect 8823 1220 8837 1254
rect 8775 1182 8837 1220
rect 8775 1148 8789 1182
rect 8823 1148 8837 1182
rect 8775 1110 8837 1148
rect 8775 1076 8789 1110
rect 8823 1076 8837 1110
rect 8109 1004 8123 1038
rect 8157 1004 8171 1038
rect 8109 966 8171 1004
rect 7443 930 7505 932
rect 8109 932 8123 966
rect 8157 932 8171 966
rect 8775 1038 8837 1076
rect 9737 1436 9751 1470
rect 9785 1436 9799 1470
rect 10403 1470 10465 1505
rect 9737 1398 9799 1436
rect 9737 1364 9751 1398
rect 9785 1364 9799 1398
rect 9737 1326 9799 1364
rect 9737 1292 9751 1326
rect 9785 1292 9799 1326
rect 9737 1254 9799 1292
rect 9737 1220 9751 1254
rect 9785 1220 9799 1254
rect 9737 1182 9799 1220
rect 9737 1148 9751 1182
rect 9785 1148 9799 1182
rect 9737 1110 9799 1148
rect 9737 1076 9751 1110
rect 9785 1076 9799 1110
rect 8775 1004 8789 1038
rect 8823 1004 8837 1038
rect 8775 966 8837 1004
rect 8109 930 8171 932
rect 8775 932 8789 966
rect 8823 932 8837 966
rect 9737 1038 9799 1076
rect 10403 1436 10417 1470
rect 10451 1436 10465 1470
rect 11365 1470 11427 1505
rect 10403 1398 10465 1436
rect 10403 1364 10417 1398
rect 10451 1364 10465 1398
rect 10403 1326 10465 1364
rect 10403 1292 10417 1326
rect 10451 1292 10465 1326
rect 10403 1254 10465 1292
rect 10403 1220 10417 1254
rect 10451 1220 10465 1254
rect 10403 1182 10465 1220
rect 10403 1148 10417 1182
rect 10451 1148 10465 1182
rect 10403 1110 10465 1148
rect 10403 1076 10417 1110
rect 10451 1076 10465 1110
rect 9737 1004 9751 1038
rect 9785 1004 9799 1038
rect 9737 966 9799 1004
rect 8775 930 8837 932
rect 9737 932 9751 966
rect 9785 932 9799 966
rect 10403 1038 10465 1076
rect 11365 1436 11379 1470
rect 11413 1436 11427 1470
rect 12327 1470 12389 1505
rect 11365 1398 11427 1436
rect 11365 1364 11379 1398
rect 11413 1364 11427 1398
rect 11365 1326 11427 1364
rect 11365 1292 11379 1326
rect 11413 1292 11427 1326
rect 11365 1254 11427 1292
rect 11365 1220 11379 1254
rect 11413 1220 11427 1254
rect 11365 1182 11427 1220
rect 11365 1148 11379 1182
rect 11413 1148 11427 1182
rect 11365 1110 11427 1148
rect 11365 1076 11379 1110
rect 11413 1076 11427 1110
rect 10403 1004 10417 1038
rect 10451 1004 10465 1038
rect 10403 966 10465 1004
rect 9737 930 9799 932
rect 10403 932 10417 966
rect 10451 932 10465 966
rect 11365 1038 11427 1076
rect 12327 1436 12341 1470
rect 12375 1436 12389 1470
rect 12993 1470 13055 1505
rect 12327 1398 12389 1436
rect 12327 1364 12341 1398
rect 12375 1364 12389 1398
rect 12327 1326 12389 1364
rect 12327 1292 12341 1326
rect 12375 1292 12389 1326
rect 12327 1254 12389 1292
rect 12327 1220 12341 1254
rect 12375 1220 12389 1254
rect 12327 1182 12389 1220
rect 12327 1148 12341 1182
rect 12375 1148 12389 1182
rect 12327 1110 12389 1148
rect 12327 1076 12341 1110
rect 12375 1076 12389 1110
rect 11365 1004 11379 1038
rect 11413 1004 11427 1038
rect 11365 966 11427 1004
rect 10403 930 10465 932
rect 11365 932 11379 966
rect 11413 932 11427 966
rect 12327 1038 12389 1076
rect 12993 1436 13007 1470
rect 13041 1436 13055 1470
rect 13659 1470 13721 1505
rect 12993 1398 13055 1436
rect 12993 1364 13007 1398
rect 13041 1364 13055 1398
rect 12993 1326 13055 1364
rect 12993 1292 13007 1326
rect 13041 1292 13055 1326
rect 12993 1254 13055 1292
rect 12993 1220 13007 1254
rect 13041 1220 13055 1254
rect 12993 1182 13055 1220
rect 12993 1148 13007 1182
rect 13041 1148 13055 1182
rect 12993 1110 13055 1148
rect 12993 1076 13007 1110
rect 13041 1076 13055 1110
rect 12327 1004 12341 1038
rect 12375 1004 12389 1038
rect 12327 966 12389 1004
rect 11365 930 11427 932
rect 12327 932 12341 966
rect 12375 932 12389 966
rect 12993 1038 13055 1076
rect 13659 1436 13673 1470
rect 13707 1436 13721 1470
rect 14621 1470 14683 1505
rect 13659 1398 13721 1436
rect 13659 1364 13673 1398
rect 13707 1364 13721 1398
rect 13659 1326 13721 1364
rect 13659 1292 13673 1326
rect 13707 1292 13721 1326
rect 13659 1254 13721 1292
rect 13659 1220 13673 1254
rect 13707 1220 13721 1254
rect 13659 1182 13721 1220
rect 13659 1148 13673 1182
rect 13707 1148 13721 1182
rect 13659 1110 13721 1148
rect 13659 1076 13673 1110
rect 13707 1076 13721 1110
rect 12993 1004 13007 1038
rect 13041 1004 13055 1038
rect 12993 966 13055 1004
rect 12327 930 12389 932
rect 12993 932 13007 966
rect 13041 932 13055 966
rect 13659 1038 13721 1076
rect 14621 1436 14635 1470
rect 14669 1436 14683 1470
rect 15287 1470 15349 1505
rect 14621 1398 14683 1436
rect 14621 1364 14635 1398
rect 14669 1364 14683 1398
rect 14621 1326 14683 1364
rect 14621 1292 14635 1326
rect 14669 1292 14683 1326
rect 14621 1254 14683 1292
rect 14621 1220 14635 1254
rect 14669 1220 14683 1254
rect 14621 1182 14683 1220
rect 14621 1148 14635 1182
rect 14669 1148 14683 1182
rect 14621 1110 14683 1148
rect 14621 1076 14635 1110
rect 14669 1076 14683 1110
rect 13659 1004 13673 1038
rect 13707 1004 13721 1038
rect 13659 966 13721 1004
rect 12993 930 13055 932
rect 13659 932 13673 966
rect 13707 932 13721 966
rect 14621 1038 14683 1076
rect 15287 1436 15301 1470
rect 15335 1436 15349 1470
rect 15953 1470 16015 1505
rect 15287 1398 15349 1436
rect 15287 1364 15301 1398
rect 15335 1364 15349 1398
rect 15287 1326 15349 1364
rect 15287 1292 15301 1326
rect 15335 1292 15349 1326
rect 15287 1254 15349 1292
rect 15287 1220 15301 1254
rect 15335 1220 15349 1254
rect 15287 1182 15349 1220
rect 15287 1148 15301 1182
rect 15335 1148 15349 1182
rect 15287 1110 15349 1148
rect 15287 1076 15301 1110
rect 15335 1076 15349 1110
rect 14621 1004 14635 1038
rect 14669 1004 14683 1038
rect 14621 966 14683 1004
rect 13659 930 13721 932
rect 14621 932 14635 966
rect 14669 932 14683 966
rect 15287 1038 15349 1076
rect 15953 1436 15967 1470
rect 16001 1436 16015 1470
rect 16619 1470 16681 1505
rect 15953 1398 16015 1436
rect 15953 1364 15967 1398
rect 16001 1364 16015 1398
rect 15953 1326 16015 1364
rect 15953 1292 15967 1326
rect 16001 1292 16015 1326
rect 15953 1254 16015 1292
rect 15953 1220 15967 1254
rect 16001 1220 16015 1254
rect 15953 1182 16015 1220
rect 15953 1148 15967 1182
rect 16001 1148 16015 1182
rect 15953 1110 16015 1148
rect 15953 1076 15967 1110
rect 16001 1076 16015 1110
rect 15287 1004 15301 1038
rect 15335 1004 15349 1038
rect 15287 966 15349 1004
rect 14621 930 14683 932
rect 15287 932 15301 966
rect 15335 932 15349 966
rect 15953 1038 16015 1076
rect 16619 1436 16633 1470
rect 16667 1436 16681 1470
rect 16619 1398 16681 1436
rect 16619 1364 16633 1398
rect 16667 1364 16681 1398
rect 16619 1326 16681 1364
rect 16619 1292 16633 1326
rect 16667 1292 16681 1326
rect 16619 1254 16681 1292
rect 16619 1220 16633 1254
rect 16667 1220 16681 1254
rect 16619 1182 16681 1220
rect 16619 1148 16633 1182
rect 16667 1148 16681 1182
rect 16619 1110 16681 1148
rect 16619 1076 16633 1110
rect 16667 1076 16681 1110
rect 15953 1004 15967 1038
rect 16001 1004 16015 1038
rect 15953 966 16015 1004
rect 15287 930 15349 932
rect 15953 932 15967 966
rect 16001 932 16015 966
rect 16619 1038 16681 1076
rect 16619 1004 16633 1038
rect 16667 1004 16681 1038
rect 16619 966 16681 1004
rect 15953 930 16015 932
rect 16619 932 16633 966
rect 16667 932 16681 966
rect 16619 930 16681 932
rect -31 868 16681 930
<< psubdiffcont >>
rect -17 512 17 546
rect 649 512 683 546
rect 1611 512 1645 546
rect 2573 512 2607 546
rect 3239 512 3273 546
rect 3905 512 3939 546
rect 4867 512 4901 546
rect 5533 512 5567 546
rect 6495 512 6529 546
rect 7457 512 7491 546
rect 8123 512 8157 546
rect 8789 512 8823 546
rect 9751 512 9785 546
rect 10417 512 10451 546
rect 11379 512 11413 546
rect 12341 512 12375 546
rect 13007 512 13041 546
rect 13673 512 13707 546
rect 14635 512 14669 546
rect 15301 512 15335 546
rect 15967 512 16001 546
rect 16633 512 16667 546
rect -17 440 17 474
rect -17 368 17 402
rect 649 440 683 474
rect -17 296 17 330
rect -17 224 17 258
rect -17 152 17 186
rect -17 80 17 114
rect 649 368 683 402
rect 1611 440 1645 474
rect 649 296 683 330
rect 649 224 683 258
rect 649 152 683 186
rect 649 80 683 114
rect 1611 368 1645 402
rect 2573 440 2607 474
rect 1611 296 1645 330
rect 1611 224 1645 258
rect 1611 152 1645 186
rect 1611 80 1645 114
rect 2573 368 2607 402
rect 3239 440 3273 474
rect 2573 296 2607 330
rect 2573 224 2607 258
rect 2573 152 2607 186
rect 2573 80 2607 114
rect 3239 368 3273 402
rect 3905 440 3939 474
rect 3239 296 3273 330
rect 3239 224 3273 258
rect 3239 152 3273 186
rect 3239 80 3273 114
rect 3905 368 3939 402
rect 4867 440 4901 474
rect 3905 296 3939 330
rect 3905 224 3939 258
rect 3905 152 3939 186
rect 3905 80 3939 114
rect 4867 368 4901 402
rect 5533 440 5567 474
rect 4867 296 4901 330
rect 4867 224 4901 258
rect 4867 152 4901 186
rect 4867 80 4901 114
rect 5533 368 5567 402
rect 6495 440 6529 474
rect 5533 296 5567 330
rect 5533 224 5567 258
rect 5533 152 5567 186
rect 5533 80 5567 114
rect 6495 368 6529 402
rect 7457 440 7491 474
rect 6495 296 6529 330
rect 6495 224 6529 258
rect 6495 152 6529 186
rect 6495 80 6529 114
rect 7457 368 7491 402
rect 8123 440 8157 474
rect 7457 296 7491 330
rect 7457 224 7491 258
rect 7457 152 7491 186
rect 7457 80 7491 114
rect 8123 368 8157 402
rect 8789 440 8823 474
rect 8123 296 8157 330
rect 8123 224 8157 258
rect 8123 152 8157 186
rect 8123 80 8157 114
rect 8789 368 8823 402
rect 9751 440 9785 474
rect 8789 296 8823 330
rect 8789 224 8823 258
rect 8789 152 8823 186
rect 8789 80 8823 114
rect 9751 368 9785 402
rect 10417 440 10451 474
rect 9751 296 9785 330
rect 9751 224 9785 258
rect 9751 152 9785 186
rect 9751 80 9785 114
rect 10417 368 10451 402
rect 11379 440 11413 474
rect 10417 296 10451 330
rect 10417 224 10451 258
rect 10417 152 10451 186
rect 10417 80 10451 114
rect 11379 368 11413 402
rect 12341 440 12375 474
rect 11379 296 11413 330
rect 11379 224 11413 258
rect 11379 152 11413 186
rect 11379 80 11413 114
rect 12341 368 12375 402
rect 13007 440 13041 474
rect 12341 296 12375 330
rect 12341 224 12375 258
rect 12341 152 12375 186
rect 12341 80 12375 114
rect 13007 368 13041 402
rect 13673 440 13707 474
rect 13007 296 13041 330
rect 13007 224 13041 258
rect 13007 152 13041 186
rect 13007 80 13041 114
rect 13673 368 13707 402
rect 14635 440 14669 474
rect 15301 440 15335 474
rect 13673 296 13707 330
rect 13673 224 13707 258
rect 13673 152 13707 186
rect 13673 80 13707 114
rect 14635 368 14669 402
rect 14635 296 14669 330
rect 14635 224 14669 258
rect 14635 152 14669 186
rect 14635 80 14669 114
rect 15301 368 15335 402
rect 15967 440 16001 474
rect 16633 440 16667 474
rect 15301 296 15335 330
rect 15301 224 15335 258
rect 15301 152 15335 186
rect 15301 80 15335 114
rect 15967 368 16001 402
rect 15967 296 16001 330
rect 15967 224 16001 258
rect 15967 152 16001 186
rect 15967 80 16001 114
rect 16633 368 16667 402
rect 16633 296 16667 330
rect 16633 224 16667 258
rect 16633 152 16667 186
rect 16633 80 16667 114
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 361 13 395 47
rect 433 13 467 47
rect 505 13 539 47
rect 577 13 611 47
rect 721 13 755 47
rect 793 13 827 47
rect 865 13 899 47
rect 937 13 971 47
rect 1009 13 1043 47
rect 1081 13 1115 47
rect 1179 13 1213 47
rect 1251 13 1285 47
rect 1323 13 1357 47
rect 1395 13 1429 47
rect 1467 13 1501 47
rect 1539 13 1573 47
rect 1683 13 1717 47
rect 1755 13 1789 47
rect 1827 13 1861 47
rect 1899 13 1933 47
rect 1971 13 2005 47
rect 2043 13 2077 47
rect 2141 13 2175 47
rect 2213 13 2247 47
rect 2285 13 2319 47
rect 2357 13 2391 47
rect 2429 13 2463 47
rect 2501 13 2535 47
rect 2645 13 2679 47
rect 2717 13 2751 47
rect 2789 13 2823 47
rect 2861 13 2895 47
rect 2951 13 2985 47
rect 3023 13 3057 47
rect 3095 13 3129 47
rect 3167 13 3201 47
rect 3311 13 3345 47
rect 3383 13 3417 47
rect 3455 13 3489 47
rect 3527 13 3561 47
rect 3617 13 3651 47
rect 3689 13 3723 47
rect 3761 13 3795 47
rect 3833 13 3867 47
rect 3977 13 4011 47
rect 4049 13 4083 47
rect 4121 13 4155 47
rect 4193 13 4227 47
rect 4265 13 4299 47
rect 4337 13 4371 47
rect 4435 13 4469 47
rect 4507 13 4541 47
rect 4579 13 4613 47
rect 4651 13 4685 47
rect 4723 13 4757 47
rect 4795 13 4829 47
rect 4939 13 4973 47
rect 5011 13 5045 47
rect 5083 13 5117 47
rect 5155 13 5189 47
rect 5245 13 5279 47
rect 5317 13 5351 47
rect 5389 13 5423 47
rect 5461 13 5495 47
rect 5605 13 5639 47
rect 5677 13 5711 47
rect 5749 13 5783 47
rect 5821 13 5855 47
rect 5893 13 5927 47
rect 5965 13 5999 47
rect 6063 13 6097 47
rect 6135 13 6169 47
rect 6207 13 6241 47
rect 6279 13 6313 47
rect 6351 13 6385 47
rect 6423 13 6457 47
rect 6567 13 6601 47
rect 6639 13 6673 47
rect 6711 13 6745 47
rect 6783 13 6817 47
rect 6855 13 6889 47
rect 6927 13 6961 47
rect 7025 13 7059 47
rect 7097 13 7131 47
rect 7169 13 7203 47
rect 7241 13 7275 47
rect 7313 13 7347 47
rect 7385 13 7419 47
rect 7529 13 7563 47
rect 7601 13 7635 47
rect 7673 13 7707 47
rect 7745 13 7779 47
rect 7835 13 7869 47
rect 7907 13 7941 47
rect 7979 13 8013 47
rect 8051 13 8085 47
rect 8195 13 8229 47
rect 8267 13 8301 47
rect 8339 13 8373 47
rect 8411 13 8445 47
rect 8501 13 8535 47
rect 8573 13 8607 47
rect 8645 13 8679 47
rect 8717 13 8751 47
rect 8861 13 8895 47
rect 8933 13 8967 47
rect 9005 13 9039 47
rect 9077 13 9111 47
rect 9149 13 9183 47
rect 9221 13 9255 47
rect 9319 13 9353 47
rect 9391 13 9425 47
rect 9463 13 9497 47
rect 9535 13 9569 47
rect 9607 13 9641 47
rect 9679 13 9713 47
rect 9823 13 9857 47
rect 9895 13 9929 47
rect 9967 13 10001 47
rect 10039 13 10073 47
rect 10129 13 10163 47
rect 10201 13 10235 47
rect 10273 13 10307 47
rect 10345 13 10379 47
rect 10489 13 10523 47
rect 10561 13 10595 47
rect 10633 13 10667 47
rect 10705 13 10739 47
rect 10777 13 10811 47
rect 10849 13 10883 47
rect 10947 13 10981 47
rect 11019 13 11053 47
rect 11091 13 11125 47
rect 11163 13 11197 47
rect 11235 13 11269 47
rect 11307 13 11341 47
rect 11451 13 11485 47
rect 11523 13 11557 47
rect 11595 13 11629 47
rect 11667 13 11701 47
rect 11739 13 11773 47
rect 11811 13 11845 47
rect 11909 13 11943 47
rect 11981 13 12015 47
rect 12053 13 12087 47
rect 12125 13 12159 47
rect 12197 13 12231 47
rect 12269 13 12303 47
rect 12413 13 12447 47
rect 12485 13 12519 47
rect 12557 13 12591 47
rect 12629 13 12663 47
rect 12719 13 12753 47
rect 12791 13 12825 47
rect 12863 13 12897 47
rect 12935 13 12969 47
rect 13079 13 13113 47
rect 13151 13 13185 47
rect 13223 13 13257 47
rect 13295 13 13329 47
rect 13385 13 13419 47
rect 13457 13 13491 47
rect 13529 13 13563 47
rect 13601 13 13635 47
rect 13745 13 13779 47
rect 13817 13 13851 47
rect 13889 13 13923 47
rect 13961 13 13995 47
rect 14033 13 14067 47
rect 14105 13 14139 47
rect 14203 13 14237 47
rect 14275 13 14309 47
rect 14347 13 14381 47
rect 14419 13 14453 47
rect 14491 13 14525 47
rect 14563 13 14597 47
rect 14707 13 14741 47
rect 14779 13 14813 47
rect 14851 13 14885 47
rect 14923 13 14957 47
rect 15013 13 15047 47
rect 15085 13 15119 47
rect 15157 13 15191 47
rect 15229 13 15263 47
rect 15373 13 15407 47
rect 15445 13 15479 47
rect 15517 13 15551 47
rect 15589 13 15623 47
rect 15679 13 15713 47
rect 15751 13 15785 47
rect 15823 13 15857 47
rect 15895 13 15929 47
rect 16039 13 16073 47
rect 16111 13 16145 47
rect 16183 13 16217 47
rect 16255 13 16289 47
rect 16345 13 16379 47
rect 16417 13 16451 47
rect 16489 13 16523 47
rect 16561 13 16595 47
<< nsubdiffcont >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 361 1505 395 1539
rect 433 1505 467 1539
rect 505 1505 539 1539
rect 577 1505 611 1539
rect 721 1505 755 1539
rect 793 1505 827 1539
rect 865 1505 899 1539
rect 937 1505 971 1539
rect 1009 1505 1043 1539
rect 1081 1505 1115 1539
rect 1179 1505 1213 1539
rect 1251 1505 1285 1539
rect 1323 1505 1357 1539
rect 1395 1505 1429 1539
rect 1467 1505 1501 1539
rect 1539 1505 1573 1539
rect 1683 1505 1717 1539
rect 1755 1505 1789 1539
rect 1827 1505 1861 1539
rect 1899 1505 1933 1539
rect 1971 1505 2005 1539
rect 2043 1505 2077 1539
rect 2141 1505 2175 1539
rect 2213 1505 2247 1539
rect 2285 1505 2319 1539
rect 2357 1505 2391 1539
rect 2429 1505 2463 1539
rect 2501 1505 2535 1539
rect 2645 1505 2679 1539
rect 2717 1505 2751 1539
rect 2789 1505 2823 1539
rect 2861 1505 2895 1539
rect 2951 1505 2985 1539
rect 3023 1505 3057 1539
rect 3095 1505 3129 1539
rect 3167 1505 3201 1539
rect 3311 1505 3345 1539
rect 3383 1505 3417 1539
rect 3455 1505 3489 1539
rect 3527 1505 3561 1539
rect 3617 1505 3651 1539
rect 3689 1505 3723 1539
rect 3761 1505 3795 1539
rect 3833 1505 3867 1539
rect 3977 1505 4011 1539
rect 4049 1505 4083 1539
rect 4121 1505 4155 1539
rect 4193 1505 4227 1539
rect 4265 1505 4299 1539
rect 4337 1505 4371 1539
rect 4435 1505 4469 1539
rect 4507 1505 4541 1539
rect 4579 1505 4613 1539
rect 4651 1505 4685 1539
rect 4723 1505 4757 1539
rect 4795 1505 4829 1539
rect 4939 1505 4973 1539
rect 5011 1505 5045 1539
rect 5083 1505 5117 1539
rect 5155 1505 5189 1539
rect 5245 1505 5279 1539
rect 5317 1505 5351 1539
rect 5389 1505 5423 1539
rect 5461 1505 5495 1539
rect 5605 1505 5639 1539
rect 5677 1505 5711 1539
rect 5749 1505 5783 1539
rect 5821 1505 5855 1539
rect 5893 1505 5927 1539
rect 5965 1505 5999 1539
rect 6063 1505 6097 1539
rect 6135 1505 6169 1539
rect 6207 1505 6241 1539
rect 6279 1505 6313 1539
rect 6351 1505 6385 1539
rect 6423 1505 6457 1539
rect 6567 1505 6601 1539
rect 6639 1505 6673 1539
rect 6711 1505 6745 1539
rect 6783 1505 6817 1539
rect 6855 1505 6889 1539
rect 6927 1505 6961 1539
rect 7025 1505 7059 1539
rect 7097 1505 7131 1539
rect 7169 1505 7203 1539
rect 7241 1505 7275 1539
rect 7313 1505 7347 1539
rect 7385 1505 7419 1539
rect 7529 1505 7563 1539
rect 7601 1505 7635 1539
rect 7673 1505 7707 1539
rect 7745 1505 7779 1539
rect 7835 1505 7869 1539
rect 7907 1505 7941 1539
rect 7979 1505 8013 1539
rect 8051 1505 8085 1539
rect 8195 1505 8229 1539
rect 8267 1505 8301 1539
rect 8339 1505 8373 1539
rect 8411 1505 8445 1539
rect 8501 1505 8535 1539
rect 8573 1505 8607 1539
rect 8645 1505 8679 1539
rect 8717 1505 8751 1539
rect 8861 1505 8895 1539
rect 8933 1505 8967 1539
rect 9005 1505 9039 1539
rect 9077 1505 9111 1539
rect 9149 1505 9183 1539
rect 9221 1505 9255 1539
rect 9319 1505 9353 1539
rect 9391 1505 9425 1539
rect 9463 1505 9497 1539
rect 9535 1505 9569 1539
rect 9607 1505 9641 1539
rect 9679 1505 9713 1539
rect 9823 1505 9857 1539
rect 9895 1505 9929 1539
rect 9967 1505 10001 1539
rect 10039 1505 10073 1539
rect 10129 1505 10163 1539
rect 10201 1505 10235 1539
rect 10273 1505 10307 1539
rect 10345 1505 10379 1539
rect 10489 1505 10523 1539
rect 10561 1505 10595 1539
rect 10633 1505 10667 1539
rect 10705 1505 10739 1539
rect 10777 1505 10811 1539
rect 10849 1505 10883 1539
rect 10947 1505 10981 1539
rect 11019 1505 11053 1539
rect 11091 1505 11125 1539
rect 11163 1505 11197 1539
rect 11235 1505 11269 1539
rect 11307 1505 11341 1539
rect 11451 1505 11485 1539
rect 11523 1505 11557 1539
rect 11595 1505 11629 1539
rect 11667 1505 11701 1539
rect 11739 1505 11773 1539
rect 11811 1505 11845 1539
rect 11909 1505 11943 1539
rect 11981 1505 12015 1539
rect 12053 1505 12087 1539
rect 12125 1505 12159 1539
rect 12197 1505 12231 1539
rect 12269 1505 12303 1539
rect 12413 1505 12447 1539
rect 12485 1505 12519 1539
rect 12557 1505 12591 1539
rect 12629 1505 12663 1539
rect 12719 1505 12753 1539
rect 12791 1505 12825 1539
rect 12863 1505 12897 1539
rect 12935 1505 12969 1539
rect 13079 1505 13113 1539
rect 13151 1505 13185 1539
rect 13223 1505 13257 1539
rect 13295 1505 13329 1539
rect 13385 1505 13419 1539
rect 13457 1505 13491 1539
rect 13529 1505 13563 1539
rect 13601 1505 13635 1539
rect 13745 1505 13779 1539
rect 13817 1505 13851 1539
rect 13889 1505 13923 1539
rect 13961 1505 13995 1539
rect 14033 1505 14067 1539
rect 14105 1505 14139 1539
rect 14203 1505 14237 1539
rect 14275 1505 14309 1539
rect 14347 1505 14381 1539
rect 14419 1505 14453 1539
rect 14491 1505 14525 1539
rect 14563 1505 14597 1539
rect 14707 1505 14741 1539
rect 14779 1505 14813 1539
rect 14851 1505 14885 1539
rect 14923 1505 14957 1539
rect 15013 1505 15047 1539
rect 15085 1505 15119 1539
rect 15157 1505 15191 1539
rect 15229 1505 15263 1539
rect 15373 1505 15407 1539
rect 15445 1505 15479 1539
rect 15517 1505 15551 1539
rect 15589 1505 15623 1539
rect 15679 1505 15713 1539
rect 15751 1505 15785 1539
rect 15823 1505 15857 1539
rect 15895 1505 15929 1539
rect 16039 1505 16073 1539
rect 16111 1505 16145 1539
rect 16183 1505 16217 1539
rect 16255 1505 16289 1539
rect 16345 1505 16379 1539
rect 16417 1505 16451 1539
rect 16489 1505 16523 1539
rect 16561 1505 16595 1539
rect -17 1436 17 1470
rect -17 1364 17 1398
rect -17 1292 17 1326
rect -17 1220 17 1254
rect -17 1148 17 1182
rect -17 1076 17 1110
rect 649 1436 683 1470
rect 649 1364 683 1398
rect 649 1292 683 1326
rect 649 1220 683 1254
rect 649 1148 683 1182
rect 649 1076 683 1110
rect -17 1004 17 1038
rect -17 932 17 966
rect 1611 1436 1645 1470
rect 1611 1364 1645 1398
rect 1611 1292 1645 1326
rect 1611 1220 1645 1254
rect 1611 1148 1645 1182
rect 1611 1076 1645 1110
rect 649 1004 683 1038
rect 649 932 683 966
rect 2573 1436 2607 1470
rect 2573 1364 2607 1398
rect 2573 1292 2607 1326
rect 2573 1220 2607 1254
rect 2573 1148 2607 1182
rect 2573 1076 2607 1110
rect 1611 1004 1645 1038
rect 1611 932 1645 966
rect 3239 1436 3273 1470
rect 3239 1364 3273 1398
rect 3239 1292 3273 1326
rect 3239 1220 3273 1254
rect 3239 1148 3273 1182
rect 3239 1076 3273 1110
rect 2573 1004 2607 1038
rect 2573 932 2607 966
rect 3905 1436 3939 1470
rect 3905 1364 3939 1398
rect 3905 1292 3939 1326
rect 3905 1220 3939 1254
rect 3905 1148 3939 1182
rect 3905 1076 3939 1110
rect 3239 1004 3273 1038
rect 3239 932 3273 966
rect 4867 1436 4901 1470
rect 4867 1364 4901 1398
rect 4867 1292 4901 1326
rect 4867 1220 4901 1254
rect 4867 1148 4901 1182
rect 4867 1076 4901 1110
rect 3905 1004 3939 1038
rect 3905 932 3939 966
rect 5533 1436 5567 1470
rect 5533 1364 5567 1398
rect 5533 1292 5567 1326
rect 5533 1220 5567 1254
rect 5533 1148 5567 1182
rect 5533 1076 5567 1110
rect 4867 1004 4901 1038
rect 4867 932 4901 966
rect 6495 1436 6529 1470
rect 6495 1364 6529 1398
rect 6495 1292 6529 1326
rect 6495 1220 6529 1254
rect 6495 1148 6529 1182
rect 6495 1076 6529 1110
rect 5533 1004 5567 1038
rect 5533 932 5567 966
rect 7457 1436 7491 1470
rect 7457 1364 7491 1398
rect 7457 1292 7491 1326
rect 7457 1220 7491 1254
rect 7457 1148 7491 1182
rect 7457 1076 7491 1110
rect 6495 1004 6529 1038
rect 6495 932 6529 966
rect 8123 1436 8157 1470
rect 8123 1364 8157 1398
rect 8123 1292 8157 1326
rect 8123 1220 8157 1254
rect 8123 1148 8157 1182
rect 8123 1076 8157 1110
rect 7457 1004 7491 1038
rect 7457 932 7491 966
rect 8789 1436 8823 1470
rect 8789 1364 8823 1398
rect 8789 1292 8823 1326
rect 8789 1220 8823 1254
rect 8789 1148 8823 1182
rect 8789 1076 8823 1110
rect 8123 1004 8157 1038
rect 8123 932 8157 966
rect 9751 1436 9785 1470
rect 9751 1364 9785 1398
rect 9751 1292 9785 1326
rect 9751 1220 9785 1254
rect 9751 1148 9785 1182
rect 9751 1076 9785 1110
rect 8789 1004 8823 1038
rect 8789 932 8823 966
rect 10417 1436 10451 1470
rect 10417 1364 10451 1398
rect 10417 1292 10451 1326
rect 10417 1220 10451 1254
rect 10417 1148 10451 1182
rect 10417 1076 10451 1110
rect 9751 1004 9785 1038
rect 9751 932 9785 966
rect 11379 1436 11413 1470
rect 11379 1364 11413 1398
rect 11379 1292 11413 1326
rect 11379 1220 11413 1254
rect 11379 1148 11413 1182
rect 11379 1076 11413 1110
rect 10417 1004 10451 1038
rect 10417 932 10451 966
rect 12341 1436 12375 1470
rect 12341 1364 12375 1398
rect 12341 1292 12375 1326
rect 12341 1220 12375 1254
rect 12341 1148 12375 1182
rect 12341 1076 12375 1110
rect 11379 1004 11413 1038
rect 11379 932 11413 966
rect 13007 1436 13041 1470
rect 13007 1364 13041 1398
rect 13007 1292 13041 1326
rect 13007 1220 13041 1254
rect 13007 1148 13041 1182
rect 13007 1076 13041 1110
rect 12341 1004 12375 1038
rect 12341 932 12375 966
rect 13673 1436 13707 1470
rect 13673 1364 13707 1398
rect 13673 1292 13707 1326
rect 13673 1220 13707 1254
rect 13673 1148 13707 1182
rect 13673 1076 13707 1110
rect 13007 1004 13041 1038
rect 13007 932 13041 966
rect 14635 1436 14669 1470
rect 14635 1364 14669 1398
rect 14635 1292 14669 1326
rect 14635 1220 14669 1254
rect 14635 1148 14669 1182
rect 14635 1076 14669 1110
rect 13673 1004 13707 1038
rect 13673 932 13707 966
rect 15301 1436 15335 1470
rect 15301 1364 15335 1398
rect 15301 1292 15335 1326
rect 15301 1220 15335 1254
rect 15301 1148 15335 1182
rect 15301 1076 15335 1110
rect 14635 1004 14669 1038
rect 14635 932 14669 966
rect 15967 1436 16001 1470
rect 15967 1364 16001 1398
rect 15967 1292 16001 1326
rect 15967 1220 16001 1254
rect 15967 1148 16001 1182
rect 15967 1076 16001 1110
rect 15301 1004 15335 1038
rect 15301 932 15335 966
rect 16633 1436 16667 1470
rect 16633 1364 16667 1398
rect 16633 1292 16667 1326
rect 16633 1220 16667 1254
rect 16633 1148 16667 1182
rect 16633 1076 16667 1110
rect 15967 1004 16001 1038
rect 15967 932 16001 966
rect 16633 1004 16667 1038
rect 16633 932 16667 966
<< poly >>
rect 187 1450 217 1476
rect 275 1450 305 1476
rect 363 1450 393 1476
rect 451 1450 481 1476
rect 913 1450 943 1476
rect 1001 1450 1031 1476
rect 1089 1450 1119 1476
rect 1177 1450 1207 1476
rect 1265 1450 1295 1476
rect 1353 1450 1383 1476
rect 187 1019 217 1050
rect 275 1019 305 1050
rect 363 1019 393 1050
rect 451 1019 481 1050
rect 187 1003 305 1019
rect 187 989 205 1003
rect 195 969 205 989
rect 239 989 305 1003
rect 349 1003 481 1019
rect 239 969 249 989
rect 195 953 249 969
rect 349 969 359 1003
rect 393 989 481 1003
rect 1875 1450 1905 1476
rect 1963 1450 1993 1476
rect 2051 1450 2081 1476
rect 2139 1450 2169 1476
rect 2227 1450 2257 1476
rect 2315 1450 2345 1476
rect 913 1019 943 1050
rect 1001 1019 1031 1050
rect 1089 1019 1119 1050
rect 1177 1019 1207 1050
rect 393 969 403 989
rect 349 953 403 969
rect 861 1003 1031 1019
rect 861 969 871 1003
rect 905 989 1031 1003
rect 1083 1003 1207 1019
rect 905 969 915 989
rect 861 953 915 969
rect 1083 969 1093 1003
rect 1127 989 1207 1003
rect 1265 1019 1295 1050
rect 1353 1019 1383 1050
rect 1265 1003 1383 1019
rect 1265 989 1315 1003
rect 1127 969 1137 989
rect 1083 953 1137 969
rect 1305 969 1315 989
rect 1349 989 1383 1003
rect 2777 1450 2807 1476
rect 2865 1450 2895 1476
rect 2953 1450 2983 1476
rect 3041 1450 3071 1476
rect 1875 1019 1905 1050
rect 1963 1019 1993 1050
rect 2051 1019 2081 1050
rect 2139 1019 2169 1050
rect 1349 969 1359 989
rect 1305 953 1359 969
rect 1823 1003 1993 1019
rect 1823 969 1833 1003
rect 1867 989 1993 1003
rect 2045 1003 2169 1019
rect 1867 969 1877 989
rect 1823 953 1877 969
rect 2045 969 2055 1003
rect 2089 989 2169 1003
rect 2227 1019 2257 1050
rect 2315 1019 2345 1050
rect 2227 1003 2345 1019
rect 2227 989 2277 1003
rect 2089 969 2099 989
rect 2045 953 2099 969
rect 2267 969 2277 989
rect 2311 989 2345 1003
rect 3443 1450 3473 1476
rect 3531 1450 3561 1476
rect 3619 1450 3649 1476
rect 3707 1450 3737 1476
rect 2311 969 2321 989
rect 2267 953 2321 969
rect 2777 1019 2807 1050
rect 2865 1019 2895 1050
rect 2953 1019 2983 1050
rect 3041 1019 3071 1050
rect 2777 1003 2895 1019
rect 2777 989 2795 1003
rect 2785 969 2795 989
rect 2829 989 2895 1003
rect 2939 1003 3071 1019
rect 2829 969 2839 989
rect 2785 953 2839 969
rect 2939 969 2949 1003
rect 2983 989 3071 1003
rect 4169 1450 4199 1476
rect 4257 1450 4287 1476
rect 4345 1450 4375 1476
rect 4433 1450 4463 1476
rect 4521 1450 4551 1476
rect 4609 1450 4639 1476
rect 2983 969 2993 989
rect 2939 953 2993 969
rect 3443 1019 3473 1050
rect 3531 1019 3561 1050
rect 3619 1019 3649 1050
rect 3707 1019 3737 1050
rect 3443 1003 3561 1019
rect 3443 989 3461 1003
rect 3451 969 3461 989
rect 3495 989 3561 1003
rect 3605 1003 3737 1019
rect 3495 969 3505 989
rect 3451 953 3505 969
rect 3605 969 3615 1003
rect 3649 989 3737 1003
rect 5071 1450 5101 1476
rect 5159 1450 5189 1476
rect 5247 1450 5277 1476
rect 5335 1450 5365 1476
rect 4169 1019 4199 1050
rect 4257 1019 4287 1050
rect 4345 1019 4375 1050
rect 4433 1019 4463 1050
rect 3649 969 3659 989
rect 3605 953 3659 969
rect 4117 1003 4287 1019
rect 4117 969 4127 1003
rect 4161 989 4287 1003
rect 4339 1003 4463 1019
rect 4161 969 4171 989
rect 4117 953 4171 969
rect 4339 969 4349 1003
rect 4383 989 4463 1003
rect 4521 1019 4551 1050
rect 4609 1019 4639 1050
rect 4521 1003 4639 1019
rect 4521 989 4571 1003
rect 4383 969 4393 989
rect 4339 953 4393 969
rect 4561 969 4571 989
rect 4605 989 4639 1003
rect 5797 1450 5827 1476
rect 5885 1450 5915 1476
rect 5973 1450 6003 1476
rect 6061 1450 6091 1476
rect 6149 1450 6179 1476
rect 6237 1450 6267 1476
rect 4605 969 4615 989
rect 4561 953 4615 969
rect 5071 1019 5101 1050
rect 5159 1019 5189 1050
rect 5247 1019 5277 1050
rect 5335 1019 5365 1050
rect 5071 1003 5189 1019
rect 5071 989 5089 1003
rect 5079 969 5089 989
rect 5123 989 5189 1003
rect 5233 1003 5365 1019
rect 5123 969 5133 989
rect 5079 953 5133 969
rect 5233 969 5243 1003
rect 5277 989 5365 1003
rect 6759 1450 6789 1476
rect 6847 1450 6877 1476
rect 6935 1450 6965 1476
rect 7023 1450 7053 1476
rect 7111 1450 7141 1476
rect 7199 1450 7229 1476
rect 5797 1019 5827 1050
rect 5885 1019 5915 1050
rect 5973 1019 6003 1050
rect 6061 1019 6091 1050
rect 5277 969 5287 989
rect 5233 953 5287 969
rect 5745 1003 5915 1019
rect 5745 969 5755 1003
rect 5789 989 5915 1003
rect 5967 1003 6091 1019
rect 5789 969 5799 989
rect 5745 953 5799 969
rect 5967 969 5977 1003
rect 6011 989 6091 1003
rect 6149 1019 6179 1050
rect 6237 1019 6267 1050
rect 6149 1003 6267 1019
rect 6149 989 6199 1003
rect 6011 969 6021 989
rect 5967 953 6021 969
rect 6189 969 6199 989
rect 6233 989 6267 1003
rect 7661 1450 7691 1476
rect 7749 1450 7779 1476
rect 7837 1450 7867 1476
rect 7925 1450 7955 1476
rect 6759 1019 6789 1050
rect 6847 1019 6877 1050
rect 6935 1019 6965 1050
rect 7023 1019 7053 1050
rect 6233 969 6243 989
rect 6189 953 6243 969
rect 6707 1003 6877 1019
rect 6707 969 6717 1003
rect 6751 989 6877 1003
rect 6929 1003 7053 1019
rect 6751 969 6761 989
rect 6707 953 6761 969
rect 6929 969 6939 1003
rect 6973 989 7053 1003
rect 7111 1019 7141 1050
rect 7199 1019 7229 1050
rect 7111 1003 7229 1019
rect 7111 989 7161 1003
rect 6973 969 6983 989
rect 6929 953 6983 969
rect 7151 969 7161 989
rect 7195 989 7229 1003
rect 8327 1450 8357 1476
rect 8415 1450 8445 1476
rect 8503 1450 8533 1476
rect 8591 1450 8621 1476
rect 7195 969 7205 989
rect 7151 953 7205 969
rect 7661 1019 7691 1050
rect 7749 1019 7779 1050
rect 7837 1019 7867 1050
rect 7925 1019 7955 1050
rect 7661 1003 7779 1019
rect 7661 989 7679 1003
rect 7669 969 7679 989
rect 7713 989 7779 1003
rect 7823 1003 7955 1019
rect 7713 969 7723 989
rect 7669 953 7723 969
rect 7823 969 7833 1003
rect 7867 989 7955 1003
rect 9053 1450 9083 1476
rect 9141 1450 9171 1476
rect 9229 1450 9259 1476
rect 9317 1450 9347 1476
rect 9405 1450 9435 1476
rect 9493 1450 9523 1476
rect 7867 969 7877 989
rect 7823 953 7877 969
rect 8327 1019 8357 1050
rect 8415 1019 8445 1050
rect 8503 1019 8533 1050
rect 8591 1019 8621 1050
rect 8327 1003 8445 1019
rect 8327 989 8345 1003
rect 8335 969 8345 989
rect 8379 989 8445 1003
rect 8489 1003 8621 1019
rect 8379 969 8389 989
rect 8335 953 8389 969
rect 8489 969 8499 1003
rect 8533 989 8621 1003
rect 9955 1450 9985 1476
rect 10043 1450 10073 1476
rect 10131 1450 10161 1476
rect 10219 1450 10249 1476
rect 9053 1019 9083 1050
rect 9141 1019 9171 1050
rect 9229 1019 9259 1050
rect 9317 1019 9347 1050
rect 8533 969 8543 989
rect 8489 953 8543 969
rect 9001 1003 9171 1019
rect 9001 969 9011 1003
rect 9045 989 9171 1003
rect 9223 1003 9347 1019
rect 9045 969 9055 989
rect 9001 953 9055 969
rect 9223 969 9233 1003
rect 9267 989 9347 1003
rect 9405 1019 9435 1050
rect 9493 1019 9523 1050
rect 9405 1003 9523 1019
rect 9405 989 9455 1003
rect 9267 969 9277 989
rect 9223 953 9277 969
rect 9445 969 9455 989
rect 9489 989 9523 1003
rect 10681 1450 10711 1476
rect 10769 1450 10799 1476
rect 10857 1450 10887 1476
rect 10945 1450 10975 1476
rect 11033 1450 11063 1476
rect 11121 1450 11151 1476
rect 9489 969 9499 989
rect 9445 953 9499 969
rect 9955 1019 9985 1050
rect 10043 1019 10073 1050
rect 10131 1019 10161 1050
rect 10219 1019 10249 1050
rect 9955 1003 10073 1019
rect 9955 989 9973 1003
rect 9963 969 9973 989
rect 10007 989 10073 1003
rect 10117 1003 10249 1019
rect 10007 969 10017 989
rect 9963 953 10017 969
rect 10117 969 10127 1003
rect 10161 989 10249 1003
rect 11643 1450 11673 1476
rect 11731 1450 11761 1476
rect 11819 1450 11849 1476
rect 11907 1450 11937 1476
rect 11995 1450 12025 1476
rect 12083 1450 12113 1476
rect 10681 1019 10711 1050
rect 10769 1019 10799 1050
rect 10857 1019 10887 1050
rect 10945 1019 10975 1050
rect 10161 969 10171 989
rect 10117 953 10171 969
rect 10629 1003 10799 1019
rect 10629 969 10639 1003
rect 10673 989 10799 1003
rect 10851 1003 10975 1019
rect 10673 969 10683 989
rect 10629 953 10683 969
rect 10851 969 10861 1003
rect 10895 989 10975 1003
rect 11033 1019 11063 1050
rect 11121 1019 11151 1050
rect 11033 1003 11151 1019
rect 11033 989 11083 1003
rect 10895 969 10905 989
rect 10851 953 10905 969
rect 11073 969 11083 989
rect 11117 989 11151 1003
rect 12545 1450 12575 1476
rect 12633 1450 12663 1476
rect 12721 1450 12751 1476
rect 12809 1450 12839 1476
rect 11643 1019 11673 1050
rect 11731 1019 11761 1050
rect 11819 1019 11849 1050
rect 11907 1019 11937 1050
rect 11117 969 11127 989
rect 11073 953 11127 969
rect 11591 1003 11761 1019
rect 11591 969 11601 1003
rect 11635 989 11761 1003
rect 11813 1003 11937 1019
rect 11635 969 11645 989
rect 11591 953 11645 969
rect 11813 969 11823 1003
rect 11857 989 11937 1003
rect 11995 1019 12025 1050
rect 12083 1019 12113 1050
rect 11995 1003 12113 1019
rect 11995 989 12045 1003
rect 11857 969 11867 989
rect 11813 953 11867 969
rect 12035 969 12045 989
rect 12079 989 12113 1003
rect 13211 1450 13241 1476
rect 13299 1450 13329 1476
rect 13387 1450 13417 1476
rect 13475 1450 13505 1476
rect 12079 969 12089 989
rect 12035 953 12089 969
rect 12545 1019 12575 1050
rect 12633 1019 12663 1050
rect 12721 1019 12751 1050
rect 12809 1019 12839 1050
rect 12545 1003 12663 1019
rect 12545 989 12563 1003
rect 12553 969 12563 989
rect 12597 989 12663 1003
rect 12707 1003 12839 1019
rect 12597 969 12607 989
rect 12553 953 12607 969
rect 12707 969 12717 1003
rect 12751 989 12839 1003
rect 13937 1450 13967 1476
rect 14025 1450 14055 1476
rect 14113 1450 14143 1476
rect 14201 1450 14231 1476
rect 14289 1450 14319 1476
rect 14377 1450 14407 1476
rect 12751 969 12761 989
rect 12707 953 12761 969
rect 13211 1019 13241 1050
rect 13299 1019 13329 1050
rect 13387 1019 13417 1050
rect 13475 1019 13505 1050
rect 13211 1003 13329 1019
rect 13211 989 13229 1003
rect 13219 969 13229 989
rect 13263 989 13329 1003
rect 13373 1003 13505 1019
rect 13263 969 13273 989
rect 13219 953 13273 969
rect 13373 969 13383 1003
rect 13417 989 13505 1003
rect 14839 1451 14869 1477
rect 14927 1451 14957 1477
rect 15015 1451 15045 1477
rect 15103 1451 15133 1477
rect 13937 1019 13967 1050
rect 14025 1019 14055 1050
rect 14113 1019 14143 1050
rect 14201 1019 14231 1050
rect 13417 969 13427 989
rect 13373 953 13427 969
rect 13885 1003 14055 1019
rect 13885 969 13895 1003
rect 13929 989 14055 1003
rect 14107 1003 14231 1019
rect 13929 969 13939 989
rect 13885 953 13939 969
rect 14107 969 14117 1003
rect 14151 989 14231 1003
rect 14289 1019 14319 1050
rect 14377 1019 14407 1050
rect 14289 1003 14407 1019
rect 14289 989 14339 1003
rect 14151 969 14161 989
rect 14107 953 14161 969
rect 14329 969 14339 989
rect 14373 989 14407 1003
rect 15503 1451 15533 1477
rect 15591 1451 15621 1477
rect 15679 1451 15709 1477
rect 15767 1451 15797 1477
rect 14839 1020 14869 1051
rect 14927 1020 14957 1051
rect 15015 1020 15045 1051
rect 15103 1020 15133 1051
rect 14373 969 14383 989
rect 14329 953 14383 969
rect 14773 1004 14957 1020
rect 14773 970 14783 1004
rect 14817 990 14957 1004
rect 15003 1004 15133 1020
rect 14817 970 14827 990
rect 14773 954 14827 970
rect 15003 970 15013 1004
rect 15047 990 15133 1004
rect 16171 1451 16201 1477
rect 16259 1451 16289 1477
rect 16347 1451 16377 1477
rect 16435 1451 16465 1477
rect 15047 970 15057 990
rect 15003 954 15057 970
rect 15503 1020 15533 1051
rect 15591 1020 15621 1051
rect 15503 1004 15621 1020
rect 15503 990 15523 1004
rect 15513 970 15523 990
rect 15557 990 15621 1004
rect 15679 1020 15709 1051
rect 15767 1020 15797 1051
rect 15679 1004 15863 1020
rect 15679 990 15819 1004
rect 15557 970 15567 990
rect 15513 954 15567 970
rect 15809 970 15819 990
rect 15853 970 15863 1004
rect 15809 954 15863 970
rect 16171 1020 16201 1051
rect 16259 1020 16289 1051
rect 16347 1020 16377 1051
rect 16435 1020 16465 1051
rect 16105 1004 16289 1020
rect 16105 970 16115 1004
rect 16149 990 16289 1004
rect 16331 1004 16465 1020
rect 16149 970 16159 990
rect 16105 954 16159 970
rect 16331 970 16341 1004
rect 16375 990 16465 1004
rect 16375 970 16385 990
rect 16331 954 16385 970
rect 195 461 249 477
rect 195 441 205 461
rect 168 427 205 441
rect 239 427 249 461
rect 168 411 249 427
rect 343 461 397 477
rect 343 427 353 461
rect 387 427 397 461
rect 343 411 397 427
rect 861 461 915 477
rect 861 441 871 461
rect 168 377 198 411
rect 362 377 392 411
rect 813 427 871 441
rect 905 427 915 461
rect 813 411 915 427
rect 1083 461 1137 477
rect 1083 427 1093 461
rect 1127 441 1137 461
rect 1305 461 1359 477
rect 1127 427 1143 441
rect 1083 411 1143 427
rect 1305 427 1315 461
rect 1349 427 1359 461
rect 1305 411 1359 427
rect 1823 461 1877 477
rect 1823 441 1833 461
rect 813 379 843 411
rect 1113 379 1143 411
rect 1315 379 1345 411
rect 1775 427 1833 441
rect 1867 427 1877 461
rect 1775 411 1877 427
rect 2045 461 2099 477
rect 2045 427 2055 461
rect 2089 441 2099 461
rect 2267 461 2321 477
rect 2089 427 2105 441
rect 2045 411 2105 427
rect 2267 427 2277 461
rect 2311 427 2321 461
rect 2267 411 2321 427
rect 2785 461 2839 477
rect 2785 441 2795 461
rect 1775 379 1805 411
rect 2075 379 2105 411
rect 2277 379 2307 411
rect 2758 427 2795 441
rect 2829 427 2839 461
rect 2758 411 2839 427
rect 2933 461 2987 477
rect 2933 427 2943 461
rect 2977 427 2987 461
rect 2933 411 2987 427
rect 3451 461 3505 477
rect 3451 441 3461 461
rect 2758 377 2788 411
rect 2952 377 2982 411
rect 3424 427 3461 441
rect 3495 427 3505 461
rect 3424 411 3505 427
rect 3599 461 3653 477
rect 3599 427 3609 461
rect 3643 427 3653 461
rect 3599 411 3653 427
rect 4117 461 4171 477
rect 4117 441 4127 461
rect 3424 377 3454 411
rect 3618 377 3648 411
rect 4069 427 4127 441
rect 4161 427 4171 461
rect 4069 411 4171 427
rect 4339 461 4393 477
rect 4339 427 4349 461
rect 4383 441 4393 461
rect 4561 461 4615 477
rect 4383 427 4399 441
rect 4339 411 4399 427
rect 4561 427 4571 461
rect 4605 427 4615 461
rect 4561 411 4615 427
rect 5079 461 5133 477
rect 5079 441 5089 461
rect 4069 379 4099 411
rect 4369 379 4399 411
rect 4571 379 4601 411
rect 5052 427 5089 441
rect 5123 427 5133 461
rect 5052 411 5133 427
rect 5227 461 5281 477
rect 5227 427 5237 461
rect 5271 427 5281 461
rect 5227 411 5281 427
rect 5745 461 5799 477
rect 5745 441 5755 461
rect 5052 377 5082 411
rect 5246 377 5276 411
rect 5697 427 5755 441
rect 5789 427 5799 461
rect 5697 411 5799 427
rect 5967 461 6021 477
rect 5967 427 5977 461
rect 6011 441 6021 461
rect 6189 461 6243 477
rect 6011 427 6027 441
rect 5967 411 6027 427
rect 6189 427 6199 461
rect 6233 427 6243 461
rect 6189 411 6243 427
rect 6707 461 6761 477
rect 6707 441 6717 461
rect 5697 379 5727 411
rect 5997 379 6027 411
rect 6199 379 6229 411
rect 6659 427 6717 441
rect 6751 427 6761 461
rect 6659 411 6761 427
rect 6929 461 6983 477
rect 6929 427 6939 461
rect 6973 441 6983 461
rect 7151 461 7205 477
rect 6973 427 6989 441
rect 6929 411 6989 427
rect 7151 427 7161 461
rect 7195 427 7205 461
rect 7151 411 7205 427
rect 7669 461 7723 477
rect 7669 441 7679 461
rect 6659 379 6689 411
rect 6959 379 6989 411
rect 7161 379 7191 411
rect 7642 427 7679 441
rect 7713 427 7723 461
rect 7642 411 7723 427
rect 7817 461 7871 477
rect 7817 427 7827 461
rect 7861 427 7871 461
rect 7817 411 7871 427
rect 8335 461 8389 477
rect 8335 441 8345 461
rect 7642 377 7672 411
rect 7836 377 7866 411
rect 8308 427 8345 441
rect 8379 427 8389 461
rect 8308 411 8389 427
rect 8483 461 8537 477
rect 8483 427 8493 461
rect 8527 427 8537 461
rect 8483 411 8537 427
rect 9001 461 9055 477
rect 9001 441 9011 461
rect 8308 377 8338 411
rect 8502 377 8532 411
rect 8953 427 9011 441
rect 9045 427 9055 461
rect 8953 411 9055 427
rect 9223 461 9277 477
rect 9223 427 9233 461
rect 9267 441 9277 461
rect 9445 461 9499 477
rect 9267 427 9283 441
rect 9223 411 9283 427
rect 9445 427 9455 461
rect 9489 427 9499 461
rect 9445 411 9499 427
rect 9963 461 10017 477
rect 9963 441 9973 461
rect 8953 379 8983 411
rect 9253 379 9283 411
rect 9455 379 9485 411
rect 9936 427 9973 441
rect 10007 427 10017 461
rect 9936 411 10017 427
rect 10111 461 10165 477
rect 10111 427 10121 461
rect 10155 427 10165 461
rect 10111 411 10165 427
rect 10629 461 10683 477
rect 10629 441 10639 461
rect 9936 377 9966 411
rect 10130 377 10160 411
rect 10581 427 10639 441
rect 10673 427 10683 461
rect 10581 411 10683 427
rect 10851 461 10905 477
rect 10851 427 10861 461
rect 10895 441 10905 461
rect 11073 461 11127 477
rect 10895 427 10911 441
rect 10851 411 10911 427
rect 11073 427 11083 461
rect 11117 427 11127 461
rect 11073 411 11127 427
rect 11591 461 11645 477
rect 11591 441 11601 461
rect 10581 379 10611 411
rect 10881 379 10911 411
rect 11083 379 11113 411
rect 11543 427 11601 441
rect 11635 427 11645 461
rect 11543 411 11645 427
rect 11813 461 11867 477
rect 11813 427 11823 461
rect 11857 441 11867 461
rect 12035 461 12089 477
rect 11857 427 11873 441
rect 11813 411 11873 427
rect 12035 427 12045 461
rect 12079 427 12089 461
rect 12035 411 12089 427
rect 12553 461 12607 477
rect 12553 441 12563 461
rect 11543 379 11573 411
rect 11843 379 11873 411
rect 12045 379 12075 411
rect 12526 427 12563 441
rect 12597 427 12607 461
rect 12526 411 12607 427
rect 12701 461 12755 477
rect 12701 427 12711 461
rect 12745 427 12755 461
rect 12701 411 12755 427
rect 13219 461 13273 477
rect 13219 441 13229 461
rect 12526 377 12556 411
rect 12720 377 12750 411
rect 13192 427 13229 441
rect 13263 427 13273 461
rect 13192 411 13273 427
rect 13367 461 13421 477
rect 13367 427 13377 461
rect 13411 427 13421 461
rect 13367 411 13421 427
rect 13885 461 13939 477
rect 13885 441 13895 461
rect 13192 377 13222 411
rect 13386 377 13416 411
rect 13837 427 13895 441
rect 13929 427 13939 461
rect 13837 411 13939 427
rect 14107 461 14161 477
rect 14107 427 14117 461
rect 14151 441 14161 461
rect 14329 461 14383 477
rect 14151 427 14167 441
rect 14107 411 14167 427
rect 14329 427 14339 461
rect 14373 427 14383 461
rect 14329 411 14383 427
rect 13837 379 13867 411
rect 14137 379 14167 411
rect 14339 379 14369 411
rect 14773 461 14827 477
rect 14773 427 14783 461
rect 14817 441 14827 461
rect 14995 461 15049 477
rect 14817 427 14850 441
rect 14773 411 14850 427
rect 14995 427 15005 461
rect 15039 427 15049 461
rect 14995 411 15049 427
rect 15513 461 15567 477
rect 15513 441 15523 461
rect 14820 377 14850 411
rect 15014 377 15044 411
rect 15486 427 15523 441
rect 15557 427 15567 461
rect 15809 461 15863 477
rect 15809 441 15819 461
rect 15486 411 15567 427
rect 15786 427 15819 441
rect 15853 427 15863 461
rect 15786 411 15863 427
rect 15486 377 15516 411
rect 15786 377 15816 411
rect 16105 461 16159 477
rect 16105 427 16115 461
rect 16149 441 16159 461
rect 16327 461 16381 477
rect 16149 427 16182 441
rect 16105 411 16182 427
rect 16327 427 16337 461
rect 16371 427 16381 461
rect 16327 411 16381 427
rect 16152 377 16182 411
rect 16346 377 16376 411
<< polycont >>
rect 205 969 239 1003
rect 359 969 393 1003
rect 871 969 905 1003
rect 1093 969 1127 1003
rect 1315 969 1349 1003
rect 1833 969 1867 1003
rect 2055 969 2089 1003
rect 2277 969 2311 1003
rect 2795 969 2829 1003
rect 2949 969 2983 1003
rect 3461 969 3495 1003
rect 3615 969 3649 1003
rect 4127 969 4161 1003
rect 4349 969 4383 1003
rect 4571 969 4605 1003
rect 5089 969 5123 1003
rect 5243 969 5277 1003
rect 5755 969 5789 1003
rect 5977 969 6011 1003
rect 6199 969 6233 1003
rect 6717 969 6751 1003
rect 6939 969 6973 1003
rect 7161 969 7195 1003
rect 7679 969 7713 1003
rect 7833 969 7867 1003
rect 8345 969 8379 1003
rect 8499 969 8533 1003
rect 9011 969 9045 1003
rect 9233 969 9267 1003
rect 9455 969 9489 1003
rect 9973 969 10007 1003
rect 10127 969 10161 1003
rect 10639 969 10673 1003
rect 10861 969 10895 1003
rect 11083 969 11117 1003
rect 11601 969 11635 1003
rect 11823 969 11857 1003
rect 12045 969 12079 1003
rect 12563 969 12597 1003
rect 12717 969 12751 1003
rect 13229 969 13263 1003
rect 13383 969 13417 1003
rect 13895 969 13929 1003
rect 14117 969 14151 1003
rect 14339 969 14373 1003
rect 14783 970 14817 1004
rect 15013 970 15047 1004
rect 15523 970 15557 1004
rect 15819 970 15853 1004
rect 16115 970 16149 1004
rect 16341 970 16375 1004
rect 205 427 239 461
rect 353 427 387 461
rect 871 427 905 461
rect 1093 427 1127 461
rect 1315 427 1349 461
rect 1833 427 1867 461
rect 2055 427 2089 461
rect 2277 427 2311 461
rect 2795 427 2829 461
rect 2943 427 2977 461
rect 3461 427 3495 461
rect 3609 427 3643 461
rect 4127 427 4161 461
rect 4349 427 4383 461
rect 4571 427 4605 461
rect 5089 427 5123 461
rect 5237 427 5271 461
rect 5755 427 5789 461
rect 5977 427 6011 461
rect 6199 427 6233 461
rect 6717 427 6751 461
rect 6939 427 6973 461
rect 7161 427 7195 461
rect 7679 427 7713 461
rect 7827 427 7861 461
rect 8345 427 8379 461
rect 8493 427 8527 461
rect 9011 427 9045 461
rect 9233 427 9267 461
rect 9455 427 9489 461
rect 9973 427 10007 461
rect 10121 427 10155 461
rect 10639 427 10673 461
rect 10861 427 10895 461
rect 11083 427 11117 461
rect 11601 427 11635 461
rect 11823 427 11857 461
rect 12045 427 12079 461
rect 12563 427 12597 461
rect 12711 427 12745 461
rect 13229 427 13263 461
rect 13377 427 13411 461
rect 13895 427 13929 461
rect 14117 427 14151 461
rect 14339 427 14373 461
rect 14783 427 14817 461
rect 15005 427 15039 461
rect 15523 427 15557 461
rect 15819 427 15853 461
rect 16115 427 16149 461
rect 16337 427 16371 461
<< locali >>
rect -31 1539 16681 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 361 1539
rect 395 1505 433 1539
rect 467 1505 505 1539
rect 539 1505 577 1539
rect 611 1505 721 1539
rect 755 1505 793 1539
rect 827 1505 865 1539
rect 899 1505 937 1539
rect 971 1505 1009 1539
rect 1043 1505 1081 1539
rect 1115 1505 1179 1539
rect 1213 1505 1251 1539
rect 1285 1505 1323 1539
rect 1357 1505 1395 1539
rect 1429 1505 1467 1539
rect 1501 1505 1539 1539
rect 1573 1505 1683 1539
rect 1717 1505 1755 1539
rect 1789 1505 1827 1539
rect 1861 1505 1899 1539
rect 1933 1505 1971 1539
rect 2005 1505 2043 1539
rect 2077 1505 2141 1539
rect 2175 1505 2213 1539
rect 2247 1505 2285 1539
rect 2319 1505 2357 1539
rect 2391 1505 2429 1539
rect 2463 1505 2501 1539
rect 2535 1505 2645 1539
rect 2679 1505 2717 1539
rect 2751 1505 2789 1539
rect 2823 1505 2861 1539
rect 2895 1505 2951 1539
rect 2985 1505 3023 1539
rect 3057 1505 3095 1539
rect 3129 1505 3167 1539
rect 3201 1505 3311 1539
rect 3345 1505 3383 1539
rect 3417 1505 3455 1539
rect 3489 1505 3527 1539
rect 3561 1505 3617 1539
rect 3651 1505 3689 1539
rect 3723 1505 3761 1539
rect 3795 1505 3833 1539
rect 3867 1505 3977 1539
rect 4011 1505 4049 1539
rect 4083 1505 4121 1539
rect 4155 1505 4193 1539
rect 4227 1505 4265 1539
rect 4299 1505 4337 1539
rect 4371 1505 4435 1539
rect 4469 1505 4507 1539
rect 4541 1505 4579 1539
rect 4613 1505 4651 1539
rect 4685 1505 4723 1539
rect 4757 1505 4795 1539
rect 4829 1505 4939 1539
rect 4973 1505 5011 1539
rect 5045 1505 5083 1539
rect 5117 1505 5155 1539
rect 5189 1505 5245 1539
rect 5279 1505 5317 1539
rect 5351 1505 5389 1539
rect 5423 1505 5461 1539
rect 5495 1505 5605 1539
rect 5639 1505 5677 1539
rect 5711 1505 5749 1539
rect 5783 1505 5821 1539
rect 5855 1505 5893 1539
rect 5927 1505 5965 1539
rect 5999 1505 6063 1539
rect 6097 1505 6135 1539
rect 6169 1505 6207 1539
rect 6241 1505 6279 1539
rect 6313 1505 6351 1539
rect 6385 1505 6423 1539
rect 6457 1505 6567 1539
rect 6601 1505 6639 1539
rect 6673 1505 6711 1539
rect 6745 1505 6783 1539
rect 6817 1505 6855 1539
rect 6889 1505 6927 1539
rect 6961 1505 7025 1539
rect 7059 1505 7097 1539
rect 7131 1505 7169 1539
rect 7203 1505 7241 1539
rect 7275 1505 7313 1539
rect 7347 1505 7385 1539
rect 7419 1505 7529 1539
rect 7563 1505 7601 1539
rect 7635 1505 7673 1539
rect 7707 1505 7745 1539
rect 7779 1505 7835 1539
rect 7869 1505 7907 1539
rect 7941 1505 7979 1539
rect 8013 1505 8051 1539
rect 8085 1505 8195 1539
rect 8229 1505 8267 1539
rect 8301 1505 8339 1539
rect 8373 1505 8411 1539
rect 8445 1505 8501 1539
rect 8535 1505 8573 1539
rect 8607 1505 8645 1539
rect 8679 1505 8717 1539
rect 8751 1505 8861 1539
rect 8895 1505 8933 1539
rect 8967 1505 9005 1539
rect 9039 1505 9077 1539
rect 9111 1505 9149 1539
rect 9183 1505 9221 1539
rect 9255 1505 9319 1539
rect 9353 1505 9391 1539
rect 9425 1505 9463 1539
rect 9497 1505 9535 1539
rect 9569 1505 9607 1539
rect 9641 1505 9679 1539
rect 9713 1505 9823 1539
rect 9857 1505 9895 1539
rect 9929 1505 9967 1539
rect 10001 1505 10039 1539
rect 10073 1505 10129 1539
rect 10163 1505 10201 1539
rect 10235 1505 10273 1539
rect 10307 1505 10345 1539
rect 10379 1505 10489 1539
rect 10523 1505 10561 1539
rect 10595 1505 10633 1539
rect 10667 1505 10705 1539
rect 10739 1505 10777 1539
rect 10811 1505 10849 1539
rect 10883 1505 10947 1539
rect 10981 1505 11019 1539
rect 11053 1505 11091 1539
rect 11125 1505 11163 1539
rect 11197 1505 11235 1539
rect 11269 1505 11307 1539
rect 11341 1505 11451 1539
rect 11485 1505 11523 1539
rect 11557 1505 11595 1539
rect 11629 1505 11667 1539
rect 11701 1505 11739 1539
rect 11773 1505 11811 1539
rect 11845 1505 11909 1539
rect 11943 1505 11981 1539
rect 12015 1505 12053 1539
rect 12087 1505 12125 1539
rect 12159 1505 12197 1539
rect 12231 1505 12269 1539
rect 12303 1505 12413 1539
rect 12447 1505 12485 1539
rect 12519 1505 12557 1539
rect 12591 1505 12629 1539
rect 12663 1505 12719 1539
rect 12753 1505 12791 1539
rect 12825 1505 12863 1539
rect 12897 1505 12935 1539
rect 12969 1505 13079 1539
rect 13113 1505 13151 1539
rect 13185 1505 13223 1539
rect 13257 1505 13295 1539
rect 13329 1505 13385 1539
rect 13419 1505 13457 1539
rect 13491 1505 13529 1539
rect 13563 1505 13601 1539
rect 13635 1505 13745 1539
rect 13779 1505 13817 1539
rect 13851 1505 13889 1539
rect 13923 1505 13961 1539
rect 13995 1505 14033 1539
rect 14067 1505 14105 1539
rect 14139 1505 14203 1539
rect 14237 1505 14275 1539
rect 14309 1505 14347 1539
rect 14381 1505 14419 1539
rect 14453 1505 14491 1539
rect 14525 1505 14563 1539
rect 14597 1505 14707 1539
rect 14741 1505 14779 1539
rect 14813 1505 14851 1539
rect 14885 1505 14923 1539
rect 14957 1505 15013 1539
rect 15047 1505 15085 1539
rect 15119 1505 15157 1539
rect 15191 1505 15229 1539
rect 15263 1505 15373 1539
rect 15407 1505 15445 1539
rect 15479 1505 15517 1539
rect 15551 1505 15589 1539
rect 15623 1505 15679 1539
rect 15713 1505 15751 1539
rect 15785 1505 15823 1539
rect 15857 1505 15895 1539
rect 15929 1505 16039 1539
rect 16073 1505 16111 1539
rect 16145 1505 16183 1539
rect 16217 1505 16255 1539
rect 16289 1505 16345 1539
rect 16379 1505 16417 1539
rect 16451 1505 16489 1539
rect 16523 1505 16561 1539
rect 16595 1505 16681 1539
rect -31 1492 16681 1505
rect -31 1470 31 1492
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect -31 1038 31 1076
rect 141 1412 175 1492
rect 141 1344 175 1378
rect 141 1276 175 1310
rect 141 1208 175 1242
rect 141 1139 175 1174
rect 141 1073 175 1105
rect 229 1412 263 1450
rect 229 1344 263 1378
rect 229 1276 263 1310
rect 229 1208 263 1242
rect 229 1139 263 1174
rect 317 1412 351 1492
rect 317 1344 351 1378
rect 317 1276 351 1310
rect 317 1208 351 1242
rect 317 1157 351 1174
rect 405 1412 439 1450
rect 405 1344 439 1378
rect 405 1276 439 1310
rect 405 1208 439 1242
rect 229 1103 263 1105
rect 405 1139 439 1174
rect 493 1412 527 1492
rect 493 1344 527 1378
rect 493 1276 527 1310
rect 493 1208 527 1242
rect 493 1157 527 1174
rect 635 1470 697 1492
rect 635 1436 649 1470
rect 683 1436 697 1470
rect 635 1398 697 1436
rect 635 1364 649 1398
rect 683 1364 697 1398
rect 635 1326 697 1364
rect 635 1292 649 1326
rect 683 1292 697 1326
rect 635 1254 697 1292
rect 635 1220 649 1254
rect 683 1220 697 1254
rect 635 1182 697 1220
rect 405 1103 439 1105
rect 635 1148 649 1182
rect 683 1148 697 1182
rect 635 1110 697 1148
rect 229 1069 535 1103
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect -31 868 31 932
rect 205 1003 239 1019
rect 359 1003 393 1019
rect -31 546 31 572
rect -31 512 -17 546
rect 17 512 31 546
rect -31 474 31 512
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect 205 461 239 969
rect 205 411 239 427
rect 353 969 359 988
rect 353 953 393 969
rect 353 905 387 953
rect 353 461 387 871
rect 353 411 387 427
rect 501 609 535 1069
rect 635 1076 649 1110
rect 683 1076 697 1110
rect 867 1412 901 1492
rect 867 1344 901 1378
rect 867 1276 901 1310
rect 867 1208 901 1242
rect 867 1139 901 1174
rect 867 1089 901 1105
rect 955 1412 989 1450
rect 955 1344 989 1378
rect 955 1276 989 1310
rect 955 1208 989 1242
rect 955 1139 989 1174
rect 1043 1412 1077 1492
rect 1043 1344 1077 1378
rect 1043 1276 1077 1310
rect 1043 1208 1077 1242
rect 1043 1157 1077 1174
rect 1131 1412 1165 1450
rect 1131 1344 1165 1378
rect 1131 1276 1165 1310
rect 1131 1208 1165 1242
rect 955 1094 989 1105
rect 1131 1139 1165 1174
rect 1219 1412 1253 1492
rect 1219 1344 1253 1378
rect 1219 1276 1253 1310
rect 1219 1208 1253 1242
rect 1219 1157 1253 1174
rect 1307 1412 1341 1450
rect 1307 1344 1341 1378
rect 1307 1276 1341 1310
rect 1307 1208 1341 1242
rect 1131 1094 1165 1105
rect 1307 1139 1341 1174
rect 1395 1412 1429 1492
rect 1395 1344 1429 1378
rect 1395 1276 1429 1310
rect 1395 1208 1429 1242
rect 1395 1157 1429 1174
rect 1597 1470 1659 1492
rect 1597 1436 1611 1470
rect 1645 1436 1659 1470
rect 1597 1398 1659 1436
rect 1597 1364 1611 1398
rect 1645 1364 1659 1398
rect 1597 1326 1659 1364
rect 1597 1292 1611 1326
rect 1645 1292 1659 1326
rect 1597 1254 1659 1292
rect 1597 1220 1611 1254
rect 1645 1220 1659 1254
rect 1597 1182 1659 1220
rect 1307 1094 1341 1105
rect 1597 1148 1611 1182
rect 1645 1148 1659 1182
rect 1597 1110 1659 1148
rect 635 1038 697 1076
rect 955 1060 1497 1094
rect 635 1004 649 1038
rect 683 1004 697 1038
rect 635 966 697 1004
rect 635 932 649 966
rect 683 932 697 966
rect 635 868 697 932
rect 871 1003 905 1019
rect -31 368 -17 402
rect 17 368 31 402
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect 122 361 156 377
rect 316 361 350 377
rect 501 376 535 575
rect 871 608 905 969
rect 156 327 219 361
rect 253 327 316 361
rect 122 289 156 327
rect 122 221 156 255
rect 316 289 350 327
rect 122 151 156 187
rect 122 101 156 117
rect 219 236 253 252
rect -31 62 31 80
rect 219 62 253 202
rect 316 221 350 255
rect 413 342 535 376
rect 635 546 697 572
rect 635 512 649 546
rect 683 512 697 546
rect 635 474 697 512
rect 635 440 649 474
rect 683 440 697 474
rect 635 402 697 440
rect 871 461 905 574
rect 871 411 905 427
rect 1093 1003 1127 1019
rect 1093 461 1127 945
rect 1093 411 1127 427
rect 1315 1003 1349 1019
rect 1315 831 1349 969
rect 1463 921 1497 1060
rect 1462 905 1497 921
rect 1496 871 1497 905
rect 1462 855 1497 871
rect 1597 1076 1611 1110
rect 1645 1076 1659 1110
rect 1829 1412 1863 1492
rect 1829 1344 1863 1378
rect 1829 1276 1863 1310
rect 1829 1208 1863 1242
rect 1829 1139 1863 1174
rect 1829 1089 1863 1105
rect 1917 1412 1951 1450
rect 1917 1344 1951 1378
rect 1917 1276 1951 1310
rect 1917 1208 1951 1242
rect 1917 1139 1951 1174
rect 2005 1412 2039 1492
rect 2005 1344 2039 1378
rect 2005 1276 2039 1310
rect 2005 1208 2039 1242
rect 2005 1157 2039 1174
rect 2093 1412 2127 1450
rect 2093 1344 2127 1378
rect 2093 1276 2127 1310
rect 2093 1208 2127 1242
rect 1917 1094 1951 1105
rect 2093 1139 2127 1174
rect 2181 1412 2215 1492
rect 2181 1344 2215 1378
rect 2181 1276 2215 1310
rect 2181 1208 2215 1242
rect 2181 1157 2215 1174
rect 2269 1412 2303 1450
rect 2269 1344 2303 1378
rect 2269 1276 2303 1310
rect 2269 1208 2303 1242
rect 2093 1094 2127 1105
rect 2269 1139 2303 1174
rect 2357 1412 2391 1492
rect 2357 1344 2391 1378
rect 2357 1276 2391 1310
rect 2357 1208 2391 1242
rect 2357 1157 2391 1174
rect 2559 1470 2621 1492
rect 2559 1436 2573 1470
rect 2607 1436 2621 1470
rect 2559 1398 2621 1436
rect 2559 1364 2573 1398
rect 2607 1364 2621 1398
rect 2559 1326 2621 1364
rect 2559 1292 2573 1326
rect 2607 1292 2621 1326
rect 2559 1254 2621 1292
rect 2559 1220 2573 1254
rect 2607 1220 2621 1254
rect 2559 1182 2621 1220
rect 2269 1094 2303 1105
rect 2559 1148 2573 1182
rect 2607 1148 2621 1182
rect 2559 1110 2621 1148
rect 1597 1038 1659 1076
rect 1917 1060 2459 1094
rect 1597 1004 1611 1038
rect 1645 1004 1659 1038
rect 1597 966 1659 1004
rect 1597 932 1611 966
rect 1645 932 1659 966
rect 1597 868 1659 932
rect 1833 1003 1867 1019
rect 1315 461 1349 797
rect 1315 411 1349 427
rect 635 368 649 402
rect 683 368 697 402
rect 413 245 447 342
rect 635 330 697 368
rect 413 195 447 211
rect 510 289 544 305
rect 510 221 544 255
rect 316 151 350 187
rect 510 151 544 187
rect 350 117 413 151
rect 447 117 510 151
rect 316 101 350 117
rect 510 101 544 117
rect 635 296 649 330
rect 683 296 697 330
rect 635 258 697 296
rect 635 224 649 258
rect 683 224 697 258
rect 635 186 697 224
rect 635 152 649 186
rect 683 152 697 186
rect 635 114 697 152
rect 635 80 649 114
rect 683 80 697 114
rect 767 363 801 379
rect 961 363 995 379
rect 1155 363 1189 379
rect 801 329 864 363
rect 898 329 961 363
rect 995 329 1058 363
rect 1092 329 1155 363
rect 767 291 801 329
rect 767 223 801 257
rect 961 291 995 329
rect 1155 313 1189 329
rect 1269 363 1303 379
rect 1463 378 1497 855
rect 1833 609 1867 969
rect 1269 291 1303 329
rect 767 153 801 189
rect 767 103 801 119
rect 864 238 898 254
rect 635 62 697 80
rect 864 62 898 204
rect 961 223 995 257
rect 1059 244 1093 260
rect 1269 244 1303 257
rect 1093 223 1303 244
rect 1093 210 1269 223
rect 1059 194 1093 210
rect 961 153 995 189
rect 1366 344 1497 378
rect 1597 546 1659 572
rect 1597 512 1611 546
rect 1645 512 1659 546
rect 1597 474 1659 512
rect 1597 440 1611 474
rect 1645 440 1659 474
rect 1597 402 1659 440
rect 1833 461 1867 575
rect 1833 411 1867 427
rect 2055 1003 2089 1019
rect 2055 535 2089 969
rect 2055 461 2089 501
rect 2055 411 2089 427
rect 2277 1003 2311 1019
rect 2277 831 2311 969
rect 2277 461 2311 797
rect 2277 411 2311 427
rect 2425 609 2459 1060
rect 2559 1076 2573 1110
rect 2607 1076 2621 1110
rect 2559 1038 2621 1076
rect 2731 1412 2765 1492
rect 2731 1344 2765 1378
rect 2731 1276 2765 1310
rect 2731 1208 2765 1242
rect 2731 1139 2765 1174
rect 2731 1073 2765 1105
rect 2819 1412 2853 1450
rect 2819 1344 2853 1378
rect 2819 1276 2853 1310
rect 2819 1208 2853 1242
rect 2819 1139 2853 1174
rect 2907 1412 2941 1492
rect 2907 1344 2941 1378
rect 2907 1276 2941 1310
rect 2907 1208 2941 1242
rect 2907 1157 2941 1174
rect 2995 1412 3029 1450
rect 2995 1344 3029 1378
rect 2995 1276 3029 1310
rect 2995 1208 3029 1242
rect 2819 1103 2853 1105
rect 2995 1139 3029 1174
rect 3083 1412 3117 1492
rect 3083 1344 3117 1378
rect 3083 1276 3117 1310
rect 3083 1208 3117 1242
rect 3083 1157 3117 1174
rect 3225 1470 3287 1492
rect 3225 1436 3239 1470
rect 3273 1436 3287 1470
rect 3225 1398 3287 1436
rect 3225 1364 3239 1398
rect 3273 1364 3287 1398
rect 3225 1326 3287 1364
rect 3225 1292 3239 1326
rect 3273 1292 3287 1326
rect 3225 1254 3287 1292
rect 3225 1220 3239 1254
rect 3273 1220 3287 1254
rect 3225 1182 3287 1220
rect 2995 1103 3029 1105
rect 3225 1148 3239 1182
rect 3273 1148 3287 1182
rect 3225 1110 3287 1148
rect 2819 1069 3125 1103
rect 2559 1004 2573 1038
rect 2607 1004 2621 1038
rect 2559 966 2621 1004
rect 2559 932 2573 966
rect 2607 932 2621 966
rect 2559 868 2621 932
rect 2795 1003 2829 1019
rect 2949 1003 2983 1019
rect 1597 368 1611 402
rect 1645 368 1659 402
rect 1366 247 1400 344
rect 1597 330 1659 368
rect 1366 197 1400 213
rect 1463 291 1497 307
rect 1463 223 1497 257
rect 1155 153 1189 169
rect 995 119 1058 153
rect 1092 119 1155 153
rect 961 103 995 119
rect 1155 103 1189 119
rect 1269 153 1303 189
rect 1463 153 1497 189
rect 1303 119 1366 153
rect 1400 119 1463 153
rect 1269 103 1303 119
rect 1463 103 1497 119
rect 1597 296 1611 330
rect 1645 296 1659 330
rect 1597 258 1659 296
rect 1597 224 1611 258
rect 1645 224 1659 258
rect 1597 186 1659 224
rect 1597 152 1611 186
rect 1645 152 1659 186
rect 1597 114 1659 152
rect 1597 80 1611 114
rect 1645 80 1659 114
rect 1729 363 1763 379
rect 1923 363 1957 379
rect 2117 363 2151 379
rect 1763 329 1826 363
rect 1860 329 1923 363
rect 1957 329 2020 363
rect 2054 329 2117 363
rect 1729 291 1763 329
rect 1729 223 1763 257
rect 1923 291 1957 329
rect 2117 313 2151 329
rect 2231 363 2265 379
rect 2425 378 2459 575
rect 2795 609 2829 969
rect 2231 291 2265 329
rect 1729 153 1763 189
rect 1729 103 1763 119
rect 1826 238 1860 254
rect 1597 62 1659 80
rect 1826 62 1860 204
rect 1923 223 1957 257
rect 2021 244 2055 260
rect 2231 244 2265 257
rect 2055 223 2265 244
rect 2055 210 2231 223
rect 2021 194 2055 210
rect 1923 153 1957 189
rect 2328 344 2459 378
rect 2559 546 2621 572
rect 2559 512 2573 546
rect 2607 512 2621 546
rect 2559 474 2621 512
rect 2559 440 2573 474
rect 2607 440 2621 474
rect 2559 402 2621 440
rect 2795 461 2829 575
rect 2795 411 2829 427
rect 2943 979 2949 995
rect 2977 953 2983 969
rect 2943 461 2977 945
rect 2943 411 2977 427
rect 3091 831 3125 1069
rect 3225 1076 3239 1110
rect 3273 1076 3287 1110
rect 3225 1038 3287 1076
rect 3397 1412 3431 1492
rect 3397 1344 3431 1378
rect 3397 1276 3431 1310
rect 3397 1208 3431 1242
rect 3397 1139 3431 1174
rect 3397 1073 3431 1105
rect 3485 1412 3519 1450
rect 3485 1344 3519 1378
rect 3485 1276 3519 1310
rect 3485 1208 3519 1242
rect 3485 1139 3519 1174
rect 3573 1412 3607 1492
rect 3573 1344 3607 1378
rect 3573 1276 3607 1310
rect 3573 1208 3607 1242
rect 3573 1157 3607 1174
rect 3661 1412 3695 1450
rect 3661 1344 3695 1378
rect 3661 1276 3695 1310
rect 3661 1208 3695 1242
rect 3485 1103 3519 1105
rect 3661 1139 3695 1174
rect 3749 1412 3783 1492
rect 3749 1344 3783 1378
rect 3749 1276 3783 1310
rect 3749 1208 3783 1242
rect 3749 1157 3783 1174
rect 3891 1470 3953 1492
rect 3891 1436 3905 1470
rect 3939 1436 3953 1470
rect 3891 1398 3953 1436
rect 3891 1364 3905 1398
rect 3939 1364 3953 1398
rect 3891 1326 3953 1364
rect 3891 1292 3905 1326
rect 3939 1292 3953 1326
rect 3891 1254 3953 1292
rect 3891 1220 3905 1254
rect 3939 1220 3953 1254
rect 3891 1182 3953 1220
rect 3661 1103 3695 1105
rect 3891 1148 3905 1182
rect 3939 1148 3953 1182
rect 3891 1110 3953 1148
rect 3485 1069 3791 1103
rect 3225 1004 3239 1038
rect 3273 1004 3287 1038
rect 3225 966 3287 1004
rect 3225 932 3239 966
rect 3273 932 3287 966
rect 3225 868 3287 932
rect 3461 1003 3495 1019
rect 3615 1003 3649 1019
rect 3461 905 3495 969
rect 2559 368 2573 402
rect 2607 368 2621 402
rect 2328 247 2362 344
rect 2559 330 2621 368
rect 2328 197 2362 213
rect 2425 291 2459 307
rect 2425 223 2459 257
rect 2117 153 2151 169
rect 1957 119 2020 153
rect 2054 119 2117 153
rect 1923 103 1957 119
rect 2117 103 2151 119
rect 2231 153 2265 189
rect 2425 153 2459 189
rect 2265 119 2328 153
rect 2362 119 2425 153
rect 2231 103 2265 119
rect 2425 103 2459 119
rect 2559 296 2573 330
rect 2607 296 2621 330
rect 2559 258 2621 296
rect 2559 224 2573 258
rect 2607 224 2621 258
rect 2559 186 2621 224
rect 2559 152 2573 186
rect 2607 152 2621 186
rect 2559 114 2621 152
rect 2559 80 2573 114
rect 2607 80 2621 114
rect 2712 361 2746 377
rect 2906 361 2940 377
rect 3091 376 3125 797
rect 2746 327 2809 361
rect 2843 327 2906 361
rect 2712 289 2746 327
rect 2712 221 2746 255
rect 2906 289 2940 327
rect 2712 151 2746 187
rect 2712 101 2746 117
rect 2809 236 2843 252
rect 2559 62 2621 80
rect 2809 62 2843 202
rect 2906 221 2940 255
rect 3003 342 3125 376
rect 3225 546 3287 572
rect 3225 512 3239 546
rect 3273 512 3287 546
rect 3225 474 3287 512
rect 3225 440 3239 474
rect 3273 440 3287 474
rect 3225 402 3287 440
rect 3461 461 3495 871
rect 3461 411 3495 427
rect 3609 969 3615 988
rect 3609 953 3649 969
rect 3609 683 3643 953
rect 3609 461 3643 649
rect 3609 411 3643 427
rect 3757 905 3791 1069
rect 3225 368 3239 402
rect 3273 368 3287 402
rect 3003 245 3037 342
rect 3225 330 3287 368
rect 3003 195 3037 211
rect 3100 289 3134 305
rect 3100 221 3134 255
rect 2906 151 2940 187
rect 3100 151 3134 187
rect 2940 117 3003 151
rect 3037 117 3100 151
rect 2906 101 2940 117
rect 3100 101 3134 117
rect 3225 296 3239 330
rect 3273 296 3287 330
rect 3225 258 3287 296
rect 3225 224 3239 258
rect 3273 224 3287 258
rect 3225 186 3287 224
rect 3225 152 3239 186
rect 3273 152 3287 186
rect 3225 114 3287 152
rect 3225 80 3239 114
rect 3273 80 3287 114
rect 3378 361 3412 377
rect 3572 361 3606 377
rect 3757 376 3791 871
rect 3891 1076 3905 1110
rect 3939 1076 3953 1110
rect 4123 1412 4157 1492
rect 4123 1344 4157 1378
rect 4123 1276 4157 1310
rect 4123 1208 4157 1242
rect 4123 1139 4157 1174
rect 4123 1089 4157 1105
rect 4211 1412 4245 1450
rect 4211 1344 4245 1378
rect 4211 1276 4245 1310
rect 4211 1208 4245 1242
rect 4211 1139 4245 1174
rect 4299 1412 4333 1492
rect 4299 1344 4333 1378
rect 4299 1276 4333 1310
rect 4299 1208 4333 1242
rect 4299 1157 4333 1174
rect 4387 1412 4421 1450
rect 4387 1344 4421 1378
rect 4387 1276 4421 1310
rect 4387 1208 4421 1242
rect 4211 1094 4245 1105
rect 4387 1139 4421 1174
rect 4475 1412 4509 1492
rect 4475 1344 4509 1378
rect 4475 1276 4509 1310
rect 4475 1208 4509 1242
rect 4475 1157 4509 1174
rect 4563 1412 4597 1450
rect 4563 1344 4597 1378
rect 4563 1276 4597 1310
rect 4563 1208 4597 1242
rect 4387 1094 4421 1105
rect 4563 1139 4597 1174
rect 4651 1412 4685 1492
rect 4651 1344 4685 1378
rect 4651 1276 4685 1310
rect 4651 1208 4685 1242
rect 4651 1157 4685 1174
rect 4853 1470 4915 1492
rect 4853 1436 4867 1470
rect 4901 1436 4915 1470
rect 4853 1398 4915 1436
rect 4853 1364 4867 1398
rect 4901 1364 4915 1398
rect 4853 1326 4915 1364
rect 4853 1292 4867 1326
rect 4901 1292 4915 1326
rect 4853 1254 4915 1292
rect 4853 1220 4867 1254
rect 4901 1220 4915 1254
rect 4853 1182 4915 1220
rect 4563 1094 4597 1105
rect 4853 1148 4867 1182
rect 4901 1148 4915 1182
rect 4853 1110 4915 1148
rect 3891 1038 3953 1076
rect 4211 1060 4753 1094
rect 3891 1004 3905 1038
rect 3939 1004 3953 1038
rect 3891 966 3953 1004
rect 3891 932 3905 966
rect 3939 932 3953 966
rect 3891 868 3953 932
rect 4127 1003 4161 1019
rect 4127 905 4161 969
rect 3412 327 3475 361
rect 3509 327 3572 361
rect 3378 289 3412 327
rect 3378 221 3412 255
rect 3572 289 3606 327
rect 3378 151 3412 187
rect 3378 101 3412 117
rect 3475 236 3509 252
rect 3225 62 3287 80
rect 3475 62 3509 202
rect 3572 221 3606 255
rect 3669 342 3791 376
rect 3891 546 3953 572
rect 3891 512 3905 546
rect 3939 512 3953 546
rect 3891 474 3953 512
rect 3891 440 3905 474
rect 3939 440 3953 474
rect 3891 402 3953 440
rect 4127 461 4161 871
rect 4127 411 4161 427
rect 4349 1003 4383 1019
rect 4349 535 4383 969
rect 4349 461 4383 501
rect 4349 411 4383 427
rect 4571 1003 4605 1019
rect 4571 831 4605 969
rect 4571 461 4605 797
rect 4571 411 4605 427
rect 4719 683 4753 1060
rect 4853 1076 4867 1110
rect 4901 1076 4915 1110
rect 4853 1038 4915 1076
rect 5025 1412 5059 1492
rect 5025 1344 5059 1378
rect 5025 1276 5059 1310
rect 5025 1208 5059 1242
rect 5025 1139 5059 1174
rect 5025 1073 5059 1105
rect 5113 1412 5147 1450
rect 5113 1344 5147 1378
rect 5113 1276 5147 1310
rect 5113 1208 5147 1242
rect 5113 1139 5147 1174
rect 5201 1412 5235 1492
rect 5201 1344 5235 1378
rect 5201 1276 5235 1310
rect 5201 1208 5235 1242
rect 5201 1157 5235 1174
rect 5289 1412 5323 1450
rect 5289 1344 5323 1378
rect 5289 1276 5323 1310
rect 5289 1208 5323 1242
rect 5113 1103 5147 1105
rect 5289 1139 5323 1174
rect 5377 1412 5411 1492
rect 5377 1344 5411 1378
rect 5377 1276 5411 1310
rect 5377 1208 5411 1242
rect 5377 1157 5411 1174
rect 5519 1470 5581 1492
rect 5519 1436 5533 1470
rect 5567 1436 5581 1470
rect 5519 1398 5581 1436
rect 5519 1364 5533 1398
rect 5567 1364 5581 1398
rect 5519 1326 5581 1364
rect 5519 1292 5533 1326
rect 5567 1292 5581 1326
rect 5519 1254 5581 1292
rect 5519 1220 5533 1254
rect 5567 1220 5581 1254
rect 5519 1182 5581 1220
rect 5289 1103 5323 1105
rect 5519 1148 5533 1182
rect 5567 1148 5581 1182
rect 5519 1110 5581 1148
rect 5113 1069 5419 1103
rect 4853 1004 4867 1038
rect 4901 1004 4915 1038
rect 4853 966 4915 1004
rect 4853 932 4867 966
rect 4901 932 4915 966
rect 4853 868 4915 932
rect 5089 1003 5123 1019
rect 5243 1003 5277 1019
rect 3891 368 3905 402
rect 3939 368 3953 402
rect 3669 245 3703 342
rect 3891 330 3953 368
rect 3669 195 3703 211
rect 3766 289 3800 305
rect 3766 221 3800 255
rect 3572 151 3606 187
rect 3766 151 3800 187
rect 3606 117 3669 151
rect 3703 117 3766 151
rect 3572 101 3606 117
rect 3766 101 3800 117
rect 3891 296 3905 330
rect 3939 296 3953 330
rect 3891 258 3953 296
rect 3891 224 3905 258
rect 3939 224 3953 258
rect 3891 186 3953 224
rect 3891 152 3905 186
rect 3939 152 3953 186
rect 3891 114 3953 152
rect 3891 80 3905 114
rect 3939 80 3953 114
rect 4023 363 4057 379
rect 4217 363 4251 379
rect 4411 363 4445 379
rect 4057 329 4120 363
rect 4154 329 4217 363
rect 4251 329 4314 363
rect 4348 329 4411 363
rect 4023 291 4057 329
rect 4023 223 4057 257
rect 4217 291 4251 329
rect 4411 313 4445 329
rect 4525 363 4559 379
rect 4719 378 4753 649
rect 4525 291 4559 329
rect 4023 153 4057 189
rect 4023 103 4057 119
rect 4120 238 4154 254
rect 3891 62 3953 80
rect 4120 62 4154 204
rect 4217 223 4251 257
rect 4315 244 4349 260
rect 4525 244 4559 257
rect 4349 223 4559 244
rect 4349 210 4525 223
rect 4315 194 4349 210
rect 4217 153 4251 189
rect 4622 344 4753 378
rect 4853 546 4915 572
rect 4853 512 4867 546
rect 4901 512 4915 546
rect 4853 474 4915 512
rect 4853 440 4867 474
rect 4901 440 4915 474
rect 4853 402 4915 440
rect 5089 461 5123 969
rect 5089 411 5123 427
rect 5237 969 5243 988
rect 5237 953 5277 969
rect 5237 905 5271 953
rect 5237 461 5271 871
rect 5237 411 5271 427
rect 5385 609 5419 1069
rect 5519 1076 5533 1110
rect 5567 1076 5581 1110
rect 5751 1412 5785 1492
rect 5751 1344 5785 1378
rect 5751 1276 5785 1310
rect 5751 1208 5785 1242
rect 5751 1139 5785 1174
rect 5751 1089 5785 1105
rect 5839 1412 5873 1450
rect 5839 1344 5873 1378
rect 5839 1276 5873 1310
rect 5839 1208 5873 1242
rect 5839 1139 5873 1174
rect 5927 1412 5961 1492
rect 5927 1344 5961 1378
rect 5927 1276 5961 1310
rect 5927 1208 5961 1242
rect 5927 1157 5961 1174
rect 6015 1412 6049 1450
rect 6015 1344 6049 1378
rect 6015 1276 6049 1310
rect 6015 1208 6049 1242
rect 5839 1094 5873 1105
rect 6015 1139 6049 1174
rect 6103 1412 6137 1492
rect 6103 1344 6137 1378
rect 6103 1276 6137 1310
rect 6103 1208 6137 1242
rect 6103 1157 6137 1174
rect 6191 1412 6225 1450
rect 6191 1344 6225 1378
rect 6191 1276 6225 1310
rect 6191 1208 6225 1242
rect 6015 1094 6049 1105
rect 6191 1139 6225 1174
rect 6279 1412 6313 1492
rect 6279 1344 6313 1378
rect 6279 1276 6313 1310
rect 6279 1208 6313 1242
rect 6279 1157 6313 1174
rect 6481 1470 6543 1492
rect 6481 1436 6495 1470
rect 6529 1436 6543 1470
rect 6481 1398 6543 1436
rect 6481 1364 6495 1398
rect 6529 1364 6543 1398
rect 6481 1326 6543 1364
rect 6481 1292 6495 1326
rect 6529 1292 6543 1326
rect 6481 1254 6543 1292
rect 6481 1220 6495 1254
rect 6529 1220 6543 1254
rect 6481 1182 6543 1220
rect 6191 1094 6225 1105
rect 6481 1148 6495 1182
rect 6529 1148 6543 1182
rect 6481 1110 6543 1148
rect 5519 1038 5581 1076
rect 5839 1060 6381 1094
rect 5519 1004 5533 1038
rect 5567 1004 5581 1038
rect 5519 966 5581 1004
rect 5519 932 5533 966
rect 5567 932 5581 966
rect 5519 868 5581 932
rect 5755 1003 5789 1019
rect 4853 368 4867 402
rect 4901 368 4915 402
rect 4622 247 4656 344
rect 4853 330 4915 368
rect 4622 197 4656 213
rect 4719 291 4753 307
rect 4719 223 4753 257
rect 4411 153 4445 169
rect 4251 119 4314 153
rect 4348 119 4411 153
rect 4217 103 4251 119
rect 4411 103 4445 119
rect 4525 153 4559 189
rect 4719 153 4753 189
rect 4559 119 4622 153
rect 4656 119 4719 153
rect 4525 103 4559 119
rect 4719 103 4753 119
rect 4853 296 4867 330
rect 4901 296 4915 330
rect 4853 258 4915 296
rect 4853 224 4867 258
rect 4901 224 4915 258
rect 4853 186 4915 224
rect 4853 152 4867 186
rect 4901 152 4915 186
rect 4853 114 4915 152
rect 4853 80 4867 114
rect 4901 80 4915 114
rect 5006 361 5040 377
rect 5200 361 5234 377
rect 5385 376 5419 575
rect 5755 608 5789 969
rect 5040 327 5103 361
rect 5137 327 5200 361
rect 5006 289 5040 327
rect 5006 221 5040 255
rect 5200 289 5234 327
rect 5006 151 5040 187
rect 5006 101 5040 117
rect 5103 236 5137 252
rect 4853 62 4915 80
rect 5103 62 5137 202
rect 5200 221 5234 255
rect 5297 342 5419 376
rect 5519 546 5581 572
rect 5519 512 5533 546
rect 5567 512 5581 546
rect 5519 474 5581 512
rect 5519 440 5533 474
rect 5567 440 5581 474
rect 5519 402 5581 440
rect 5755 461 5789 574
rect 5755 411 5789 427
rect 5977 1003 6011 1019
rect 5977 461 6011 945
rect 5977 411 6011 427
rect 6199 1003 6233 1019
rect 6199 831 6233 969
rect 6347 921 6381 1060
rect 6346 905 6381 921
rect 6380 871 6381 905
rect 6346 855 6381 871
rect 6481 1076 6495 1110
rect 6529 1076 6543 1110
rect 6713 1412 6747 1492
rect 6713 1344 6747 1378
rect 6713 1276 6747 1310
rect 6713 1208 6747 1242
rect 6713 1139 6747 1174
rect 6713 1089 6747 1105
rect 6801 1412 6835 1450
rect 6801 1344 6835 1378
rect 6801 1276 6835 1310
rect 6801 1208 6835 1242
rect 6801 1139 6835 1174
rect 6889 1412 6923 1492
rect 6889 1344 6923 1378
rect 6889 1276 6923 1310
rect 6889 1208 6923 1242
rect 6889 1157 6923 1174
rect 6977 1412 7011 1450
rect 6977 1344 7011 1378
rect 6977 1276 7011 1310
rect 6977 1208 7011 1242
rect 6801 1094 6835 1105
rect 6977 1139 7011 1174
rect 7065 1412 7099 1492
rect 7065 1344 7099 1378
rect 7065 1276 7099 1310
rect 7065 1208 7099 1242
rect 7065 1157 7099 1174
rect 7153 1412 7187 1450
rect 7153 1344 7187 1378
rect 7153 1276 7187 1310
rect 7153 1208 7187 1242
rect 6977 1094 7011 1105
rect 7153 1139 7187 1174
rect 7241 1412 7275 1492
rect 7241 1344 7275 1378
rect 7241 1276 7275 1310
rect 7241 1208 7275 1242
rect 7241 1157 7275 1174
rect 7443 1470 7505 1492
rect 7443 1436 7457 1470
rect 7491 1436 7505 1470
rect 7443 1398 7505 1436
rect 7443 1364 7457 1398
rect 7491 1364 7505 1398
rect 7443 1326 7505 1364
rect 7443 1292 7457 1326
rect 7491 1292 7505 1326
rect 7443 1254 7505 1292
rect 7443 1220 7457 1254
rect 7491 1220 7505 1254
rect 7443 1182 7505 1220
rect 7153 1094 7187 1105
rect 7443 1148 7457 1182
rect 7491 1148 7505 1182
rect 7443 1110 7505 1148
rect 6481 1038 6543 1076
rect 6801 1060 7343 1094
rect 6481 1004 6495 1038
rect 6529 1004 6543 1038
rect 6481 966 6543 1004
rect 6481 932 6495 966
rect 6529 932 6543 966
rect 6481 868 6543 932
rect 6717 1003 6751 1019
rect 6199 461 6233 797
rect 6199 411 6233 427
rect 5519 368 5533 402
rect 5567 368 5581 402
rect 5297 245 5331 342
rect 5519 330 5581 368
rect 5297 195 5331 211
rect 5394 289 5428 305
rect 5394 221 5428 255
rect 5200 151 5234 187
rect 5394 151 5428 187
rect 5234 117 5297 151
rect 5331 117 5394 151
rect 5200 101 5234 117
rect 5394 101 5428 117
rect 5519 296 5533 330
rect 5567 296 5581 330
rect 5519 258 5581 296
rect 5519 224 5533 258
rect 5567 224 5581 258
rect 5519 186 5581 224
rect 5519 152 5533 186
rect 5567 152 5581 186
rect 5519 114 5581 152
rect 5519 80 5533 114
rect 5567 80 5581 114
rect 5651 363 5685 379
rect 5845 363 5879 379
rect 6039 363 6073 379
rect 5685 329 5748 363
rect 5782 329 5845 363
rect 5879 329 5942 363
rect 5976 329 6039 363
rect 5651 291 5685 329
rect 5651 223 5685 257
rect 5845 291 5879 329
rect 6039 313 6073 329
rect 6153 363 6187 379
rect 6347 378 6381 855
rect 6717 609 6751 969
rect 6153 291 6187 329
rect 5651 153 5685 189
rect 5651 103 5685 119
rect 5748 238 5782 254
rect 5519 62 5581 80
rect 5748 62 5782 204
rect 5845 223 5879 257
rect 5943 244 5977 260
rect 6153 244 6187 257
rect 5977 223 6187 244
rect 5977 210 6153 223
rect 5943 194 5977 210
rect 5845 153 5879 189
rect 6250 344 6381 378
rect 6481 546 6543 572
rect 6481 512 6495 546
rect 6529 512 6543 546
rect 6481 474 6543 512
rect 6481 440 6495 474
rect 6529 440 6543 474
rect 6481 402 6543 440
rect 6717 461 6751 575
rect 6717 411 6751 427
rect 6939 1003 6973 1019
rect 6939 535 6973 969
rect 6939 461 6973 501
rect 6939 411 6973 427
rect 7161 1003 7195 1019
rect 7161 831 7195 969
rect 7161 461 7195 797
rect 7161 411 7195 427
rect 7309 609 7343 1060
rect 7443 1076 7457 1110
rect 7491 1076 7505 1110
rect 7443 1038 7505 1076
rect 7615 1412 7649 1492
rect 7615 1344 7649 1378
rect 7615 1276 7649 1310
rect 7615 1208 7649 1242
rect 7615 1139 7649 1174
rect 7615 1073 7649 1105
rect 7703 1412 7737 1450
rect 7703 1344 7737 1378
rect 7703 1276 7737 1310
rect 7703 1208 7737 1242
rect 7703 1139 7737 1174
rect 7791 1412 7825 1492
rect 7791 1344 7825 1378
rect 7791 1276 7825 1310
rect 7791 1208 7825 1242
rect 7791 1157 7825 1174
rect 7879 1412 7913 1450
rect 7879 1344 7913 1378
rect 7879 1276 7913 1310
rect 7879 1208 7913 1242
rect 7703 1103 7737 1105
rect 7879 1139 7913 1174
rect 7967 1412 8001 1492
rect 7967 1344 8001 1378
rect 7967 1276 8001 1310
rect 7967 1208 8001 1242
rect 7967 1157 8001 1174
rect 8109 1470 8171 1492
rect 8109 1436 8123 1470
rect 8157 1436 8171 1470
rect 8109 1398 8171 1436
rect 8109 1364 8123 1398
rect 8157 1364 8171 1398
rect 8109 1326 8171 1364
rect 8109 1292 8123 1326
rect 8157 1292 8171 1326
rect 8109 1254 8171 1292
rect 8109 1220 8123 1254
rect 8157 1220 8171 1254
rect 8109 1182 8171 1220
rect 7879 1103 7913 1105
rect 8109 1148 8123 1182
rect 8157 1148 8171 1182
rect 8109 1110 8171 1148
rect 7703 1069 8009 1103
rect 7443 1004 7457 1038
rect 7491 1004 7505 1038
rect 7443 966 7505 1004
rect 7443 932 7457 966
rect 7491 932 7505 966
rect 7443 868 7505 932
rect 7679 1003 7713 1019
rect 7833 1003 7867 1019
rect 6481 368 6495 402
rect 6529 368 6543 402
rect 6250 247 6284 344
rect 6481 330 6543 368
rect 6250 197 6284 213
rect 6347 291 6381 307
rect 6347 223 6381 257
rect 6039 153 6073 169
rect 5879 119 5942 153
rect 5976 119 6039 153
rect 5845 103 5879 119
rect 6039 103 6073 119
rect 6153 153 6187 189
rect 6347 153 6381 189
rect 6187 119 6250 153
rect 6284 119 6347 153
rect 6153 103 6187 119
rect 6347 103 6381 119
rect 6481 296 6495 330
rect 6529 296 6543 330
rect 6481 258 6543 296
rect 6481 224 6495 258
rect 6529 224 6543 258
rect 6481 186 6543 224
rect 6481 152 6495 186
rect 6529 152 6543 186
rect 6481 114 6543 152
rect 6481 80 6495 114
rect 6529 80 6543 114
rect 6613 363 6647 379
rect 6807 363 6841 379
rect 7001 363 7035 379
rect 6647 329 6710 363
rect 6744 329 6807 363
rect 6841 329 6904 363
rect 6938 329 7001 363
rect 6613 291 6647 329
rect 6613 223 6647 257
rect 6807 291 6841 329
rect 7001 313 7035 329
rect 7115 363 7149 379
rect 7309 378 7343 575
rect 7679 609 7713 969
rect 7115 291 7149 329
rect 6613 153 6647 189
rect 6613 103 6647 119
rect 6710 238 6744 254
rect 6481 62 6543 80
rect 6710 62 6744 204
rect 6807 223 6841 257
rect 6905 244 6939 260
rect 7115 244 7149 257
rect 6939 223 7149 244
rect 6939 210 7115 223
rect 6905 194 6939 210
rect 6807 153 6841 189
rect 7212 344 7343 378
rect 7443 546 7505 572
rect 7443 512 7457 546
rect 7491 512 7505 546
rect 7443 474 7505 512
rect 7443 440 7457 474
rect 7491 440 7505 474
rect 7443 402 7505 440
rect 7679 461 7713 575
rect 7679 411 7713 427
rect 7827 979 7833 995
rect 7861 953 7867 969
rect 7827 461 7861 945
rect 7827 411 7861 427
rect 7975 831 8009 1069
rect 8109 1076 8123 1110
rect 8157 1076 8171 1110
rect 8109 1038 8171 1076
rect 8281 1412 8315 1492
rect 8281 1344 8315 1378
rect 8281 1276 8315 1310
rect 8281 1208 8315 1242
rect 8281 1139 8315 1174
rect 8281 1073 8315 1105
rect 8369 1412 8403 1450
rect 8369 1344 8403 1378
rect 8369 1276 8403 1310
rect 8369 1208 8403 1242
rect 8369 1139 8403 1174
rect 8457 1412 8491 1492
rect 8457 1344 8491 1378
rect 8457 1276 8491 1310
rect 8457 1208 8491 1242
rect 8457 1157 8491 1174
rect 8545 1412 8579 1450
rect 8545 1344 8579 1378
rect 8545 1276 8579 1310
rect 8545 1208 8579 1242
rect 8369 1103 8403 1105
rect 8545 1139 8579 1174
rect 8633 1412 8667 1492
rect 8633 1344 8667 1378
rect 8633 1276 8667 1310
rect 8633 1208 8667 1242
rect 8633 1157 8667 1174
rect 8775 1470 8837 1492
rect 8775 1436 8789 1470
rect 8823 1436 8837 1470
rect 8775 1398 8837 1436
rect 8775 1364 8789 1398
rect 8823 1364 8837 1398
rect 8775 1326 8837 1364
rect 8775 1292 8789 1326
rect 8823 1292 8837 1326
rect 8775 1254 8837 1292
rect 8775 1220 8789 1254
rect 8823 1220 8837 1254
rect 8775 1182 8837 1220
rect 8545 1103 8579 1105
rect 8775 1148 8789 1182
rect 8823 1148 8837 1182
rect 8775 1110 8837 1148
rect 8369 1069 8675 1103
rect 8109 1004 8123 1038
rect 8157 1004 8171 1038
rect 8109 966 8171 1004
rect 8109 932 8123 966
rect 8157 932 8171 966
rect 8109 868 8171 932
rect 8345 1003 8379 1019
rect 8499 1003 8533 1019
rect 8345 905 8379 969
rect 7443 368 7457 402
rect 7491 368 7505 402
rect 7212 247 7246 344
rect 7443 330 7505 368
rect 7212 197 7246 213
rect 7309 291 7343 307
rect 7309 223 7343 257
rect 7001 153 7035 169
rect 6841 119 6904 153
rect 6938 119 7001 153
rect 6807 103 6841 119
rect 7001 103 7035 119
rect 7115 153 7149 189
rect 7309 153 7343 189
rect 7149 119 7212 153
rect 7246 119 7309 153
rect 7115 103 7149 119
rect 7309 103 7343 119
rect 7443 296 7457 330
rect 7491 296 7505 330
rect 7443 258 7505 296
rect 7443 224 7457 258
rect 7491 224 7505 258
rect 7443 186 7505 224
rect 7443 152 7457 186
rect 7491 152 7505 186
rect 7443 114 7505 152
rect 7443 80 7457 114
rect 7491 80 7505 114
rect 7596 361 7630 377
rect 7790 361 7824 377
rect 7975 376 8009 797
rect 7630 327 7693 361
rect 7727 327 7790 361
rect 7596 289 7630 327
rect 7596 221 7630 255
rect 7790 289 7824 327
rect 7596 151 7630 187
rect 7596 101 7630 117
rect 7693 236 7727 252
rect 7443 62 7505 80
rect 7693 62 7727 202
rect 7790 221 7824 255
rect 7887 342 8009 376
rect 8109 546 8171 572
rect 8109 512 8123 546
rect 8157 512 8171 546
rect 8109 474 8171 512
rect 8109 440 8123 474
rect 8157 440 8171 474
rect 8109 402 8171 440
rect 8345 461 8379 871
rect 8345 411 8379 427
rect 8493 969 8499 988
rect 8493 953 8533 969
rect 8493 757 8527 953
rect 8493 461 8527 723
rect 8493 411 8527 427
rect 8641 905 8675 1069
rect 8109 368 8123 402
rect 8157 368 8171 402
rect 7887 245 7921 342
rect 8109 330 8171 368
rect 7887 195 7921 211
rect 7984 289 8018 305
rect 7984 221 8018 255
rect 7790 151 7824 187
rect 7984 151 8018 187
rect 7824 117 7887 151
rect 7921 117 7984 151
rect 7790 101 7824 117
rect 7984 101 8018 117
rect 8109 296 8123 330
rect 8157 296 8171 330
rect 8109 258 8171 296
rect 8109 224 8123 258
rect 8157 224 8171 258
rect 8109 186 8171 224
rect 8109 152 8123 186
rect 8157 152 8171 186
rect 8109 114 8171 152
rect 8109 80 8123 114
rect 8157 80 8171 114
rect 8262 361 8296 377
rect 8456 361 8490 377
rect 8641 376 8675 871
rect 8775 1076 8789 1110
rect 8823 1076 8837 1110
rect 9007 1412 9041 1492
rect 9007 1344 9041 1378
rect 9007 1276 9041 1310
rect 9007 1208 9041 1242
rect 9007 1139 9041 1174
rect 9007 1089 9041 1105
rect 9095 1412 9129 1450
rect 9095 1344 9129 1378
rect 9095 1276 9129 1310
rect 9095 1208 9129 1242
rect 9095 1139 9129 1174
rect 9183 1412 9217 1492
rect 9183 1344 9217 1378
rect 9183 1276 9217 1310
rect 9183 1208 9217 1242
rect 9183 1157 9217 1174
rect 9271 1412 9305 1450
rect 9271 1344 9305 1378
rect 9271 1276 9305 1310
rect 9271 1208 9305 1242
rect 9095 1094 9129 1105
rect 9271 1139 9305 1174
rect 9359 1412 9393 1492
rect 9359 1344 9393 1378
rect 9359 1276 9393 1310
rect 9359 1208 9393 1242
rect 9359 1157 9393 1174
rect 9447 1412 9481 1450
rect 9447 1344 9481 1378
rect 9447 1276 9481 1310
rect 9447 1208 9481 1242
rect 9271 1094 9305 1105
rect 9447 1139 9481 1174
rect 9535 1412 9569 1492
rect 9535 1344 9569 1378
rect 9535 1276 9569 1310
rect 9535 1208 9569 1242
rect 9535 1157 9569 1174
rect 9737 1470 9799 1492
rect 9737 1436 9751 1470
rect 9785 1436 9799 1470
rect 9737 1398 9799 1436
rect 9737 1364 9751 1398
rect 9785 1364 9799 1398
rect 9737 1326 9799 1364
rect 9737 1292 9751 1326
rect 9785 1292 9799 1326
rect 9737 1254 9799 1292
rect 9737 1220 9751 1254
rect 9785 1220 9799 1254
rect 9737 1182 9799 1220
rect 9447 1094 9481 1105
rect 9737 1148 9751 1182
rect 9785 1148 9799 1182
rect 9737 1110 9799 1148
rect 8775 1038 8837 1076
rect 9095 1060 9637 1094
rect 8775 1004 8789 1038
rect 8823 1004 8837 1038
rect 8775 966 8837 1004
rect 8775 932 8789 966
rect 8823 932 8837 966
rect 8775 868 8837 932
rect 9011 1003 9045 1019
rect 9011 905 9045 969
rect 8296 327 8359 361
rect 8393 327 8456 361
rect 8262 289 8296 327
rect 8262 221 8296 255
rect 8456 289 8490 327
rect 8262 151 8296 187
rect 8262 101 8296 117
rect 8359 236 8393 252
rect 8109 62 8171 80
rect 8359 62 8393 202
rect 8456 221 8490 255
rect 8553 342 8675 376
rect 8775 546 8837 572
rect 8775 512 8789 546
rect 8823 512 8837 546
rect 8775 474 8837 512
rect 8775 440 8789 474
rect 8823 440 8837 474
rect 8775 402 8837 440
rect 9011 461 9045 871
rect 9011 411 9045 427
rect 9233 1003 9267 1019
rect 9233 535 9267 969
rect 9233 461 9267 501
rect 9233 411 9267 427
rect 9455 1003 9489 1019
rect 9455 831 9489 969
rect 9455 461 9489 797
rect 9455 411 9489 427
rect 9603 757 9637 1060
rect 9737 1076 9751 1110
rect 9785 1076 9799 1110
rect 9737 1038 9799 1076
rect 9909 1412 9943 1492
rect 9909 1344 9943 1378
rect 9909 1276 9943 1310
rect 9909 1208 9943 1242
rect 9909 1139 9943 1174
rect 9909 1073 9943 1105
rect 9997 1412 10031 1450
rect 9997 1344 10031 1378
rect 9997 1276 10031 1310
rect 9997 1208 10031 1242
rect 9997 1139 10031 1174
rect 10085 1412 10119 1492
rect 10085 1344 10119 1378
rect 10085 1276 10119 1310
rect 10085 1208 10119 1242
rect 10085 1157 10119 1174
rect 10173 1412 10207 1450
rect 10173 1344 10207 1378
rect 10173 1276 10207 1310
rect 10173 1208 10207 1242
rect 9997 1103 10031 1105
rect 10173 1139 10207 1174
rect 10261 1412 10295 1492
rect 10261 1344 10295 1378
rect 10261 1276 10295 1310
rect 10261 1208 10295 1242
rect 10261 1157 10295 1174
rect 10403 1470 10465 1492
rect 10403 1436 10417 1470
rect 10451 1436 10465 1470
rect 10403 1398 10465 1436
rect 10403 1364 10417 1398
rect 10451 1364 10465 1398
rect 10403 1326 10465 1364
rect 10403 1292 10417 1326
rect 10451 1292 10465 1326
rect 10403 1254 10465 1292
rect 10403 1220 10417 1254
rect 10451 1220 10465 1254
rect 10403 1182 10465 1220
rect 10173 1103 10207 1105
rect 10403 1148 10417 1182
rect 10451 1148 10465 1182
rect 10403 1110 10465 1148
rect 9997 1069 10303 1103
rect 9737 1004 9751 1038
rect 9785 1004 9799 1038
rect 9737 966 9799 1004
rect 9737 932 9751 966
rect 9785 932 9799 966
rect 9737 868 9799 932
rect 9973 1003 10007 1019
rect 10127 1003 10161 1019
rect 8775 368 8789 402
rect 8823 368 8837 402
rect 8553 245 8587 342
rect 8775 330 8837 368
rect 8553 195 8587 211
rect 8650 289 8684 305
rect 8650 221 8684 255
rect 8456 151 8490 187
rect 8650 151 8684 187
rect 8490 117 8553 151
rect 8587 117 8650 151
rect 8456 101 8490 117
rect 8650 101 8684 117
rect 8775 296 8789 330
rect 8823 296 8837 330
rect 8775 258 8837 296
rect 8775 224 8789 258
rect 8823 224 8837 258
rect 8775 186 8837 224
rect 8775 152 8789 186
rect 8823 152 8837 186
rect 8775 114 8837 152
rect 8775 80 8789 114
rect 8823 80 8837 114
rect 8907 363 8941 379
rect 9101 363 9135 379
rect 9295 363 9329 379
rect 8941 329 9004 363
rect 9038 329 9101 363
rect 9135 329 9198 363
rect 9232 329 9295 363
rect 8907 291 8941 329
rect 8907 223 8941 257
rect 9101 291 9135 329
rect 9295 313 9329 329
rect 9409 363 9443 379
rect 9603 378 9637 723
rect 9409 291 9443 329
rect 8907 153 8941 189
rect 8907 103 8941 119
rect 9004 238 9038 254
rect 8775 62 8837 80
rect 9004 62 9038 204
rect 9101 223 9135 257
rect 9199 244 9233 260
rect 9409 244 9443 257
rect 9233 223 9443 244
rect 9233 210 9409 223
rect 9199 194 9233 210
rect 9101 153 9135 189
rect 9506 344 9637 378
rect 9737 546 9799 572
rect 9737 512 9751 546
rect 9785 512 9799 546
rect 9737 474 9799 512
rect 9737 440 9751 474
rect 9785 440 9799 474
rect 9737 402 9799 440
rect 9973 461 10007 969
rect 9973 411 10007 427
rect 10121 969 10127 988
rect 10121 953 10161 969
rect 10121 905 10155 953
rect 10121 461 10155 871
rect 10121 411 10155 427
rect 10269 609 10303 1069
rect 10403 1076 10417 1110
rect 10451 1076 10465 1110
rect 10635 1412 10669 1492
rect 10635 1344 10669 1378
rect 10635 1276 10669 1310
rect 10635 1208 10669 1242
rect 10635 1139 10669 1174
rect 10635 1089 10669 1105
rect 10723 1412 10757 1450
rect 10723 1344 10757 1378
rect 10723 1276 10757 1310
rect 10723 1208 10757 1242
rect 10723 1139 10757 1174
rect 10811 1412 10845 1492
rect 10811 1344 10845 1378
rect 10811 1276 10845 1310
rect 10811 1208 10845 1242
rect 10811 1157 10845 1174
rect 10899 1412 10933 1450
rect 10899 1344 10933 1378
rect 10899 1276 10933 1310
rect 10899 1208 10933 1242
rect 10723 1094 10757 1105
rect 10899 1139 10933 1174
rect 10987 1412 11021 1492
rect 10987 1344 11021 1378
rect 10987 1276 11021 1310
rect 10987 1208 11021 1242
rect 10987 1157 11021 1174
rect 11075 1412 11109 1450
rect 11075 1344 11109 1378
rect 11075 1276 11109 1310
rect 11075 1208 11109 1242
rect 10899 1094 10933 1105
rect 11075 1139 11109 1174
rect 11163 1412 11197 1492
rect 11163 1344 11197 1378
rect 11163 1276 11197 1310
rect 11163 1208 11197 1242
rect 11163 1157 11197 1174
rect 11365 1470 11427 1492
rect 11365 1436 11379 1470
rect 11413 1436 11427 1470
rect 11365 1398 11427 1436
rect 11365 1364 11379 1398
rect 11413 1364 11427 1398
rect 11365 1326 11427 1364
rect 11365 1292 11379 1326
rect 11413 1292 11427 1326
rect 11365 1254 11427 1292
rect 11365 1220 11379 1254
rect 11413 1220 11427 1254
rect 11365 1182 11427 1220
rect 11075 1094 11109 1105
rect 11365 1148 11379 1182
rect 11413 1148 11427 1182
rect 11365 1110 11427 1148
rect 10403 1038 10465 1076
rect 10723 1060 11265 1094
rect 10403 1004 10417 1038
rect 10451 1004 10465 1038
rect 10403 966 10465 1004
rect 10403 932 10417 966
rect 10451 932 10465 966
rect 10403 868 10465 932
rect 10639 1003 10673 1019
rect 9737 368 9751 402
rect 9785 368 9799 402
rect 9506 247 9540 344
rect 9737 330 9799 368
rect 9506 197 9540 213
rect 9603 291 9637 307
rect 9603 223 9637 257
rect 9295 153 9329 169
rect 9135 119 9198 153
rect 9232 119 9295 153
rect 9101 103 9135 119
rect 9295 103 9329 119
rect 9409 153 9443 189
rect 9603 153 9637 189
rect 9443 119 9506 153
rect 9540 119 9603 153
rect 9409 103 9443 119
rect 9603 103 9637 119
rect 9737 296 9751 330
rect 9785 296 9799 330
rect 9737 258 9799 296
rect 9737 224 9751 258
rect 9785 224 9799 258
rect 9737 186 9799 224
rect 9737 152 9751 186
rect 9785 152 9799 186
rect 9737 114 9799 152
rect 9737 80 9751 114
rect 9785 80 9799 114
rect 9890 361 9924 377
rect 10084 361 10118 377
rect 10269 376 10303 575
rect 10639 608 10673 969
rect 9924 327 9987 361
rect 10021 327 10084 361
rect 9890 289 9924 327
rect 9890 221 9924 255
rect 10084 289 10118 327
rect 9890 151 9924 187
rect 9890 101 9924 117
rect 9987 236 10021 252
rect 9737 62 9799 80
rect 9987 62 10021 202
rect 10084 221 10118 255
rect 10181 342 10303 376
rect 10403 546 10465 572
rect 10403 512 10417 546
rect 10451 512 10465 546
rect 10403 474 10465 512
rect 10403 440 10417 474
rect 10451 440 10465 474
rect 10403 402 10465 440
rect 10639 461 10673 574
rect 10639 411 10673 427
rect 10861 1003 10895 1019
rect 10861 461 10895 945
rect 10861 411 10895 427
rect 11083 1003 11117 1019
rect 11083 831 11117 969
rect 11231 921 11265 1060
rect 11230 905 11265 921
rect 11264 871 11265 905
rect 11230 855 11265 871
rect 11365 1076 11379 1110
rect 11413 1076 11427 1110
rect 11597 1412 11631 1492
rect 11597 1344 11631 1378
rect 11597 1276 11631 1310
rect 11597 1208 11631 1242
rect 11597 1139 11631 1174
rect 11597 1089 11631 1105
rect 11685 1412 11719 1450
rect 11685 1344 11719 1378
rect 11685 1276 11719 1310
rect 11685 1208 11719 1242
rect 11685 1139 11719 1174
rect 11773 1412 11807 1492
rect 11773 1344 11807 1378
rect 11773 1276 11807 1310
rect 11773 1208 11807 1242
rect 11773 1157 11807 1174
rect 11861 1412 11895 1450
rect 11861 1344 11895 1378
rect 11861 1276 11895 1310
rect 11861 1208 11895 1242
rect 11685 1094 11719 1105
rect 11861 1139 11895 1174
rect 11949 1412 11983 1492
rect 11949 1344 11983 1378
rect 11949 1276 11983 1310
rect 11949 1208 11983 1242
rect 11949 1157 11983 1174
rect 12037 1412 12071 1450
rect 12037 1344 12071 1378
rect 12037 1276 12071 1310
rect 12037 1208 12071 1242
rect 11861 1094 11895 1105
rect 12037 1139 12071 1174
rect 12125 1412 12159 1492
rect 12125 1344 12159 1378
rect 12125 1276 12159 1310
rect 12125 1208 12159 1242
rect 12125 1157 12159 1174
rect 12327 1470 12389 1492
rect 12327 1436 12341 1470
rect 12375 1436 12389 1470
rect 12327 1398 12389 1436
rect 12327 1364 12341 1398
rect 12375 1364 12389 1398
rect 12327 1326 12389 1364
rect 12327 1292 12341 1326
rect 12375 1292 12389 1326
rect 12327 1254 12389 1292
rect 12327 1220 12341 1254
rect 12375 1220 12389 1254
rect 12327 1182 12389 1220
rect 12037 1094 12071 1105
rect 12327 1148 12341 1182
rect 12375 1148 12389 1182
rect 12327 1110 12389 1148
rect 11365 1038 11427 1076
rect 11685 1060 12227 1094
rect 11365 1004 11379 1038
rect 11413 1004 11427 1038
rect 11365 966 11427 1004
rect 11365 932 11379 966
rect 11413 932 11427 966
rect 11365 868 11427 932
rect 11601 1003 11635 1019
rect 11083 461 11117 797
rect 11083 411 11117 427
rect 10403 368 10417 402
rect 10451 368 10465 402
rect 10181 245 10215 342
rect 10403 330 10465 368
rect 10181 195 10215 211
rect 10278 289 10312 305
rect 10278 221 10312 255
rect 10084 151 10118 187
rect 10278 151 10312 187
rect 10118 117 10181 151
rect 10215 117 10278 151
rect 10084 101 10118 117
rect 10278 101 10312 117
rect 10403 296 10417 330
rect 10451 296 10465 330
rect 10403 258 10465 296
rect 10403 224 10417 258
rect 10451 224 10465 258
rect 10403 186 10465 224
rect 10403 152 10417 186
rect 10451 152 10465 186
rect 10403 114 10465 152
rect 10403 80 10417 114
rect 10451 80 10465 114
rect 10535 363 10569 379
rect 10729 363 10763 379
rect 10923 363 10957 379
rect 10569 329 10632 363
rect 10666 329 10729 363
rect 10763 329 10826 363
rect 10860 329 10923 363
rect 10535 291 10569 329
rect 10535 223 10569 257
rect 10729 291 10763 329
rect 10923 313 10957 329
rect 11037 363 11071 379
rect 11231 378 11265 855
rect 11601 609 11635 969
rect 11037 291 11071 329
rect 10535 153 10569 189
rect 10535 103 10569 119
rect 10632 238 10666 254
rect 10403 62 10465 80
rect 10632 62 10666 204
rect 10729 223 10763 257
rect 10827 244 10861 260
rect 11037 244 11071 257
rect 10861 223 11071 244
rect 10861 210 11037 223
rect 10827 194 10861 210
rect 10729 153 10763 189
rect 11134 344 11265 378
rect 11365 546 11427 572
rect 11365 512 11379 546
rect 11413 512 11427 546
rect 11365 474 11427 512
rect 11365 440 11379 474
rect 11413 440 11427 474
rect 11365 402 11427 440
rect 11601 461 11635 575
rect 11601 411 11635 427
rect 11823 1003 11857 1019
rect 11823 535 11857 969
rect 11823 461 11857 501
rect 11823 411 11857 427
rect 12045 1003 12079 1019
rect 12045 831 12079 969
rect 12045 461 12079 797
rect 12045 411 12079 427
rect 12193 609 12227 1060
rect 12327 1076 12341 1110
rect 12375 1076 12389 1110
rect 12327 1038 12389 1076
rect 12499 1412 12533 1492
rect 12499 1344 12533 1378
rect 12499 1276 12533 1310
rect 12499 1208 12533 1242
rect 12499 1139 12533 1174
rect 12499 1073 12533 1105
rect 12587 1412 12621 1450
rect 12587 1344 12621 1378
rect 12587 1276 12621 1310
rect 12587 1208 12621 1242
rect 12587 1139 12621 1174
rect 12675 1412 12709 1492
rect 12675 1344 12709 1378
rect 12675 1276 12709 1310
rect 12675 1208 12709 1242
rect 12675 1157 12709 1174
rect 12763 1412 12797 1450
rect 12763 1344 12797 1378
rect 12763 1276 12797 1310
rect 12763 1208 12797 1242
rect 12587 1103 12621 1105
rect 12763 1139 12797 1174
rect 12851 1412 12885 1492
rect 12851 1344 12885 1378
rect 12851 1276 12885 1310
rect 12851 1208 12885 1242
rect 12851 1157 12885 1174
rect 12993 1470 13055 1492
rect 12993 1436 13007 1470
rect 13041 1436 13055 1470
rect 12993 1398 13055 1436
rect 12993 1364 13007 1398
rect 13041 1364 13055 1398
rect 12993 1326 13055 1364
rect 12993 1292 13007 1326
rect 13041 1292 13055 1326
rect 12993 1254 13055 1292
rect 12993 1220 13007 1254
rect 13041 1220 13055 1254
rect 12993 1182 13055 1220
rect 12763 1103 12797 1105
rect 12993 1148 13007 1182
rect 13041 1148 13055 1182
rect 12993 1110 13055 1148
rect 12587 1069 12893 1103
rect 12327 1004 12341 1038
rect 12375 1004 12389 1038
rect 12327 966 12389 1004
rect 12327 932 12341 966
rect 12375 932 12389 966
rect 12327 868 12389 932
rect 12563 1003 12597 1019
rect 12717 1003 12751 1019
rect 11365 368 11379 402
rect 11413 368 11427 402
rect 11134 247 11168 344
rect 11365 330 11427 368
rect 11134 197 11168 213
rect 11231 291 11265 307
rect 11231 223 11265 257
rect 10923 153 10957 169
rect 10763 119 10826 153
rect 10860 119 10923 153
rect 10729 103 10763 119
rect 10923 103 10957 119
rect 11037 153 11071 189
rect 11231 153 11265 189
rect 11071 119 11134 153
rect 11168 119 11231 153
rect 11037 103 11071 119
rect 11231 103 11265 119
rect 11365 296 11379 330
rect 11413 296 11427 330
rect 11365 258 11427 296
rect 11365 224 11379 258
rect 11413 224 11427 258
rect 11365 186 11427 224
rect 11365 152 11379 186
rect 11413 152 11427 186
rect 11365 114 11427 152
rect 11365 80 11379 114
rect 11413 80 11427 114
rect 11497 363 11531 379
rect 11691 363 11725 379
rect 11885 363 11919 379
rect 11531 329 11594 363
rect 11628 329 11691 363
rect 11725 329 11788 363
rect 11822 329 11885 363
rect 11497 291 11531 329
rect 11497 223 11531 257
rect 11691 291 11725 329
rect 11885 313 11919 329
rect 11999 363 12033 379
rect 12193 378 12227 575
rect 12563 609 12597 969
rect 11999 291 12033 329
rect 11497 153 11531 189
rect 11497 103 11531 119
rect 11594 238 11628 254
rect 11365 62 11427 80
rect 11594 62 11628 204
rect 11691 223 11725 257
rect 11789 244 11823 260
rect 11999 244 12033 257
rect 11823 223 12033 244
rect 11823 210 11999 223
rect 11789 194 11823 210
rect 11691 153 11725 189
rect 12096 344 12227 378
rect 12327 546 12389 572
rect 12327 512 12341 546
rect 12375 512 12389 546
rect 12327 474 12389 512
rect 12327 440 12341 474
rect 12375 440 12389 474
rect 12327 402 12389 440
rect 12563 461 12597 575
rect 12563 411 12597 427
rect 12711 979 12717 995
rect 12745 953 12751 969
rect 12711 461 12745 945
rect 12711 411 12745 427
rect 12859 831 12893 1069
rect 12993 1076 13007 1110
rect 13041 1076 13055 1110
rect 12993 1038 13055 1076
rect 13165 1412 13199 1492
rect 13165 1344 13199 1378
rect 13165 1276 13199 1310
rect 13165 1208 13199 1242
rect 13165 1139 13199 1174
rect 13165 1073 13199 1105
rect 13253 1412 13287 1450
rect 13253 1344 13287 1378
rect 13253 1276 13287 1310
rect 13253 1208 13287 1242
rect 13253 1139 13287 1174
rect 13341 1412 13375 1492
rect 13341 1344 13375 1378
rect 13341 1276 13375 1310
rect 13341 1208 13375 1242
rect 13341 1157 13375 1174
rect 13429 1412 13463 1450
rect 13429 1344 13463 1378
rect 13429 1276 13463 1310
rect 13429 1208 13463 1242
rect 13253 1103 13287 1105
rect 13429 1139 13463 1174
rect 13517 1412 13551 1492
rect 13517 1344 13551 1378
rect 13517 1276 13551 1310
rect 13517 1208 13551 1242
rect 13517 1157 13551 1174
rect 13659 1470 13721 1492
rect 13659 1436 13673 1470
rect 13707 1436 13721 1470
rect 13659 1398 13721 1436
rect 13659 1364 13673 1398
rect 13707 1364 13721 1398
rect 13659 1326 13721 1364
rect 13659 1292 13673 1326
rect 13707 1292 13721 1326
rect 13659 1254 13721 1292
rect 13659 1220 13673 1254
rect 13707 1220 13721 1254
rect 13659 1182 13721 1220
rect 13429 1103 13463 1105
rect 13659 1148 13673 1182
rect 13707 1148 13721 1182
rect 13659 1110 13721 1148
rect 13253 1069 13559 1103
rect 12993 1004 13007 1038
rect 13041 1004 13055 1038
rect 12993 966 13055 1004
rect 12993 932 13007 966
rect 13041 932 13055 966
rect 12993 868 13055 932
rect 13229 1003 13263 1019
rect 13383 1003 13417 1019
rect 13229 905 13263 969
rect 12327 368 12341 402
rect 12375 368 12389 402
rect 12096 247 12130 344
rect 12327 330 12389 368
rect 12096 197 12130 213
rect 12193 291 12227 307
rect 12193 223 12227 257
rect 11885 153 11919 169
rect 11725 119 11788 153
rect 11822 119 11885 153
rect 11691 103 11725 119
rect 11885 103 11919 119
rect 11999 153 12033 189
rect 12193 153 12227 189
rect 12033 119 12096 153
rect 12130 119 12193 153
rect 11999 103 12033 119
rect 12193 103 12227 119
rect 12327 296 12341 330
rect 12375 296 12389 330
rect 12327 258 12389 296
rect 12327 224 12341 258
rect 12375 224 12389 258
rect 12327 186 12389 224
rect 12327 152 12341 186
rect 12375 152 12389 186
rect 12327 114 12389 152
rect 12327 80 12341 114
rect 12375 80 12389 114
rect 12480 361 12514 377
rect 12674 361 12708 377
rect 12859 376 12893 797
rect 12514 327 12577 361
rect 12611 327 12674 361
rect 12480 289 12514 327
rect 12480 221 12514 255
rect 12674 289 12708 327
rect 12480 151 12514 187
rect 12480 101 12514 117
rect 12577 236 12611 252
rect 12327 62 12389 80
rect 12577 62 12611 202
rect 12674 221 12708 255
rect 12771 342 12893 376
rect 12993 546 13055 572
rect 12993 512 13007 546
rect 13041 512 13055 546
rect 12993 474 13055 512
rect 12993 440 13007 474
rect 13041 440 13055 474
rect 12993 402 13055 440
rect 13229 461 13263 871
rect 13229 411 13263 427
rect 13377 969 13383 988
rect 13377 953 13417 969
rect 13525 979 13559 1069
rect 13377 905 13411 953
rect 13377 461 13411 871
rect 13377 411 13411 427
rect 12993 368 13007 402
rect 13041 368 13055 402
rect 12771 245 12805 342
rect 12993 330 13055 368
rect 12771 195 12805 211
rect 12868 289 12902 305
rect 12868 221 12902 255
rect 12674 151 12708 187
rect 12868 151 12902 187
rect 12708 117 12771 151
rect 12805 117 12868 151
rect 12674 101 12708 117
rect 12868 101 12902 117
rect 12993 296 13007 330
rect 13041 296 13055 330
rect 12993 258 13055 296
rect 12993 224 13007 258
rect 13041 224 13055 258
rect 12993 186 13055 224
rect 12993 152 13007 186
rect 13041 152 13055 186
rect 12993 114 13055 152
rect 12993 80 13007 114
rect 13041 80 13055 114
rect 13146 361 13180 377
rect 13340 361 13374 377
rect 13525 376 13559 945
rect 13659 1076 13673 1110
rect 13707 1076 13721 1110
rect 13891 1412 13925 1492
rect 13891 1344 13925 1378
rect 13891 1276 13925 1310
rect 13891 1208 13925 1242
rect 13891 1139 13925 1174
rect 13891 1089 13925 1105
rect 13979 1412 14013 1450
rect 13979 1344 14013 1378
rect 13979 1276 14013 1310
rect 13979 1208 14013 1242
rect 13979 1139 14013 1174
rect 14067 1412 14101 1492
rect 14067 1344 14101 1378
rect 14067 1276 14101 1310
rect 14067 1208 14101 1242
rect 14067 1157 14101 1174
rect 14155 1412 14189 1450
rect 14155 1344 14189 1378
rect 14155 1276 14189 1310
rect 14155 1208 14189 1242
rect 13979 1094 14013 1105
rect 14155 1139 14189 1174
rect 14243 1412 14277 1492
rect 14243 1344 14277 1378
rect 14243 1276 14277 1310
rect 14243 1208 14277 1242
rect 14243 1157 14277 1174
rect 14331 1412 14365 1450
rect 14331 1344 14365 1378
rect 14331 1276 14365 1310
rect 14331 1208 14365 1242
rect 14155 1094 14189 1105
rect 14331 1139 14365 1174
rect 14419 1412 14453 1492
rect 14419 1344 14453 1378
rect 14419 1276 14453 1310
rect 14419 1208 14453 1242
rect 14419 1157 14453 1174
rect 14621 1470 14683 1492
rect 14621 1436 14635 1470
rect 14669 1436 14683 1470
rect 14621 1398 14683 1436
rect 14621 1364 14635 1398
rect 14669 1364 14683 1398
rect 14621 1326 14683 1364
rect 14621 1292 14635 1326
rect 14669 1292 14683 1326
rect 14621 1254 14683 1292
rect 14621 1220 14635 1254
rect 14669 1220 14683 1254
rect 14621 1182 14683 1220
rect 14331 1094 14365 1105
rect 14621 1148 14635 1182
rect 14669 1148 14683 1182
rect 14621 1110 14683 1148
rect 13659 1038 13721 1076
rect 13979 1060 14521 1094
rect 13659 1004 13673 1038
rect 13707 1004 13721 1038
rect 13659 966 13721 1004
rect 13659 932 13673 966
rect 13707 932 13721 966
rect 13659 868 13721 932
rect 13895 1003 13929 1019
rect 13180 327 13243 361
rect 13277 327 13340 361
rect 13146 289 13180 327
rect 13146 221 13180 255
rect 13340 289 13374 327
rect 13146 151 13180 187
rect 13146 101 13180 117
rect 13243 236 13277 252
rect 12993 62 13055 80
rect 13243 62 13277 202
rect 13340 221 13374 255
rect 13437 342 13559 376
rect 13659 546 13721 572
rect 13659 512 13673 546
rect 13707 512 13721 546
rect 13659 474 13721 512
rect 13659 440 13673 474
rect 13707 440 13721 474
rect 13659 402 13721 440
rect 13895 461 13929 945
rect 13895 411 13929 427
rect 14117 1003 14151 1019
rect 14117 535 14151 969
rect 14117 461 14151 501
rect 14117 411 14151 427
rect 14339 1003 14373 1019
rect 14339 831 14373 969
rect 14339 461 14373 797
rect 14339 411 14373 427
rect 14487 905 14521 1060
rect 13659 368 13673 402
rect 13707 368 13721 402
rect 13437 245 13471 342
rect 13659 330 13721 368
rect 13437 195 13471 211
rect 13534 289 13568 305
rect 13534 221 13568 255
rect 13340 151 13374 187
rect 13534 151 13568 187
rect 13374 117 13437 151
rect 13471 117 13534 151
rect 13340 101 13374 117
rect 13534 101 13568 117
rect 13659 296 13673 330
rect 13707 296 13721 330
rect 13659 258 13721 296
rect 13659 224 13673 258
rect 13707 224 13721 258
rect 13659 186 13721 224
rect 13659 152 13673 186
rect 13707 152 13721 186
rect 13659 114 13721 152
rect 13659 80 13673 114
rect 13707 80 13721 114
rect 13791 363 13825 379
rect 13985 363 14019 379
rect 14179 363 14213 379
rect 13825 329 13888 363
rect 13922 329 13985 363
rect 14019 329 14082 363
rect 14116 329 14179 363
rect 13791 291 13825 329
rect 13791 223 13825 257
rect 13985 291 14019 329
rect 14179 313 14213 329
rect 14293 363 14327 379
rect 14487 378 14521 871
rect 14621 1076 14635 1110
rect 14669 1076 14683 1110
rect 14621 1038 14683 1076
rect 14793 1411 14827 1492
rect 14793 1343 14827 1377
rect 14793 1275 14827 1309
rect 14793 1207 14827 1241
rect 14793 1139 14827 1173
rect 14793 1071 14827 1105
rect 14881 1411 14917 1445
rect 14969 1411 15003 1492
rect 14881 1343 14915 1377
rect 14881 1275 14915 1309
rect 14881 1207 14915 1241
rect 14881 1139 14915 1173
rect 14969 1343 15003 1377
rect 14969 1275 15003 1309
rect 14969 1207 15003 1241
rect 14969 1157 15003 1173
rect 15057 1411 15091 1445
rect 15057 1343 15091 1377
rect 15057 1275 15091 1309
rect 15057 1207 15091 1241
rect 15057 1105 15091 1173
rect 14881 1071 15057 1105
rect 15145 1411 15179 1492
rect 15145 1343 15179 1377
rect 15145 1275 15179 1309
rect 15145 1207 15179 1241
rect 15145 1139 15179 1173
rect 15145 1071 15179 1105
rect 15287 1470 15349 1492
rect 15287 1436 15301 1470
rect 15335 1436 15349 1470
rect 15953 1470 16015 1492
rect 15287 1398 15349 1436
rect 15287 1364 15301 1398
rect 15335 1364 15349 1398
rect 15287 1326 15349 1364
rect 15287 1292 15301 1326
rect 15335 1292 15349 1326
rect 15287 1254 15349 1292
rect 15287 1220 15301 1254
rect 15335 1220 15349 1254
rect 15287 1182 15349 1220
rect 15287 1148 15301 1182
rect 15335 1148 15349 1182
rect 15287 1110 15349 1148
rect 15287 1076 15301 1110
rect 15335 1076 15349 1110
rect 15057 1055 15091 1071
rect 14621 1004 14635 1038
rect 14669 1004 14683 1038
rect 15287 1038 15349 1076
rect 15457 1411 15843 1445
rect 15457 1343 15491 1377
rect 15457 1275 15491 1309
rect 15457 1207 15491 1241
rect 15457 1105 15491 1173
rect 15545 1343 15579 1359
rect 15545 1275 15579 1309
rect 15545 1207 15579 1241
rect 15545 1139 15579 1173
rect 15633 1343 15667 1377
rect 15633 1275 15667 1309
rect 15633 1207 15667 1241
rect 15633 1157 15667 1173
rect 15721 1343 15755 1359
rect 15721 1275 15755 1309
rect 15721 1207 15755 1241
rect 15721 1105 15755 1173
rect 15809 1343 15843 1377
rect 15809 1275 15843 1309
rect 15809 1207 15843 1241
rect 15809 1121 15843 1173
rect 15953 1436 15967 1470
rect 16001 1436 16015 1470
rect 16619 1470 16681 1492
rect 15953 1398 16015 1436
rect 15953 1364 15967 1398
rect 16001 1364 16015 1398
rect 15953 1326 16015 1364
rect 15953 1292 15967 1326
rect 16001 1292 16015 1326
rect 15953 1254 16015 1292
rect 15953 1220 15967 1254
rect 16001 1220 16015 1254
rect 15953 1182 16015 1220
rect 15953 1148 15967 1182
rect 16001 1148 16015 1182
rect 15545 1071 15721 1105
rect 15457 1055 15491 1071
rect 15721 1055 15755 1071
rect 15953 1110 16015 1148
rect 15953 1076 15967 1110
rect 16001 1076 16015 1110
rect 14621 966 14683 1004
rect 14621 932 14635 966
rect 14669 932 14683 966
rect 14621 868 14683 932
rect 14783 1004 14817 1020
rect 15013 1004 15047 1020
rect 14783 757 14817 945
rect 14293 291 14327 329
rect 13791 153 13825 189
rect 13791 103 13825 119
rect 13888 238 13922 254
rect 13659 62 13721 80
rect 13888 62 13922 204
rect 13985 223 14019 257
rect 14083 244 14117 260
rect 14293 244 14327 257
rect 14117 223 14327 244
rect 14117 210 14293 223
rect 14083 194 14117 210
rect 13985 153 14019 189
rect 14390 344 14521 378
rect 14621 546 14683 572
rect 14621 512 14635 546
rect 14669 512 14683 546
rect 14621 474 14683 512
rect 14621 440 14635 474
rect 14669 440 14683 474
rect 14621 402 14683 440
rect 14783 461 14817 723
rect 14783 411 14817 427
rect 15005 970 15013 988
rect 15005 954 15047 970
rect 15287 1004 15301 1038
rect 15335 1004 15349 1038
rect 15953 1038 16015 1076
rect 16125 1411 16511 1445
rect 16125 1343 16159 1377
rect 16125 1275 16159 1309
rect 16125 1207 16159 1241
rect 16125 1105 16159 1173
rect 16213 1343 16247 1359
rect 16213 1275 16247 1309
rect 16213 1207 16247 1241
rect 16213 1139 16247 1173
rect 16301 1343 16335 1377
rect 16301 1275 16335 1309
rect 16301 1207 16335 1241
rect 16301 1157 16335 1173
rect 16389 1343 16423 1359
rect 16389 1275 16423 1309
rect 16389 1207 16423 1241
rect 16389 1139 16423 1173
rect 16477 1343 16511 1377
rect 16477 1275 16511 1309
rect 16477 1207 16511 1241
rect 16477 1157 16511 1173
rect 16619 1436 16633 1470
rect 16667 1436 16681 1470
rect 16619 1398 16681 1436
rect 16619 1364 16633 1398
rect 16667 1364 16681 1398
rect 16619 1326 16681 1364
rect 16619 1292 16633 1326
rect 16667 1292 16681 1326
rect 16619 1254 16681 1292
rect 16619 1220 16633 1254
rect 16667 1220 16681 1254
rect 16619 1182 16681 1220
rect 16619 1148 16633 1182
rect 16667 1148 16681 1182
rect 16619 1110 16681 1148
rect 16213 1071 16519 1105
rect 16125 1055 16159 1071
rect 15287 966 15349 1004
rect 15005 905 15039 954
rect 15005 461 15039 871
rect 15287 932 15301 966
rect 15335 932 15349 966
rect 15287 868 15349 932
rect 15523 1004 15557 1020
rect 15005 411 15039 427
rect 15287 546 15349 572
rect 15287 512 15301 546
rect 15335 512 15349 546
rect 15287 474 15349 512
rect 15287 440 15301 474
rect 15335 440 15349 474
rect 14621 368 14635 402
rect 14669 368 14683 402
rect 15287 402 15349 440
rect 15523 461 15557 945
rect 15523 411 15557 427
rect 15819 1004 15853 1020
rect 15819 683 15853 970
rect 15953 1004 15967 1038
rect 16001 1004 16015 1038
rect 15953 966 16015 1004
rect 15953 932 15967 966
rect 16001 932 16015 966
rect 15953 868 16015 932
rect 16115 1004 16149 1020
rect 15819 461 15853 649
rect 15819 411 15853 427
rect 15953 546 16015 572
rect 15953 512 15967 546
rect 16001 512 16015 546
rect 15953 474 16015 512
rect 15953 440 15967 474
rect 16001 440 16015 474
rect 14390 247 14424 344
rect 14621 330 14683 368
rect 14390 197 14424 213
rect 14487 291 14521 307
rect 14487 223 14521 257
rect 14179 153 14213 169
rect 14019 119 14082 153
rect 14116 119 14179 153
rect 13985 103 14019 119
rect 14179 103 14213 119
rect 14293 153 14327 189
rect 14487 153 14521 189
rect 14327 119 14390 153
rect 14424 119 14487 153
rect 14293 103 14327 119
rect 14487 103 14521 119
rect 14621 296 14635 330
rect 14669 296 14683 330
rect 14621 258 14683 296
rect 14621 224 14635 258
rect 14669 224 14683 258
rect 14621 186 14683 224
rect 14621 152 14635 186
rect 14669 152 14683 186
rect 14621 114 14683 152
rect 14621 80 14635 114
rect 14669 80 14683 114
rect 14774 361 14808 377
rect 14968 361 15002 377
rect 14808 327 14871 361
rect 14905 327 14968 361
rect 14774 289 14808 327
rect 14774 221 14808 255
rect 14968 289 15002 327
rect 15162 361 15196 377
rect 15065 281 15099 297
rect 14774 151 14808 187
rect 14774 101 14808 117
rect 14871 236 14905 252
rect 14621 62 14683 80
rect 14871 62 14905 202
rect 14968 221 15002 255
rect 15064 247 15065 262
rect 15064 245 15099 247
rect 15098 231 15099 245
rect 15162 289 15196 327
rect 15064 195 15098 211
rect 15162 221 15196 255
rect 14968 151 15002 187
rect 15162 151 15196 187
rect 15002 117 15064 151
rect 15098 117 15162 151
rect 14968 101 15002 117
rect 15162 101 15196 117
rect 15287 368 15301 402
rect 15335 368 15349 402
rect 15953 402 16015 440
rect 16115 461 16149 970
rect 16115 411 16149 427
rect 16337 1004 16375 1020
rect 16337 970 16341 1004
rect 16337 954 16375 970
rect 16337 905 16371 954
rect 16337 461 16371 871
rect 16337 411 16371 427
rect 16485 831 16519 1071
rect 16619 1076 16633 1110
rect 16667 1076 16681 1110
rect 16619 1038 16681 1076
rect 16619 1004 16633 1038
rect 16667 1004 16681 1038
rect 16619 966 16681 1004
rect 16619 932 16633 966
rect 16667 932 16681 966
rect 16619 868 16681 932
rect 15287 330 15349 368
rect 15287 296 15301 330
rect 15335 296 15349 330
rect 15287 258 15349 296
rect 15287 224 15301 258
rect 15335 224 15349 258
rect 15287 186 15349 224
rect 15287 152 15301 186
rect 15335 152 15349 186
rect 15287 114 15349 152
rect 15287 80 15301 114
rect 15335 80 15349 114
rect 15440 361 15474 377
rect 15634 361 15668 377
rect 15474 327 15537 361
rect 15571 327 15634 361
rect 15440 289 15474 327
rect 15440 221 15474 255
rect 15634 289 15668 327
rect 15828 361 15862 377
rect 15440 151 15474 187
rect 15440 101 15474 117
rect 15537 236 15571 252
rect 15287 62 15349 80
rect 15537 62 15571 202
rect 15634 221 15668 255
rect 15731 281 15765 297
rect 15731 245 15765 247
rect 15731 195 15765 211
rect 15828 289 15862 327
rect 15828 221 15862 255
rect 15634 151 15668 187
rect 15828 151 15862 187
rect 15668 117 15731 151
rect 15765 117 15828 151
rect 15634 101 15668 117
rect 15828 101 15862 117
rect 15953 368 15967 402
rect 16001 368 16015 402
rect 15953 330 16015 368
rect 15953 296 15967 330
rect 16001 296 16015 330
rect 15953 258 16015 296
rect 15953 224 15967 258
rect 16001 224 16015 258
rect 15953 186 16015 224
rect 15953 152 15967 186
rect 16001 152 16015 186
rect 15953 114 16015 152
rect 15953 80 15967 114
rect 16001 80 16015 114
rect 16106 361 16140 377
rect 16300 361 16334 377
rect 16485 374 16519 797
rect 16140 327 16203 361
rect 16237 327 16300 361
rect 16106 289 16140 327
rect 16106 221 16140 255
rect 16300 289 16334 327
rect 16106 151 16140 187
rect 16106 101 16140 117
rect 16203 236 16237 252
rect 15953 62 16015 80
rect 16203 62 16237 202
rect 16300 221 16334 255
rect 16397 340 16519 374
rect 16619 546 16681 572
rect 16619 512 16633 546
rect 16667 512 16681 546
rect 16619 474 16681 512
rect 16619 440 16633 474
rect 16667 440 16681 474
rect 16619 402 16681 440
rect 16619 368 16633 402
rect 16667 368 16681 402
rect 16397 281 16431 340
rect 16619 330 16681 368
rect 16397 245 16431 247
rect 16397 195 16431 211
rect 16494 289 16528 306
rect 16494 221 16528 255
rect 16300 151 16334 187
rect 16494 151 16528 187
rect 16334 117 16397 151
rect 16431 117 16494 151
rect 16300 101 16334 117
rect 16494 101 16528 117
rect 16619 296 16633 330
rect 16667 296 16681 330
rect 16619 258 16681 296
rect 16619 224 16633 258
rect 16667 224 16681 258
rect 16619 186 16681 224
rect 16619 152 16633 186
rect 16667 152 16681 186
rect 16619 114 16681 152
rect 16619 80 16633 114
rect 16667 80 16681 114
rect 16619 62 16681 80
rect -31 47 15731 62
rect 15765 47 16681 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 361 47
rect 395 13 433 47
rect 467 13 505 47
rect 539 13 577 47
rect 611 13 721 47
rect 755 13 793 47
rect 827 13 865 47
rect 899 13 937 47
rect 971 13 1009 47
rect 1043 13 1081 47
rect 1115 13 1179 47
rect 1213 13 1251 47
rect 1285 13 1323 47
rect 1357 13 1395 47
rect 1429 13 1467 47
rect 1501 13 1539 47
rect 1573 13 1683 47
rect 1717 13 1755 47
rect 1789 13 1827 47
rect 1861 13 1899 47
rect 1933 13 1971 47
rect 2005 13 2043 47
rect 2077 13 2141 47
rect 2175 13 2213 47
rect 2247 13 2285 47
rect 2319 13 2357 47
rect 2391 13 2429 47
rect 2463 13 2501 47
rect 2535 13 2645 47
rect 2679 13 2717 47
rect 2751 13 2789 47
rect 2823 13 2861 47
rect 2895 13 2951 47
rect 2985 13 3023 47
rect 3057 13 3095 47
rect 3129 13 3167 47
rect 3201 13 3311 47
rect 3345 13 3383 47
rect 3417 13 3455 47
rect 3489 13 3527 47
rect 3561 13 3617 47
rect 3651 13 3689 47
rect 3723 13 3761 47
rect 3795 13 3833 47
rect 3867 13 3977 47
rect 4011 13 4049 47
rect 4083 13 4121 47
rect 4155 13 4193 47
rect 4227 13 4265 47
rect 4299 13 4337 47
rect 4371 13 4435 47
rect 4469 13 4507 47
rect 4541 13 4579 47
rect 4613 13 4651 47
rect 4685 13 4723 47
rect 4757 13 4795 47
rect 4829 13 4939 47
rect 4973 13 5011 47
rect 5045 13 5083 47
rect 5117 13 5155 47
rect 5189 13 5245 47
rect 5279 13 5317 47
rect 5351 13 5389 47
rect 5423 13 5461 47
rect 5495 13 5605 47
rect 5639 13 5677 47
rect 5711 13 5749 47
rect 5783 13 5821 47
rect 5855 13 5893 47
rect 5927 13 5965 47
rect 5999 13 6063 47
rect 6097 13 6135 47
rect 6169 13 6207 47
rect 6241 13 6279 47
rect 6313 13 6351 47
rect 6385 13 6423 47
rect 6457 13 6567 47
rect 6601 13 6639 47
rect 6673 13 6711 47
rect 6745 13 6783 47
rect 6817 13 6855 47
rect 6889 13 6927 47
rect 6961 13 7025 47
rect 7059 13 7097 47
rect 7131 13 7169 47
rect 7203 13 7241 47
rect 7275 13 7313 47
rect 7347 13 7385 47
rect 7419 13 7529 47
rect 7563 13 7601 47
rect 7635 13 7673 47
rect 7707 13 7745 47
rect 7779 13 7835 47
rect 7869 13 7907 47
rect 7941 13 7979 47
rect 8013 13 8051 47
rect 8085 13 8195 47
rect 8229 13 8267 47
rect 8301 13 8339 47
rect 8373 13 8411 47
rect 8445 13 8501 47
rect 8535 13 8573 47
rect 8607 13 8645 47
rect 8679 13 8717 47
rect 8751 13 8861 47
rect 8895 13 8933 47
rect 8967 13 9005 47
rect 9039 13 9077 47
rect 9111 13 9149 47
rect 9183 13 9221 47
rect 9255 13 9319 47
rect 9353 13 9391 47
rect 9425 13 9463 47
rect 9497 13 9535 47
rect 9569 13 9607 47
rect 9641 13 9679 47
rect 9713 13 9823 47
rect 9857 13 9895 47
rect 9929 13 9967 47
rect 10001 13 10039 47
rect 10073 13 10129 47
rect 10163 13 10201 47
rect 10235 13 10273 47
rect 10307 13 10345 47
rect 10379 13 10489 47
rect 10523 13 10561 47
rect 10595 13 10633 47
rect 10667 13 10705 47
rect 10739 13 10777 47
rect 10811 13 10849 47
rect 10883 13 10947 47
rect 10981 13 11019 47
rect 11053 13 11091 47
rect 11125 13 11163 47
rect 11197 13 11235 47
rect 11269 13 11307 47
rect 11341 13 11451 47
rect 11485 13 11523 47
rect 11557 13 11595 47
rect 11629 13 11667 47
rect 11701 13 11739 47
rect 11773 13 11811 47
rect 11845 13 11909 47
rect 11943 13 11981 47
rect 12015 13 12053 47
rect 12087 13 12125 47
rect 12159 13 12197 47
rect 12231 13 12269 47
rect 12303 13 12413 47
rect 12447 13 12485 47
rect 12519 13 12557 47
rect 12591 13 12629 47
rect 12663 13 12719 47
rect 12753 13 12791 47
rect 12825 13 12863 47
rect 12897 13 12935 47
rect 12969 13 13079 47
rect 13113 13 13151 47
rect 13185 13 13223 47
rect 13257 13 13295 47
rect 13329 13 13385 47
rect 13419 13 13457 47
rect 13491 13 13529 47
rect 13563 13 13601 47
rect 13635 13 13745 47
rect 13779 13 13817 47
rect 13851 13 13889 47
rect 13923 13 13961 47
rect 13995 13 14033 47
rect 14067 13 14105 47
rect 14139 13 14203 47
rect 14237 13 14275 47
rect 14309 13 14347 47
rect 14381 13 14419 47
rect 14453 13 14491 47
rect 14525 13 14563 47
rect 14597 13 14707 47
rect 14741 13 14779 47
rect 14813 13 14851 47
rect 14885 13 14923 47
rect 14957 13 15013 47
rect 15047 13 15085 47
rect 15119 13 15157 47
rect 15191 13 15229 47
rect 15263 13 15373 47
rect 15407 13 15445 47
rect 15479 13 15517 47
rect 15551 13 15589 47
rect 15623 13 15679 47
rect 15713 13 15751 47
rect 15785 13 15823 47
rect 15857 13 15895 47
rect 15929 13 16039 47
rect 16073 13 16111 47
rect 16145 13 16183 47
rect 16217 13 16255 47
rect 16289 13 16345 47
rect 16379 13 16417 47
rect 16451 13 16489 47
rect 16523 13 16561 47
rect 16595 13 16681 47
rect -31 0 16681 13
<< viali >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 361 1505 395 1539
rect 433 1505 467 1539
rect 505 1505 539 1539
rect 577 1505 611 1539
rect 721 1505 755 1539
rect 793 1505 827 1539
rect 865 1505 899 1539
rect 937 1505 971 1539
rect 1009 1505 1043 1539
rect 1081 1505 1115 1539
rect 1179 1505 1213 1539
rect 1251 1505 1285 1539
rect 1323 1505 1357 1539
rect 1395 1505 1429 1539
rect 1467 1505 1501 1539
rect 1539 1505 1573 1539
rect 1683 1505 1717 1539
rect 1755 1505 1789 1539
rect 1827 1505 1861 1539
rect 1899 1505 1933 1539
rect 1971 1505 2005 1539
rect 2043 1505 2077 1539
rect 2141 1505 2175 1539
rect 2213 1505 2247 1539
rect 2285 1505 2319 1539
rect 2357 1505 2391 1539
rect 2429 1505 2463 1539
rect 2501 1505 2535 1539
rect 2645 1505 2679 1539
rect 2717 1505 2751 1539
rect 2789 1505 2823 1539
rect 2861 1505 2895 1539
rect 2951 1505 2985 1539
rect 3023 1505 3057 1539
rect 3095 1505 3129 1539
rect 3167 1505 3201 1539
rect 3311 1505 3345 1539
rect 3383 1505 3417 1539
rect 3455 1505 3489 1539
rect 3527 1505 3561 1539
rect 3617 1505 3651 1539
rect 3689 1505 3723 1539
rect 3761 1505 3795 1539
rect 3833 1505 3867 1539
rect 3977 1505 4011 1539
rect 4049 1505 4083 1539
rect 4121 1505 4155 1539
rect 4193 1505 4227 1539
rect 4265 1505 4299 1539
rect 4337 1505 4371 1539
rect 4435 1505 4469 1539
rect 4507 1505 4541 1539
rect 4579 1505 4613 1539
rect 4651 1505 4685 1539
rect 4723 1505 4757 1539
rect 4795 1505 4829 1539
rect 4939 1505 4973 1539
rect 5011 1505 5045 1539
rect 5083 1505 5117 1539
rect 5155 1505 5189 1539
rect 5245 1505 5279 1539
rect 5317 1505 5351 1539
rect 5389 1505 5423 1539
rect 5461 1505 5495 1539
rect 5605 1505 5639 1539
rect 5677 1505 5711 1539
rect 5749 1505 5783 1539
rect 5821 1505 5855 1539
rect 5893 1505 5927 1539
rect 5965 1505 5999 1539
rect 6063 1505 6097 1539
rect 6135 1505 6169 1539
rect 6207 1505 6241 1539
rect 6279 1505 6313 1539
rect 6351 1505 6385 1539
rect 6423 1505 6457 1539
rect 6567 1505 6601 1539
rect 6639 1505 6673 1539
rect 6711 1505 6745 1539
rect 6783 1505 6817 1539
rect 6855 1505 6889 1539
rect 6927 1505 6961 1539
rect 7025 1505 7059 1539
rect 7097 1505 7131 1539
rect 7169 1505 7203 1539
rect 7241 1505 7275 1539
rect 7313 1505 7347 1539
rect 7385 1505 7419 1539
rect 7529 1505 7563 1539
rect 7601 1505 7635 1539
rect 7673 1505 7707 1539
rect 7745 1505 7779 1539
rect 7835 1505 7869 1539
rect 7907 1505 7941 1539
rect 7979 1505 8013 1539
rect 8051 1505 8085 1539
rect 8195 1505 8229 1539
rect 8267 1505 8301 1539
rect 8339 1505 8373 1539
rect 8411 1505 8445 1539
rect 8501 1505 8535 1539
rect 8573 1505 8607 1539
rect 8645 1505 8679 1539
rect 8717 1505 8751 1539
rect 8861 1505 8895 1539
rect 8933 1505 8967 1539
rect 9005 1505 9039 1539
rect 9077 1505 9111 1539
rect 9149 1505 9183 1539
rect 9221 1505 9255 1539
rect 9319 1505 9353 1539
rect 9391 1505 9425 1539
rect 9463 1505 9497 1539
rect 9535 1505 9569 1539
rect 9607 1505 9641 1539
rect 9679 1505 9713 1539
rect 9823 1505 9857 1539
rect 9895 1505 9929 1539
rect 9967 1505 10001 1539
rect 10039 1505 10073 1539
rect 10129 1505 10163 1539
rect 10201 1505 10235 1539
rect 10273 1505 10307 1539
rect 10345 1505 10379 1539
rect 10489 1505 10523 1539
rect 10561 1505 10595 1539
rect 10633 1505 10667 1539
rect 10705 1505 10739 1539
rect 10777 1505 10811 1539
rect 10849 1505 10883 1539
rect 10947 1505 10981 1539
rect 11019 1505 11053 1539
rect 11091 1505 11125 1539
rect 11163 1505 11197 1539
rect 11235 1505 11269 1539
rect 11307 1505 11341 1539
rect 11451 1505 11485 1539
rect 11523 1505 11557 1539
rect 11595 1505 11629 1539
rect 11667 1505 11701 1539
rect 11739 1505 11773 1539
rect 11811 1505 11845 1539
rect 11909 1505 11943 1539
rect 11981 1505 12015 1539
rect 12053 1505 12087 1539
rect 12125 1505 12159 1539
rect 12197 1505 12231 1539
rect 12269 1505 12303 1539
rect 12413 1505 12447 1539
rect 12485 1505 12519 1539
rect 12557 1505 12591 1539
rect 12629 1505 12663 1539
rect 12719 1505 12753 1539
rect 12791 1505 12825 1539
rect 12863 1505 12897 1539
rect 12935 1505 12969 1539
rect 13079 1505 13113 1539
rect 13151 1505 13185 1539
rect 13223 1505 13257 1539
rect 13295 1505 13329 1539
rect 13385 1505 13419 1539
rect 13457 1505 13491 1539
rect 13529 1505 13563 1539
rect 13601 1505 13635 1539
rect 13745 1505 13779 1539
rect 13817 1505 13851 1539
rect 13889 1505 13923 1539
rect 13961 1505 13995 1539
rect 14033 1505 14067 1539
rect 14105 1505 14139 1539
rect 14203 1505 14237 1539
rect 14275 1505 14309 1539
rect 14347 1505 14381 1539
rect 14419 1505 14453 1539
rect 14491 1505 14525 1539
rect 14563 1505 14597 1539
rect 14707 1505 14741 1539
rect 14779 1505 14813 1539
rect 14851 1505 14885 1539
rect 14923 1505 14957 1539
rect 15013 1505 15047 1539
rect 15085 1505 15119 1539
rect 15157 1505 15191 1539
rect 15229 1505 15263 1539
rect 15373 1505 15407 1539
rect 15445 1505 15479 1539
rect 15517 1505 15551 1539
rect 15589 1505 15623 1539
rect 15679 1505 15713 1539
rect 15751 1505 15785 1539
rect 15823 1505 15857 1539
rect 15895 1505 15929 1539
rect 16039 1505 16073 1539
rect 16111 1505 16145 1539
rect 16183 1505 16217 1539
rect 16255 1505 16289 1539
rect 16345 1505 16379 1539
rect 16417 1505 16451 1539
rect 16489 1505 16523 1539
rect 16561 1505 16595 1539
rect 205 427 239 461
rect 353 871 387 905
rect 501 575 535 609
rect 871 574 905 608
rect 1093 969 1127 979
rect 1093 945 1127 969
rect 1462 871 1496 905
rect 1315 797 1349 831
rect 1833 575 1867 609
rect 2055 501 2089 535
rect 2277 797 2311 831
rect 2425 575 2459 609
rect 2795 575 2829 609
rect 2943 969 2949 979
rect 2949 969 2977 979
rect 2943 945 2977 969
rect 3461 871 3495 905
rect 3091 797 3125 831
rect 3609 649 3643 683
rect 3757 871 3791 905
rect 4127 871 4161 905
rect 4349 501 4383 535
rect 4571 797 4605 831
rect 4719 649 4753 683
rect 5089 427 5123 461
rect 5237 871 5271 905
rect 5385 575 5419 609
rect 5755 574 5789 608
rect 5977 969 6011 979
rect 5977 945 6011 969
rect 6346 871 6380 905
rect 6199 797 6233 831
rect 6717 575 6751 609
rect 6939 501 6973 535
rect 7161 797 7195 831
rect 7309 575 7343 609
rect 7679 575 7713 609
rect 7827 969 7833 979
rect 7833 969 7861 979
rect 7827 945 7861 969
rect 8345 871 8379 905
rect 7975 797 8009 831
rect 8493 723 8527 757
rect 8641 871 8675 905
rect 9011 871 9045 905
rect 9233 501 9267 535
rect 9455 797 9489 831
rect 9603 723 9637 757
rect 9973 427 10007 461
rect 10121 871 10155 905
rect 10269 575 10303 609
rect 10639 574 10673 608
rect 10861 969 10895 979
rect 10861 945 10895 969
rect 11230 871 11264 905
rect 11083 797 11117 831
rect 11601 575 11635 609
rect 11823 501 11857 535
rect 12045 797 12079 831
rect 12193 575 12227 609
rect 12563 575 12597 609
rect 12711 969 12717 979
rect 12717 969 12745 979
rect 12711 945 12745 969
rect 13229 871 13263 905
rect 12859 797 12893 831
rect 13377 871 13411 905
rect 13525 945 13559 979
rect 13895 969 13929 979
rect 13895 945 13929 969
rect 14117 501 14151 535
rect 14339 797 14373 831
rect 14487 871 14521 905
rect 15057 1071 15091 1105
rect 15457 1071 15491 1105
rect 15721 1071 15755 1105
rect 14783 970 14817 979
rect 14783 945 14817 970
rect 14783 723 14817 757
rect 16125 1071 16159 1105
rect 15005 871 15039 905
rect 15523 970 15557 979
rect 15523 945 15557 970
rect 15819 649 15853 683
rect 15819 427 15853 461
rect 15065 247 15099 281
rect 16115 427 16149 461
rect 16337 871 16371 905
rect 16485 797 16519 831
rect 15731 247 15765 281
rect 16397 247 16431 281
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 361 13 395 47
rect 433 13 467 47
rect 505 13 539 47
rect 577 13 611 47
rect 721 13 755 47
rect 793 13 827 47
rect 865 13 899 47
rect 937 13 971 47
rect 1009 13 1043 47
rect 1081 13 1115 47
rect 1179 13 1213 47
rect 1251 13 1285 47
rect 1323 13 1357 47
rect 1395 13 1429 47
rect 1467 13 1501 47
rect 1539 13 1573 47
rect 1683 13 1717 47
rect 1755 13 1789 47
rect 1827 13 1861 47
rect 1899 13 1933 47
rect 1971 13 2005 47
rect 2043 13 2077 47
rect 2141 13 2175 47
rect 2213 13 2247 47
rect 2285 13 2319 47
rect 2357 13 2391 47
rect 2429 13 2463 47
rect 2501 13 2535 47
rect 2645 13 2679 47
rect 2717 13 2751 47
rect 2789 13 2823 47
rect 2861 13 2895 47
rect 2951 13 2985 47
rect 3023 13 3057 47
rect 3095 13 3129 47
rect 3167 13 3201 47
rect 3311 13 3345 47
rect 3383 13 3417 47
rect 3455 13 3489 47
rect 3527 13 3561 47
rect 3617 13 3651 47
rect 3689 13 3723 47
rect 3761 13 3795 47
rect 3833 13 3867 47
rect 3977 13 4011 47
rect 4049 13 4083 47
rect 4121 13 4155 47
rect 4193 13 4227 47
rect 4265 13 4299 47
rect 4337 13 4371 47
rect 4435 13 4469 47
rect 4507 13 4541 47
rect 4579 13 4613 47
rect 4651 13 4685 47
rect 4723 13 4757 47
rect 4795 13 4829 47
rect 4939 13 4973 47
rect 5011 13 5045 47
rect 5083 13 5117 47
rect 5155 13 5189 47
rect 5245 13 5279 47
rect 5317 13 5351 47
rect 5389 13 5423 47
rect 5461 13 5495 47
rect 5605 13 5639 47
rect 5677 13 5711 47
rect 5749 13 5783 47
rect 5821 13 5855 47
rect 5893 13 5927 47
rect 5965 13 5999 47
rect 6063 13 6097 47
rect 6135 13 6169 47
rect 6207 13 6241 47
rect 6279 13 6313 47
rect 6351 13 6385 47
rect 6423 13 6457 47
rect 6567 13 6601 47
rect 6639 13 6673 47
rect 6711 13 6745 47
rect 6783 13 6817 47
rect 6855 13 6889 47
rect 6927 13 6961 47
rect 7025 13 7059 47
rect 7097 13 7131 47
rect 7169 13 7203 47
rect 7241 13 7275 47
rect 7313 13 7347 47
rect 7385 13 7419 47
rect 7529 13 7563 47
rect 7601 13 7635 47
rect 7673 13 7707 47
rect 7745 13 7779 47
rect 7835 13 7869 47
rect 7907 13 7941 47
rect 7979 13 8013 47
rect 8051 13 8085 47
rect 8195 13 8229 47
rect 8267 13 8301 47
rect 8339 13 8373 47
rect 8411 13 8445 47
rect 8501 13 8535 47
rect 8573 13 8607 47
rect 8645 13 8679 47
rect 8717 13 8751 47
rect 8861 13 8895 47
rect 8933 13 8967 47
rect 9005 13 9039 47
rect 9077 13 9111 47
rect 9149 13 9183 47
rect 9221 13 9255 47
rect 9319 13 9353 47
rect 9391 13 9425 47
rect 9463 13 9497 47
rect 9535 13 9569 47
rect 9607 13 9641 47
rect 9679 13 9713 47
rect 9823 13 9857 47
rect 9895 13 9929 47
rect 9967 13 10001 47
rect 10039 13 10073 47
rect 10129 13 10163 47
rect 10201 13 10235 47
rect 10273 13 10307 47
rect 10345 13 10379 47
rect 10489 13 10523 47
rect 10561 13 10595 47
rect 10633 13 10667 47
rect 10705 13 10739 47
rect 10777 13 10811 47
rect 10849 13 10883 47
rect 10947 13 10981 47
rect 11019 13 11053 47
rect 11091 13 11125 47
rect 11163 13 11197 47
rect 11235 13 11269 47
rect 11307 13 11341 47
rect 11451 13 11485 47
rect 11523 13 11557 47
rect 11595 13 11629 47
rect 11667 13 11701 47
rect 11739 13 11773 47
rect 11811 13 11845 47
rect 11909 13 11943 47
rect 11981 13 12015 47
rect 12053 13 12087 47
rect 12125 13 12159 47
rect 12197 13 12231 47
rect 12269 13 12303 47
rect 12413 13 12447 47
rect 12485 13 12519 47
rect 12557 13 12591 47
rect 12629 13 12663 47
rect 12719 13 12753 47
rect 12791 13 12825 47
rect 12863 13 12897 47
rect 12935 13 12969 47
rect 13079 13 13113 47
rect 13151 13 13185 47
rect 13223 13 13257 47
rect 13295 13 13329 47
rect 13385 13 13419 47
rect 13457 13 13491 47
rect 13529 13 13563 47
rect 13601 13 13635 47
rect 13745 13 13779 47
rect 13817 13 13851 47
rect 13889 13 13923 47
rect 13961 13 13995 47
rect 14033 13 14067 47
rect 14105 13 14139 47
rect 14203 13 14237 47
rect 14275 13 14309 47
rect 14347 13 14381 47
rect 14419 13 14453 47
rect 14491 13 14525 47
rect 14563 13 14597 47
rect 14707 13 14741 47
rect 14779 13 14813 47
rect 14851 13 14885 47
rect 14923 13 14957 47
rect 15013 13 15047 47
rect 15085 13 15119 47
rect 15157 13 15191 47
rect 15229 13 15263 47
rect 15373 13 15407 47
rect 15445 13 15479 47
rect 15517 13 15551 47
rect 15589 13 15623 47
rect 15679 13 15713 47
rect 15751 13 15785 47
rect 15823 13 15857 47
rect 15895 13 15929 47
rect 16039 13 16073 47
rect 16111 13 16145 47
rect 16183 13 16217 47
rect 16255 13 16289 47
rect 16345 13 16379 47
rect 16417 13 16451 47
rect 16489 13 16523 47
rect 16561 13 16595 47
<< metal1 >>
rect -31 1539 16681 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 361 1539
rect 395 1505 433 1539
rect 467 1505 505 1539
rect 539 1505 577 1539
rect 611 1505 721 1539
rect 755 1505 793 1539
rect 827 1505 865 1539
rect 899 1505 937 1539
rect 971 1505 1009 1539
rect 1043 1505 1081 1539
rect 1115 1505 1179 1539
rect 1213 1505 1251 1539
rect 1285 1505 1323 1539
rect 1357 1505 1395 1539
rect 1429 1505 1467 1539
rect 1501 1505 1539 1539
rect 1573 1505 1683 1539
rect 1717 1505 1755 1539
rect 1789 1505 1827 1539
rect 1861 1505 1899 1539
rect 1933 1505 1971 1539
rect 2005 1505 2043 1539
rect 2077 1505 2141 1539
rect 2175 1505 2213 1539
rect 2247 1505 2285 1539
rect 2319 1505 2357 1539
rect 2391 1505 2429 1539
rect 2463 1505 2501 1539
rect 2535 1505 2645 1539
rect 2679 1505 2717 1539
rect 2751 1505 2789 1539
rect 2823 1505 2861 1539
rect 2895 1505 2951 1539
rect 2985 1505 3023 1539
rect 3057 1505 3095 1539
rect 3129 1505 3167 1539
rect 3201 1505 3311 1539
rect 3345 1505 3383 1539
rect 3417 1505 3455 1539
rect 3489 1505 3527 1539
rect 3561 1505 3617 1539
rect 3651 1505 3689 1539
rect 3723 1505 3761 1539
rect 3795 1505 3833 1539
rect 3867 1505 3977 1539
rect 4011 1505 4049 1539
rect 4083 1505 4121 1539
rect 4155 1505 4193 1539
rect 4227 1505 4265 1539
rect 4299 1505 4337 1539
rect 4371 1505 4435 1539
rect 4469 1505 4507 1539
rect 4541 1505 4579 1539
rect 4613 1505 4651 1539
rect 4685 1505 4723 1539
rect 4757 1505 4795 1539
rect 4829 1505 4939 1539
rect 4973 1505 5011 1539
rect 5045 1505 5083 1539
rect 5117 1505 5155 1539
rect 5189 1505 5245 1539
rect 5279 1505 5317 1539
rect 5351 1505 5389 1539
rect 5423 1505 5461 1539
rect 5495 1505 5605 1539
rect 5639 1505 5677 1539
rect 5711 1505 5749 1539
rect 5783 1505 5821 1539
rect 5855 1505 5893 1539
rect 5927 1505 5965 1539
rect 5999 1505 6063 1539
rect 6097 1505 6135 1539
rect 6169 1505 6207 1539
rect 6241 1505 6279 1539
rect 6313 1505 6351 1539
rect 6385 1505 6423 1539
rect 6457 1505 6567 1539
rect 6601 1505 6639 1539
rect 6673 1505 6711 1539
rect 6745 1505 6783 1539
rect 6817 1505 6855 1539
rect 6889 1505 6927 1539
rect 6961 1505 7025 1539
rect 7059 1505 7097 1539
rect 7131 1505 7169 1539
rect 7203 1505 7241 1539
rect 7275 1505 7313 1539
rect 7347 1505 7385 1539
rect 7419 1505 7529 1539
rect 7563 1505 7601 1539
rect 7635 1505 7673 1539
rect 7707 1505 7745 1539
rect 7779 1505 7835 1539
rect 7869 1505 7907 1539
rect 7941 1505 7979 1539
rect 8013 1505 8051 1539
rect 8085 1505 8195 1539
rect 8229 1505 8267 1539
rect 8301 1505 8339 1539
rect 8373 1505 8411 1539
rect 8445 1505 8501 1539
rect 8535 1505 8573 1539
rect 8607 1505 8645 1539
rect 8679 1505 8717 1539
rect 8751 1505 8861 1539
rect 8895 1505 8933 1539
rect 8967 1505 9005 1539
rect 9039 1505 9077 1539
rect 9111 1505 9149 1539
rect 9183 1505 9221 1539
rect 9255 1505 9319 1539
rect 9353 1505 9391 1539
rect 9425 1505 9463 1539
rect 9497 1505 9535 1539
rect 9569 1505 9607 1539
rect 9641 1505 9679 1539
rect 9713 1505 9823 1539
rect 9857 1505 9895 1539
rect 9929 1505 9967 1539
rect 10001 1505 10039 1539
rect 10073 1505 10129 1539
rect 10163 1505 10201 1539
rect 10235 1505 10273 1539
rect 10307 1505 10345 1539
rect 10379 1505 10489 1539
rect 10523 1505 10561 1539
rect 10595 1505 10633 1539
rect 10667 1505 10705 1539
rect 10739 1505 10777 1539
rect 10811 1505 10849 1539
rect 10883 1505 10947 1539
rect 10981 1505 11019 1539
rect 11053 1505 11091 1539
rect 11125 1505 11163 1539
rect 11197 1505 11235 1539
rect 11269 1505 11307 1539
rect 11341 1505 11451 1539
rect 11485 1505 11523 1539
rect 11557 1505 11595 1539
rect 11629 1505 11667 1539
rect 11701 1505 11739 1539
rect 11773 1505 11811 1539
rect 11845 1505 11909 1539
rect 11943 1505 11981 1539
rect 12015 1505 12053 1539
rect 12087 1505 12125 1539
rect 12159 1505 12197 1539
rect 12231 1505 12269 1539
rect 12303 1505 12413 1539
rect 12447 1505 12485 1539
rect 12519 1505 12557 1539
rect 12591 1505 12629 1539
rect 12663 1505 12719 1539
rect 12753 1505 12791 1539
rect 12825 1505 12863 1539
rect 12897 1505 12935 1539
rect 12969 1505 13079 1539
rect 13113 1505 13151 1539
rect 13185 1505 13223 1539
rect 13257 1505 13295 1539
rect 13329 1505 13385 1539
rect 13419 1505 13457 1539
rect 13491 1505 13529 1539
rect 13563 1505 13601 1539
rect 13635 1505 13745 1539
rect 13779 1505 13817 1539
rect 13851 1505 13889 1539
rect 13923 1505 13961 1539
rect 13995 1505 14033 1539
rect 14067 1505 14105 1539
rect 14139 1505 14203 1539
rect 14237 1505 14275 1539
rect 14309 1505 14347 1539
rect 14381 1505 14419 1539
rect 14453 1505 14491 1539
rect 14525 1505 14563 1539
rect 14597 1505 14707 1539
rect 14741 1505 14779 1539
rect 14813 1505 14851 1539
rect 14885 1505 14923 1539
rect 14957 1505 15013 1539
rect 15047 1505 15085 1539
rect 15119 1505 15157 1539
rect 15191 1505 15229 1539
rect 15263 1505 15373 1539
rect 15407 1505 15445 1539
rect 15479 1505 15517 1539
rect 15551 1505 15589 1539
rect 15623 1505 15679 1539
rect 15713 1505 15751 1539
rect 15785 1505 15823 1539
rect 15857 1505 15895 1539
rect 15929 1505 16039 1539
rect 16073 1505 16111 1539
rect 16145 1505 16183 1539
rect 16217 1505 16255 1539
rect 16289 1505 16345 1539
rect 16379 1505 16417 1539
rect 16451 1505 16489 1539
rect 16523 1505 16561 1539
rect 16595 1505 16681 1539
rect -31 1492 16681 1505
rect 15051 1105 15097 1111
rect 15451 1105 15497 1111
rect 15715 1105 15761 1111
rect 16119 1105 16165 1111
rect 15045 1071 15057 1105
rect 15091 1071 15457 1105
rect 15491 1071 15503 1105
rect 15709 1071 15721 1105
rect 15755 1071 16125 1105
rect 16159 1071 16171 1105
rect 15051 1065 15097 1071
rect 15451 1065 15497 1071
rect 15715 1065 15761 1071
rect 16119 1065 16165 1071
rect 1087 979 1133 985
rect 2937 979 2983 985
rect 5971 979 6017 985
rect 7821 979 7867 985
rect 10855 979 10901 985
rect 12705 979 12751 985
rect 13519 979 13565 985
rect 13889 979 13935 985
rect 14777 979 14823 985
rect 15517 979 15563 985
rect 1081 945 1093 979
rect 1127 945 2943 979
rect 2977 945 5977 979
rect 6011 945 7827 979
rect 7861 945 10861 979
rect 10895 945 12711 979
rect 12745 945 12757 979
rect 13513 945 13525 979
rect 13559 945 13895 979
rect 13929 945 13941 979
rect 14771 945 14783 979
rect 14817 945 15523 979
rect 15557 945 15569 979
rect 1087 939 1133 945
rect 2937 939 2983 945
rect 5971 939 6017 945
rect 7821 939 7867 945
rect 10855 939 10901 945
rect 12705 939 12751 945
rect 13519 939 13565 945
rect 13889 939 13935 945
rect 14777 939 14823 945
rect 15517 939 15563 945
rect 347 905 393 911
rect 1456 905 1502 911
rect 3455 905 3501 911
rect 3751 905 3797 911
rect 4121 905 4167 911
rect 5231 905 5277 911
rect 6340 905 6386 911
rect 8339 905 8385 911
rect 8635 905 8681 911
rect 9005 905 9051 911
rect 10115 905 10161 911
rect 11224 905 11270 911
rect 13223 905 13269 911
rect 13371 905 13417 911
rect 14481 905 14527 911
rect 14999 905 15045 911
rect 16331 905 16377 911
rect 341 871 353 905
rect 387 871 1462 905
rect 1496 871 3461 905
rect 3495 871 3507 905
rect 3745 871 3757 905
rect 3791 871 4127 905
rect 4161 871 4173 905
rect 5225 871 5237 905
rect 5271 871 6346 905
rect 6380 871 8345 905
rect 8379 871 8391 905
rect 8629 871 8641 905
rect 8675 871 9011 905
rect 9045 871 9057 905
rect 10109 871 10121 905
rect 10155 871 11230 905
rect 11264 871 13229 905
rect 13263 871 13275 905
rect 13365 871 13377 905
rect 13411 871 14487 905
rect 14521 871 15005 905
rect 15039 871 16337 905
rect 16371 871 16383 905
rect 347 865 393 871
rect 1456 865 1502 871
rect 3455 865 3501 871
rect 3751 865 3797 871
rect 4121 865 4167 871
rect 5231 865 5277 871
rect 6340 865 6386 871
rect 8339 865 8385 871
rect 8635 865 8681 871
rect 9005 865 9051 871
rect 10115 865 10161 871
rect 11224 865 11270 871
rect 13223 865 13269 871
rect 13371 865 13417 871
rect 14481 865 14527 871
rect 14999 865 15045 871
rect 16331 865 16377 871
rect 1309 831 1355 837
rect 2271 831 2317 837
rect 3085 831 3131 837
rect 4565 831 4611 837
rect 6193 831 6239 837
rect 7155 831 7201 837
rect 7969 831 8015 837
rect 9449 831 9495 837
rect 11077 831 11123 837
rect 12039 831 12085 837
rect 12853 831 12899 837
rect 14333 831 14379 837
rect 16479 831 16525 837
rect 1303 797 1315 831
rect 1349 797 2277 831
rect 2311 797 3091 831
rect 3125 797 4571 831
rect 4605 797 4617 831
rect 6187 797 6199 831
rect 6233 797 7161 831
rect 7195 797 7975 831
rect 8009 797 9455 831
rect 9489 797 9501 831
rect 11071 797 11083 831
rect 11117 797 12045 831
rect 12079 797 12859 831
rect 12893 797 14339 831
rect 14373 797 14385 831
rect 16473 797 16485 831
rect 16519 797 16555 831
rect 1309 791 1355 797
rect 2271 791 2317 797
rect 3085 791 3131 797
rect 4565 791 4611 797
rect 6193 791 6239 797
rect 7155 791 7201 797
rect 7969 791 8015 797
rect 9449 791 9495 797
rect 11077 791 11123 797
rect 12039 791 12085 797
rect 12853 791 12899 797
rect 14333 791 14379 797
rect 16479 791 16525 797
rect 8487 757 8533 763
rect 9597 757 9643 763
rect 14777 757 14823 763
rect 8481 723 8493 757
rect 8527 723 9603 757
rect 9637 723 14783 757
rect 14817 723 14829 757
rect 8487 717 8533 723
rect 9597 717 9643 723
rect 14777 717 14823 723
rect 3603 683 3649 689
rect 4713 683 4759 689
rect 15813 683 15859 689
rect 3597 649 3609 683
rect 3643 649 4719 683
rect 4753 649 15819 683
rect 15853 649 15865 683
rect 3603 643 3649 649
rect 4713 643 4759 649
rect 15813 643 15859 649
rect 495 609 541 615
rect 865 609 911 614
rect 1827 609 1873 615
rect 2419 609 2465 615
rect 2789 609 2835 615
rect 5379 609 5425 615
rect 5749 609 5795 614
rect 6711 609 6757 615
rect 7303 609 7349 615
rect 7673 609 7719 615
rect 10263 609 10309 615
rect 10633 609 10679 614
rect 11595 609 11641 615
rect 12187 609 12233 615
rect 12557 609 12603 615
rect 489 575 501 609
rect 535 608 1833 609
rect 535 575 871 608
rect 495 569 541 575
rect 859 574 871 575
rect 905 575 1833 608
rect 1867 575 1879 609
rect 2413 575 2425 609
rect 2459 575 2795 609
rect 2829 575 2841 609
rect 5373 575 5385 609
rect 5419 608 6717 609
rect 5419 575 5755 608
rect 905 574 941 575
rect 865 568 911 574
rect 1827 569 1873 575
rect 2419 569 2465 575
rect 2789 569 2835 575
rect 5379 569 5425 575
rect 5743 574 5755 575
rect 5789 575 6717 608
rect 6751 575 6763 609
rect 7297 575 7309 609
rect 7343 575 7679 609
rect 7713 575 7725 609
rect 10257 575 10269 609
rect 10303 608 11601 609
rect 10303 575 10639 608
rect 5789 574 5825 575
rect 5749 568 5795 574
rect 6711 569 6757 575
rect 7303 569 7349 575
rect 7673 569 7719 575
rect 10263 569 10309 575
rect 10627 574 10639 575
rect 10673 575 11601 608
rect 11635 575 11647 609
rect 12181 575 12193 609
rect 12227 575 12563 609
rect 12597 575 12609 609
rect 10673 574 10709 575
rect 10633 568 10679 574
rect 11595 569 11641 575
rect 12187 569 12233 575
rect 12557 569 12603 575
rect 2049 535 2095 541
rect 4343 535 4389 541
rect 6933 535 6979 541
rect 9227 535 9273 541
rect 11817 535 11863 541
rect 14111 535 14157 541
rect 2043 501 2055 535
rect 2089 501 4349 535
rect 4383 501 6939 535
rect 6973 501 9233 535
rect 9267 501 11823 535
rect 11857 501 14117 535
rect 14151 501 14163 535
rect 2049 495 2095 501
rect 4343 495 4389 501
rect 6933 495 6979 501
rect 9227 495 9273 501
rect 11817 495 11863 501
rect 14111 495 14157 501
rect 199 461 245 467
rect 5083 461 5129 467
rect 9967 461 10013 467
rect 15813 461 15859 467
rect 16109 461 16155 467
rect 193 427 205 461
rect 239 427 5089 461
rect 5123 427 9973 461
rect 10007 427 10019 461
rect 15807 427 15819 461
rect 15853 427 16115 461
rect 16149 427 16161 461
rect 199 421 245 427
rect 5083 421 5129 427
rect 9967 421 10013 427
rect 15813 421 15859 427
rect 16109 421 16155 427
rect 15059 281 15105 287
rect 15725 281 15771 287
rect 16391 281 16437 287
rect 15053 247 15065 281
rect 15099 247 15731 281
rect 15765 247 16397 281
rect 16431 247 16443 281
rect 15059 241 15105 247
rect 15725 241 15771 247
rect 16391 241 16437 247
rect -31 47 16681 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 361 47
rect 395 13 433 47
rect 467 13 505 47
rect 539 13 577 47
rect 611 13 721 47
rect 755 13 793 47
rect 827 13 865 47
rect 899 13 937 47
rect 971 13 1009 47
rect 1043 13 1081 47
rect 1115 13 1179 47
rect 1213 13 1251 47
rect 1285 13 1323 47
rect 1357 13 1395 47
rect 1429 13 1467 47
rect 1501 13 1539 47
rect 1573 13 1683 47
rect 1717 13 1755 47
rect 1789 13 1827 47
rect 1861 13 1899 47
rect 1933 13 1971 47
rect 2005 13 2043 47
rect 2077 13 2141 47
rect 2175 13 2213 47
rect 2247 13 2285 47
rect 2319 13 2357 47
rect 2391 13 2429 47
rect 2463 13 2501 47
rect 2535 13 2645 47
rect 2679 13 2717 47
rect 2751 13 2789 47
rect 2823 13 2861 47
rect 2895 13 2951 47
rect 2985 13 3023 47
rect 3057 13 3095 47
rect 3129 13 3167 47
rect 3201 13 3311 47
rect 3345 13 3383 47
rect 3417 13 3455 47
rect 3489 13 3527 47
rect 3561 13 3617 47
rect 3651 13 3689 47
rect 3723 13 3761 47
rect 3795 13 3833 47
rect 3867 13 3977 47
rect 4011 13 4049 47
rect 4083 13 4121 47
rect 4155 13 4193 47
rect 4227 13 4265 47
rect 4299 13 4337 47
rect 4371 13 4435 47
rect 4469 13 4507 47
rect 4541 13 4579 47
rect 4613 13 4651 47
rect 4685 13 4723 47
rect 4757 13 4795 47
rect 4829 13 4939 47
rect 4973 13 5011 47
rect 5045 13 5083 47
rect 5117 13 5155 47
rect 5189 13 5245 47
rect 5279 13 5317 47
rect 5351 13 5389 47
rect 5423 13 5461 47
rect 5495 13 5605 47
rect 5639 13 5677 47
rect 5711 13 5749 47
rect 5783 13 5821 47
rect 5855 13 5893 47
rect 5927 13 5965 47
rect 5999 13 6063 47
rect 6097 13 6135 47
rect 6169 13 6207 47
rect 6241 13 6279 47
rect 6313 13 6351 47
rect 6385 13 6423 47
rect 6457 13 6567 47
rect 6601 13 6639 47
rect 6673 13 6711 47
rect 6745 13 6783 47
rect 6817 13 6855 47
rect 6889 13 6927 47
rect 6961 13 7025 47
rect 7059 13 7097 47
rect 7131 13 7169 47
rect 7203 13 7241 47
rect 7275 13 7313 47
rect 7347 13 7385 47
rect 7419 13 7529 47
rect 7563 13 7601 47
rect 7635 13 7673 47
rect 7707 13 7745 47
rect 7779 13 7835 47
rect 7869 13 7907 47
rect 7941 13 7979 47
rect 8013 13 8051 47
rect 8085 13 8195 47
rect 8229 13 8267 47
rect 8301 13 8339 47
rect 8373 13 8411 47
rect 8445 13 8501 47
rect 8535 13 8573 47
rect 8607 13 8645 47
rect 8679 13 8717 47
rect 8751 13 8861 47
rect 8895 13 8933 47
rect 8967 13 9005 47
rect 9039 13 9077 47
rect 9111 13 9149 47
rect 9183 13 9221 47
rect 9255 13 9319 47
rect 9353 13 9391 47
rect 9425 13 9463 47
rect 9497 13 9535 47
rect 9569 13 9607 47
rect 9641 13 9679 47
rect 9713 13 9823 47
rect 9857 13 9895 47
rect 9929 13 9967 47
rect 10001 13 10039 47
rect 10073 13 10129 47
rect 10163 13 10201 47
rect 10235 13 10273 47
rect 10307 13 10345 47
rect 10379 13 10489 47
rect 10523 13 10561 47
rect 10595 13 10633 47
rect 10667 13 10705 47
rect 10739 13 10777 47
rect 10811 13 10849 47
rect 10883 13 10947 47
rect 10981 13 11019 47
rect 11053 13 11091 47
rect 11125 13 11163 47
rect 11197 13 11235 47
rect 11269 13 11307 47
rect 11341 13 11451 47
rect 11485 13 11523 47
rect 11557 13 11595 47
rect 11629 13 11667 47
rect 11701 13 11739 47
rect 11773 13 11811 47
rect 11845 13 11909 47
rect 11943 13 11981 47
rect 12015 13 12053 47
rect 12087 13 12125 47
rect 12159 13 12197 47
rect 12231 13 12269 47
rect 12303 13 12413 47
rect 12447 13 12485 47
rect 12519 13 12557 47
rect 12591 13 12629 47
rect 12663 13 12719 47
rect 12753 13 12791 47
rect 12825 13 12863 47
rect 12897 13 12935 47
rect 12969 13 13079 47
rect 13113 13 13151 47
rect 13185 13 13223 47
rect 13257 13 13295 47
rect 13329 13 13385 47
rect 13419 13 13457 47
rect 13491 13 13529 47
rect 13563 13 13601 47
rect 13635 13 13745 47
rect 13779 13 13817 47
rect 13851 13 13889 47
rect 13923 13 13961 47
rect 13995 13 14033 47
rect 14067 13 14105 47
rect 14139 13 14203 47
rect 14237 13 14275 47
rect 14309 13 14347 47
rect 14381 13 14419 47
rect 14453 13 14491 47
rect 14525 13 14563 47
rect 14597 13 14707 47
rect 14741 13 14779 47
rect 14813 13 14851 47
rect 14885 13 14923 47
rect 14957 13 15013 47
rect 15047 13 15085 47
rect 15119 13 15157 47
rect 15191 13 15229 47
rect 15263 13 15373 47
rect 15407 13 15445 47
rect 15479 13 15517 47
rect 15551 13 15589 47
rect 15623 13 15679 47
rect 15713 13 15751 47
rect 15785 13 15823 47
rect 15857 13 15895 47
rect 15929 13 16039 47
rect 16073 13 16111 47
rect 16145 13 16183 47
rect 16217 13 16255 47
rect 16289 13 16345 47
rect 16379 13 16417 47
rect 16451 13 16489 47
rect 16523 13 16561 47
rect 16595 13 16681 47
rect -31 0 16681 13
<< labels >>
rlabel metal1 16485 797 16519 831 1 QN
port 1 n
rlabel metal1 205 427 239 461 1 D
port 2 n
rlabel metal1 1093 945 1127 979 1 CLK
port 3 n
rlabel metal1 2055 501 2089 535 1 SN
port 4 n
rlabel metal1 72 1522 72 1522 1 VDD
port 5 n
rlabel metal1 72 30 72 30 1 VSS
port 6 n
<< end >>
