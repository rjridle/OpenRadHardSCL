magic
tech sky130A
magscale 1 2
timestamp 1648751721
<< nwell >>
rect -84 832 750 1575
<< nmos >>
rect 168 324 198 377
tri 198 324 214 340 sw
rect 362 324 392 377
tri 392 324 408 340 sw
rect 168 294 274 324
tri 274 294 304 324 sw
rect 168 193 198 294
tri 198 278 214 294 nw
tri 258 278 274 294 ne
tri 198 193 214 209 sw
tri 258 193 274 209 se
rect 274 193 304 294
rect 362 294 468 324
tri 468 294 498 324 sw
rect 362 279 393 294
tri 393 279 408 294 nw
tri 452 279 467 294 ne
rect 467 279 498 294
tri 168 163 198 193 ne
rect 198 163 274 193
tri 274 163 304 193 nw
rect 362 193 392 279
tri 392 193 408 209 sw
tri 452 193 468 209 se
rect 468 193 498 279
tri 362 163 392 193 ne
rect 392 163 468 193
tri 468 163 498 193 nw
<< pmos >>
rect 187 1051 217 1451
rect 275 1051 305 1451
rect 363 1051 393 1451
rect 451 1051 481 1451
<< ndiff >>
rect 112 361 168 377
rect 112 327 122 361
rect 156 327 168 361
rect 112 289 168 327
rect 198 340 362 377
tri 198 324 214 340 ne
rect 214 324 362 340
rect 392 340 554 377
tri 392 324 408 340 ne
rect 408 324 554 340
tri 274 294 304 324 ne
rect 112 255 122 289
rect 156 255 168 289
rect 112 221 168 255
rect 112 187 122 221
rect 156 187 168 221
tri 198 278 214 294 se
rect 214 278 258 294
tri 258 278 274 294 sw
rect 198 245 274 278
rect 198 211 219 245
rect 253 211 274 245
rect 198 209 274 211
tri 198 193 214 209 ne
rect 214 193 258 209
tri 258 193 274 209 nw
rect 304 289 362 324
tri 468 294 498 324 ne
rect 304 255 316 289
rect 350 255 362 289
tri 393 279 408 294 se
rect 408 279 452 294
tri 452 279 467 294 sw
rect 498 289 554 324
rect 304 221 362 255
rect 112 163 168 187
tri 168 163 198 193 sw
tri 274 163 304 193 se
rect 304 187 316 221
rect 350 187 362 221
rect 392 245 468 279
rect 392 211 413 245
rect 447 211 468 245
rect 392 209 468 211
tri 392 193 408 209 ne
rect 408 193 452 209
tri 452 193 468 209 nw
rect 498 255 510 289
rect 544 255 554 289
rect 498 221 554 255
rect 304 163 362 187
tri 362 163 392 193 sw
tri 468 163 498 193 se
rect 498 187 510 221
rect 544 187 554 221
rect 498 163 554 187
rect 112 151 554 163
rect 112 117 122 151
rect 156 117 219 151
rect 253 117 316 151
rect 350 117 413 151
rect 447 117 510 151
rect 544 117 554 151
rect 112 101 554 117
<< pdiff >>
rect 131 1411 187 1451
rect 131 1377 141 1411
rect 175 1377 187 1411
rect 131 1343 187 1377
rect 131 1309 141 1343
rect 175 1309 187 1343
rect 131 1275 187 1309
rect 131 1241 141 1275
rect 175 1241 187 1275
rect 131 1207 187 1241
rect 131 1173 141 1207
rect 175 1173 187 1207
rect 131 1139 187 1173
rect 131 1105 141 1139
rect 175 1105 187 1139
rect 131 1051 187 1105
rect 217 1411 275 1451
rect 217 1377 229 1411
rect 263 1377 275 1411
rect 217 1343 275 1377
rect 217 1309 229 1343
rect 263 1309 275 1343
rect 217 1275 275 1309
rect 217 1241 229 1275
rect 263 1241 275 1275
rect 217 1207 275 1241
rect 217 1173 229 1207
rect 263 1173 275 1207
rect 217 1051 275 1173
rect 305 1411 363 1451
rect 305 1377 317 1411
rect 351 1377 363 1411
rect 305 1343 363 1377
rect 305 1309 317 1343
rect 351 1309 363 1343
rect 305 1275 363 1309
rect 305 1241 317 1275
rect 351 1241 363 1275
rect 305 1207 363 1241
rect 305 1173 317 1207
rect 351 1173 363 1207
rect 305 1139 363 1173
rect 305 1105 317 1139
rect 351 1105 363 1139
rect 305 1051 363 1105
rect 393 1343 451 1451
rect 393 1309 405 1343
rect 439 1309 451 1343
rect 393 1275 451 1309
rect 393 1241 405 1275
rect 439 1241 451 1275
rect 393 1207 451 1241
rect 393 1173 405 1207
rect 439 1173 451 1207
rect 393 1139 451 1173
rect 393 1105 405 1139
rect 439 1105 451 1139
rect 393 1051 451 1105
rect 481 1411 535 1451
rect 481 1377 493 1411
rect 527 1377 535 1411
rect 481 1343 535 1377
rect 481 1309 493 1343
rect 527 1309 535 1343
rect 481 1275 535 1309
rect 481 1241 493 1275
rect 527 1241 535 1275
rect 481 1207 535 1241
rect 481 1173 493 1207
rect 527 1173 535 1207
rect 481 1051 535 1173
<< ndiffc >>
rect 122 327 156 361
rect 122 255 156 289
rect 122 187 156 221
rect 219 211 253 245
rect 316 255 350 289
rect 316 187 350 221
rect 413 211 447 245
rect 510 255 544 289
rect 510 187 544 221
rect 122 117 156 151
rect 219 117 253 151
rect 316 117 350 151
rect 413 117 447 151
rect 510 117 544 151
<< pdiffc >>
rect 141 1377 175 1411
rect 141 1309 175 1343
rect 141 1241 175 1275
rect 141 1173 175 1207
rect 141 1105 175 1139
rect 229 1377 263 1411
rect 229 1309 263 1343
rect 229 1241 263 1275
rect 229 1173 263 1207
rect 317 1377 351 1411
rect 317 1309 351 1343
rect 317 1241 351 1275
rect 317 1173 351 1207
rect 317 1105 351 1139
rect 405 1309 439 1343
rect 405 1241 439 1275
rect 405 1173 439 1207
rect 405 1105 439 1139
rect 493 1377 527 1411
rect 493 1309 527 1343
rect 493 1241 527 1275
rect 493 1173 527 1207
<< psubdiff >>
rect -31 546 697 572
rect -31 512 -17 546
rect 17 512 649 546
rect 683 512 697 546
rect -31 510 697 512
rect -31 474 31 510
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect -31 368 -17 402
rect 17 368 31 402
rect 635 474 697 510
rect 635 440 649 474
rect 683 440 697 474
rect 635 402 697 440
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect 635 368 649 402
rect 683 368 697 402
rect 635 330 697 368
rect 635 296 649 330
rect 683 296 697 330
rect 635 258 697 296
rect 635 224 649 258
rect 683 224 697 258
rect 635 186 697 224
rect 635 152 649 186
rect 683 152 697 186
rect 635 114 697 152
rect -31 47 31 80
rect 635 80 649 114
rect 683 80 697 114
rect 635 47 697 80
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 361 47
rect 395 13 433 47
rect 467 13 505 47
rect 539 13 577 47
rect 611 13 697 47
rect -31 11 31 13
rect 635 11 697 13
<< nsubdiff >>
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 361 1539
rect 395 1505 433 1539
rect 467 1505 505 1539
rect 539 1505 577 1539
rect 611 1505 697 1539
rect -31 1470 31 1505
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect 635 1470 697 1505
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect -31 1038 31 1076
rect 635 1436 649 1470
rect 683 1436 697 1470
rect 635 1398 697 1436
rect 635 1364 649 1398
rect 683 1364 697 1398
rect 635 1326 697 1364
rect 635 1292 649 1326
rect 683 1292 697 1326
rect 635 1254 697 1292
rect 635 1220 649 1254
rect 683 1220 697 1254
rect 635 1182 697 1220
rect 635 1148 649 1182
rect 683 1148 697 1182
rect 635 1110 697 1148
rect 635 1076 649 1110
rect 683 1076 697 1110
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect 635 1038 697 1076
rect 635 1004 649 1038
rect 683 1004 697 1038
rect 635 966 697 1004
rect -31 930 31 932
rect 635 932 649 966
rect 683 932 697 966
rect 635 930 697 932
rect -31 868 697 930
<< psubdiffcont >>
rect -17 512 17 546
rect 649 512 683 546
rect -17 440 17 474
rect -17 368 17 402
rect 649 440 683 474
rect -17 296 17 330
rect -17 224 17 258
rect -17 152 17 186
rect -17 80 17 114
rect 649 368 683 402
rect 649 296 683 330
rect 649 224 683 258
rect 649 152 683 186
rect 649 80 683 114
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 361 13 395 47
rect 433 13 467 47
rect 505 13 539 47
rect 577 13 611 47
<< nsubdiffcont >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 361 1505 395 1539
rect 433 1505 467 1539
rect 505 1505 539 1539
rect 577 1505 611 1539
rect -17 1436 17 1470
rect -17 1364 17 1398
rect -17 1292 17 1326
rect -17 1220 17 1254
rect -17 1148 17 1182
rect -17 1076 17 1110
rect 649 1436 683 1470
rect 649 1364 683 1398
rect 649 1292 683 1326
rect 649 1220 683 1254
rect 649 1148 683 1182
rect 649 1076 683 1110
rect -17 1004 17 1038
rect -17 932 17 966
rect 649 1004 683 1038
rect 649 932 683 966
<< poly >>
rect 187 1451 217 1477
rect 275 1451 305 1477
rect 363 1451 393 1477
rect 451 1451 481 1477
rect 187 1020 217 1051
rect 275 1020 305 1051
rect 363 1020 393 1051
rect 451 1020 481 1051
rect 164 1004 305 1020
rect 164 970 174 1004
rect 208 990 305 1004
rect 350 1004 481 1020
rect 208 970 218 990
rect 164 954 218 970
rect 350 970 360 1004
rect 394 990 481 1004
rect 394 970 404 990
rect 350 954 404 970
rect 195 461 249 477
rect 195 441 205 461
rect 168 427 205 441
rect 239 427 249 461
rect 168 411 249 427
rect 343 461 397 477
rect 343 427 353 461
rect 387 427 397 461
rect 343 411 397 427
rect 168 377 198 411
rect 362 377 392 411
<< polycont >>
rect 174 970 208 1004
rect 360 970 394 1004
rect 205 427 239 461
rect 353 427 387 461
<< locali >>
rect -31 1539 697 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 361 1539
rect 395 1505 433 1539
rect 467 1505 505 1539
rect 539 1505 577 1539
rect 611 1505 697 1539
rect -31 1492 697 1505
rect -31 1470 31 1492
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect -31 1038 31 1076
rect 141 1411 175 1451
rect 141 1343 175 1377
rect 141 1275 175 1309
rect 141 1207 175 1241
rect 141 1139 175 1173
rect 229 1411 263 1492
rect 635 1470 697 1492
rect 229 1343 263 1377
rect 229 1275 263 1309
rect 229 1207 263 1241
rect 229 1157 263 1173
rect 317 1411 527 1445
rect 317 1343 351 1377
rect 317 1275 351 1309
rect 317 1207 351 1241
rect 317 1139 351 1173
rect 141 1071 351 1105
rect 405 1343 439 1359
rect 405 1275 439 1309
rect 405 1207 439 1241
rect 405 1139 439 1173
rect 493 1343 527 1377
rect 493 1275 527 1309
rect 493 1207 527 1241
rect 493 1157 527 1173
rect 635 1436 649 1470
rect 683 1436 697 1470
rect 635 1398 697 1436
rect 635 1364 649 1398
rect 683 1364 697 1398
rect 635 1326 697 1364
rect 635 1292 649 1326
rect 683 1292 697 1326
rect 635 1254 697 1292
rect 635 1220 649 1254
rect 683 1220 697 1254
rect 635 1182 697 1220
rect 635 1148 649 1182
rect 683 1148 697 1182
rect 635 1110 697 1148
rect 405 1071 535 1105
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect 174 1004 208 1020
rect 360 1004 394 1020
rect 208 970 239 988
rect 174 954 239 970
rect -31 868 31 932
rect 205 831 239 954
rect -31 546 31 572
rect -31 512 -17 546
rect 17 512 31 546
rect -31 474 31 512
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect 205 461 239 797
rect 205 411 239 427
rect 353 970 360 988
rect 353 954 394 970
rect 353 757 387 954
rect 501 773 535 1071
rect 635 1076 649 1110
rect 683 1076 697 1110
rect 635 1038 697 1076
rect 635 1004 649 1038
rect 683 1004 697 1038
rect 635 966 697 1004
rect 635 932 649 966
rect 683 932 697 966
rect 635 868 697 932
rect 353 461 387 723
rect 500 757 535 773
rect 534 723 535 757
rect 500 707 535 723
rect 353 411 387 427
rect -31 368 -17 402
rect 17 368 31 402
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect -31 62 31 80
rect 122 361 156 377
rect 501 376 535 707
rect 122 289 156 327
rect 122 221 156 255
rect 219 342 535 376
rect 635 546 697 572
rect 635 512 649 546
rect 683 512 697 546
rect 635 474 697 512
rect 635 440 649 474
rect 683 440 697 474
rect 635 402 697 440
rect 635 368 649 402
rect 683 368 697 402
rect 219 245 253 342
rect 219 195 253 211
rect 316 289 350 306
rect 316 221 350 255
rect 122 151 156 187
rect 413 245 447 342
rect 635 330 697 368
rect 413 195 447 211
rect 510 289 544 306
rect 510 221 544 255
rect 316 151 350 187
rect 510 151 544 187
rect 156 117 219 151
rect 253 117 316 151
rect 350 117 413 151
rect 447 117 510 151
rect 122 62 156 117
rect 219 62 253 117
rect 316 62 350 117
rect 413 62 447 117
rect 510 62 544 117
rect 635 296 649 330
rect 683 296 697 330
rect 635 258 697 296
rect 635 224 649 258
rect 683 224 697 258
rect 635 186 697 224
rect 635 152 649 186
rect 683 152 697 186
rect 635 114 697 152
rect 635 80 649 114
rect 683 80 697 114
rect 635 62 697 80
rect -31 47 697 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 361 47
rect 395 13 433 47
rect 467 13 505 47
rect 539 13 577 47
rect 611 13 697 47
rect -31 0 697 13
<< viali >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 361 1505 395 1539
rect 433 1505 467 1539
rect 505 1505 539 1539
rect 577 1505 611 1539
rect 205 797 239 831
rect 353 723 387 757
rect 500 723 534 757
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 361 13 395 47
rect 433 13 467 47
rect 505 13 539 47
rect 577 13 611 47
<< metal1 >>
rect -31 1539 697 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 361 1539
rect 395 1505 433 1539
rect 467 1505 505 1539
rect 539 1505 577 1539
rect 611 1505 697 1539
rect -31 1492 697 1505
rect 199 831 245 837
rect 169 797 205 831
rect 239 797 251 831
rect 199 791 245 797
rect 347 757 393 763
rect 494 757 540 763
rect 317 723 353 757
rect 387 723 399 757
rect 488 723 500 757
rect 534 723 570 757
rect 347 717 393 723
rect 494 717 540 723
rect -31 47 697 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 361 47
rect 395 13 433 47
rect 467 13 505 47
rect 539 13 577 47
rect 611 13 697 47
rect -31 0 697 13
<< labels >>
rlabel metal1 500 723 534 757 1 Y
port 1 n
rlabel metal1 205 797 239 831 1 A
port 2 n
rlabel metal1 353 723 387 757 1 B
port 3 n
rlabel metal1 55 1505 89 1539 1 VDD
port 4 n
rlabel metal1 55 13 89 47 1 VSS
port 5 n
<< end >>
