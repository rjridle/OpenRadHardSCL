* HSPICE file created from tmp.ext - technology: sky130A

.option scale=5000u

.subckt tmp Y A B C VDD VSS
X0 a_277_1051 C VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=67200 ps=2736 w=400 l=30 M=2
X1 VDD a_277_1051 Y VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=11600 ps=458 w=400 l=30 M=2
X2 VDD A a_277_1051 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=400 l=30 M=2
X3 a_277_1051 C a_372_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=598 l=30
X4 VDD B a_277_1051 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=400 l=30 M=2
X5 Y a_277_1051 VSS VSS sky130_fd_pr__nfet_01v8 ad=7088 pd=312 as=53378 ps=1936 w=598 l=30
X6 a_372_210 B a_91_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=600 l=30
X7 VSS A a_91_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=598 l=30
C0 VDD a_277_1051 2.89fF
.ends

** hspice subcircuit dictionary
