magic
tech sky130
magscale 1 2
timestamp 1651259629
<< metal1 >>
rect 1377 945 3313 979
rect 1660 797 5490 831
rect 716 723 4024 757
rect 831 576 2174 610
rect 2757 575 3055 609
rect 426 501 4265 535
rect 2351 427 5210 461
use nand3x1_pcell  nand3x1_pcell_1
timestamp 1651259484
transform 1 0 962 0 1 0
box -84 0 1046 1575
use nand3x1_pcell  nand3x1_pcell_0
timestamp 1651259484
transform 1 0 0 0 1 0
box -84 0 1046 1575
use li1_M1_contact  li1_M1_contact_2
timestamp 1648061256
transform -1 0 444 0 -1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform -1 0 666 0 -1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_3
timestamp 1648061256
transform -1 0 814 0 -1 593
box -53 -33 29 33
use nand3x1_pcell  nand3x1_pcell_2
timestamp 1651259484
transform 1 0 1924 0 1 0
box -84 0 1046 1575
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform -1 0 1405 0 -1 962
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_7
timestamp 1648061256
transform -1 0 1776 0 -1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_8
timestamp 1648061256
transform 1 0 2146 0 1 593
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_5
timestamp 1648061256
transform -1 0 1184 0 -1 593
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_4
timestamp 1648061256
transform -1 0 1627 0 -1 814
box -53 -33 29 33
use nand3x1_pcell  nand3x1_pcell_3
timestamp 1651259484
transform 1 0 2886 0 1 0
box -84 0 1046 1575
use li1_M1_contact  li1_M1_contact_6
timestamp 1648061256
transform 1 0 3330 0 1 962
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_10
timestamp 1648061256
transform -1 0 2368 0 -1 445
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_17
timestamp 1648061256
transform 1 0 3108 0 1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_11
timestamp 1648061256
transform -1 0 2738 0 -1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_9
timestamp 1648061256
transform 1 0 2590 0 1 814
box -53 -33 29 33
use nand3x1_pcell  nand3x1_pcell_4
timestamp 1651259484
transform 1 0 3848 0 1 0
box -84 0 1046 1575
use li1_M1_contact  li1_M1_contact_12
timestamp 1648061256
transform -1 0 3552 0 -1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_18
timestamp 1648061256
transform 1 0 4292 0 1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_19
timestamp 1648061256
transform 1 0 4070 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_13
timestamp 1648061256
transform -1 0 3700 0 -1 814
box -53 -33 29 33
use nand3x1_pcell  nand3x1_pcell_5
timestamp 1651259484
transform 1 0 4810 0 1 0
box -84 0 1046 1575
use li1_M1_contact  li1_M1_contact_22
timestamp 1648061256
transform 1 0 5254 0 1 444
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_20
timestamp 1648061256
transform 1 0 5476 0 1 814
box -53 -33 29 33
<< end >>
