magic
tech sky130A
magscale 1 2
timestamp 1643175030
<< nmos >>
rect 56 202 86 270
rect 56 172 152 202
tri 152 172 182 202 sw
rect 56 80 86 172
tri 86 156 102 172 nw
tri 136 156 152 172 ne
tri 86 80 102 96 sw
tri 136 80 152 96 se
rect 152 80 182 172
tri 56 50 86 80 ne
rect 86 50 152 80
tri 152 50 182 80 nw
<< ndiff >>
rect 0 254 56 270
rect 0 220 10 254
rect 44 220 56 254
rect 0 186 56 220
rect 86 254 238 270
rect 86 220 126 254
rect 160 220 194 254
rect 228 220 238 254
rect 86 202 238 220
rect 0 152 10 186
rect 44 152 56 186
tri 152 172 182 202 ne
rect 182 186 238 202
rect 0 118 56 152
rect 0 84 10 118
rect 44 84 56 118
rect 0 50 56 84
tri 86 156 102 172 se
rect 102 156 136 172
tri 136 156 152 172 sw
rect 86 143 152 156
rect 86 109 102 143
rect 136 109 152 143
rect 86 96 152 109
tri 86 80 102 96 ne
rect 102 80 136 96
tri 136 80 152 96 nw
rect 182 152 194 186
rect 228 152 238 186
rect 182 118 238 152
rect 182 84 194 118
rect 228 84 238 118
tri 56 50 86 80 sw
tri 152 50 182 80 se
rect 182 50 238 84
rect 0 16 10 50
rect 44 16 194 50
rect 228 16 238 50
rect 0 0 238 16
<< ndiffc >>
rect 10 220 44 254
rect 126 220 160 254
rect 194 220 228 254
rect 10 152 44 186
rect 10 84 44 118
rect 102 109 136 143
rect 194 152 228 186
rect 194 84 228 118
rect 10 16 44 50
rect 194 16 228 50
<< poly >>
rect 56 270 86 296
<< locali >>
rect 10 254 44 270
rect 194 254 228 270
rect 44 220 126 254
rect 160 220 194 254
rect 10 186 44 220
rect 194 186 228 220
rect 10 118 44 152
rect 10 50 44 84
rect 10 0 44 16
rect 102 143 136 159
rect 102 0 136 109
rect 194 118 228 152
rect 194 50 228 84
rect 194 0 228 16
<< end >>
