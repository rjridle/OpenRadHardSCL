* SPICE3 file created from MUX2X1.ext - technology: sky130A

.subckt MUX2X1 Y A0 A1 S VDD VSS
X0 VDD a_185_209 a_1327_1050 VDD sky130_fd_pr__pfet_01v8 ad=6.14p pd=5.014u as=0p ps=0u w=2u l=0.15u M=2
X1 a_185_209 S VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X2 Y a_1327_1050 a_1888_101 VSS sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=0p ps=0u w=3u l=0.15u
X3 a_661_1050 A0 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X4 VSS S a_556_101 VSS sky130_fd_pr__nfet_01v8 ad=1.6781p pd=1.281u as=0p ps=0u w=3u l=0.15u
X5 VDD A1 a_1327_1050 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X6 a_185_209 S VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X7 a_661_1050 S VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X8 a_1327_1050 A1 a_1222_101 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X9 VDD a_1327_1050 Y VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.16p ps=9.16u w=2u l=0.15u M=2
X10 a_661_1050 A0 a_556_101 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X11 VDD a_661_1050 Y VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X12 VSS a_661_1050 a_1888_101 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X13 VSS a_185_209 a_1222_101 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
C0 VDD a_661_1050 2.21fF
C1 VDD a_1327_1050 2.21fF
C2 VDD VSS 3.98fF
.ends
