magic
tech sky130
magscale 1 2
timestamp 1651259543
<< metal1 >>
rect 537 501 841 535
rect 1203 501 1512 535
use nand2x1_pcell  nand2x1_pcell_1
timestamp 1651259477
transform 1 0 1332 0 1 0
box -84 0 750 1575
use nand2x1_pcell  nand2x1_pcell_0
timestamp 1651259477
transform 1 0 0 0 1 0
box -84 0 750 1575
use nor2x1_pcell  nor2x1_pcell_0
timestamp 1651259490
transform 1 0 666 0 1 0
box -84 0 750 1575
use li1_M1_contact  li1_M1_contact_3
timestamp 1648061256
transform 1 0 1554 0 1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_2
timestamp 1648061256
transform -1 0 1184 0 -1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform 1 0 888 0 1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform -1 0 518 0 -1 518
box -53 -33 29 33
<< end >>
