magic
tech sky130
magscale 1 2
timestamp 1651260992
<< nwell >>
rect 55 1505 89 1539
<< pwell >>
rect 55 13 89 47
<< metal1 >>
rect -31 1492 697 1554
rect 205 797 239 831
rect 353 723 387 757
rect 500 723 534 757
rect -31 0 697 62
use nor2x1_pcell  nor2x1_pcell_0 pcells
timestamp 1651259490
transform 1 0 0 0 1 0
box -84 0 750 1575
use li1_M1_contact  li1_M1_contact_2 pcells
timestamp 1648061256
transform -1 0 517 0 -1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform 1 0 370 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform 1 0 222 0 1 814
box -53 -33 29 33
<< labels >>
rlabel metal1 500 723 534 757 1 Y
port 1 nsew signal output
rlabel metal1 205 797 239 831 1 A
port 2 nsew signal input
rlabel metal1 353 723 387 757 1 B
port 3 nsew signal input
rlabel metal1 -31 1492 697 1554 1 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 -31 0 697 62 1 VGND
port 5 nsew ground bidirectional abutment
rlabel nwell 55 1505 89 1539 1 VPB
port 6 nsew power bidirectional
rlabel pwell 55 13 89 47 1 VNB
port 7 nsew ground bidirectional
<< end >>
