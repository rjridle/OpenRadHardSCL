* SPICE3 file created from NOR2X1.ext - technology: sky130A

.subckt NOR2X1 Y A B VDD GND
X0 Y A.t1 GND.t0 GND sky130_fd_pr__nfet_01v8 ad=3.582p pd=3.15u as=0p ps=0u w=0u l=0u
X1 a_131_1051.t2 A.t0 VDD.t4 VDD.t3 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X2 Y A GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.9366p ps=1.294u w=3u l=0.15u
X3 a_131_1051.t0 B.t0 Y.t0  �4�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X4 Y B.t1 GND.t1 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X5 Y B GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X6 VDD.t2 A.t2 a_131_1051.t1 �4�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X7 Y.t3 B.t2 a_131_1051.t3  �4�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
C0 Y VDD 0.50fF
C1 B VDD 0.32fF
C2 Y B 0.29fF
C3 A VDD 0.36fF
C4 Y A 0.11fF
C5 B A 0.26fF
R0 A.n0 A.t0 486.819
R1 A.n0 A.t2 384.527
R2 A.n1 A.t1 378.637
R3 A.n1 A.n0 151.269
R4 A.n2 A.n1 4.65
R5 A.n2 A 0.046
R6 VDD.n64 VDD.n63 129.849
R7 VDD.n44 VDD.n43 92.5
R8 VDD.n42 VDD.n41 92.5
R9 VDD.n40 VDD.n39 92.5
R10 VDD.n38 VDD.n37 92.5
R11 VDD.n46 VDD.n45 92.5
R12 VDD.n14 VDD.n1 92.5
R13 VDD.n5 VDD.n4 92.5
R14 VDD.n7 VDD.n6 92.5
R15 VDD.n9 VDD.n8 92.5
R16 VDD.n11 VDD.n10 92.5
R17 VDD.n13 VDD.n12 92.5
R18 VDD.n21 VDD.n20 92.059
R19 VDD.n55 VDD.n54 92.059
R20 VDD.n20 VDD.n16 67.194
R21 VDD.n20 VDD.n17 67.194
R22 VDD.n20 VDD.n18 67.194
R23 VDD.n20 VDD.n19 67.194
R24 VDD.n5 VDD.n3 44.141
R25 VDD.n3 VDD.n2 44.107
R26 VDD.n20 VDD.n15 41.052
R27 VDD.n53 VDD.n51 39.742
R28 VDD.n53 VDD.n52 39.742
R29 VDD.n50 VDD.n49 39.742
R30 VDD.n1 VDD.n0 30.923
R31 VDD.n54 VDD.n53 26.38
R32 VDD.n54 VDD.n50 26.38
R33 VDD.n54 VDD.n48 26.38
R34 VDD.n54 VDD.n47 26.38
R35 VDD.n57 VDD.n46 22.915
R36 VDD.n23 VDD.n14 22.915
R37 VDD.n28  �4�� 20.457
R38 VDD.n65 �4�� 17.9
R39 VDD.n46 VDD.n44 14.864
R40 VDD.n44 VDD.n42 14.864
R41 VDD.n42 VDD.n40 14.864
R42 VDD.n40 VDD.n38 14.864
R43 VDD.n38 VDD.n36 14.864
R44 VDD.n36 VDD.n35 14.864
R45 VDD.n14 VDD.n13 14.864
R46 VDD.n13 VDD.n11 14.864
R47 VDD.n11 VDD.n9 14.864
R48 VDD.n9 VDD.n7 14.864
R49 VDD.n7 VDD.n5 14.864
R50 VDD.n63 VDD.t4 14.282
R51 VDD.n63 VDD.t2 14.282
R52 VDD.n23 VDD.n22 8.855
R53 VDD.n22 VDD.n21 8.855
R54 VDD.n26 VDD.n25 8.855
R55 VDD.n25 VDD.n24 8.855
R56 VDD.n30 VDD.n29 8.855
R57 VDD.n29 VDD.n28 8.855
R58 VDD.n33 VDD.n32 8.855
R59 VDD.n32  �4�� 8.855
R60 VDD.n71 VDD.n70 8.855
R61 VDD.n70 VDD.n69 8.855
R62 VDD.n67 VDD.n66 8.855
R63 VDD.n66 VDD.n65 8.855
R64 VDD.n61 VDD.n60 8.855
R65 VDD.n60 VDD.n59 8.855
R66 VDD.n57 VDD.n56 8.855
R67 VDD.n56 VDD.n55 8.855
R68 VDD.n67 VDD.n64 6.193
R69 VDD.n31 VDD.n30 4.65
R70 VDD.n34 VDD.n33 4.65
R71 VDD.n72 VDD.n71 4.65
R72 VDD.n68 VDD.n67 4.65
R73 VDD.n62 VDD.n61 4.65
R74 VDD.n58 VDD.n57 4.65
R75 VDD.n27 VDD.n23 2.933
R76 VDD.n27 VDD.n26 2.844
R77 VDD.n69 VDD.t3 2.557
R78 VDD.n31 VDD.n27 1.063
R79 VDD.n58 VDD 0.207
R80 VDD.n34 VDD.n31 0.145
R81 VDD.n72 VDD.n68 0.145
R82 VDD.n68 VDD.n62 0.145
R83 VDD.n62 VDD.n58 0.145
R84 VDD VDD.n34 0.09
R85 VDD VDD.n72 0.09
R86 a_131_1051.n0 a_131_1051.t0 228.369
R87 a_131_1051.n0 a_131_1051.t1 219.778
R88 a_131_1051.n1 a_131_1051.n0 42.29
R89 a_131_1051.n1 a_131_1051.t3 14.282
R90 a_131_1051.t2 a_131_1051.n1 14.282
R91 GND.n11 GND.n10 92.5
R92 GND.n29 GND.n28 92.5
R93 GND.n23 GND.t0 45.413
R94 GND.n37 GND.n36 40.431
R95 GND.n23 GND.n22 39.307
R96 GND.n3 GND.n2 35.865
R97 GND.n4 GND.n3 28.503
R98 GND.n24 GND.n23 23.77
R99 GND.n30 GND.n29 20.705
R100 GND.n38 GND.n37 20.705
R101 GND.n12 GND.n11 20.705
R102 GND.n5 GND.n4 20.705
R103 GND.n25 GND.n24 20.705
R104 GND.n36 GND.t1 13.654
R105 GND.n36 GND.n35 13.654
R106 GND.n40 GND.n38 9.29
R107 GND.n26 GND.n21 9.154
R108 GND.n32 GND.n31 9.154
R109 GND.n40 GND.n39 9.154
R110 GND.n16 GND.n15 9.154
R111 GND.n13 GND.n9 9.154
R112 GND.n7 GND.n6 9.154
R113 GND.t1 GND.n34 7.04
R114 GND.n8 GND.n1 4.795
R115 GND.n20 GND.n19 4.65
R116 GND.n8 GND.n7 4.65
R117 GND.n14 GND.n13 4.65
R118 GND.n17 GND.n16 4.65
R119 GND.n41 GND.n40 4.65
R120 GND.n33 GND.n32 4.65