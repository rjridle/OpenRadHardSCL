magic
tech sky130A
magscale 1 2
timestamp 1643653892
<< nwell >>
rect 492 1323 1114 1353
rect 492 1319 1111 1323
rect 492 1281 520 1319
rect 564 1318 1111 1319
rect 564 1317 1102 1318
rect 564 1281 1111 1317
rect 492 1279 1111 1281
rect 492 794 1114 1279
rect 492 770 1129 794
rect 1135 770 1202 794
rect 492 759 1216 770
<< ndiff >>
rect 727 272 761 346
<< psubdiff >>
rect 571 490 1101 552
rect 509 13 516 47
rect 563 13 591 47
rect 625 13 659 47
rect 693 13 727 47
rect 761 13 819 47
rect 853 13 911 47
rect 945 13 979 47
rect 1013 13 1047 47
rect 1081 13 1101 47
<< nsubdiff >>
rect 509 1283 520 1317
rect 564 1283 592 1317
rect 627 1283 661 1317
rect 696 1283 730 1317
rect 765 1283 819 1317
rect 854 1283 908 1317
rect 943 1283 977 1317
rect 1012 1283 1046 1317
rect 1081 1283 1111 1317
rect 509 795 1163 857
<< psubdiffcont >>
rect 591 13 625 47
rect 659 13 693 47
rect 727 13 761 47
rect 819 13 853 47
rect 911 13 945 47
rect 979 13 1013 47
rect 1047 13 1081 47
<< nsubdiffcont >>
rect 592 1283 627 1317
rect 661 1283 696 1317
rect 730 1283 765 1317
rect 819 1283 854 1317
rect 908 1283 943 1317
rect 977 1283 1012 1317
rect 1046 1283 1081 1317
<< poly >>
rect 681 916 685 946
rect 681 403 711 465
<< locali >>
rect 509 1319 1101 1332
rect 509 1281 520 1319
rect 564 1317 1101 1319
rect 564 1283 592 1317
rect 627 1283 661 1317
rect 696 1283 730 1317
rect 765 1283 819 1317
rect 854 1283 908 1317
rect 943 1283 977 1317
rect 1012 1283 1046 1317
rect 1081 1283 1111 1317
rect 564 1281 1101 1283
rect 509 1270 1101 1281
rect 727 1036 761 1060
rect 727 272 761 1002
rect 903 1035 937 1041
rect 903 995 937 1001
rect 509 55 1101 62
rect 509 7 516 55
rect 563 47 1101 55
rect 563 13 591 47
rect 625 13 659 47
rect 693 13 727 47
rect 761 13 819 47
rect 853 13 911 47
rect 945 13 979 47
rect 1013 13 1047 47
rect 1081 13 1101 47
rect 563 7 1101 13
rect 509 0 1101 7
<< viali >>
rect 592 1283 627 1317
rect 661 1283 696 1317
rect 730 1283 765 1317
rect 819 1283 854 1317
rect 908 1283 943 1317
rect 977 1283 1012 1317
rect 1046 1283 1081 1317
rect 727 1002 761 1036
rect 903 1001 937 1035
rect 591 13 625 47
rect 659 13 693 47
rect 727 13 761 47
rect 819 13 853 47
rect 911 13 945 47
rect 979 13 1013 47
rect 1047 13 1081 47
<< metal1 >>
rect 509 1319 1101 1332
rect 509 1281 520 1319
rect 564 1317 1101 1319
rect 564 1283 592 1317
rect 627 1283 661 1317
rect 696 1283 730 1317
rect 765 1283 819 1317
rect 854 1283 908 1317
rect 943 1283 977 1317
rect 1012 1283 1046 1317
rect 1081 1283 1111 1317
rect 564 1281 1101 1283
rect 509 1270 1101 1281
rect 721 1036 767 1042
rect 897 1036 943 1041
rect 715 1002 727 1036
rect 761 1035 943 1036
rect 761 1002 903 1035
rect 721 1001 903 1002
rect 937 1001 949 1035
rect 721 996 767 1001
rect 897 995 943 1001
rect 637 473 671 874
rect 871 473 905 936
rect 509 55 1101 62
rect 509 7 516 55
rect 563 47 1101 55
rect 563 13 591 47
rect 625 13 659 47
rect 693 13 727 47
rect 761 13 819 47
rect 853 13 911 47
rect 945 13 979 47
rect 1013 13 1047 47
rect 1081 13 1101 47
rect 563 7 1101 13
rect 509 0 1101 7
use nmos_bottom_left  nmos_bottom_left_0 pcells
timestamp 1643178650
transform 1 0 854 0 1 165
box -45 -64 193 238
use diff_ring_side  diff_ring_side_1 pcells
timestamp 1643181737
transform 1 0 1207 0 1 0
box -159 0 9 1353
use pmos  pmos_1 pcells
timestamp 1643179034
transform 1 0 805 0 1 1228
box -36 -312 264 42
use M1_M2_contact  M1_M2_contact_3 pcells
timestamp 1643652910
transform 1 0 791 0 1 481
box 64 391 130 473
use M1_M2_contact  M1_M2_contact_1
timestamp 1643652910
transform 1 0 791 0 1 0
box 64 391 130 473
use diff_ring_side  diff_ring_side_0
timestamp 1643181737
transform 1 0 615 0 1 0
box -159 0 9 1353
use nmos_top_left  nmos_top_left_0 pcells
timestamp 1643177486
transform 1 0 670 0 1 165
box -45 -64 193 238
use M1_M2_contact  M1_M2_contact_0
timestamp 1643652910
transform 1 0 557 0 1 0
box 64 391 130 473
use M1_M2_contact  M1_M2_contact_2
timestamp 1643652910
transform 1 0 557 0 1 481
box 64 391 130 473
use pmos  pmos_0
timestamp 1643179034
transform 1 0 629 0 1 1228
box -36 -312 264 42
<< labels >>
rlabel metal1 727 1002 761 1036 1 YN
port 1 n
rlabel nwell 637 896 671 930 1 A
port 2 n
rlabel metal1 871 896 905 930 1 B
port 3 n
<< end >>
