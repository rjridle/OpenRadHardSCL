magic
tech sky130A
magscale 1 2
timestamp 1649549313
<< nwell >>
rect -84 832 2526 1575
<< nmos >>
rect 155 324 185 377
tri 185 324 201 340 sw
rect 155 294 261 324
tri 261 294 291 324 sw
rect 155 193 185 294
tri 185 278 201 294 nw
tri 245 278 261 294 ne
tri 185 193 201 209 sw
tri 245 193 261 209 se
rect 261 193 291 294
tri 155 163 185 193 ne
rect 185 163 261 193
tri 261 163 291 193 nw
rect 612 316 642 377
tri 642 316 658 332 sw
rect 806 324 836 377
tri 836 324 852 340 sw
rect 612 286 718 316
tri 718 286 748 316 sw
rect 806 294 912 324
tri 912 294 942 324 sw
rect 612 185 642 286
tri 642 270 658 286 nw
tri 702 270 718 286 ne
tri 642 185 658 201 sw
tri 702 185 718 201 se
rect 718 185 748 286
rect 806 193 836 294
tri 836 278 852 294 nw
tri 896 278 912 294 ne
tri 836 193 852 209 sw
tri 896 193 912 209 se
rect 912 193 942 294
tri 612 155 642 185 ne
rect 642 155 718 185
tri 718 155 748 185 nw
tri 806 163 836 193 ne
rect 836 163 912 193
tri 912 163 942 193 nw
rect 1278 316 1308 377
tri 1308 316 1324 332 sw
rect 1472 324 1502 377
tri 1502 324 1518 340 sw
rect 1278 286 1384 316
tri 1384 286 1414 316 sw
rect 1472 294 1578 324
tri 1578 294 1608 324 sw
rect 1278 185 1308 286
tri 1308 270 1324 286 nw
tri 1368 270 1384 286 ne
tri 1308 185 1324 201 sw
tri 1368 185 1384 201 se
rect 1384 185 1414 286
rect 1472 193 1502 294
tri 1502 278 1518 294 nw
tri 1562 278 1578 294 ne
tri 1502 193 1518 209 sw
tri 1562 193 1578 209 se
rect 1578 193 1608 294
tri 1278 155 1308 185 ne
rect 1308 155 1384 185
tri 1384 155 1414 185 nw
tri 1472 163 1502 193 ne
rect 1502 163 1578 193
tri 1578 163 1608 193 nw
rect 1944 316 1974 377
tri 1974 316 1990 332 sw
rect 2138 324 2168 377
tri 2168 324 2184 340 sw
rect 1944 286 2050 316
tri 2050 286 2080 316 sw
rect 2138 294 2244 324
tri 2244 294 2274 324 sw
rect 1944 185 1974 286
tri 1974 270 1990 286 nw
tri 2034 270 2050 286 ne
tri 1974 185 1990 201 sw
tri 2034 185 2050 201 se
rect 2050 185 2080 286
rect 2138 193 2168 294
tri 2168 278 2184 294 nw
tri 2228 278 2244 294 ne
tri 2168 193 2184 209 sw
tri 2228 193 2244 209 se
rect 2244 193 2274 294
tri 1944 155 1974 185 ne
rect 1974 155 2050 185
tri 2050 155 2080 185 nw
tri 2138 163 2168 193 ne
rect 2168 163 2244 193
tri 2244 163 2274 193 nw
<< pmos >>
rect 163 1050 193 1450
rect 251 1050 281 1450
rect 631 1050 661 1450
rect 719 1050 749 1450
rect 807 1050 837 1450
rect 895 1050 925 1450
rect 1297 1050 1327 1450
rect 1385 1050 1415 1450
rect 1473 1050 1503 1450
rect 1561 1050 1591 1450
rect 1963 1050 1993 1450
rect 2051 1050 2081 1450
rect 2139 1050 2169 1450
rect 2227 1050 2257 1450
<< ndiff >>
rect 99 361 155 377
rect 99 327 109 361
rect 143 327 155 361
rect 99 289 155 327
rect 185 361 345 377
rect 185 340 303 361
tri 185 324 201 340 ne
rect 201 327 303 340
rect 337 327 345 361
rect 201 324 345 327
tri 261 294 291 324 ne
rect 99 255 109 289
rect 143 255 155 289
rect 99 221 155 255
rect 99 187 109 221
rect 143 187 155 221
tri 185 278 201 294 se
rect 201 278 245 294
tri 245 278 261 294 sw
rect 185 245 261 278
rect 185 211 205 245
rect 239 211 261 245
rect 185 209 261 211
tri 185 193 201 209 ne
rect 201 193 245 209
tri 245 193 261 209 nw
rect 291 289 345 324
rect 291 255 303 289
rect 337 255 345 289
rect 291 221 345 255
rect 99 163 155 187
tri 155 163 185 193 sw
tri 261 163 291 193 se
rect 291 187 303 221
rect 337 187 345 221
rect 291 163 345 187
rect 99 151 345 163
rect 99 117 109 151
rect 143 117 205 151
rect 239 117 303 151
rect 337 117 345 151
rect 99 101 345 117
rect 556 361 612 377
rect 556 327 566 361
rect 600 327 612 361
rect 556 289 612 327
rect 642 361 806 377
rect 642 332 663 361
tri 642 316 658 332 ne
rect 658 327 663 332
rect 697 327 760 361
rect 794 327 806 361
rect 658 316 806 327
rect 836 340 998 377
tri 836 324 852 340 ne
rect 852 324 998 340
rect 556 255 566 289
rect 600 255 612 289
tri 718 286 748 316 ne
rect 748 289 806 316
tri 912 294 942 324 ne
rect 556 221 612 255
rect 556 187 566 221
rect 600 187 612 221
rect 556 155 612 187
tri 642 270 658 286 se
rect 658 270 702 286
tri 702 270 718 286 sw
rect 642 236 718 270
rect 642 202 663 236
rect 697 202 718 236
rect 642 201 718 202
tri 642 185 658 201 ne
rect 658 185 702 201
tri 702 185 718 201 nw
rect 748 255 760 289
rect 794 255 806 289
rect 748 221 806 255
rect 748 187 760 221
rect 794 187 806 221
tri 836 278 852 294 se
rect 852 278 896 294
tri 896 278 912 294 sw
rect 836 245 912 278
rect 836 211 857 245
rect 891 211 912 245
rect 836 209 912 211
tri 836 193 852 209 ne
rect 852 193 896 209
tri 896 193 912 209 nw
rect 942 289 998 324
rect 942 255 954 289
rect 988 255 998 289
rect 942 221 998 255
tri 612 155 642 185 sw
tri 718 155 748 185 se
rect 748 163 806 187
tri 806 163 836 193 sw
tri 912 163 942 193 se
rect 942 187 954 221
rect 988 187 998 221
rect 942 163 998 187
rect 748 155 998 163
rect 556 151 998 155
rect 556 117 566 151
rect 600 117 760 151
rect 794 117 857 151
rect 891 117 954 151
rect 988 117 998 151
rect 556 101 998 117
rect 1222 361 1278 377
rect 1222 327 1232 361
rect 1266 327 1278 361
rect 1222 289 1278 327
rect 1308 361 1472 377
rect 1308 332 1329 361
tri 1308 316 1324 332 ne
rect 1324 327 1329 332
rect 1363 327 1426 361
rect 1460 327 1472 361
rect 1324 316 1472 327
rect 1502 340 1664 377
tri 1502 324 1518 340 ne
rect 1518 324 1664 340
rect 1222 255 1232 289
rect 1266 255 1278 289
tri 1384 286 1414 316 ne
rect 1414 289 1472 316
tri 1578 294 1608 324 ne
rect 1222 221 1278 255
rect 1222 187 1232 221
rect 1266 187 1278 221
rect 1222 155 1278 187
tri 1308 270 1324 286 se
rect 1324 270 1368 286
tri 1368 270 1384 286 sw
rect 1308 236 1384 270
rect 1308 202 1329 236
rect 1363 202 1384 236
rect 1308 201 1384 202
tri 1308 185 1324 201 ne
rect 1324 185 1368 201
tri 1368 185 1384 201 nw
rect 1414 255 1426 289
rect 1460 255 1472 289
rect 1414 221 1472 255
rect 1414 187 1426 221
rect 1460 187 1472 221
tri 1502 278 1518 294 se
rect 1518 278 1562 294
tri 1562 278 1578 294 sw
rect 1502 245 1578 278
rect 1502 211 1523 245
rect 1557 211 1578 245
rect 1502 209 1578 211
tri 1502 193 1518 209 ne
rect 1518 193 1562 209
tri 1562 193 1578 209 nw
rect 1608 289 1664 324
rect 1608 255 1620 289
rect 1654 255 1664 289
rect 1608 221 1664 255
tri 1278 155 1308 185 sw
tri 1384 155 1414 185 se
rect 1414 163 1472 187
tri 1472 163 1502 193 sw
tri 1578 163 1608 193 se
rect 1608 187 1620 221
rect 1654 187 1664 221
rect 1608 163 1664 187
rect 1414 155 1664 163
rect 1222 151 1664 155
rect 1222 117 1232 151
rect 1266 117 1426 151
rect 1460 117 1523 151
rect 1557 117 1620 151
rect 1654 117 1664 151
rect 1222 101 1664 117
rect 1888 361 1944 377
rect 1888 327 1898 361
rect 1932 327 1944 361
rect 1888 289 1944 327
rect 1974 361 2138 377
rect 1974 332 1995 361
tri 1974 316 1990 332 ne
rect 1990 327 1995 332
rect 2029 327 2092 361
rect 2126 327 2138 361
rect 1990 316 2138 327
rect 2168 340 2330 377
tri 2168 324 2184 340 ne
rect 2184 324 2330 340
rect 1888 255 1898 289
rect 1932 255 1944 289
tri 2050 286 2080 316 ne
rect 2080 289 2138 316
tri 2244 294 2274 324 ne
rect 1888 221 1944 255
rect 1888 187 1898 221
rect 1932 187 1944 221
rect 1888 155 1944 187
tri 1974 270 1990 286 se
rect 1990 270 2034 286
tri 2034 270 2050 286 sw
rect 1974 236 2050 270
rect 1974 202 1995 236
rect 2029 202 2050 236
rect 1974 201 2050 202
tri 1974 185 1990 201 ne
rect 1990 185 2034 201
tri 2034 185 2050 201 nw
rect 2080 255 2092 289
rect 2126 255 2138 289
rect 2080 221 2138 255
rect 2080 187 2092 221
rect 2126 187 2138 221
tri 2168 278 2184 294 se
rect 2184 278 2228 294
tri 2228 278 2244 294 sw
rect 2168 245 2244 278
rect 2168 211 2189 245
rect 2223 211 2244 245
rect 2168 209 2244 211
tri 2168 193 2184 209 ne
rect 2184 193 2228 209
tri 2228 193 2244 209 nw
rect 2274 289 2330 324
rect 2274 255 2286 289
rect 2320 255 2330 289
rect 2274 221 2330 255
tri 1944 155 1974 185 sw
tri 2050 155 2080 185 se
rect 2080 163 2138 187
tri 2138 163 2168 193 sw
tri 2244 163 2274 193 se
rect 2274 187 2286 221
rect 2320 187 2330 221
rect 2274 163 2330 187
rect 2080 155 2330 163
rect 1888 151 2330 155
rect 1888 117 1898 151
rect 1932 117 2092 151
rect 2126 117 2189 151
rect 2223 117 2286 151
rect 2320 117 2330 151
rect 1888 101 2330 117
<< pdiff >>
rect 107 1412 163 1450
rect 107 1378 117 1412
rect 151 1378 163 1412
rect 107 1344 163 1378
rect 107 1310 117 1344
rect 151 1310 163 1344
rect 107 1276 163 1310
rect 107 1242 117 1276
rect 151 1242 163 1276
rect 107 1208 163 1242
rect 107 1174 117 1208
rect 151 1174 163 1208
rect 107 1139 163 1174
rect 107 1105 117 1139
rect 151 1105 163 1139
rect 107 1050 163 1105
rect 193 1412 251 1450
rect 193 1378 205 1412
rect 239 1378 251 1412
rect 193 1344 251 1378
rect 193 1310 205 1344
rect 239 1310 251 1344
rect 193 1276 251 1310
rect 193 1242 205 1276
rect 239 1242 251 1276
rect 193 1208 251 1242
rect 193 1174 205 1208
rect 239 1174 251 1208
rect 193 1139 251 1174
rect 193 1105 205 1139
rect 239 1105 251 1139
rect 193 1050 251 1105
rect 281 1412 335 1450
rect 281 1378 293 1412
rect 327 1378 335 1412
rect 281 1344 335 1378
rect 281 1310 293 1344
rect 327 1310 335 1344
rect 281 1276 335 1310
rect 281 1242 293 1276
rect 327 1242 335 1276
rect 281 1208 335 1242
rect 281 1174 293 1208
rect 327 1174 335 1208
rect 281 1139 335 1174
rect 281 1105 293 1139
rect 327 1105 335 1139
rect 281 1050 335 1105
rect 575 1412 631 1450
rect 575 1378 585 1412
rect 619 1378 631 1412
rect 575 1344 631 1378
rect 575 1310 585 1344
rect 619 1310 631 1344
rect 575 1276 631 1310
rect 575 1242 585 1276
rect 619 1242 631 1276
rect 575 1208 631 1242
rect 575 1174 585 1208
rect 619 1174 631 1208
rect 575 1139 631 1174
rect 575 1105 585 1139
rect 619 1105 631 1139
rect 575 1050 631 1105
rect 661 1412 719 1450
rect 661 1378 673 1412
rect 707 1378 719 1412
rect 661 1344 719 1378
rect 661 1310 673 1344
rect 707 1310 719 1344
rect 661 1276 719 1310
rect 661 1242 673 1276
rect 707 1242 719 1276
rect 661 1208 719 1242
rect 661 1174 673 1208
rect 707 1174 719 1208
rect 661 1139 719 1174
rect 661 1105 673 1139
rect 707 1105 719 1139
rect 661 1050 719 1105
rect 749 1412 807 1450
rect 749 1378 761 1412
rect 795 1378 807 1412
rect 749 1344 807 1378
rect 749 1310 761 1344
rect 795 1310 807 1344
rect 749 1276 807 1310
rect 749 1242 761 1276
rect 795 1242 807 1276
rect 749 1208 807 1242
rect 749 1174 761 1208
rect 795 1174 807 1208
rect 749 1050 807 1174
rect 837 1412 895 1450
rect 837 1378 849 1412
rect 883 1378 895 1412
rect 837 1344 895 1378
rect 837 1310 849 1344
rect 883 1310 895 1344
rect 837 1276 895 1310
rect 837 1242 849 1276
rect 883 1242 895 1276
rect 837 1208 895 1242
rect 837 1174 849 1208
rect 883 1174 895 1208
rect 837 1139 895 1174
rect 837 1105 849 1139
rect 883 1105 895 1139
rect 837 1050 895 1105
rect 925 1412 979 1450
rect 925 1378 937 1412
rect 971 1378 979 1412
rect 925 1344 979 1378
rect 925 1310 937 1344
rect 971 1310 979 1344
rect 925 1276 979 1310
rect 925 1242 937 1276
rect 971 1242 979 1276
rect 925 1208 979 1242
rect 925 1174 937 1208
rect 971 1174 979 1208
rect 925 1050 979 1174
rect 1241 1412 1297 1450
rect 1241 1378 1251 1412
rect 1285 1378 1297 1412
rect 1241 1344 1297 1378
rect 1241 1310 1251 1344
rect 1285 1310 1297 1344
rect 1241 1276 1297 1310
rect 1241 1242 1251 1276
rect 1285 1242 1297 1276
rect 1241 1208 1297 1242
rect 1241 1174 1251 1208
rect 1285 1174 1297 1208
rect 1241 1139 1297 1174
rect 1241 1105 1251 1139
rect 1285 1105 1297 1139
rect 1241 1050 1297 1105
rect 1327 1412 1385 1450
rect 1327 1378 1339 1412
rect 1373 1378 1385 1412
rect 1327 1344 1385 1378
rect 1327 1310 1339 1344
rect 1373 1310 1385 1344
rect 1327 1276 1385 1310
rect 1327 1242 1339 1276
rect 1373 1242 1385 1276
rect 1327 1208 1385 1242
rect 1327 1174 1339 1208
rect 1373 1174 1385 1208
rect 1327 1139 1385 1174
rect 1327 1105 1339 1139
rect 1373 1105 1385 1139
rect 1327 1050 1385 1105
rect 1415 1412 1473 1450
rect 1415 1378 1427 1412
rect 1461 1378 1473 1412
rect 1415 1344 1473 1378
rect 1415 1310 1427 1344
rect 1461 1310 1473 1344
rect 1415 1276 1473 1310
rect 1415 1242 1427 1276
rect 1461 1242 1473 1276
rect 1415 1208 1473 1242
rect 1415 1174 1427 1208
rect 1461 1174 1473 1208
rect 1415 1050 1473 1174
rect 1503 1412 1561 1450
rect 1503 1378 1515 1412
rect 1549 1378 1561 1412
rect 1503 1344 1561 1378
rect 1503 1310 1515 1344
rect 1549 1310 1561 1344
rect 1503 1276 1561 1310
rect 1503 1242 1515 1276
rect 1549 1242 1561 1276
rect 1503 1208 1561 1242
rect 1503 1174 1515 1208
rect 1549 1174 1561 1208
rect 1503 1139 1561 1174
rect 1503 1105 1515 1139
rect 1549 1105 1561 1139
rect 1503 1050 1561 1105
rect 1591 1412 1645 1450
rect 1591 1378 1603 1412
rect 1637 1378 1645 1412
rect 1591 1344 1645 1378
rect 1591 1310 1603 1344
rect 1637 1310 1645 1344
rect 1591 1276 1645 1310
rect 1591 1242 1603 1276
rect 1637 1242 1645 1276
rect 1591 1208 1645 1242
rect 1591 1174 1603 1208
rect 1637 1174 1645 1208
rect 1591 1050 1645 1174
rect 1907 1412 1963 1450
rect 1907 1378 1917 1412
rect 1951 1378 1963 1412
rect 1907 1344 1963 1378
rect 1907 1310 1917 1344
rect 1951 1310 1963 1344
rect 1907 1276 1963 1310
rect 1907 1242 1917 1276
rect 1951 1242 1963 1276
rect 1907 1208 1963 1242
rect 1907 1174 1917 1208
rect 1951 1174 1963 1208
rect 1907 1139 1963 1174
rect 1907 1105 1917 1139
rect 1951 1105 1963 1139
rect 1907 1050 1963 1105
rect 1993 1412 2051 1450
rect 1993 1378 2005 1412
rect 2039 1378 2051 1412
rect 1993 1344 2051 1378
rect 1993 1310 2005 1344
rect 2039 1310 2051 1344
rect 1993 1276 2051 1310
rect 1993 1242 2005 1276
rect 2039 1242 2051 1276
rect 1993 1208 2051 1242
rect 1993 1174 2005 1208
rect 2039 1174 2051 1208
rect 1993 1139 2051 1174
rect 1993 1105 2005 1139
rect 2039 1105 2051 1139
rect 1993 1050 2051 1105
rect 2081 1412 2139 1450
rect 2081 1378 2093 1412
rect 2127 1378 2139 1412
rect 2081 1344 2139 1378
rect 2081 1310 2093 1344
rect 2127 1310 2139 1344
rect 2081 1276 2139 1310
rect 2081 1242 2093 1276
rect 2127 1242 2139 1276
rect 2081 1208 2139 1242
rect 2081 1174 2093 1208
rect 2127 1174 2139 1208
rect 2081 1050 2139 1174
rect 2169 1412 2227 1450
rect 2169 1378 2181 1412
rect 2215 1378 2227 1412
rect 2169 1344 2227 1378
rect 2169 1310 2181 1344
rect 2215 1310 2227 1344
rect 2169 1276 2227 1310
rect 2169 1242 2181 1276
rect 2215 1242 2227 1276
rect 2169 1208 2227 1242
rect 2169 1174 2181 1208
rect 2215 1174 2227 1208
rect 2169 1139 2227 1174
rect 2169 1105 2181 1139
rect 2215 1105 2227 1139
rect 2169 1050 2227 1105
rect 2257 1412 2311 1450
rect 2257 1378 2269 1412
rect 2303 1378 2311 1412
rect 2257 1344 2311 1378
rect 2257 1310 2269 1344
rect 2303 1310 2311 1344
rect 2257 1276 2311 1310
rect 2257 1242 2269 1276
rect 2303 1242 2311 1276
rect 2257 1208 2311 1242
rect 2257 1174 2269 1208
rect 2303 1174 2311 1208
rect 2257 1050 2311 1174
<< ndiffc >>
rect 109 327 143 361
rect 303 327 337 361
rect 109 255 143 289
rect 109 187 143 221
rect 205 211 239 245
rect 303 255 337 289
rect 303 187 337 221
rect 109 117 143 151
rect 205 117 239 151
rect 303 117 337 151
rect 566 327 600 361
rect 663 327 697 361
rect 760 327 794 361
rect 566 255 600 289
rect 566 187 600 221
rect 663 202 697 236
rect 760 255 794 289
rect 760 187 794 221
rect 857 211 891 245
rect 954 255 988 289
rect 954 187 988 221
rect 566 117 600 151
rect 760 117 794 151
rect 857 117 891 151
rect 954 117 988 151
rect 1232 327 1266 361
rect 1329 327 1363 361
rect 1426 327 1460 361
rect 1232 255 1266 289
rect 1232 187 1266 221
rect 1329 202 1363 236
rect 1426 255 1460 289
rect 1426 187 1460 221
rect 1523 211 1557 245
rect 1620 255 1654 289
rect 1620 187 1654 221
rect 1232 117 1266 151
rect 1426 117 1460 151
rect 1523 117 1557 151
rect 1620 117 1654 151
rect 1898 327 1932 361
rect 1995 327 2029 361
rect 2092 327 2126 361
rect 1898 255 1932 289
rect 1898 187 1932 221
rect 1995 202 2029 236
rect 2092 255 2126 289
rect 2092 187 2126 221
rect 2189 211 2223 245
rect 2286 255 2320 289
rect 2286 187 2320 221
rect 1898 117 1932 151
rect 2092 117 2126 151
rect 2189 117 2223 151
rect 2286 117 2320 151
<< pdiffc >>
rect 117 1378 151 1412
rect 117 1310 151 1344
rect 117 1242 151 1276
rect 117 1174 151 1208
rect 117 1105 151 1139
rect 205 1378 239 1412
rect 205 1310 239 1344
rect 205 1242 239 1276
rect 205 1174 239 1208
rect 205 1105 239 1139
rect 293 1378 327 1412
rect 293 1310 327 1344
rect 293 1242 327 1276
rect 293 1174 327 1208
rect 293 1105 327 1139
rect 585 1378 619 1412
rect 585 1310 619 1344
rect 585 1242 619 1276
rect 585 1174 619 1208
rect 585 1105 619 1139
rect 673 1378 707 1412
rect 673 1310 707 1344
rect 673 1242 707 1276
rect 673 1174 707 1208
rect 673 1105 707 1139
rect 761 1378 795 1412
rect 761 1310 795 1344
rect 761 1242 795 1276
rect 761 1174 795 1208
rect 849 1378 883 1412
rect 849 1310 883 1344
rect 849 1242 883 1276
rect 849 1174 883 1208
rect 849 1105 883 1139
rect 937 1378 971 1412
rect 937 1310 971 1344
rect 937 1242 971 1276
rect 937 1174 971 1208
rect 1251 1378 1285 1412
rect 1251 1310 1285 1344
rect 1251 1242 1285 1276
rect 1251 1174 1285 1208
rect 1251 1105 1285 1139
rect 1339 1378 1373 1412
rect 1339 1310 1373 1344
rect 1339 1242 1373 1276
rect 1339 1174 1373 1208
rect 1339 1105 1373 1139
rect 1427 1378 1461 1412
rect 1427 1310 1461 1344
rect 1427 1242 1461 1276
rect 1427 1174 1461 1208
rect 1515 1378 1549 1412
rect 1515 1310 1549 1344
rect 1515 1242 1549 1276
rect 1515 1174 1549 1208
rect 1515 1105 1549 1139
rect 1603 1378 1637 1412
rect 1603 1310 1637 1344
rect 1603 1242 1637 1276
rect 1603 1174 1637 1208
rect 1917 1378 1951 1412
rect 1917 1310 1951 1344
rect 1917 1242 1951 1276
rect 1917 1174 1951 1208
rect 1917 1105 1951 1139
rect 2005 1378 2039 1412
rect 2005 1310 2039 1344
rect 2005 1242 2039 1276
rect 2005 1174 2039 1208
rect 2005 1105 2039 1139
rect 2093 1378 2127 1412
rect 2093 1310 2127 1344
rect 2093 1242 2127 1276
rect 2093 1174 2127 1208
rect 2181 1378 2215 1412
rect 2181 1310 2215 1344
rect 2181 1242 2215 1276
rect 2181 1174 2215 1208
rect 2181 1105 2215 1139
rect 2269 1378 2303 1412
rect 2269 1310 2303 1344
rect 2269 1242 2303 1276
rect 2269 1174 2303 1208
<< psubdiff >>
rect -31 546 2473 572
rect -31 512 -17 546
rect 17 512 427 546
rect 461 512 1093 546
rect 1127 512 1759 546
rect 1793 512 2425 546
rect 2459 512 2473 546
rect -31 510 2473 512
rect -31 474 31 510
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect 413 474 475 510
rect -31 368 -17 402
rect 17 368 31 402
rect 413 440 427 474
rect 461 440 475 474
rect 413 402 475 440
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect 413 368 427 402
rect 461 368 475 402
rect 1079 474 1141 510
rect 1079 440 1093 474
rect 1127 440 1141 474
rect 1079 402 1141 440
rect 413 330 475 368
rect 413 296 427 330
rect 461 296 475 330
rect 413 258 475 296
rect 413 224 427 258
rect 461 224 475 258
rect 413 186 475 224
rect 413 152 427 186
rect 461 152 475 186
rect 413 114 475 152
rect -31 47 31 80
rect 413 80 427 114
rect 461 80 475 114
rect 1079 368 1093 402
rect 1127 368 1141 402
rect 1745 474 1807 510
rect 1745 440 1759 474
rect 1793 440 1807 474
rect 1745 402 1807 440
rect 1079 330 1141 368
rect 1079 296 1093 330
rect 1127 296 1141 330
rect 1079 258 1141 296
rect 1079 224 1093 258
rect 1127 224 1141 258
rect 1079 186 1141 224
rect 1079 152 1093 186
rect 1127 152 1141 186
rect 1079 114 1141 152
rect 413 47 475 80
rect 1079 80 1093 114
rect 1127 80 1141 114
rect 1745 368 1759 402
rect 1793 368 1807 402
rect 2411 474 2473 510
rect 2411 440 2425 474
rect 2459 440 2473 474
rect 2411 402 2473 440
rect 1745 330 1807 368
rect 1745 296 1759 330
rect 1793 296 1807 330
rect 1745 258 1807 296
rect 1745 224 1759 258
rect 1793 224 1807 258
rect 1745 186 1807 224
rect 1745 152 1759 186
rect 1793 152 1807 186
rect 1745 114 1807 152
rect 1079 47 1141 80
rect 1745 80 1759 114
rect 1793 80 1807 114
rect 2411 368 2425 402
rect 2459 368 2473 402
rect 2411 330 2473 368
rect 2411 296 2425 330
rect 2459 296 2473 330
rect 2411 258 2473 296
rect 2411 224 2425 258
rect 2459 224 2473 258
rect 2411 186 2473 224
rect 2411 152 2425 186
rect 2459 152 2473 186
rect 2411 114 2473 152
rect 1745 47 1807 80
rect 2411 80 2425 114
rect 2459 80 2473 114
rect 2411 47 2473 80
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 205 47
rect 239 13 283 47
rect 317 13 355 47
rect 389 13 499 47
rect 533 13 571 47
rect 605 13 643 47
rect 677 13 715 47
rect 749 13 805 47
rect 839 13 877 47
rect 911 13 949 47
rect 983 13 1021 47
rect 1055 13 1165 47
rect 1199 13 1237 47
rect 1271 13 1309 47
rect 1343 13 1381 47
rect 1415 13 1471 47
rect 1505 13 1543 47
rect 1577 13 1615 47
rect 1649 13 1687 47
rect 1721 13 1831 47
rect 1865 13 1903 47
rect 1937 13 1975 47
rect 2009 13 2047 47
rect 2081 13 2137 47
rect 2171 13 2209 47
rect 2243 13 2281 47
rect 2315 13 2353 47
rect 2387 13 2473 47
rect -31 11 31 13
rect 413 11 475 13
rect 1079 11 1141 13
rect 1745 11 1807 13
rect 2411 11 2473 13
<< nsubdiff >>
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 205 1539
rect 239 1505 283 1539
rect 317 1505 355 1539
rect 389 1505 499 1539
rect 533 1505 571 1539
rect 605 1505 643 1539
rect 677 1505 715 1539
rect 749 1505 805 1539
rect 839 1505 877 1539
rect 911 1505 949 1539
rect 983 1505 1021 1539
rect 1055 1505 1165 1539
rect 1199 1505 1237 1539
rect 1271 1505 1309 1539
rect 1343 1505 1381 1539
rect 1415 1505 1471 1539
rect 1505 1505 1543 1539
rect 1577 1505 1615 1539
rect 1649 1505 1687 1539
rect 1721 1505 1831 1539
rect 1865 1505 1903 1539
rect 1937 1505 1975 1539
rect 2009 1505 2047 1539
rect 2081 1505 2137 1539
rect 2171 1505 2209 1539
rect 2243 1505 2281 1539
rect 2315 1505 2353 1539
rect 2387 1505 2473 1539
rect -31 1470 31 1505
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect 413 1470 475 1505
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect -31 1038 31 1076
rect 413 1436 427 1470
rect 461 1436 475 1470
rect 1079 1470 1141 1505
rect 413 1398 475 1436
rect 413 1364 427 1398
rect 461 1364 475 1398
rect 413 1326 475 1364
rect 413 1292 427 1326
rect 461 1292 475 1326
rect 413 1254 475 1292
rect 413 1220 427 1254
rect 461 1220 475 1254
rect 413 1182 475 1220
rect 413 1148 427 1182
rect 461 1148 475 1182
rect 413 1110 475 1148
rect 413 1076 427 1110
rect 461 1076 475 1110
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect 413 1038 475 1076
rect 1079 1436 1093 1470
rect 1127 1436 1141 1470
rect 1745 1470 1807 1505
rect 1079 1398 1141 1436
rect 1079 1364 1093 1398
rect 1127 1364 1141 1398
rect 1079 1326 1141 1364
rect 1079 1292 1093 1326
rect 1127 1292 1141 1326
rect 1079 1254 1141 1292
rect 1079 1220 1093 1254
rect 1127 1220 1141 1254
rect 1079 1182 1141 1220
rect 1079 1148 1093 1182
rect 1127 1148 1141 1182
rect 1079 1110 1141 1148
rect 1079 1076 1093 1110
rect 1127 1076 1141 1110
rect 413 1004 427 1038
rect 461 1004 475 1038
rect 413 966 475 1004
rect -31 930 31 932
rect 413 932 427 966
rect 461 932 475 966
rect 1079 1038 1141 1076
rect 1745 1436 1759 1470
rect 1793 1436 1807 1470
rect 2411 1470 2473 1505
rect 1745 1398 1807 1436
rect 1745 1364 1759 1398
rect 1793 1364 1807 1398
rect 1745 1326 1807 1364
rect 1745 1292 1759 1326
rect 1793 1292 1807 1326
rect 1745 1254 1807 1292
rect 1745 1220 1759 1254
rect 1793 1220 1807 1254
rect 1745 1182 1807 1220
rect 1745 1148 1759 1182
rect 1793 1148 1807 1182
rect 1745 1110 1807 1148
rect 1745 1076 1759 1110
rect 1793 1076 1807 1110
rect 1079 1004 1093 1038
rect 1127 1004 1141 1038
rect 1079 966 1141 1004
rect 413 930 475 932
rect 1079 932 1093 966
rect 1127 932 1141 966
rect 1745 1038 1807 1076
rect 2411 1436 2425 1470
rect 2459 1436 2473 1470
rect 2411 1398 2473 1436
rect 2411 1364 2425 1398
rect 2459 1364 2473 1398
rect 2411 1326 2473 1364
rect 2411 1292 2425 1326
rect 2459 1292 2473 1326
rect 2411 1254 2473 1292
rect 2411 1220 2425 1254
rect 2459 1220 2473 1254
rect 2411 1182 2473 1220
rect 2411 1148 2425 1182
rect 2459 1148 2473 1182
rect 2411 1110 2473 1148
rect 2411 1076 2425 1110
rect 2459 1076 2473 1110
rect 1745 1004 1759 1038
rect 1793 1004 1807 1038
rect 1745 966 1807 1004
rect 1079 930 1141 932
rect 1745 932 1759 966
rect 1793 932 1807 966
rect 2411 1038 2473 1076
rect 2411 1004 2425 1038
rect 2459 1004 2473 1038
rect 2411 966 2473 1004
rect 1745 930 1807 932
rect 2411 932 2425 966
rect 2459 932 2473 966
rect 2411 930 2473 932
rect -31 868 2473 930
<< psubdiffcont >>
rect -17 512 17 546
rect 427 512 461 546
rect 1093 512 1127 546
rect 1759 512 1793 546
rect 2425 512 2459 546
rect -17 440 17 474
rect -17 368 17 402
rect 427 440 461 474
rect -17 296 17 330
rect -17 224 17 258
rect -17 152 17 186
rect -17 80 17 114
rect 427 368 461 402
rect 1093 440 1127 474
rect 427 296 461 330
rect 427 224 461 258
rect 427 152 461 186
rect 427 80 461 114
rect 1093 368 1127 402
rect 1759 440 1793 474
rect 1093 296 1127 330
rect 1093 224 1127 258
rect 1093 152 1127 186
rect 1093 80 1127 114
rect 1759 368 1793 402
rect 2425 440 2459 474
rect 1759 296 1793 330
rect 1759 224 1793 258
rect 1759 152 1793 186
rect 1759 80 1793 114
rect 2425 368 2459 402
rect 2425 296 2459 330
rect 2425 224 2459 258
rect 2425 152 2459 186
rect 2425 80 2459 114
rect 55 13 89 47
rect 127 13 161 47
rect 205 13 239 47
rect 283 13 317 47
rect 355 13 389 47
rect 499 13 533 47
rect 571 13 605 47
rect 643 13 677 47
rect 715 13 749 47
rect 805 13 839 47
rect 877 13 911 47
rect 949 13 983 47
rect 1021 13 1055 47
rect 1165 13 1199 47
rect 1237 13 1271 47
rect 1309 13 1343 47
rect 1381 13 1415 47
rect 1471 13 1505 47
rect 1543 13 1577 47
rect 1615 13 1649 47
rect 1687 13 1721 47
rect 1831 13 1865 47
rect 1903 13 1937 47
rect 1975 13 2009 47
rect 2047 13 2081 47
rect 2137 13 2171 47
rect 2209 13 2243 47
rect 2281 13 2315 47
rect 2353 13 2387 47
<< nsubdiffcont >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 205 1505 239 1539
rect 283 1505 317 1539
rect 355 1505 389 1539
rect 499 1505 533 1539
rect 571 1505 605 1539
rect 643 1505 677 1539
rect 715 1505 749 1539
rect 805 1505 839 1539
rect 877 1505 911 1539
rect 949 1505 983 1539
rect 1021 1505 1055 1539
rect 1165 1505 1199 1539
rect 1237 1505 1271 1539
rect 1309 1505 1343 1539
rect 1381 1505 1415 1539
rect 1471 1505 1505 1539
rect 1543 1505 1577 1539
rect 1615 1505 1649 1539
rect 1687 1505 1721 1539
rect 1831 1505 1865 1539
rect 1903 1505 1937 1539
rect 1975 1505 2009 1539
rect 2047 1505 2081 1539
rect 2137 1505 2171 1539
rect 2209 1505 2243 1539
rect 2281 1505 2315 1539
rect 2353 1505 2387 1539
rect -17 1436 17 1470
rect -17 1364 17 1398
rect -17 1292 17 1326
rect -17 1220 17 1254
rect -17 1148 17 1182
rect -17 1076 17 1110
rect 427 1436 461 1470
rect 427 1364 461 1398
rect 427 1292 461 1326
rect 427 1220 461 1254
rect 427 1148 461 1182
rect 427 1076 461 1110
rect -17 1004 17 1038
rect -17 932 17 966
rect 1093 1436 1127 1470
rect 1093 1364 1127 1398
rect 1093 1292 1127 1326
rect 1093 1220 1127 1254
rect 1093 1148 1127 1182
rect 1093 1076 1127 1110
rect 427 1004 461 1038
rect 427 932 461 966
rect 1759 1436 1793 1470
rect 1759 1364 1793 1398
rect 1759 1292 1793 1326
rect 1759 1220 1793 1254
rect 1759 1148 1793 1182
rect 1759 1076 1793 1110
rect 1093 1004 1127 1038
rect 1093 932 1127 966
rect 2425 1436 2459 1470
rect 2425 1364 2459 1398
rect 2425 1292 2459 1326
rect 2425 1220 2459 1254
rect 2425 1148 2459 1182
rect 2425 1076 2459 1110
rect 1759 1004 1793 1038
rect 1759 932 1793 966
rect 2425 1004 2459 1038
rect 2425 932 2459 966
<< poly >>
rect 163 1450 193 1476
rect 251 1450 281 1476
rect 631 1450 661 1476
rect 719 1450 749 1476
rect 807 1450 837 1476
rect 895 1450 925 1476
rect 163 1019 193 1050
rect 251 1019 281 1050
rect 121 1003 281 1019
rect 121 969 131 1003
rect 165 989 281 1003
rect 1297 1450 1327 1476
rect 1385 1450 1415 1476
rect 1473 1450 1503 1476
rect 1561 1450 1591 1476
rect 165 969 175 989
rect 121 953 175 969
rect 631 1019 661 1050
rect 719 1019 749 1050
rect 807 1019 837 1050
rect 895 1019 925 1050
rect 631 1003 749 1019
rect 631 989 649 1003
rect 639 969 649 989
rect 683 989 749 1003
rect 793 1003 925 1019
rect 683 969 693 989
rect 639 953 693 969
rect 793 969 803 1003
rect 837 989 925 1003
rect 1963 1450 1993 1476
rect 2051 1450 2081 1476
rect 2139 1450 2169 1476
rect 2227 1450 2257 1476
rect 837 969 847 989
rect 793 953 847 969
rect 1297 1019 1327 1050
rect 1385 1019 1415 1050
rect 1473 1019 1503 1050
rect 1561 1019 1591 1050
rect 1297 1003 1415 1019
rect 1297 989 1315 1003
rect 1305 969 1315 989
rect 1349 989 1415 1003
rect 1459 1003 1591 1019
rect 1349 969 1359 989
rect 1305 953 1359 969
rect 1459 969 1469 1003
rect 1503 989 1591 1003
rect 1503 969 1513 989
rect 1459 953 1513 969
rect 1963 1019 1993 1050
rect 2051 1019 2081 1050
rect 2139 1019 2169 1050
rect 2227 1019 2257 1050
rect 1963 1003 2081 1019
rect 1963 989 1981 1003
rect 1971 969 1981 989
rect 2015 989 2081 1003
rect 2125 1003 2257 1019
rect 2015 969 2025 989
rect 1971 953 2025 969
rect 2125 969 2135 1003
rect 2169 989 2257 1003
rect 2169 969 2179 989
rect 2125 953 2179 969
rect 121 461 175 477
rect 121 427 131 461
rect 165 441 175 461
rect 165 427 185 441
rect 121 411 185 427
rect 155 377 185 411
rect 639 461 693 477
rect 639 441 649 461
rect 612 427 649 441
rect 683 427 693 461
rect 612 411 693 427
rect 787 461 841 477
rect 787 427 797 461
rect 831 427 841 461
rect 787 411 841 427
rect 1305 461 1359 477
rect 1305 441 1315 461
rect 612 377 642 411
rect 806 377 836 411
rect 1278 427 1315 441
rect 1349 427 1359 461
rect 1278 411 1359 427
rect 1453 461 1507 477
rect 1453 427 1463 461
rect 1497 427 1507 461
rect 1453 411 1507 427
rect 1971 461 2025 477
rect 1971 441 1981 461
rect 1278 377 1308 411
rect 1472 377 1502 411
rect 1944 427 1981 441
rect 2015 427 2025 461
rect 1944 411 2025 427
rect 2119 461 2173 477
rect 2119 427 2129 461
rect 2163 427 2173 461
rect 2119 411 2173 427
rect 1944 377 1974 411
rect 2138 377 2168 411
<< polycont >>
rect 131 969 165 1003
rect 649 969 683 1003
rect 803 969 837 1003
rect 1315 969 1349 1003
rect 1469 969 1503 1003
rect 1981 969 2015 1003
rect 2135 969 2169 1003
rect 131 427 165 461
rect 649 427 683 461
rect 797 427 831 461
rect 1315 427 1349 461
rect 1463 427 1497 461
rect 1981 427 2015 461
rect 2129 427 2163 461
<< locali >>
rect -31 1539 2473 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 205 1539
rect 239 1505 283 1539
rect 317 1505 355 1539
rect 389 1505 499 1539
rect 533 1505 571 1539
rect 605 1505 643 1539
rect 677 1505 715 1539
rect 749 1505 805 1539
rect 839 1505 877 1539
rect 911 1505 949 1539
rect 983 1505 1021 1539
rect 1055 1505 1165 1539
rect 1199 1505 1237 1539
rect 1271 1505 1309 1539
rect 1343 1505 1381 1539
rect 1415 1505 1471 1539
rect 1505 1505 1543 1539
rect 1577 1505 1615 1539
rect 1649 1505 1687 1539
rect 1721 1505 1831 1539
rect 1865 1505 1903 1539
rect 1937 1505 1975 1539
rect 2009 1505 2047 1539
rect 2081 1505 2137 1539
rect 2171 1505 2209 1539
rect 2243 1505 2281 1539
rect 2315 1505 2353 1539
rect 2387 1505 2473 1539
rect -31 1492 2473 1505
rect -31 1470 31 1492
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect 117 1412 151 1492
rect 117 1344 151 1378
rect 117 1276 151 1310
rect 117 1208 151 1242
rect 117 1139 151 1174
rect 117 1083 151 1105
rect 205 1412 239 1450
rect 205 1344 239 1378
rect 205 1276 239 1310
rect 205 1208 239 1242
rect 205 1139 239 1174
rect -31 1038 31 1076
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect -31 868 31 932
rect 131 1003 165 1019
rect 131 609 165 969
rect 205 979 239 1105
rect 293 1412 327 1492
rect 293 1344 327 1378
rect 293 1276 327 1310
rect 293 1208 327 1242
rect 293 1139 327 1174
rect 293 1083 327 1105
rect 413 1470 475 1492
rect 413 1436 427 1470
rect 461 1436 475 1470
rect 413 1398 475 1436
rect 413 1364 427 1398
rect 461 1364 475 1398
rect 413 1326 475 1364
rect 413 1292 427 1326
rect 461 1292 475 1326
rect 413 1254 475 1292
rect 413 1220 427 1254
rect 461 1220 475 1254
rect 413 1182 475 1220
rect 413 1148 427 1182
rect 461 1148 475 1182
rect 413 1110 475 1148
rect 413 1076 427 1110
rect 461 1076 475 1110
rect 413 1038 475 1076
rect 585 1412 619 1492
rect 585 1344 619 1378
rect 585 1276 619 1310
rect 585 1208 619 1242
rect 585 1139 619 1174
rect 585 1073 619 1105
rect 673 1412 707 1450
rect 673 1344 707 1378
rect 673 1276 707 1310
rect 673 1208 707 1242
rect 673 1139 707 1174
rect 761 1412 795 1492
rect 761 1344 795 1378
rect 761 1276 795 1310
rect 761 1208 795 1242
rect 761 1157 795 1174
rect 849 1412 883 1450
rect 849 1344 883 1378
rect 849 1276 883 1310
rect 849 1208 883 1242
rect 673 1103 707 1105
rect 849 1139 883 1174
rect 937 1412 971 1492
rect 937 1344 971 1378
rect 937 1276 971 1310
rect 937 1208 971 1242
rect 937 1157 971 1174
rect 1079 1470 1141 1492
rect 1079 1436 1093 1470
rect 1127 1436 1141 1470
rect 1079 1398 1141 1436
rect 1079 1364 1093 1398
rect 1127 1364 1141 1398
rect 1079 1326 1141 1364
rect 1079 1292 1093 1326
rect 1127 1292 1141 1326
rect 1079 1254 1141 1292
rect 1079 1220 1093 1254
rect 1127 1220 1141 1254
rect 1079 1182 1141 1220
rect 849 1103 883 1105
rect 1079 1148 1093 1182
rect 1127 1148 1141 1182
rect 1079 1110 1141 1148
rect 673 1069 979 1103
rect 413 1004 427 1038
rect 461 1004 475 1038
rect 205 945 313 979
rect -31 546 31 572
rect -31 512 -17 546
rect 17 512 31 546
rect -31 474 31 512
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect 131 461 165 575
rect 279 683 313 945
rect 413 966 475 1004
rect 413 932 427 966
rect 461 932 475 966
rect 413 868 475 932
rect 649 1003 683 1019
rect 803 1003 837 1019
rect 279 461 313 649
rect 649 609 683 969
rect 131 411 165 427
rect 205 427 313 461
rect 413 546 475 572
rect 413 512 427 546
rect 461 512 475 546
rect 413 474 475 512
rect 413 440 427 474
rect 461 440 475 474
rect -31 368 -17 402
rect 17 368 31 402
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect -31 62 31 80
rect 109 361 143 377
rect 109 289 143 327
rect 109 221 143 255
rect 205 245 239 427
rect 413 402 475 440
rect 649 461 683 575
rect 649 411 683 427
rect 797 969 803 988
rect 797 953 837 969
rect 797 757 831 953
rect 797 461 831 723
rect 797 411 831 427
rect 945 609 979 1069
rect 1079 1076 1093 1110
rect 1127 1076 1141 1110
rect 1079 1038 1141 1076
rect 1251 1412 1285 1492
rect 1251 1344 1285 1378
rect 1251 1276 1285 1310
rect 1251 1208 1285 1242
rect 1251 1139 1285 1174
rect 1251 1073 1285 1105
rect 1339 1412 1373 1450
rect 1339 1344 1373 1378
rect 1339 1276 1373 1310
rect 1339 1208 1373 1242
rect 1339 1139 1373 1174
rect 1427 1412 1461 1492
rect 1427 1344 1461 1378
rect 1427 1276 1461 1310
rect 1427 1208 1461 1242
rect 1427 1157 1461 1174
rect 1515 1412 1549 1450
rect 1515 1344 1549 1378
rect 1515 1276 1549 1310
rect 1515 1208 1549 1242
rect 1339 1103 1373 1105
rect 1515 1139 1549 1174
rect 1603 1412 1637 1492
rect 1603 1344 1637 1378
rect 1603 1276 1637 1310
rect 1603 1208 1637 1242
rect 1603 1157 1637 1174
rect 1745 1470 1807 1492
rect 1745 1436 1759 1470
rect 1793 1436 1807 1470
rect 1745 1398 1807 1436
rect 1745 1364 1759 1398
rect 1793 1364 1807 1398
rect 1745 1326 1807 1364
rect 1745 1292 1759 1326
rect 1793 1292 1807 1326
rect 1745 1254 1807 1292
rect 1745 1220 1759 1254
rect 1793 1220 1807 1254
rect 1745 1182 1807 1220
rect 1515 1103 1549 1105
rect 1745 1148 1759 1182
rect 1793 1148 1807 1182
rect 1745 1110 1807 1148
rect 1339 1069 1645 1103
rect 1079 1004 1093 1038
rect 1127 1004 1141 1038
rect 1079 966 1141 1004
rect 1079 932 1093 966
rect 1127 932 1141 966
rect 1079 868 1141 932
rect 1315 1003 1349 1019
rect 1469 1003 1503 1019
rect 205 195 239 211
rect 303 361 337 377
rect 303 289 337 327
rect 303 221 337 255
rect 109 151 143 187
rect 303 151 337 187
rect 143 117 205 151
rect 239 117 303 151
rect 109 62 143 117
rect 206 62 240 117
rect 303 62 337 117
rect 413 368 427 402
rect 461 368 475 402
rect 413 330 475 368
rect 413 296 427 330
rect 461 296 475 330
rect 413 258 475 296
rect 413 224 427 258
rect 461 224 475 258
rect 413 186 475 224
rect 413 152 427 186
rect 461 152 475 186
rect 413 114 475 152
rect 413 80 427 114
rect 461 80 475 114
rect 566 361 600 377
rect 760 361 794 377
rect 945 376 979 575
rect 1315 683 1349 969
rect 600 327 663 361
rect 697 327 760 361
rect 566 289 600 327
rect 566 221 600 255
rect 760 289 794 327
rect 566 151 600 187
rect 566 101 600 117
rect 663 236 697 252
rect 413 62 475 80
rect 663 62 697 202
rect 760 221 794 255
rect 857 342 979 376
rect 1079 546 1141 572
rect 1079 512 1093 546
rect 1127 512 1141 546
rect 1079 474 1141 512
rect 1079 440 1093 474
rect 1127 440 1141 474
rect 1079 402 1141 440
rect 1315 461 1349 649
rect 1315 411 1349 427
rect 1463 969 1469 988
rect 1463 953 1503 969
rect 1463 831 1497 953
rect 1463 461 1497 797
rect 1463 411 1497 427
rect 1611 683 1645 1069
rect 1745 1076 1759 1110
rect 1793 1076 1807 1110
rect 1745 1038 1807 1076
rect 1917 1412 1951 1492
rect 1917 1344 1951 1378
rect 1917 1276 1951 1310
rect 1917 1208 1951 1242
rect 1917 1139 1951 1174
rect 1917 1073 1951 1105
rect 2005 1412 2039 1450
rect 2005 1344 2039 1378
rect 2005 1276 2039 1310
rect 2005 1208 2039 1242
rect 2005 1139 2039 1174
rect 2093 1412 2127 1492
rect 2093 1344 2127 1378
rect 2093 1276 2127 1310
rect 2093 1208 2127 1242
rect 2093 1157 2127 1174
rect 2181 1412 2215 1450
rect 2181 1344 2215 1378
rect 2181 1276 2215 1310
rect 2181 1208 2215 1242
rect 2005 1103 2039 1105
rect 2181 1139 2215 1174
rect 2269 1412 2303 1492
rect 2269 1344 2303 1378
rect 2269 1276 2303 1310
rect 2269 1208 2303 1242
rect 2269 1157 2303 1174
rect 2411 1470 2473 1492
rect 2411 1436 2425 1470
rect 2459 1436 2473 1470
rect 2411 1398 2473 1436
rect 2411 1364 2425 1398
rect 2459 1364 2473 1398
rect 2411 1326 2473 1364
rect 2411 1292 2425 1326
rect 2459 1292 2473 1326
rect 2411 1254 2473 1292
rect 2411 1220 2425 1254
rect 2459 1220 2473 1254
rect 2411 1182 2473 1220
rect 2181 1103 2215 1105
rect 2411 1148 2425 1182
rect 2459 1148 2473 1182
rect 2411 1110 2473 1148
rect 2005 1069 2311 1103
rect 1745 1004 1759 1038
rect 1793 1004 1807 1038
rect 1745 966 1807 1004
rect 1745 932 1759 966
rect 1793 932 1807 966
rect 1745 868 1807 932
rect 1981 1003 2015 1019
rect 2135 1003 2169 1019
rect 1079 368 1093 402
rect 1127 368 1141 402
rect 857 245 891 342
rect 1079 330 1141 368
rect 857 195 891 211
rect 954 289 988 305
rect 954 221 988 255
rect 760 151 794 187
rect 954 151 988 187
rect 794 117 857 151
rect 891 117 954 151
rect 760 101 794 117
rect 954 101 988 117
rect 1079 296 1093 330
rect 1127 296 1141 330
rect 1079 258 1141 296
rect 1079 224 1093 258
rect 1127 224 1141 258
rect 1079 186 1141 224
rect 1079 152 1093 186
rect 1127 152 1141 186
rect 1079 114 1141 152
rect 1079 80 1093 114
rect 1127 80 1141 114
rect 1232 361 1266 377
rect 1426 361 1460 377
rect 1611 376 1645 649
rect 1981 609 2015 969
rect 1266 327 1329 361
rect 1363 327 1426 361
rect 1232 289 1266 327
rect 1232 221 1266 255
rect 1426 289 1460 327
rect 1232 151 1266 187
rect 1232 101 1266 117
rect 1329 236 1363 252
rect 1079 62 1141 80
rect 1329 62 1363 202
rect 1426 221 1460 255
rect 1523 342 1645 376
rect 1745 546 1807 572
rect 1745 512 1759 546
rect 1793 512 1807 546
rect 1745 474 1807 512
rect 1745 440 1759 474
rect 1793 440 1807 474
rect 1745 402 1807 440
rect 1981 461 2015 575
rect 1981 411 2015 427
rect 2129 969 2135 988
rect 2129 953 2169 969
rect 2129 683 2163 953
rect 2129 461 2163 649
rect 2129 411 2163 427
rect 2277 683 2311 1069
rect 2411 1076 2425 1110
rect 2459 1076 2473 1110
rect 2411 1038 2473 1076
rect 2411 1004 2425 1038
rect 2459 1004 2473 1038
rect 2411 966 2473 1004
rect 2411 932 2425 966
rect 2459 932 2473 966
rect 2411 868 2473 932
rect 1745 368 1759 402
rect 1793 368 1807 402
rect 1523 245 1557 342
rect 1745 330 1807 368
rect 1523 195 1557 211
rect 1620 289 1654 305
rect 1620 221 1654 255
rect 1426 151 1460 187
rect 1620 151 1654 187
rect 1460 117 1523 151
rect 1557 117 1620 151
rect 1426 101 1460 117
rect 1620 101 1654 117
rect 1745 296 1759 330
rect 1793 296 1807 330
rect 1745 258 1807 296
rect 1745 224 1759 258
rect 1793 224 1807 258
rect 1745 186 1807 224
rect 1745 152 1759 186
rect 1793 152 1807 186
rect 1745 114 1807 152
rect 1745 80 1759 114
rect 1793 80 1807 114
rect 1898 361 1932 377
rect 2092 361 2126 377
rect 2277 376 2311 649
rect 1932 327 1995 361
rect 2029 327 2092 361
rect 1898 289 1932 327
rect 1898 221 1932 255
rect 2092 289 2126 327
rect 1898 151 1932 187
rect 1898 101 1932 117
rect 1995 236 2029 252
rect 1745 62 1807 80
rect 1995 62 2029 202
rect 2092 221 2126 255
rect 2189 342 2311 376
rect 2411 546 2473 572
rect 2411 512 2425 546
rect 2459 512 2473 546
rect 2411 474 2473 512
rect 2411 440 2425 474
rect 2459 440 2473 474
rect 2411 402 2473 440
rect 2411 368 2425 402
rect 2459 368 2473 402
rect 2189 245 2223 342
rect 2411 330 2473 368
rect 2189 195 2223 211
rect 2286 289 2320 305
rect 2286 221 2320 255
rect 2092 151 2126 187
rect 2286 151 2320 187
rect 2126 117 2189 151
rect 2223 117 2286 151
rect 2092 101 2126 117
rect 2286 101 2320 117
rect 2411 296 2425 330
rect 2459 296 2473 330
rect 2411 258 2473 296
rect 2411 224 2425 258
rect 2459 224 2473 258
rect 2411 186 2473 224
rect 2411 152 2425 186
rect 2459 152 2473 186
rect 2411 114 2473 152
rect 2411 80 2425 114
rect 2459 80 2473 114
rect 2411 62 2473 80
rect -31 47 2473 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 205 47
rect 239 13 283 47
rect 317 13 355 47
rect 389 13 499 47
rect 533 13 571 47
rect 605 13 643 47
rect 677 13 715 47
rect 749 13 805 47
rect 839 13 877 47
rect 911 13 949 47
rect 983 13 1021 47
rect 1055 13 1165 47
rect 1199 13 1237 47
rect 1271 13 1309 47
rect 1343 13 1381 47
rect 1415 13 1471 47
rect 1505 13 1543 47
rect 1577 13 1615 47
rect 1649 13 1687 47
rect 1721 13 1831 47
rect 1865 13 1903 47
rect 1937 13 1975 47
rect 2009 13 2047 47
rect 2081 13 2137 47
rect 2171 13 2209 47
rect 2243 13 2281 47
rect 2315 13 2353 47
rect 2387 13 2473 47
rect -31 0 2473 13
<< viali >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 205 1505 239 1539
rect 283 1505 317 1539
rect 355 1505 389 1539
rect 499 1505 533 1539
rect 571 1505 605 1539
rect 643 1505 677 1539
rect 715 1505 749 1539
rect 805 1505 839 1539
rect 877 1505 911 1539
rect 949 1505 983 1539
rect 1021 1505 1055 1539
rect 1165 1505 1199 1539
rect 1237 1505 1271 1539
rect 1309 1505 1343 1539
rect 1381 1505 1415 1539
rect 1471 1505 1505 1539
rect 1543 1505 1577 1539
rect 1615 1505 1649 1539
rect 1687 1505 1721 1539
rect 1831 1505 1865 1539
rect 1903 1505 1937 1539
rect 1975 1505 2009 1539
rect 2047 1505 2081 1539
rect 2137 1505 2171 1539
rect 2209 1505 2243 1539
rect 2281 1505 2315 1539
rect 2353 1505 2387 1539
rect 131 575 165 609
rect 279 649 313 683
rect 649 575 683 609
rect 797 723 831 757
rect 945 575 979 609
rect 1315 649 1349 683
rect 1463 797 1497 831
rect 1611 649 1645 683
rect 1981 575 2015 609
rect 2129 649 2163 683
rect 2277 649 2311 683
rect 55 13 89 47
rect 127 13 161 47
rect 205 13 239 47
rect 283 13 317 47
rect 355 13 389 47
rect 499 13 533 47
rect 571 13 605 47
rect 643 13 677 47
rect 715 13 749 47
rect 805 13 839 47
rect 877 13 911 47
rect 949 13 983 47
rect 1021 13 1055 47
rect 1165 13 1199 47
rect 1237 13 1271 47
rect 1309 13 1343 47
rect 1381 13 1415 47
rect 1471 13 1505 47
rect 1543 13 1577 47
rect 1615 13 1649 47
rect 1687 13 1721 47
rect 1831 13 1865 47
rect 1903 13 1937 47
rect 1975 13 2009 47
rect 2047 13 2081 47
rect 2137 13 2171 47
rect 2209 13 2243 47
rect 2281 13 2315 47
rect 2353 13 2387 47
<< metal1 >>
rect -31 1539 2473 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 205 1539
rect 239 1505 283 1539
rect 317 1505 355 1539
rect 389 1505 499 1539
rect 533 1505 571 1539
rect 605 1505 643 1539
rect 677 1505 715 1539
rect 749 1505 805 1539
rect 839 1505 877 1539
rect 911 1505 949 1539
rect 983 1505 1021 1539
rect 1055 1505 1165 1539
rect 1199 1505 1237 1539
rect 1271 1505 1309 1539
rect 1343 1505 1381 1539
rect 1415 1505 1471 1539
rect 1505 1505 1543 1539
rect 1577 1505 1615 1539
rect 1649 1505 1687 1539
rect 1721 1505 1831 1539
rect 1865 1505 1903 1539
rect 1937 1505 1975 1539
rect 2009 1505 2047 1539
rect 2081 1505 2137 1539
rect 2171 1505 2209 1539
rect 2243 1505 2281 1539
rect 2315 1505 2353 1539
rect 2387 1505 2473 1539
rect -31 1492 2473 1505
rect 1457 831 1503 837
rect 1427 797 1463 831
rect 1497 797 1509 831
rect 1457 791 1503 797
rect 791 757 837 763
rect 761 723 797 757
rect 831 723 843 757
rect 791 717 837 723
rect 273 683 319 689
rect 1309 683 1355 689
rect 1605 683 1651 689
rect 2123 683 2169 689
rect 2271 683 2317 689
rect 267 649 279 683
rect 313 649 1315 683
rect 1349 649 1361 683
rect 1599 649 1611 683
rect 1645 649 2129 683
rect 2163 649 2175 683
rect 2265 649 2277 683
rect 2311 649 2347 683
rect 273 643 319 649
rect 1309 643 1355 649
rect 1605 643 1651 649
rect 2123 643 2169 649
rect 2271 643 2317 649
rect 125 609 171 615
rect 643 609 689 615
rect 939 609 985 615
rect 1975 609 2021 615
rect 95 575 131 609
rect 165 575 649 609
rect 683 575 695 609
rect 933 575 945 609
rect 979 575 1981 609
rect 2015 575 2027 609
rect 125 569 171 575
rect 643 569 689 575
rect 939 569 985 575
rect 1975 569 2021 575
rect -31 47 2473 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 205 47
rect 239 13 283 47
rect 317 13 355 47
rect 389 13 499 47
rect 533 13 571 47
rect 605 13 643 47
rect 677 13 715 47
rect 749 13 805 47
rect 839 13 877 47
rect 911 13 949 47
rect 983 13 1021 47
rect 1055 13 1165 47
rect 1199 13 1237 47
rect 1271 13 1309 47
rect 1343 13 1381 47
rect 1415 13 1471 47
rect 1505 13 1543 47
rect 1577 13 1615 47
rect 1649 13 1687 47
rect 1721 13 1831 47
rect 1865 13 1903 47
rect 1937 13 1975 47
rect 2009 13 2047 47
rect 2081 13 2137 47
rect 2171 13 2209 47
rect 2243 13 2281 47
rect 2315 13 2353 47
rect 2387 13 2473 47
rect -31 0 2473 13
<< labels >>
rlabel metal1 2277 649 2311 683 1 Y
port 1 n
rlabel metal1 797 723 831 757 1 A0
port 2 n
rlabel metal1 1463 797 1497 831 1 A1
port 3 n
rlabel metal1 131 575 165 609 1 S
port 4 n
rlabel metal1 72 1522 72 1522 1 VDD
port 5 n
rlabel metal1 72 30 72 30 1 VSS
port 6 n
<< end >>
