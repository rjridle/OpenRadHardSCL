* SPICE3 file created from DFFRNQNX1.ext - technology: sky130A

.subckt DFFRNQNX1 QN D CLK RN VDD GND
X0 a_599_989.t3 D.t0 VDD.t43 0��&�U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X1 VDD.t37 CLK.t0 a_277_1050.t6  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X2 VDD.t13 a_599_989.t7 a_2141_1050.t3 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X3 VDD.t47 a_277_1050.t7 QN.t2  �O� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X4 a_599_989.t1 RN.t0 VDD.t39 ��O� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X5 a_147_187.t3 CLK.t1 VDD.t19  �O� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X6 QN.t0 a_4151_989.t5 VDD.t27 ��O� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X7 a_4151_989.t4 QN.t7 VDD.t29  �O� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X8 VDD.t9 a_599_989.t8 a_277_1050.t3 ��O� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X9 VDD.t49 a_147_187.t9 a_2141_1050.t4  �O� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X10 VDD.t53 a_2141_1050.t5 a_147_187.t1 ��O� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X11 a_147_187.t4 RN.t1 VDD.t59  �O� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X12 GND a_147_187.t12 a_91_103.t0 GND sky130_fd_pr__nfet_01v8 ad=1.0746p pd=9.42u as=0p ps=0u w=0u l=0u
X13 a_4151_989.t1 a_147_187.t10 VDD.t35 ��O� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X14 QN a_4151_989.t7 a_3924_210.t0 GND sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=0p ps=0u w=0u l=0u
X15 a_277_1050.t0 a_147_187.t11 VDD.t5  �O� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X16 VDD.t3 a_277_1050.t8 a_599_989.t0 ��O� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X17 VDD.t61 RN.t3 a_599_989.t6  �O� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X18 VDD.t51 a_4151_989.t6 QN.t4 ��O� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X19 GND a_277_1050.t11 a_3643_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X20 a_277_1050.t5 CLK.t2 VDD.t25  �O� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X21 a_2141_1050.t2 a_599_989.t10 VDD.t15 ��O� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X22 QN.t1 a_277_1050.t9 VDD.t7  �O� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X23 GND QN.t8 a_4626_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X24 VDD.t57 RN.t4 QN.t6 ��O� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X25 GND a_599_989.t12 a_2036_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X26 VDD.t41 D.t2 a_599_989.t2  �O� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X27 GND a_2141_1050.t7 a_2681_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X28 a_599_989.t4 a_277_1050.t10 VDD.t45 ��O� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X29 a_277_1050.t2 a_599_989.t11 VDD.t23  �O� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X30 a_2141_1050.t1 a_147_187.t13 VDD.t31 ��O� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X31 QN.t5 RN.t5 VDD.t55  �O� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X32 a_147_187.t0 a_2141_1050.t6 VDD.t21 ��O� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X33 VDD.t1 CLK.t4 a_147_187.t2  �O� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X34 VDD.t11 QN.t9 a_4151_989.t3 ��O� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X35 GND a_277_1050.t12 a_1053_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X36 VDD.t63 RN.t8 a_147_187.t6  �O� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X37 VDD.t33 a_147_187.t14 a_4151_989.t0 ��O� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X38 VDD.t17 a_147_187.t15 a_277_1050.t1  �O� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
C0 QN VDD 2.82fF
C1 RN VDD 0.89fF
C2 QN RN 0.12fF
C3 D VDD 0.29fF
C4 D RN 0.18fF
C5 CLK VDD 1.98fF
C6 CLK RN 0.28fF
C7 CLK D 0.07fF
R0 D.n0 D.t2 479.223
R1 D.n0 D.t0 375.52
R2 D.n1 D.t1 287.572
R3 D.n1 D.n0 196.47
R4 D.n2 D.n1 4.65
R5 D.n2 D 0.046
R6 VDD.n307 VDD.n296 144.705
R7 VDD.n430 VDD.n428 144.705
R8 VDD.n382 VDD.n375 144.705
R9 VDD.n154 VDD.n147 144.705
R10 VDD.n79 VDD.n68 144.705
R11 VDD.n273 VDD.t9 143.754
R12 VDD.n349 VDD.t61 143.754
R13 VDD.n163 VDD.t63 143.754
R14 VDD.n88 VDD.t51 143.754
R15 VDD.n407 VDD.t49 143.754
R16 VDD.n24 VDD.t33 143.754
R17 VDD.n238 VDD.t5 135.17
R18 VDD.n314 VDD.t45 135.17
R19 VDD.n385 VDD.t15 135.17
R20 VDD.n193 VDD.t21 135.17
R21 VDD.n118 VDD.t7 135.17
R22 VDD.n46 VDD.t29 135.17
R23 VDD.n248 VDD.n247 129.472
R24 VDD.n264 VDD.n263 129.472
R25 VDD.n324 VDD.n323 129.472
R26 VDD.n340 VDD.n339 129.472
R27 VDD.n399 VDD.n398 129.472
R28 VDD.n184 VDD.n183 129.472
R29 VDD.n172 VDD.n171 129.472
R30 VDD.n109 VDD.n108 129.472
R31 VDD.n97 VDD.n96 129.472
R32 VDD.n34 VDD.n33 129.472
R33 VDD.n64 VDD.n63 92.5
R34 VDD.n62 VDD.n61 92.5
R35 VDD.n60 VDD.n59 92.5
R36 VDD.n58 VDD.n57 92.5
R37 VDD.n66 VDD.n65 92.5
R38 VDD.n143 VDD.n142 92.5
R39 VDD.n141 VDD.n140 92.5
R40 VDD.n139 VDD.n138 92.5
R41 VDD.n137 VDD.n136 92.5
R42 VDD.n145 VDD.n144 92.5
R43 VDD.n424 VDD.n423 92.5
R44 VDD.n422 VDD.n421 92.5
R45 VDD.n420 VDD.n419 92.5
R46 VDD.n418 VDD.n417 92.5
R47 VDD.n426 VDD.n425 92.5
R48 VDD.n371 VDD.n370 92.5
R49 VDD.n369 VDD.n368 92.5
R50 VDD.n367 VDD.n366 92.5
R51 VDD.n365 VDD.n364 92.5
R52 VDD.n373 VDD.n372 92.5
R53 VDD.n292 VDD.n291 92.5
R54 VDD.n290 VDD.n289 92.5
R55 VDD.n288 VDD.n287 92.5
R56 VDD.n286 VDD.n285 92.5
R57 VDD.n294 VDD.n293 92.5
R58 VDD.n222 VDD.n221 92.5
R59 VDD.n220 VDD.n219 92.5
R60 VDD.n218 VDD.n217 92.5
R61 VDD.n216 VDD.n215 92.5
R62 VDD.n224 VDD.n223 92.5
R63 VDD.n14 VDD.n1 92.5
R64 VDD.n5 VDD.n4 92.5
R65 VDD.n7 VDD.n6 92.5
R66 VDD.n9 VDD.n8 92.5
R67 VDD.n11 VDD.n10 92.5
R68 VDD.n13 VDD.n12 92.5
R69 VDD.n21 VDD.n20 92.059
R70 VDD.n78 VDD.n77 92.059
R71 VDD.n153 VDD.n152 92.059
R72 VDD.n207 VDD.n206 92.059
R73 VDD.n381 VDD.n380 92.059
R74 VDD.n306 VDD.n305 92.059
R75 VDD.n230 VDD.n229 92.059
R76 VDD.n20 VDD.n16 67.194
R77 VDD.n20 VDD.n17 67.194
R78 VDD.n20 VDD.n18 67.194
R79 VDD.n20 VDD.n19 67.194
R80 VDD.n214 VDD.n213 44.141
R81 VDD.n363 VDD.n362 44.141
R82 VDD.n416 VDD.n415 44.141
R83 VDD.n135 VDD.n134 44.141
R84 VDD.n5 VDD.n3 44.141
R85 VDD.n362 VDD.n360 44.107
R86 VDD.n415 VDD.n413 44.107
R87 VDD.n134 VDD.n132 44.107
R88 VDD.n213 VDD.n211 44.107
R89 VDD.n3 VDD.n2 44.107
R90 VDD.n20 VDD.n15 41.052
R91 VDD.n72 VDD.n70 39.742
R92 VDD.n72 VDD.n71 39.742
R93 VDD.n74 VDD.n73 39.742
R94 VDD.n149 VDD.n148 39.742
R95 VDD.n203 VDD.n202 39.742
R96 VDD.n377 VDD.n376 39.742
R97 VDD.n226 VDD.n225 39.742
R98 VDD.n304 VDD.n301 39.742
R99 VDD.n304 VDD.n303 39.742
R100 VDD.n300 VDD.n299 39.742
R101 VDD.n134 VDD.n133 38
R102 VDD.n415 VDD.n414 38
R103 VDD.n362 VDD.n361 38
R104 VDD.n213 VDD.n212 38
R105 VDD.n360 VDD.n359 36.774
R106 VDD.n413 VDD.n412 36.774
R107 VDD.n132 VDD.n131 36.774
R108 VDD.n70 VDD.n69 36.774
R109 VDD.n303 VDD.n302 36.774
R110 VDD.n90 ��O� 35.8
R111 VDD.n165  �O� 35.8
R112 VDD.n343  �O� 35.8
R113 VDD.n267 ��O� 35.8
R114 VDD.n114  �O� 33.243
R115 VDD.n189 ��O� 33.243
R116 VDD.n319 ��O� 33.243
R117 VDD.n243  �O� 33.243
R118 VDD.n1 VDD.n0 30.923
R119 VDD.n77 VDD.n75 26.38
R120 VDD.n77 VDD.n74 26.38
R121 VDD.n77 VDD.n72 26.38
R122 VDD.n77 VDD.n76 26.38
R123 VDD.n152 VDD.n150 26.38
R124 VDD.n152 VDD.n149 26.38
R125 VDD.n152 VDD.n151 26.38
R126 VDD.n206 VDD.n204 26.38
R127 VDD.n206 VDD.n203 26.38
R128 VDD.n206 VDD.n205 26.38
R129 VDD.n380 VDD.n378 26.38
R130 VDD.n380 VDD.n377 26.38
R131 VDD.n380 VDD.n379 26.38
R132 VDD.n229 VDD.n227 26.38
R133 VDD.n229 VDD.n226 26.38
R134 VDD.n229 VDD.n228 26.38
R135 VDD.n305 VDD.n304 26.38
R136 VDD.n305 VDD.n300 26.38
R137 VDD.n305 VDD.n298 26.38
R138 VDD.n305 VDD.n297 26.38
R139 VDD.n232 VDD.n224 22.915
R140 VDD.n23 VDD.n14 22.915
R141 VDD.n29 ��O� 20.457
R142 VDD.n403  �O� 20.457
R143 VDD.n42  �O� 17.9
R144 VDD.n390 ��O� 17.9
R145 VDD.n94 ��O� 15.343
R146 VDD.n169  �O� 15.343
R147 VDD.n337 ��O� 15.343
R148 VDD.n261  �O� 15.343
R149 VDD.n224 VDD.n222 14.864
R150 VDD.n222 VDD.n220 14.864
R151 VDD.n220 VDD.n218 14.864
R152 VDD.n218 VDD.n216 14.864
R153 VDD.n216 VDD.n214 14.864
R154 VDD.n373 VDD.n371 14.864
R155 VDD.n371 VDD.n369 14.864
R156 VDD.n369 VDD.n367 14.864
R157 VDD.n367 VDD.n365 14.864
R158 VDD.n365 VDD.n363 14.864
R159 VDD.n426 VDD.n424 14.864
R160 VDD.n424 VDD.n422 14.864
R161 VDD.n422 VDD.n420 14.864
R162 VDD.n420 VDD.n418 14.864
R163 VDD.n418 VDD.n416 14.864
R164 VDD.n145 VDD.n143 14.864
R165 VDD.n143 VDD.n141 14.864
R166 VDD.n141 VDD.n139 14.864
R167 VDD.n139 VDD.n137 14.864
R168 VDD.n137 VDD.n135 14.864
R169 VDD.n66 VDD.n64 14.864
R170 VDD.n64 VDD.n62 14.864
R171 VDD.n62 VDD.n60 14.864
R172 VDD.n60 VDD.n58 14.864
R173 VDD.n58 VDD.n56 14.864
R174 VDD.n56 VDD.n55 14.864
R175 VDD.n294 VDD.n292 14.864
R176 VDD.n292 VDD.n290 14.864
R177 VDD.n290 VDD.n288 14.864
R178 VDD.n288 VDD.n286 14.864
R179 VDD.n286 VDD.n284 14.864
R180 VDD.n284 VDD.n283 14.864
R181 VDD.n14 VDD.n13 14.864
R182 VDD.n13 VDD.n11 14.864
R183 VDD.n11 VDD.n9 14.864
R184 VDD.n9 VDD.n7 14.864
R185 VDD.n7 VDD.n5 14.864
R186 VDD.n80 VDD.n67 14.864
R187 VDD.n155 VDD.n146 14.864
R188 VDD.n431 VDD.n427 14.864
R189 VDD.n383 VDD.n374 14.864
R190 VDD.n308 VDD.n295 14.864
R191 VDD.n247 VDD.t25 14.282
R192 VDD.n247 VDD.t17 14.282
R193 VDD.n263 VDD.t23 14.282
R194 VDD.n263 VDD.t37 14.282
R195 VDD.n323 VDD.t43 14.282
R196 VDD.n323 VDD.t3 14.282
R197 VDD.n339 VDD.t39 14.282
R198 VDD.n339 VDD.t41 14.282
R199 VDD.n398 VDD.t31 14.282
R200 VDD.n398 VDD.t13 14.282
R201 VDD.n183 VDD.t19 14.282
R202 VDD.n183 VDD.t53 14.282
R203 VDD.n171 VDD.t59 14.282
R204 VDD.n171 VDD.t1 14.282
R205 VDD.n108 VDD.t55 14.282
R206 VDD.n108 VDD.t47 14.282
R207 VDD.n96 VDD.t27 14.282
R208 VDD.n96 VDD.t57 14.282
R209 VDD.n33 VDD.t35 14.282
R210 VDD.n33 VDD.t11 14.282
R211 VDD.n110  �O� 12.786
R212 VDD.n185 ��O� 12.786
R213 VDD.n325 ��O� 12.786
R214 VDD.n249  �O� 12.786
R215 VDD.n36 VDD.n34 9.083
R216 VDD.n401 VDD.n399 9.083
R217 VDD.n23 VDD.n22 8.855
R218 VDD.n22 VDD.n21 8.855
R219 VDD.n27 VDD.n26 8.855
R220 VDD.n26 VDD.n25 8.855
R221 VDD.n31 VDD.n30 8.855
R222 VDD.n30 VDD.n29 8.855
R223 VDD.n36 VDD.n35 8.855
R224 VDD.n35 ��O� 8.855
R225 VDD.n40 VDD.n39 8.855
R226 VDD.n39 VDD.n38 8.855
R227 VDD.n44 VDD.n43 8.855
R228 VDD.n43 VDD.n42 8.855
R229 VDD.n49 VDD.n48 8.855
R230 VDD.n48 VDD.n47 8.855
R231 VDD.n53 VDD.n52 8.855
R232 VDD.n52 VDD.n51 8.855
R233 VDD.n80 VDD.n79 8.855
R234 VDD.n79 VDD.n78 8.855
R235 VDD.n84 VDD.n83 8.855
R236 VDD.n83 VDD.n82 8.855
R237 VDD.n88 VDD.n87 8.855
R238 VDD.n87 VDD.n86 8.855
R239 VDD.n92 VDD.n91 8.855
R240 VDD.n91 VDD.n90 8.855
R241 VDD.n98 VDD.n95 8.855
R242 VDD.n95 VDD.n94 8.855
R243 VDD.n102 VDD.n101 8.855
R244 VDD.n101 VDD.n100 8.855
R245 VDD.n106 VDD.n105 8.855
R246 VDD.n105 VDD.n104 8.855
R247 VDD.n112 VDD.n111 8.855
R248 VDD.n111 VDD.n110 8.855
R249 VDD.n116 VDD.n115 8.855
R250 VDD.n115 VDD.n114 8.855
R251 VDD.n121 VDD.n120 8.855
R252 VDD.n120 VDD.n119 8.855
R253 VDD.n125 VDD.n124 8.855
R254 VDD.n124 VDD.n123 8.855
R255 VDD.n129 VDD.n128 8.855
R256 VDD.n128 VDD.n127 8.855
R257 VDD.n155 VDD.n154 8.855
R258 VDD.n154 VDD.n153 8.855
R259 VDD.n159 VDD.n158 8.855
R260 VDD.n158 VDD.n157 8.855
R261 VDD.n163 VDD.n162 8.855
R262 VDD.n162 VDD.n161 8.855
R263 VDD.n167 VDD.n166 8.855
R264 VDD.n166 VDD.n165 8.855
R265 VDD.n173 VDD.n170 8.855
R266 VDD.n170 VDD.n169 8.855
R267 VDD.n177 VDD.n176 8.855
R268 VDD.n176 VDD.n175 8.855
R269 VDD.n181 VDD.n180 8.855
R270 VDD.n180 VDD.n179 8.855
R271 VDD.n187 VDD.n186 8.855
R272 VDD.n186 VDD.n185 8.855
R273 VDD.n191 VDD.n190 8.855
R274 VDD.n190 VDD.n189 8.855
R275 VDD.n196 VDD.n195 8.855
R276 VDD.n195 VDD.n194 8.855
R277 VDD.n200 VDD.n199 8.855
R278 VDD.n199 VDD.n198 8.855
R279 VDD.n209 VDD.n208 8.855
R280 VDD.n208 VDD.n207 8.855
R281 VDD.n431 VDD.n430 8.855
R282 VDD.n430 VDD.n429 8.855
R283 VDD.n410 VDD.n409 8.855
R284 VDD.n409 VDD.n408 8.855
R285 VDD.n405 VDD.n404 8.855
R286 VDD.n404 VDD.n403 8.855
R287 VDD.n401 VDD.n400 8.855
R288 VDD.n400 ��O� 8.855
R289 VDD.n396 VDD.n395 8.855
R290 VDD.n395 VDD.n394 8.855
R291 VDD.n392 VDD.n391 8.855
R292 VDD.n391 VDD.n390 8.855
R293 VDD.n388 VDD.n387 8.855
R294 VDD.n387 VDD.n386 8.855
R295 VDD.n383 VDD.n382 8.855
R296 VDD.n382 VDD.n381 8.855
R297 VDD.n357 VDD.n356 8.855
R298 VDD.n356 VDD.n355 8.855
R299 VDD.n353 VDD.n352 8.855
R300 VDD.n352 VDD.n351 8.855
R301 VDD.n349 VDD.n348 8.855
R302 VDD.n348 VDD.n347 8.855
R303 VDD.n345 VDD.n344 8.855
R304 VDD.n344 VDD.n343 8.855
R305 VDD.n341 VDD.n338 8.855
R306 VDD.n338 VDD.n337 8.855
R307 VDD.n335 VDD.n334 8.855
R308 VDD.n334 VDD.n333 8.855
R309 VDD.n331 VDD.n330 8.855
R310 VDD.n330 VDD.n329 8.855
R311 VDD.n327 VDD.n326 8.855
R312 VDD.n326 VDD.n325 8.855
R313 VDD.n321 VDD.n320 8.855
R314 VDD.n320 VDD.n319 8.855
R315 VDD.n317 VDD.n316 8.855
R316 VDD.n316 VDD.n315 8.855
R317 VDD.n312 VDD.n311 8.855
R318 VDD.n311 VDD.n310 8.855
R319 VDD.n308 VDD.n307 8.855
R320 VDD.n307 VDD.n306 8.855
R321 VDD.n281 VDD.n280 8.855
R322 VDD.n280 VDD.n279 8.855
R323 VDD.n277 VDD.n276 8.855
R324 VDD.n276 VDD.n275 8.855
R325 VDD.n273 VDD.n272 8.855
R326 VDD.n272 VDD.n271 8.855
R327 VDD.n269 VDD.n268 8.855
R328 VDD.n268 VDD.n267 8.855
R329 VDD.n265 VDD.n262 8.855
R330 VDD.n262 VDD.n261 8.855
R331 VDD.n259 VDD.n258 8.855
R332 VDD.n258 VDD.n257 8.855
R333 VDD.n255 VDD.n254 8.855
R334 VDD.n254 VDD.n253 8.855
R335 VDD.n251 VDD.n250 8.855
R336 VDD.n250 VDD.n249 8.855
R337 VDD.n245 VDD.n244 8.855
R338 VDD.n244 VDD.n243 8.855
R339 VDD.n241 VDD.n240 8.855
R340 VDD.n240 VDD.n239 8.855
R341 VDD.n236 VDD.n235 8.855
R342 VDD.n235 VDD.n234 8.855
R343 VDD.n232 VDD.n231 8.855
R344 VDD.n231 VDD.n230 8.855
R345 VDD.n374 VDD.n373 8.051
R346 VDD.n427 VDD.n426 8.051
R347 VDD.n146 VDD.n145 8.051
R348 VDD.n67 VDD.n66 8.051
R349 VDD.n295 VDD.n294 8.051
R350 VDD.n104  �O� 7.671
R351 VDD.n179  �O� 7.671
R352 VDD.n329 0��&�U 7.671
R353 VDD.n253  �O� 7.671
R354 VDD.n112 VDD.n109 7.019
R355 VDD.n187 VDD.n184 7.019
R356 VDD.n327 VDD.n324 7.019
R357 VDD.n251 VDD.n248 7.019
R358 VDD.n98 VDD.n97 6.606
R359 VDD.n173 VDD.n172 6.606
R360 VDD.n341 VDD.n340 6.606
R361 VDD.n265 VDD.n264 6.606
R362 VDD.n100 ��O� 5.114
R363 VDD.n175  �O� 5.114
R364 VDD.n333  �O� 5.114
R365 VDD.n257 ���&�U 5.114
R366 VDD.n32 VDD.n31 4.65
R367 VDD.n37 VDD.n36 4.65
R368 VDD.n41 VDD.n40 4.65
R369 VDD.n45 VDD.n44 4.65
R370 VDD.n50 VDD.n49 4.65
R371 VDD.n54 VDD.n53 4.65
R372 VDD.n81 VDD.n80 4.65
R373 VDD.n85 VDD.n84 4.65
R374 VDD.n89 VDD.n88 4.65
R375 VDD.n93 VDD.n92 4.65
R376 VDD.n99 VDD.n98 4.65
R377 VDD.n103 VDD.n102 4.65
R378 VDD.n107 VDD.n106 4.65
R379 VDD.n113 VDD.n112 4.65
R380 VDD.n117 VDD.n116 4.65
R381 VDD.n122 VDD.n121 4.65
R382 VDD.n126 VDD.n125 4.65
R383 VDD.n130 VDD.n129 4.65
R384 VDD.n156 VDD.n155 4.65
R385 VDD.n160 VDD.n159 4.65
R386 VDD.n164 VDD.n163 4.65
R387 VDD.n168 VDD.n167 4.65
R388 VDD.n174 VDD.n173 4.65
R389 VDD.n178 VDD.n177 4.65
R390 VDD.n182 VDD.n181 4.65
R391 VDD.n188 VDD.n187 4.65
R392 VDD.n192 VDD.n191 4.65
R393 VDD.n197 VDD.n196 4.65
R394 VDD.n201 VDD.n200 4.65
R395 VDD.n210 VDD.n209 4.65
R396 VDD.n432 VDD.n431 4.65
R397 VDD.n411 VDD.n410 4.65
R398 VDD.n406 VDD.n405 4.65
R399 VDD.n402 VDD.n401 4.65
R400 VDD.n397 VDD.n396 4.65
R401 VDD.n393 VDD.n392 4.65
R402 VDD.n389 VDD.n388 4.65
R403 VDD.n384 VDD.n383 4.65
R404 VDD.n358 VDD.n357 4.65
R405 VDD.n354 VDD.n353 4.65
R406 VDD.n350 VDD.n349 4.65
R407 VDD.n346 VDD.n345 4.65
R408 VDD.n342 VDD.n341 4.65
R409 VDD.n336 VDD.n335 4.65
R410 VDD.n332 VDD.n331 4.65
R411 VDD.n328 VDD.n327 4.65
R412 VDD.n322 VDD.n321 4.65
R413 VDD.n318 VDD.n317 4.65
R414 VDD.n313 VDD.n312 4.65
R415 VDD.n309 VDD.n308 4.65
R416 VDD.n282 VDD.n281 4.65
R417 VDD.n278 VDD.n277 4.65
R418 VDD.n274 VDD.n273 4.65
R419 VDD.n270 VDD.n269 4.65
R420 VDD.n266 VDD.n265 4.65
R421 VDD.n260 VDD.n259 4.65
R422 VDD.n256 VDD.n255 4.65
R423 VDD.n252 VDD.n251 4.65
R424 VDD.n246 VDD.n245 4.65
R425 VDD.n242 VDD.n241 4.65
R426 VDD.n237 VDD.n236 4.65
R427 VDD.n233 VDD.n232 4.65
R428 VDD.n28 VDD.n23 2.933
R429 VDD.n49 VDD.n46 2.89
R430 VDD.n388 VDD.n385 2.89
R431 VDD.n28 VDD.n27 2.844
R432 VDD.n38 ��O� 2.557
R433 VDD.n394 VDD.t12 2.557
R434 VDD.n27 VDD.n24 2.477
R435 VDD.n410 VDD.n407 2.477
R436 VDD.n32 VDD.n28 1.063
R437 VDD.n121 VDD.n118 0.412
R438 VDD.n196 VDD.n193 0.412
R439 VDD.n317 VDD.n314 0.412
R440 VDD.n241 VDD.n238 0.412
R441 VDD.n81 VDD.n54 0.29
R442 VDD.n156 VDD.n130 0.29
R443 VDD.n384 VDD.n358 0.29
R444 VDD.n309 VDD.n282 0.29
R445 VDD.n233 VDD 0.207
R446 VDD.n107 VDD.n103 0.197
R447 VDD.n182 VDD.n178 0.197
R448 VDD.n336 VDD.n332 0.197
R449 VDD.n260 VDD.n256 0.197
R450 VDD.n41 VDD.n37 0.181
R451 VDD.n402 VDD.n397 0.181
R452 VDD.n37 VDD.n32 0.145
R453 VDD.n45 VDD.n41 0.145
R454 VDD.n50 VDD.n45 0.145
R455 VDD.n54 VDD.n50 0.145
R456 VDD.n85 VDD.n81 0.145
R457 VDD.n89 VDD.n85 0.145
R458 VDD.n93 VDD.n89 0.145
R459 VDD.n99 VDD.n93 0.145
R460 VDD.n103 VDD.n99 0.145
R461 VDD.n113 VDD.n107 0.145
R462 VDD.n117 VDD.n113 0.145
R463 VDD.n122 VDD.n117 0.145
R464 VDD.n126 VDD.n122 0.145
R465 VDD.n130 VDD.n126 0.145
R466 VDD.n160 VDD.n156 0.145
R467 VDD.n164 VDD.n160 0.145
R468 VDD.n168 VDD.n164 0.145
R469 VDD.n174 VDD.n168 0.145
R470 VDD.n178 VDD.n174 0.145
R471 VDD.n188 VDD.n182 0.145
R472 VDD.n192 VDD.n188 0.145
R473 VDD.n197 VDD.n192 0.145
R474 VDD.n201 VDD.n197 0.145
R475 VDD.n210 VDD.n201 0.145
R476 VDD VDD.n210 0.145
R477 VDD VDD.n432 0.145
R478 VDD.n432 VDD.n411 0.145
R479 VDD.n411 VDD.n406 0.145
R480 VDD.n406 VDD.n402 0.145
R481 VDD.n397 VDD.n393 0.145
R482 VDD.n393 VDD.n389 0.145
R483 VDD.n389 VDD.n384 0.145
R484 VDD.n358 VDD.n354 0.145
R485 VDD.n354 VDD.n350 0.145
R486 VDD.n350 VDD.n346 0.145
R487 VDD.n346 VDD.n342 0.145
R488 VDD.n342 VDD.n336 0.145
R489 VDD.n332 VDD.n328 0.145
R490 VDD.n328 VDD.n322 0.145
R491 VDD.n322 VDD.n318 0.145
R492 VDD.n318 VDD.n313 0.145
R493 VDD.n313 VDD.n309 0.145
R494 VDD.n282 VDD.n278 0.145
R495 VDD.n278 VDD.n274 0.145
R496 VDD.n274 VDD.n270 0.145
R497 VDD.n270 VDD.n266 0.145
R498 VDD.n266 VDD.n260 0.145
R499 VDD.n256 VDD.n252 0.145
R500 VDD.n252 VDD.n246 0.145
R501 VDD.n246 VDD.n242 0.145
R502 VDD.n242 VDD.n237 0.145
R503 VDD.n237 VDD.n233 0.145
R504 a_599_989.n1 a_599_989.t7 480.392
R505 a_599_989.n3 a_599_989.t11 454.685
R506 a_599_989.n3 a_599_989.t8 428.979
R507 a_599_989.n1 a_599_989.t10 403.272
R508 a_599_989.n2 a_599_989.t12 357.204
R509 a_599_989.n4 a_599_989.t9 311.683
R510 a_599_989.n10 a_599_989.n9 308.216
R511 a_599_989.n11 a_599_989.n10 179.199
R512 a_599_989.n4 a_599_989.n3 171.288
R513 a_599_989.n2 a_599_989.n1 171.288
R514 a_599_989.n13 a_599_989.n12 161.352
R515 a_599_989.n11 a_599_989.n0 95.095
R516 a_599_989.n14 a_599_989.n13 95.094
R517 a_599_989.n13 a_599_989.n11 66.258
R518 a_599_989.n9 a_599_989.n8 30
R519 a_599_989.n7 a_599_989.n6 24.383
R520 a_599_989.n9 a_599_989.n7 23.684
R521 a_599_989.n0 a_599_989.t6 14.282
R522 a_599_989.n0 a_599_989.t1 14.282
R523 a_599_989.n12 a_599_989.t0 14.282
R524 a_599_989.n12 a_599_989.t4 14.282
R525 a_599_989.n14 a_599_989.t2 14.282
R526 a_599_989.t3 a_599_989.n14 14.282
R527 a_599_989.n5 a_599_989.n4 8.685
R528 a_599_989.n5 a_599_989.n2 5.965
R529 a_599_989.n10 a_599_989.n5 4.65
R530 CLK.n2 CLK.t0 459.505
R531 CLK.n0 CLK.t4 459.505
R532 CLK.n3 CLK.t3 399.181
R533 CLK.n1 CLK.t5 399.181
R534 CLK.n2 CLK.t2 384.527
R535 CLK.n0 CLK.t1 384.527
R536 CLK.n3 CLK.n2 33.832
R537 CLK.n1 CLK.n0 33.832
R538 CLK.n4 CLK.n1 11.555
R539 CLK.n4 CLK.n3 2.079
R540 CLK.n4 CLK 0.046
R541 a_277_1050.n2 a_277_1050.t8 512.525
R542 a_277_1050.n0 a_277_1050.t7 512.525
R543 a_277_1050.n3 a_277_1050.t12 389.251
R544 a_277_1050.n1 a_277_1050.t11 389.251
R545 a_277_1050.n2 a_277_1050.t10 371.139
R546 a_277_1050.n0 a_277_1050.t9 371.139
R547 a_277_1050.n9 a_277_1050.n8 336.075
R548 a_277_1050.n3 a_277_1050.n2 207.695
R549 a_277_1050.n1 a_277_1050.n0 207.695
R550 a_277_1050.n12 a_277_1050.n11 161.352
R551 a_277_1050.n13 a_277_1050.n9 151.34
R552 a_277_1050.n12 a_277_1050.n10 95.095
R553 a_277_1050.n14 a_277_1050.n13 95.094
R554 a_277_1050.n13 a_277_1050.n12 66.258
R555 a_277_1050.n8 a_277_1050.n7 30
R556 a_277_1050.n6 a_277_1050.n5 24.383
R557 a_277_1050.n8 a_277_1050.n6 23.684
R558 a_277_1050.n10 a_277_1050.t6 14.282
R559 a_277_1050.n10 a_277_1050.t5 14.282
R560 a_277_1050.n11 a_277_1050.t1 14.282
R561 a_277_1050.n11 a_277_1050.t0 14.282
R562 a_277_1050.t3 a_277_1050.n14 14.282
R563 a_277_1050.n14 a_277_1050.t2 14.282
R564 a_277_1050.n4 a_277_1050.n1 14.126
R565 a_277_1050.n9 a_277_1050.n4 5.965
R566 a_277_1050.n4 a_277_1050.n3 4.65
R567 a_2141_1050.n1 a_2141_1050.t5 512.525
R568 a_2141_1050.n1 a_2141_1050.t6 371.139
R569 a_2141_1050.n2 a_2141_1050.t7 361.392
R570 a_2141_1050.n4 a_2141_1050.n3 327.32
R571 a_2141_1050.n2 a_2141_1050.n1 235.554
R572 a_2141_1050.n5 a_2141_1050.n4 159.999
R573 a_2141_1050.n6 a_2141_1050.n5 157.963
R574 a_2141_1050.n5 a_2141_1050.n0 91.706
R575 a_2141_1050.n0 a_2141_1050.t4 14.282
R576 a_2141_1050.n0 a_2141_1050.t1 14.282
R577 a_2141_1050.t3 a_2141_1050.n6 14.282
R578 a_2141_1050.n6 a_2141_1050.t2 14.282
R579 a_2141_1050.n4 a_2141_1050.n2 10.615
R580 QN.n0 QN.t9 480.392
R581 QN.n0 QN.t7 403.272
R582 QN.n1 QN.t8 357.204
R583 QN.n8 QN.n7 329.955
R584 QN.n8 QN.n6 179.199
R585 QN.n1 QN.n0 171.288
R586 QN.n5 QN.n4 161.352
R587 QN.n6 QN.n2 95.095
R588 QN.n5 QN.n3 95.095
R589 QN.n6 QN.n5 66.258
R590 QN.n2 QN.t4 14.282
R591 QN.n2 QN.t0 14.282
R592 QN.n3 QN.t6 14.282
R593 QN.n3 QN.t5 14.282
R594 QN.n4 QN.t2 14.282
R595 QN.n4 QN.t1 14.282
R596 QN.n9 QN.n1 5.965
R597 QN.n9 QN.n8 4.65
R598 QN.n9 QN 0.046
R599 a_1053_103.t0 a_1053_103.n3 117.777
R600 a_1053_103.n6 a_1053_103.n4 55.785
R601 a_1053_103.n6 a_1053_103.n5 51.696
R602 a_1053_103.t0 a_1053_103.n6 39.361
R603 a_1053_103.n2 a_1053_103.n0 32.662
R604 a_1053_103.t0 a_1053_103.n2 3.034
R605 a_1053_103.n2 a_1053_103.n1 0.443
R606 a_1334_210.n10 a_1334_210.n8 171.558
R607 a_1334_210.n8 a_1334_210.t1 75.764
R608 a_1334_210.n11 a_1334_210.n0 49.6
R609 a_1334_210.n3 a_1334_210.n2 27.476
R610 a_1334_210.n10 a_1334_210.n9 27.2
R611 a_1334_210.n11 a_1334_210.n10 22.4
R612 a_1334_210.t1 a_1334_210.n5 20.241
R613 a_1334_210.n7 a_1334_210.n6 19.952
R614 a_1334_210.t1 a_1334_210.n3 13.984
R615 a_1334_210.n5 a_1334_210.n4 13.494
R616 a_1334_210.t1 a_1334_210.n1 7.04
R617 a_1334_210.n8 a_1334_210.n7 1.505
R618 GND.n156 GND.n155 237.558
R619 GND.n231 GND.n230 237.558
R620 GND.n198 GND.n197 237.558
R621 GND.n76 GND.n75 237.558
R622 GND.n31 GND.n30 237.558
R623 GND.n28 GND.n27 210.82
R624 GND.n158 GND.n157 210.82
R625 GND.n200 GND.n199 210.82
R626 GND.n228 GND.n227 210.82
R627 GND.n73 GND.n72 210.82
R628 GND.n167 GND.n166 173.365
R629 GND.n125 GND.n124 173.365
R630 GND.n63 GND.n62 152.358
R631 GND.n108 GND.n107 152.358
R632 GND.n17 GND.n16 151.605
R633 GND.n211 GND.n210 151.605
R634 GND.n16 GND.n15 28.421
R635 GND.n62 GND.n61 28.421
R636 GND.n107 GND.n106 28.421
R637 GND.n210 GND.n209 28.421
R638 GND.n16 GND.n14 25.263
R639 GND.n62 GND.n60 25.263
R640 GND.n107 GND.n105 25.263
R641 GND.n210 GND.n208 25.263
R642 GND.n14 GND.n13 24.383
R643 GND.n60 GND.n59 24.383
R644 GND.n105 GND.n104 24.383
R645 GND.n208 GND.n207 24.383
R646 GND.n29 GND.n28 18.953
R647 GND.n159 GND.n158 18.953
R648 GND.n201 GND.n200 18.953
R649 GND.n229 GND.n228 18.953
R650 GND.n74 GND.n73 18.953
R651 GND.n32 GND.n29 14.864
R652 GND.n77 GND.n74 14.864
R653 GND.n232 GND.n229 14.864
R654 GND.n202 GND.n201 14.864
R655 GND.n160 GND.n159 14.864
R656 GND.n121 GND.n120 9.154
R657 GND.n126 GND.n123 9.154
R658 GND.n129 GND.n128 9.154
R659 GND.n132 GND.n131 9.154
R660 GND.n135 GND.n134 9.154
R661 GND.n138 GND.n137 9.154
R662 GND.n141 GND.n140 9.154
R663 GND.n144 GND.n143 9.154
R664 GND.n147 GND.n146 9.154
R665 GND.n150 GND.n149 9.154
R666 GND.n153 GND.n152 9.154
R667 GND.n160 GND.n156 9.154
R668 GND.n163 GND.n162 9.154
R669 GND.n168 GND.n165 9.154
R670 GND.n171 GND.n170 9.154
R671 GND.n174 GND.n173 9.154
R672 GND.n177 GND.n176 9.154
R673 GND.n180 GND.n179 9.154
R674 GND.n183 GND.n182 9.154
R675 GND.n186 GND.n185 9.154
R676 GND.n189 GND.n188 9.154
R677 GND.n192 GND.n191 9.154
R678 GND.n195 GND.n194 9.154
R679 GND.n202 GND.n198 9.154
R680 GND.n205 GND.n204 9.154
R681 GND.n213 GND.n212 9.154
R682 GND.n216 GND.n215 9.154
R683 GND.n219 GND.n218 9.154
R684 GND.n222 GND.n221 9.154
R685 GND.n225 GND.n224 9.154
R686 GND.n232 GND.n231 9.154
R687 GND.n115 GND.n114 9.154
R688 GND.n112 GND.n111 9.154
R689 GND.n109 GND.n103 9.154
R690 GND.n101 GND.n100 9.154
R691 GND.n98 GND.n97 9.154
R692 GND.n95 GND.n94 9.154
R693 GND.n92 GND.n91 9.154
R694 GND.n89 GND.n88 9.154
R695 GND.n86 GND.n85 9.154
R696 GND.n83 GND.n82 9.154
R697 GND.n80 GND.n79 9.154
R698 GND.n77 GND.n76 9.154
R699 GND.n70 GND.n69 9.154
R700 GND.n67 GND.n66 9.154
R701 GND.n64 GND.n58 9.154
R702 GND.n56 GND.n55 9.154
R703 GND.n53 GND.n52 9.154
R704 GND.n50 GND.n49 9.154
R705 GND.n47 GND.n46 9.154
R706 GND.n44 GND.n43 9.154
R707 GND.n41 GND.n40 9.154
R708 GND.n38 GND.n37 9.154
R709 GND.n35 GND.n34 9.154
R710 GND.n32 GND.n31 9.154
R711 GND.n25 GND.n24 9.154
R712 GND.n22 GND.n21 9.154
R713 GND.n19 GND.n18 9.154
R714 GND.n11 GND.n10 9.154
R715 GND.n8 GND.n7 9.154
R716 GND.n5 GND.n4 9.154
R717 GND.n2 GND.n1 9.154
R718 GND.n119 GND.n118 4.65
R719 GND.n6 GND.n5 4.65
R720 GND.n9 GND.n8 4.65
R721 GND.n12 GND.n11 4.65
R722 GND.n20 GND.n19 4.65
R723 GND.n23 GND.n22 4.65
R724 GND.n26 GND.n25 4.65
R725 GND.n33 GND.n32 4.65
R726 GND.n36 GND.n35 4.65
R727 GND.n39 GND.n38 4.65
R728 GND.n42 GND.n41 4.65
R729 GND.n45 GND.n44 4.65
R730 GND.n48 GND.n47 4.65
R731 GND.n51 GND.n50 4.65
R732 GND.n54 GND.n53 4.65
R733 GND.n57 GND.n56 4.65
R734 GND.n65 GND.n64 4.65
R735 GND.n68 GND.n67 4.65
R736 GND.n71 GND.n70 4.65
R737 GND.n78 GND.n77 4.65
R738 GND.n81 GND.n80 4.65
R739 GND.n84 GND.n83 4.65
R740 GND.n87 GND.n86 4.65
R741 GND.n90 GND.n89 4.65
R742 GND.n93 GND.n92 4.65
R743 GND.n96 GND.n95 4.65
R744 GND.n99 GND.n98 4.65
R745 GND.n102 GND.n101 4.65
R746 GND.n110 GND.n109 4.65
R747 GND.n113 GND.n112 4.65
R748 GND.n116 GND.n115 4.65
R749 GND.n233 GND.n232 4.65
R750 GND.n226 GND.n225 4.65
R751 GND.n223 GND.n222 4.65
R752 GND.n220 GND.n219 4.65
R753 GND.n217 GND.n216 4.65
R754 GND.n214 GND.n213 4.65
R755 GND.n206 GND.n205 4.65
R756 GND.n203 GND.n202 4.65
R757 GND.n196 GND.n195 4.65
R758 GND.n193 GND.n192 4.65
R759 GND.n190 GND.n189 4.65
R760 GND.n187 GND.n186 4.65
R761 GND.n184 GND.n183 4.65
R762 GND.n181 GND.n180 4.65
R763 GND.n178 GND.n177 4.65
R764 GND.n175 GND.n174 4.65
R765 GND.n172 GND.n171 4.65
R766 GND.n169 GND.n168 4.65
R767 GND.n164 GND.n163 4.65
R768 GND.n161 GND.n160 4.65
R769 GND.n154 GND.n153 4.65
R770 GND.n151 GND.n150 4.65
R771 GND.n148 GND.n147 4.65
R772 GND.n145 GND.n144 4.65
R773 GND.n142 GND.n141 4.65
R774 GND.n139 GND.n138 4.65
R775 GND.n136 GND.n135 4.65
R776 GND.n133 GND.n132 4.65
R777 GND.n130 GND.n129 4.65
R778 GND.n127 GND.n126 4.65
R779 GND.n122 GND.n121 4.65
R780 GND.n19 GND.n17 4.129
R781 GND.n213 GND.n211 4.129
R782 GND.n3 GND.n0 3.407
R783 GND.n3 GND.n2 2.844
R784 GND.n6 GND.n3 1.063
R785 GND.n118 GND.n117 0.474
R786 GND.n33 GND.n26 0.29
R787 GND.n78 GND.n71 0.29
R788 GND.n203 GND.n196 0.29
R789 GND.n161 GND.n154 0.29
R790 GND.n119 GND 0.207
R791 GND.n64 GND.n63 0.206
R792 GND.n109 GND.n108 0.206
R793 GND.n168 GND.n167 0.206
R794 GND.n126 GND.n125 0.206
R795 GND.n51 GND.n48 0.197
R796 GND.n96 GND.n93 0.197
R797 GND.n181 GND.n178 0.197
R798 GND.n139 GND.n136 0.197
R799 GND.n12 GND.n9 0.181
R800 GND.n220 GND.n217 0.181
R801 GND.n9 GND.n6 0.145
R802 GND.n20 GND.n12 0.145
R803 GND.n23 GND.n20 0.145
R804 GND.n26 GND.n23 0.145
R805 GND.n36 GND.n33 0.145
R806 GND.n39 GND.n36 0.145
R807 GND.n42 GND.n39 0.145
R808 GND.n45 GND.n42 0.145
R809 GND.n48 GND.n45 0.145
R810 GND.n54 GND.n51 0.145
R811 GND.n57 GND.n54 0.145
R812 GND.n65 GND.n57 0.145
R813 GND.n68 GND.n65 0.145
R814 GND.n71 GND.n68 0.145
R815 GND.n81 GND.n78 0.145
R816 GND.n84 GND.n81 0.145
R817 GND.n87 GND.n84 0.145
R818 GND.n90 GND.n87 0.145
R819 GND.n93 GND.n90 0.145
R820 GND.n99 GND.n96 0.145
R821 GND.n102 GND.n99 0.145
R822 GND.n110 GND.n102 0.145
R823 GND.n113 GND.n110 0.145
R824 GND.n116 GND.n113 0.145
R825 GND GND.n116 0.145
R826 GND GND.n233 0.145
R827 GND.n233 GND.n226 0.145
R828 GND.n226 GND.n223 0.145
R829 GND.n223 GND.n220 0.145
R830 GND.n217 GND.n214 0.145
R831 GND.n214 GND.n206 0.145
R832 GND.n206 GND.n203 0.145
R833 GND.n196 GND.n193 0.145
R834 GND.n193 GND.n190 0.145
R835 GND.n190 GND.n187 0.145
R836 GND.n187 GND.n184 0.145
R837 GND.n184 GND.n181 0.145
R838 GND.n178 GND.n175 0.145
R839 GND.n175 GND.n172 0.145
R840 GND.n172 GND.n169 0.145
R841 GND.n169 GND.n164 0.145
R842 GND.n164 GND.n161 0.145
R843 GND.n154 GND.n151 0.145
R844 GND.n151 GND.n148 0.145
R845 GND.n148 GND.n145 0.145
R846 GND.n145 GND.n142 0.145
R847 GND.n142 GND.n139 0.145
R848 GND.n136 GND.n133 0.145
R849 GND.n133 GND.n130 0.145
R850 GND.n130 GND.n127 0.145
R851 GND.n127 GND.n122 0.145
R852 GND.n122 GND.n119 0.145
R853 a_147_187.n6 a_147_187.t15 512.525
R854 a_147_187.n4 a_147_187.t9 472.359
R855 a_147_187.n2 a_147_187.t14 472.359
R856 a_147_187.n7 a_147_187.t12 417.109
R857 a_147_187.n4 a_147_187.t13 384.527
R858 a_147_187.n2 a_147_187.t10 384.527
R859 a_147_187.n13 a_147_187.n12 379.457
R860 a_147_187.n6 a_147_187.t11 371.139
R861 a_147_187.n5 a_147_187.t8 370.613
R862 a_147_187.n3 a_147_187.t7 370.613
R863 a_147_187.n7 a_147_187.n6 179.837
R864 a_147_187.n16 a_147_187.n15 161.352
R865 a_147_187.n5 a_147_187.n4 127.096
R866 a_147_187.n3 a_147_187.n2 127.096
R867 a_147_187.n14 a_147_187.n13 123.481
R868 a_147_187.n14 a_147_187.n1 95.095
R869 a_147_187.n15 a_147_187.n0 95.095
R870 a_147_187.n15 a_147_187.n14 66.258
R871 a_147_187.n12 a_147_187.n11 22.578
R872 a_147_187.n1 a_147_187.t6 14.282
R873 a_147_187.n1 a_147_187.t4 14.282
R874 a_147_187.n0 a_147_187.t2 14.282
R875 a_147_187.n0 a_147_187.t3 14.282
R876 a_147_187.t1 a_147_187.n16 14.282
R877 a_147_187.n16 a_147_187.t0 14.282
R878 a_147_187.n8 a_147_187.n7 12.222
R879 a_147_187.n9 a_147_187.n3 10.046
R880 a_147_187.n12 a_147_187.n10 8.58
R881 a_147_187.n8 a_147_187.n5 4.65
R882 a_147_187.n13 a_147_187.n9 4.65
R883 a_147_187.n9 a_147_187.n8 4.035
R884 a_4626_101.n3 a_4626_101.n1 42.788
R885 a_4626_101.t0 a_4626_101.n0 8.137
R886 a_4626_101.n3 a_4626_101.n2 4.665
R887 a_4626_101.t0 a_4626_101.n3 0.06
R888 a_4151_989.n0 a_4151_989.t5 454.685
R889 a_4151_989.n0 a_4151_989.t6 428.979
R890 a_4151_989.n3 a_4151_989.n2 355.179
R891 a_4151_989.n1 a_4151_989.t7 339.542
R892 a_4151_989.n5 a_4151_989.n4 157.964
R893 a_4151_989.n1 a_4151_989.n0 143.429
R894 a_4151_989.n5 a_4151_989.n3 132.141
R895 a_4151_989.n6 a_4151_989.n5 91.705
R896 a_4151_989.n4 a_4151_989.t3 14.282
R897 a_4151_989.n4 a_4151_989.t4 14.282
R898 a_4151_989.n6 a_4151_989.t0 14.282
R899 a_4151_989.t1 a_4151_989.n6 14.282
R900 a_4151_989.n3 a_4151_989.n1 12.247
R901 a_2036_101.n11 a_2036_101.n10 68.43
R902 a_2036_101.n3 a_2036_101.n2 62.817
R903 a_2036_101.n7 a_2036_101.n6 38.626
R904 a_2036_101.n6 a_2036_101.n5 35.955
R905 a_2036_101.n3 a_2036_101.n1 26.202
R906 a_2036_101.t0 a_2036_101.n3 19.737
R907 a_2036_101.t1 a_2036_101.n8 8.137
R908 a_2036_101.t0 a_2036_101.n4 7.273
R909 a_2036_101.t0 a_2036_101.n0 6.109
R910 a_2036_101.t1 a_2036_101.n7 4.864
R911 a_2036_101.t0 a_2036_101.n12 2.074
R912 a_2036_101.n12 a_2036_101.t1 0.937
R913 a_2036_101.t1 a_2036_101.n11 0.763
R914 a_2036_101.n11 a_2036_101.n9 0.185
R915 RN.n0 RN.t4 479.223
R916 RN.n5 RN.t0 454.685
R917 RN.n2 RN.t1 454.685
R918 RN.n5 RN.t3 428.979
R919 RN.n2 RN.t8 428.979
R920 RN.n0 RN.t5 375.52
R921 RN.n6 RN.n5 254.865
R922 RN.n3 RN.n2 254.865
R923 RN.n1 RN.n0 252.188
R924 RN.n1 RN.t7 231.854
R925 RN.n6 RN.t6 228.106
R926 RN.n3 RN.t2 228.106
R927 RN.n4 RN.n1 7.325
R928 RN.n7 RN.n4 5.94
R929 RN.n4 RN.n3 4.65
R930 RN.n7 RN.n6 4.65
R931 RN.n7 RN 0.046
R932 a_372_210.n9 a_372_210.n7 171.558
R933 a_372_210.t0 a_372_210.n9 75.765
R934 a_372_210.n3 a_372_210.n1 74.827
R935 a_372_210.n3 a_372_210.n2 27.476
R936 a_372_210.n7 a_372_210.n6 27.2
R937 a_372_210.n5 a_372_210.n4 23.498
R938 a_372_210.n7 a_372_210.n5 22.4
R939 a_372_210.t0 a_372_210.n11 20.241
R940 a_372_210.t0 a_372_210.n3 13.984
R941 a_372_210.n11 a_372_210.n10 13.494
R942 a_372_210.t0 a_372_210.n0 8.137
R943 a_372_210.n9 a_372_210.n8 1.505
R944 a_2962_210.n9 a_2962_210.n7 171.558
R945 a_2962_210.t0 a_2962_210.n9 75.765
R946 a_2962_210.n3 a_2962_210.n1 74.827
R947 a_2962_210.n3 a_2962_210.n2 27.476
R948 a_2962_210.n7 a_2962_210.n6 27.2
R949 a_2962_210.n5 a_2962_210.n4 23.498
R950 a_2962_210.n7 a_2962_210.n5 22.4
R951 a_2962_210.t0 a_2962_210.n11 20.241
R952 a_2962_210.t0 a_2962_210.n3 13.984
R953 a_2962_210.n11 a_2962_210.n10 13.494
R954 a_2962_210.t0 a_2962_210.n0 8.137
R955 a_2962_210.n9 a_2962_210.n8 1.505
R956 a_91_103.t0 a_91_103.n7 59.616
R957 a_91_103.n4 a_91_103.n2 54.496
R958 a_91_103.n4 a_91_103.n3 54.496
R959 a_91_103.n1 a_91_103.n0 24.679
R960 a_91_103.t0 a_91_103.n1 7.505
R961 a_91_103.n6 a_91_103.n5 2.455
R962 a_91_103.n6 a_91_103.n4 0.636
R963 a_91_103.t0 a_91_103.n6 0.246
R964 a_3924_210.n9 a_3924_210.n7 171.558
R965 a_3924_210.t0 a_3924_210.n9 75.765
R966 a_3924_210.n3 a_3924_210.n1 74.827
R967 a_3924_210.n3 a_3924_210.n2 27.476
R968 a_3924_210.n7 a_3924_210.n6 27.2
R969 a_3924_210.n5 a_3924_210.n4 23.498
R970 a_3924_210.n7 a_3924_210.n5 22.4
R971 a_3924_210.t0 a_3924_210.n11 20.241
R972 a_3924_210.t0 a_3924_210.n3 13.984
R973 a_3924_210.n11 a_3924_210.n10 13.494
R974 a_3924_210.t0 a_3924_210.n0 8.137
R975 a_3924_210.n9 a_3924_210.n8 1.505
R976 a_3643_103.t0 a_3643_103.n7 59.616
R977 a_3643_103.n4 a_3643_103.n2 54.496
R978 a_3643_103.n4 a_3643_103.n3 54.496
R979 a_3643_103.n1 a_3643_103.n0 24.679
R980 a_3643_103.t0 a_3643_103.n1 7.505
R981 a_3643_103.n6 a_3643_103.n5 2.455
R982 a_3643_103.n6 a_3643_103.n4 0.636
R983 a_3643_103.t0 a_3643_103.n6 0.246
R984 a_2681_103.n5 a_2681_103.n4 66.708
R985 a_2681_103.n2 a_2681_103.n0 25.439
R986 a_2681_103.n5 a_2681_103.n3 19.496
R987 a_2681_103.t0 a_2681_103.n5 13.756
R988 a_2681_103.n2 a_2681_103.n1 2.455
R989 a_2681_103.t0 a_2681_103.n2 0.246
C8 RN GND 1.72fF
C9 VDD GND 8.55fF
C10 a_2681_103.n0 GND 0.11fF
C11 a_2681_103.n1 GND 0.04fF
C12 a_2681_103.n2 GND 0.03fF
C13 a_2681_103.n3 GND 0.07fF
C14 a_2681_103.n4 GND 0.08fF
C15 a_2681_103.n5 GND 0.03fF
C16 a_3643_103.n0 GND 0.08fF
C17 a_3643_103.n1 GND 0.07fF
C18 a_3643_103.n2 GND 0.04fF
C19 a_3643_103.n3 GND 0.06fF
C20 a_3643_103.n4 GND 0.03fF
C21 a_3643_103.n5 GND 0.04fF
C22 a_3643_103.n7 GND 0.08fF
C23 a_3924_210.n0 GND 0.07fF
C24 a_3924_210.n1 GND 0.09fF
C25 a_3924_210.n2 GND 0.12fF
C26 a_3924_210.n3 GND 0.08fF
C27 a_3924_210.n4 GND 0.02fF
C28 a_3924_210.n5 GND 0.03fF
C29 a_3924_210.n6 GND 0.02fF
C30 a_3924_210.n7 GND 0.03fF
C31 a_3924_210.n8 GND 0.02fF
C32 a_3924_210.n9 GND 0.13fF
C33 a_3924_210.n10 GND 0.08fF
C34 a_3924_210.n11 GND 0.02fF
C35 a_91_103.n0 GND 0.08fF
C36 a_91_103.n1 GND 0.07fF
C37 a_91_103.n2 GND 0.04fF
C38 a_91_103.n3 GND 0.06fF
C39 a_91_103.n4 GND 0.03fF
C40 a_91_103.n5 GND 0.03fF
C41 a_91_103.n7 GND 0.08fF
C42 a_2962_210.n0 GND 0.07fF
C43 a_2962_210.n1 GND 0.09fF
C44 a_2962_210.n2 GND 0.12fF
C45 a_2962_210.n3 GND 0.08fF
C46 a_2962_210.n4 GND 0.02fF
C47 a_2962_210.n5 GND 0.03fF
C48 a_2962_210.n6 GND 0.02fF
C49 a_2962_210.n7 GND 0.03fF
C50 a_2962_210.n8 GND 0.02fF
C51 a_2962_210.n9 GND 0.13fF
C52 a_2962_210.n10 GND 0.08fF
C53 a_2962_210.n11 GND 0.02fF
C54 a_2962_210.t0 GND 0.31fF
C55 a_372_210.n0 GND 0.07fF
C56 a_372_210.n1 GND 0.09fF
C57 a_372_210.n2 GND 0.12fF
C58 a_372_210.n3 GND 0.08fF
C59 a_372_210.n4 GND 0.02fF
C60 a_372_210.n5 GND 0.03fF
C61 a_372_210.n6 GND 0.02fF
C62 a_372_210.n7 GND 0.03fF
C63 a_372_210.n8 GND 0.02fF
C64 a_372_210.n9 GND 0.13fF
C65 a_372_210.n10 GND 0.08fF
C66 a_372_210.n11 GND 0.02fF
C67 a_372_210.t0 GND 0.31fF
C68 RN.n0 GND 0.33fF
C69 RN.t7 GND 0.36fF
C70 RN.n1 GND 0.40fF
C71 RN.n2 GND 0.32fF
C72 RN.t2 GND 0.36fF
C73 RN.n3 GND 0.30fF
C74 RN.n4 GND 0.92fF
C75 RN.n5 GND 0.32fF
C76 RN.t6 GND 0.37fF
C77 RN.n6 GND 0.30fF
C78 RN.n7 GND 0.53fF
C79 a_2036_101.n0 GND 0.02fF
C80 a_2036_101.n1 GND 0.09fF
C81 a_2036_101.n2 GND 0.08fF
C82 a_2036_101.n3 GND 0.03fF
C83 a_2036_101.n4 GND 0.01fF
C84 a_2036_101.n5 GND 0.04fF
C85 a_2036_101.n6 GND 0.04fF
C86 a_2036_101.n7 GND 0.02fF
C87 a_2036_101.n8 GND 0.05fF
C88 a_2036_101.n9 GND 0.15fF
C89 a_2036_101.n10 GND 0.08fF
C90 a_2036_101.n11 GND 0.08fF
C91 a_2036_101.t1 GND 0.23fF
C92 a_2036_101.n12 GND 0.01fF
C93 a_4151_989.n0 GND 0.30fF
C94 a_4151_989.n1 GND 0.76fF
C95 a_4151_989.n2 GND 0.36fF
C96 a_4151_989.n3 GND 0.86fF
C97 a_4151_989.n4 GND 0.48fF
C98 a_4151_989.n5 GND 0.54fF
C99 a_4151_989.n6 GND 0.38fF
C100 a_4626_101.n0 GND 0.05fF
C101 a_4626_101.n1 GND 0.12fF
C102 a_4626_101.n2 GND 0.04fF
C103 a_4626_101.n3 GND 0.16fF
C104 a_147_187.n0 GND 0.58fF
C105 a_147_187.n1 GND 0.58fF
C106 a_147_187.n2 GND 0.41fF
C107 a_147_187.t7 GND 0.86fF
C108 a_147_187.n3 GND 1.08fF
C109 a_147_187.n4 GND 0.41fF
C110 a_147_187.t8 GND 0.86fF
C111 a_147_187.n5 GND 0.58fF
C112 a_147_187.n6 GND 0.42fF
C113 a_147_187.n7 GND 1.51fF
C114 a_147_187.n8 GND 2.43fF
C115 a_147_187.n9 GND 2.02fF
C116 a_147_187.n10 GND 0.06fF
C117 a_147_187.n11 GND 0.08fF
C118 a_147_187.n12 GND 0.45fF
C119 a_147_187.n13 GND 0.80fF
C120 a_147_187.n14 GND 0.58fF
C121 a_147_187.n15 GND 0.70fF
C122 a_147_187.n16 GND 0.74fF
C123 a_1334_210.n0 GND 0.02fF
C124 a_1334_210.n1 GND 0.09fF
C125 a_1334_210.n2 GND 0.12fF
C126 a_1334_210.n3 GND 0.08fF
C127 a_1334_210.n4 GND 0.08fF
C128 a_1334_210.n5 GND 0.02fF
C129 a_1334_210.t1 GND 0.29fF
C130 a_1334_210.n6 GND 0.09fF
C131 a_1334_210.n7 GND 0.02fF
C132 a_1334_210.n8 GND 0.13fF
C133 a_1334_210.n9 GND 0.02fF
C134 a_1334_210.n10 GND 0.03fF
C135 a_1334_210.n11 GND 0.02fF
C136 a_1053_103.n0 GND 0.13fF
C137 a_1053_103.n1 GND 0.04fF
C138 a_1053_103.n2 GND 0.09fF
C139 a_1053_103.n3 GND 0.03fF
C140 a_1053_103.n4 GND 0.08fF
C141 a_1053_103.n5 GND 0.07fF
C142 a_1053_103.n6 GND 0.04fF
C143 QN.n0 GND 0.27fF
C144 QN.n1 GND 0.39fF
C145 QN.n2 GND 0.32fF
C146 QN.n3 GND 0.32fF
C147 QN.n4 GND 0.41fF
C148 QN.n5 GND 0.39fF
C149 QN.n6 GND 0.37fF
C150 QN.n7 GND 0.28fF
C151 QN.n8 GND 0.44fF
C152 QN.n9 GND 0.25fF
C153 a_2141_1050.n0 GND 0.36fF
C154 a_2141_1050.n1 GND 0.31fF
C155 a_2141_1050.n2 GND 0.62fF
C156 a_2141_1050.n3 GND 0.31fF
C157 a_2141_1050.n4 GND 0.65fF
C158 a_2141_1050.n5 GND 0.54fF
C159 a_2141_1050.n6 GND 0.46fF
C160 a_277_1050.n0 GND 0.41fF
C161 a_277_1050.n1 GND 1.62fF
C162 a_277_1050.n2 GND 0.41fF
C163 a_277_1050.n3 GND 0.65fF
C164 a_277_1050.n4 GND 2.31fF
C165 a_277_1050.n5 GND 0.05fF
C166 a_277_1050.n6 GND 0.07fF
C167 a_277_1050.n7 GND 0.05fF
C168 a_277_1050.n8 GND 0.35fF
C169 a_277_1050.n9 GND 0.76fF
C170 a_277_1050.n10 GND 0.53fF
C171 a_277_1050.n11 GND 0.67fF
C172 a_277_1050.n12 GND 0.64fF
C173 a_277_1050.n13 GND 0.56fF
C174 a_277_1050.n14 GND 0.53fF
C175 a_599_989.n0 GND 0.40fF
C176 a_599_989.n1 GND 0.34fF
C177 a_599_989.n2 GND 0.48fF
C178 a_599_989.n3 GND 0.34fF
C179 a_599_989.t9 GND 0.55fF
C180 a_599_989.n4 GND 0.65fF
C181 a_599_989.n5 GND 1.04fF
C182 a_599_989.n6 GND 0.04fF
C183 a_599_989.n7 GND 0.06fF
C184 a_599_989.n8 GND 0.04fF
C185 a_599_989.n9 GND 0.23fF
C186 a_599_989.n10 GND 0.54fF
C187 a_599_989.n11 GND 0.46fF
C188 a_599_989.n12 GND 0.51fF
C189 a_599_989.n13 GND 0.49fF
C190 a_599_989.n14 GND 0.40fF
C191 VDD.n1 GND 0.03fF
C192 VDD.n2 GND 0.14fF
C193 VDD.n3 GND 0.03fF
C194 VDD.n4 GND 0.02fF
C195 VDD.n5 GND 0.06fF
C196 VDD.n6 GND 0.02fF
C197 VDD.n7 GND 0.02fF
C198 VDD.n8 GND 0.02fF
C199 VDD.n9 GND 0.02fF
C200 VDD.n10 GND 0.02fF
C201 VDD.n11 GND 0.02fF
C202 VDD.n12 GND 0.02fF
C203 VDD.n13 GND 0.02fF
C204 VDD.n14 GND 0.04fF
C205 VDD.n15 GND 0.01fF
C206 VDD.n20 GND 0.46fF
C207 VDD.n21 GND 0.27fF
C208 VDD.n22 GND 0.02fF
C209 VDD.n23 GND 0.03fF
C210 VDD.n24 GND 0.06fF
C211 VDD.n25 GND 0.24fF
C212 VDD.n26 GND 0.01fF
C213 VDD.n27 GND 0.01fF
C214 VDD.n28 GND 0.01fF
C215 VDD.n29 GND 0.17fF
C216 VDD.n30 GND 0.01fF
C217 VDD.n31 GND 0.02fF
C218 VDD.n32 GND 0.08fF
C219 VDD.n33 GND 0.08fF
C220 VDD.n34 GND 0.05fF
C221 VDD.n35 GND 0.01fF
C222 VDD.n36 GND 0.02fF
C223 VDD.n37 GND 0.03fF
C224 VDD.n38 GND 0.14fF
C225 VDD.n39 GND 0.01fF
C226 VDD.n40 GND 0.02fF
C227 VDD.n41 GND 0.03fF
C228 VDD.n42 GND 0.16fF
C229 VDD.n43 GND 0.01fF
C230 VDD.n44 GND 0.02fF
C231 VDD.n45 GND 0.02fF
C232 VDD.n46 GND 0.06fF
C233 VDD.n47 GND 0.25fF
C234 VDD.n48 GND 0.01fF
C235 VDD.n49 GND 0.01fF
C236 VDD.n50 GND 0.02fF
C237 VDD.n51 GND 0.27fF
C238 VDD.n52 GND 0.01fF
C239 VDD.n53 GND 0.02fF
C240 VDD.n54 GND 0.03fF
C241 VDD.n55 GND 0.05fF
C242 VDD.n56 GND 0.02fF
C243 VDD.n57 GND 0.02fF
C244 VDD.n58 GND 0.02fF
C245 VDD.n59 GND 0.02fF
C246 VDD.n60 GND 0.02fF
C247 VDD.n61 GND 0.02fF
C248 VDD.n62 GND 0.02fF
C249 VDD.n63 GND 0.02fF
C250 VDD.n64 GND 0.02fF
C251 VDD.n65 GND 0.02fF
C252 VDD.n66 GND 0.02fF
C253 VDD.n67 GND 0.03fF
C254 VDD.n68 GND 0.02fF
C255 VDD.n69 GND 0.27fF
C256 VDD.n70 GND 0.02fF
C257 VDD.n71 GND 0.02fF
C258 VDD.n73 GND 0.02fF
C259 VDD.n77 GND 0.27fF
C260 VDD.n78 GND 0.27fF
C261 VDD.n79 GND 0.01fF
C262 VDD.n80 GND 0.02fF
C263 VDD.n81 GND 0.03fF
C264 VDD.n82 GND 0.27fF
C265 VDD.n83 GND 0.01fF
C266 VDD.n84 GND 0.02fF
C267 VDD.n85 GND 0.02fF
C268 VDD.n86 GND 0.22fF
C269 VDD.n87 GND 0.01fF
C270 VDD.n88 GND 0.07fF
C271 VDD.n89 GND 0.02fF
C272 VDD.n90 GND 0.17fF
C273 VDD.n91 GND 0.01fF
C274 VDD.n92 GND 0.02fF
C275 VDD.n93 GND 0.02fF
C276 VDD.n94 GND 0.16fF
C277 VDD.n95 GND 0.01fF
C278 VDD.n96 GND 0.08fF
C279 VDD.n97 GND 0.05fF
C280 VDD.n98 GND 0.02fF
C281 VDD.n99 GND 0.02fF
C282 VDD.n100 GND 0.14fF
C283 VDD.n101 GND 0.01fF
C284 VDD.n102 GND 0.02fF
C285 VDD.n103 GND 0.03fF
C286 VDD.n104 GND 0.15fF
C287 VDD.n105 GND 0.01fF
C288 VDD.n106 GND 0.02fF
C289 VDD.n107 GND 0.03fF
C290 VDD.n108 GND 0.08fF
C291 VDD.n109 GND 0.05fF
C292 VDD.n110 GND 0.16fF
C293 VDD.n111 GND 0.01fF
C294 VDD.n112 GND 0.02fF
C295 VDD.n113 GND 0.02fF
C296 VDD.n114 GND 0.17fF
C297 VDD.n115 GND 0.01fF
C298 VDD.n116 GND 0.02fF
C299 VDD.n117 GND 0.02fF
C300 VDD.n118 GND 0.06fF
C301 VDD.n119 GND 0.22fF
C302 VDD.n120 GND 0.01fF
C303 VDD.n121 GND 0.01fF
C304 VDD.n122 GND 0.02fF
C305 VDD.n123 GND 0.27fF
C306 VDD.n124 GND 0.01fF
C307 VDD.n125 GND 0.02fF
C308 VDD.n126 GND 0.02fF
C309 VDD.n127 GND 0.27fF
C310 VDD.n128 GND 0.01fF
C311 VDD.n129 GND 0.02fF
C312 VDD.n130 GND 0.03fF
C313 VDD.n131 GND 0.31fF
C314 VDD.n132 GND 0.02fF
C315 VDD.n133 GND 0.02fF
C316 VDD.n134 GND 0.02fF
C317 VDD.n135 GND 0.06fF
C318 VDD.n136 GND 0.02fF
C319 VDD.n137 GND 0.02fF
C320 VDD.n138 GND 0.02fF
C321 VDD.n139 GND 0.02fF
C322 VDD.n140 GND 0.02fF
C323 VDD.n141 GND 0.02fF
C324 VDD.n142 GND 0.02fF
C325 VDD.n143 GND 0.02fF
C326 VDD.n144 GND 0.02fF
C327 VDD.n145 GND 0.02fF
C328 VDD.n146 GND 0.03fF
C329 VDD.n147 GND 0.02fF
C330 VDD.n148 GND 0.02fF
C331 VDD.n152 GND 0.27fF
C332 VDD.n153 GND 0.27fF
C333 VDD.n154 GND 0.01fF
C334 VDD.n155 GND 0.02fF
C335 VDD.n156 GND 0.03fF
C336 VDD.n157 GND 0.27fF
C337 VDD.n158 GND 0.01fF
C338 VDD.n159 GND 0.02fF
C339 VDD.n160 GND 0.02fF
C340 VDD.n161 GND 0.22fF
C341 VDD.n162 GND 0.01fF
C342 VDD.n163 GND 0.07fF
C343 VDD.n164 GND 0.02fF
C344 VDD.n165 GND 0.17fF
C345 VDD.n166 GND 0.01fF
C346 VDD.n167 GND 0.02fF
C347 VDD.n168 GND 0.02fF
C348 VDD.n169 GND 0.16fF
C349 VDD.n170 GND 0.01fF
C350 VDD.n171 GND 0.08fF
C351 VDD.n172 GND 0.05fF
C352 VDD.n173 GND 0.02fF
C353 VDD.n174 GND 0.02fF
C354 VDD.n175 GND 0.14fF
C355 VDD.n176 GND 0.01fF
C356 VDD.n177 GND 0.02fF
C357 VDD.n178 GND 0.03fF
C358 VDD.n179 GND 0.15fF
C359 VDD.n180 GND 0.01fF
C360 VDD.n181 GND 0.02fF
C361 VDD.n182 GND 0.03fF
C362 VDD.n183 GND 0.08fF
C363 VDD.n184 GND 0.05fF
C364 VDD.n185 GND 0.16fF
C365 VDD.n186 GND 0.01fF
C366 VDD.n187 GND 0.02fF
C367 VDD.n188 GND 0.02fF
C368 VDD.n189 GND 0.17fF
C369 VDD.n190 GND 0.01fF
C370 VDD.n191 GND 0.02fF
C371 VDD.n192 GND 0.02fF
C372 VDD.n193 GND 0.06fF
C373 VDD.n194 GND 0.22fF
C374 VDD.n195 GND 0.01fF
C375 VDD.n196 GND 0.01fF
C376 VDD.n197 GND 0.02fF
C377 VDD.n198 GND 0.27fF
C378 VDD.n199 GND 0.01fF
C379 VDD.n200 GND 0.02fF
C380 VDD.n201 GND 0.02fF
C381 VDD.n202 GND 0.02fF
C382 VDD.n206 GND 0.27fF
C383 VDD.n207 GND 0.27fF
C384 VDD.n208 GND 0.01fF
C385 VDD.n209 GND 0.02fF
C386 VDD.n210 GND 0.02fF
C387 VDD.n211 GND 0.18fF
C388 VDD.n212 GND 0.02fF
C389 VDD.n213 GND 0.02fF
C390 VDD.n214 GND 0.06fF
C391 VDD.n215 GND 0.02fF
C392 VDD.n216 GND 0.02fF
C393 VDD.n217 GND 0.02fF
C394 VDD.n218 GND 0.02fF
C395 VDD.n219 GND 0.02fF
C396 VDD.n220 GND 0.02fF
C397 VDD.n221 GND 0.02fF
C398 VDD.n222 GND 0.02fF
C399 VDD.n223 GND 0.03fF
C400 VDD.n224 GND 0.04fF
C401 VDD.n225 GND 0.02fF
C402 VDD.n229 GND 0.46fF
C403 VDD.n230 GND 0.27fF
C404 VDD.n231 GND 0.02fF
C405 VDD.n232 GND 0.03fF
C406 VDD.n233 GND 0.03fF
C407 VDD.n234 GND 0.27fF
C408 VDD.n235 GND 0.01fF
C409 VDD.n236 GND 0.02fF
C410 VDD.n237 GND 0.02fF
C411 VDD.n238 GND 0.06fF
C412 VDD.n239 GND 0.22fF
C413 VDD.n240 GND 0.01fF
C414 VDD.n241 GND 0.01fF
C415 VDD.n242 GND 0.02fF
C416 VDD.n243 GND 0.17fF
C417 VDD.n244 GND 0.01fF
C418 VDD.n245 GND 0.02fF
C419 VDD.n246 GND 0.02fF
C420 VDD.n247 GND 0.08fF
C421 VDD.n248 GND 0.05fF
C422 VDD.n249 GND 0.16fF
C423 VDD.n250 GND 0.01fF
C424 VDD.n251 GND 0.02fF
C425 VDD.n252 GND 0.02fF
C426 VDD.n253 GND 0.15fF
C427 VDD.n254 GND 0.01fF
C428 VDD.n255 GND 0.02fF
C429 VDD.n256 GND 0.03fF
C430 VDD.n257 GND 0.14fF
C431 VDD.n258 GND 0.01fF
C432 VDD.n259 GND 0.02fF
C433 VDD.n260 GND 0.03fF
C434 VDD.n261 GND 0.16fF
C435 VDD.n262 GND 0.01fF
C436 VDD.n263 GND 0.08fF
C437 VDD.n264 GND 0.05fF
C438 VDD.n265 GND 0.02fF
C439 VDD.n266 GND 0.02fF
C440 VDD.n267 GND 0.17fF
C441 VDD.n268 GND 0.01fF
C442 VDD.n269 GND 0.02fF
C443 VDD.n270 GND 0.02fF
C444 VDD.n271 GND 0.22fF
C445 VDD.n272 GND 0.01fF
C446 VDD.n273 GND 0.07fF
C447 VDD.n274 GND 0.02fF
C448 VDD.n275 GND 0.27fF
C449 VDD.n276 GND 0.01fF
C450 VDD.n277 GND 0.02fF
C451 VDD.n278 GND 0.02fF
C452 VDD.n279 GND 0.27fF
C453 VDD.n280 GND 0.01fF
C454 VDD.n281 GND 0.02fF
C455 VDD.n282 GND 0.03fF
C456 VDD.n283 GND 0.05fF
C457 VDD.n284 GND 0.02fF
C458 VDD.n285 GND 0.02fF
C459 VDD.n286 GND 0.02fF
C460 VDD.n287 GND 0.02fF
C461 VDD.n288 GND 0.02fF
C462 VDD.n289 GND 0.02fF
C463 VDD.n290 GND 0.02fF
C464 VDD.n291 GND 0.02fF
C465 VDD.n292 GND 0.02fF
C466 VDD.n293 GND 0.02fF
C467 VDD.n294 GND 0.02fF
C468 VDD.n295 GND 0.03fF
C469 VDD.n296 GND 0.02fF
C470 VDD.n299 GND 0.02fF
C471 VDD.n301 GND 0.02fF
C472 VDD.n302 GND 0.31fF
C473 VDD.n303 GND 0.02fF
C474 VDD.n305 GND 0.27fF
C475 VDD.n306 GND 0.27fF
C476 VDD.n307 GND 0.01fF
C477 VDD.n308 GND 0.02fF
C478 VDD.n309 GND 0.03fF
C479 VDD.n310 GND 0.27fF
C480 VDD.n311 GND 0.01fF
C481 VDD.n312 GND 0.02fF
C482 VDD.n313 GND 0.02fF
C483 VDD.n314 GND 0.06fF
C484 VDD.n315 GND 0.22fF
C485 VDD.n316 GND 0.01fF
C486 VDD.n317 GND 0.01fF
C487 VDD.n318 GND 0.02fF
C488 VDD.n319 GND 0.17fF
C489 VDD.n320 GND 0.01fF
C490 VDD.n321 GND 0.02fF
C491 VDD.n322 GND 0.02fF
C492 VDD.n323 GND 0.08fF
C493 VDD.n324 GND 0.05fF
C494 VDD.n325 GND 0.16fF
C495 VDD.n326 GND 0.01fF
C496 VDD.n327 GND 0.02fF
C497 VDD.n328 GND 0.02fF
C498 VDD.n329 GND 0.15fF
C499 VDD.n330 GND 0.01fF
C500 VDD.n331 GND 0.02fF
C501 VDD.n332 GND 0.03fF
C502 VDD.n333 GND 0.14fF
C503 VDD.n334 GND 0.01fF
C504 VDD.n335 GND 0.02fF
C505 VDD.n336 GND 0.03fF
C506 VDD.n337 GND 0.16fF
C507 VDD.n338 GND 0.01fF
C508 VDD.n339 GND 0.08fF
C509 VDD.n340 GND 0.05fF
C510 VDD.n341 GND 0.02fF
C511 VDD.n342 GND 0.02fF
C512 VDD.n343 GND 0.17fF
C513 VDD.n344 GND 0.01fF
C514 VDD.n345 GND 0.02fF
C515 VDD.n346 GND 0.02fF
C516 VDD.n347 GND 0.22fF
C517 VDD.n348 GND 0.01fF
C518 VDD.n349 GND 0.07fF
C519 VDD.n350 GND 0.02fF
C520 VDD.n351 GND 0.27fF
C521 VDD.n352 GND 0.01fF
C522 VDD.n353 GND 0.02fF
C523 VDD.n354 GND 0.02fF
C524 VDD.n355 GND 0.27fF
C525 VDD.n356 GND 0.01fF
C526 VDD.n357 GND 0.02fF
C527 VDD.n358 GND 0.03fF
C528 VDD.n359 GND 0.26fF
C529 VDD.n360 GND 0.02fF
C530 VDD.n361 GND 0.02fF
C531 VDD.n362 GND 0.02fF
C532 VDD.n363 GND 0.06fF
C533 VDD.n364 GND 0.02fF
C534 VDD.n365 GND 0.02fF
C535 VDD.n366 GND 0.02fF
C536 VDD.n367 GND 0.02fF
C537 VDD.n368 GND 0.02fF
C538 VDD.n369 GND 0.02fF
C539 VDD.n370 GND 0.02fF
C540 VDD.n371 GND 0.02fF
C541 VDD.n372 GND 0.02fF
C542 VDD.n373 GND 0.02fF
C543 VDD.n374 GND 0.03fF
C544 VDD.n375 GND 0.02fF
C545 VDD.n376 GND 0.02fF
C546 VDD.n380 GND 0.27fF
C547 VDD.n381 GND 0.27fF
C548 VDD.n382 GND 0.01fF
C549 VDD.n383 GND 0.02fF
C550 VDD.n384 GND 0.03fF
C551 VDD.n385 GND 0.06fF
C552 VDD.n386 GND 0.25fF
C553 VDD.n387 GND 0.01fF
C554 VDD.n388 GND 0.01fF
C555 VDD.n389 GND 0.02fF
C556 VDD.n390 GND 0.16fF
C557 VDD.n391 GND 0.01fF
C558 VDD.n392 GND 0.02fF
C559 VDD.n393 GND 0.02fF
C560 VDD.n394 GND 0.14fF
C561 VDD.n395 GND 0.01fF
C562 VDD.n396 GND 0.02fF
C563 VDD.n397 GND 0.03fF
C564 VDD.n398 GND 0.08fF
C565 VDD.n399 GND 0.05fF
C566 VDD.n400 GND 0.01fF
C567 VDD.n401 GND 0.02fF
C568 VDD.n402 GND 0.03fF
C569 VDD.n403 GND 0.17fF
C570 VDD.n404 GND 0.01fF
C571 VDD.n405 GND 0.02fF
C572 VDD.n406 GND 0.02fF
C573 VDD.n407 GND 0.06fF
C574 VDD.n408 GND 0.24fF
C575 VDD.n409 GND 0.01fF
C576 VDD.n410 GND 0.01fF
C577 VDD.n411 GND 0.02fF
C578 VDD.n412 GND 0.26fF
C579 VDD.n413 GND 0