magic
tech sky130A
magscale 1 2
timestamp 1645652543
<< poly >>
rect -33 17 33 27
rect -33 -17 -17 17
rect 17 -17 33 17
rect -33 -27 33 -17
<< polycont >>
rect -17 -17 17 17
<< locali >>
rect -33 -17 -17 17
rect 17 -17 33 17
<< end >>
