* SPICE3 file created from AND2X2.ext - technology: sky130A

.subckt AND2X2 A B Y VSS VDD
M1000 VSS B a_36_101# VSS nshort w=3u l=0.15u
+  ad=1.23735p pd=9.4u as=1.85625p ps=12.67u
M1001 Y a_128_200# VDD VDD pshort w=3u l=0.15u
+  ad=0.87p pd=6.58u as=4.29p ps=32.86u
M1002 Y a_128_200# VSS VSS nshort w=3u l=0.15u
+  ad=0.1588p pd=1.5u as=0p ps=0u
M1003 VDD B a_128_200# VDD pshort w=3u l=0.15u
+  ad=0p pd=0u as=1.74p ps=13.16u
M1004 a_128_200# A VDD VDD pshort w=3u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 VDD a_128_200# Y VDD pshort w=3u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_128_200# A a_36_101# VSS nshort w=3u l=0.15u
+  ad=0.1588p pd=1.5u as=0p ps=0u
M1007 a_128_200# B VDD VDD pshort w=3u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 VDD A a_128_200# VDD pshort w=3u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
.ends
