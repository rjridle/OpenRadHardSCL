magic
tech sky130A
magscale 1 2
timestamp 1649544039
<< nwell >>
rect -84 832 3414 1575
<< nmos >>
rect 168 316 198 377
tri 198 316 214 332 sw
rect 362 324 392 377
tri 392 324 408 340 sw
rect 168 286 274 316
tri 274 286 304 316 sw
rect 362 294 468 324
tri 468 294 498 324 sw
rect 168 185 198 286
tri 198 270 214 286 nw
tri 258 270 274 286 ne
tri 198 185 214 201 sw
tri 258 185 274 201 se
rect 274 185 304 286
rect 362 193 392 294
tri 392 278 408 294 nw
tri 452 278 468 294 ne
tri 392 193 408 209 sw
tri 452 193 468 209 se
rect 468 193 498 294
tri 168 155 198 185 ne
rect 198 155 274 185
tri 274 155 304 185 nw
tri 362 163 392 193 ne
rect 392 163 468 193
tri 468 163 498 193 nw
rect 821 324 851 377
tri 851 324 867 340 sw
rect 821 294 927 324
tri 927 294 957 324 sw
rect 821 193 851 294
tri 851 278 867 294 nw
tri 911 278 927 294 ne
tri 851 193 867 209 sw
tri 911 193 927 209 se
rect 927 193 957 294
tri 821 163 851 193 ne
rect 851 163 927 193
tri 927 163 957 193 nw
rect 1265 324 1295 377
tri 1295 324 1311 340 sw
rect 1265 294 1371 324
tri 1371 294 1401 324 sw
rect 1265 193 1295 294
tri 1295 278 1311 294 nw
tri 1355 278 1371 294 ne
tri 1295 193 1311 209 sw
tri 1355 193 1371 209 se
rect 1371 193 1401 294
tri 1265 163 1295 193 ne
rect 1295 163 1371 193
tri 1371 163 1401 193 nw
rect 1722 316 1752 377
tri 1752 316 1768 332 sw
rect 1916 324 1946 377
tri 1946 324 1962 340 sw
rect 1722 286 1828 316
tri 1828 286 1858 316 sw
rect 1916 294 2022 324
tri 2022 294 2052 324 sw
rect 1722 185 1752 286
tri 1752 270 1768 286 nw
tri 1812 270 1828 286 ne
tri 1752 185 1768 201 sw
tri 1812 185 1828 201 se
rect 1828 185 1858 286
rect 1916 193 1946 294
tri 1946 278 1962 294 nw
tri 2006 278 2022 294 ne
tri 1946 193 1962 209 sw
tri 2006 193 2022 209 se
rect 2022 193 2052 294
tri 1722 155 1752 185 ne
rect 1752 155 1828 185
tri 1828 155 1858 185 nw
tri 1916 163 1946 193 ne
rect 1946 163 2022 193
tri 2022 163 2052 193 nw
rect 2388 316 2418 377
tri 2418 316 2434 332 sw
rect 2582 324 2612 377
tri 2612 324 2628 340 sw
rect 2388 286 2494 316
tri 2494 286 2524 316 sw
rect 2582 294 2688 324
tri 2688 294 2718 324 sw
rect 2388 185 2418 286
tri 2418 270 2434 286 nw
tri 2478 270 2494 286 ne
tri 2418 185 2434 201 sw
tri 2478 185 2494 201 se
rect 2494 185 2524 286
rect 2582 193 2612 294
tri 2612 278 2628 294 nw
tri 2672 278 2688 294 ne
tri 2612 193 2628 209 sw
tri 2672 193 2688 209 se
rect 2688 193 2718 294
tri 2388 155 2418 185 ne
rect 2418 155 2494 185
tri 2494 155 2524 185 nw
tri 2582 163 2612 193 ne
rect 2612 163 2688 193
tri 2688 163 2718 193 nw
tri 3129 324 3145 340 se
rect 3145 324 3175 377
tri 3039 294 3069 324 se
rect 3069 294 3175 324
rect 3039 193 3069 294
tri 3069 278 3085 294 nw
tri 3129 278 3145 294 ne
tri 3069 193 3085 209 sw
tri 3129 193 3145 209 se
rect 3145 193 3175 294
tri 3039 163 3069 193 ne
rect 3069 163 3145 193
tri 3145 163 3175 193 nw
<< pmos >>
rect 187 1050 217 1450
rect 275 1050 305 1450
rect 363 1050 393 1450
rect 451 1050 481 1450
rect 829 1050 859 1450
rect 917 1050 947 1450
rect 1273 1050 1303 1450
rect 1361 1050 1391 1450
rect 1741 1051 1771 1451
rect 1829 1051 1859 1451
rect 1917 1051 1947 1451
rect 2005 1051 2035 1451
rect 2407 1051 2437 1451
rect 2495 1051 2525 1451
rect 2583 1051 2613 1451
rect 2671 1051 2701 1451
rect 3049 1050 3079 1450
rect 3137 1050 3167 1450
<< ndiff >>
rect 112 361 168 377
rect 112 327 122 361
rect 156 327 168 361
rect 112 289 168 327
rect 198 361 362 377
rect 198 332 219 361
tri 198 316 214 332 ne
rect 214 327 219 332
rect 253 327 316 361
rect 350 327 362 361
rect 214 316 362 327
rect 392 340 554 377
tri 392 324 408 340 ne
rect 408 324 554 340
rect 112 255 122 289
rect 156 255 168 289
tri 274 286 304 316 ne
rect 304 289 362 316
tri 468 294 498 324 ne
rect 112 221 168 255
rect 112 187 122 221
rect 156 187 168 221
rect 112 155 168 187
tri 198 270 214 286 se
rect 214 270 258 286
tri 258 270 274 286 sw
rect 198 236 274 270
rect 198 202 219 236
rect 253 202 274 236
rect 198 201 274 202
tri 198 185 214 201 ne
rect 214 185 258 201
tri 258 185 274 201 nw
rect 304 255 316 289
rect 350 255 362 289
rect 304 221 362 255
rect 304 187 316 221
rect 350 187 362 221
tri 392 278 408 294 se
rect 408 278 452 294
tri 452 278 468 294 sw
rect 392 245 468 278
rect 392 211 413 245
rect 447 211 468 245
rect 392 209 468 211
tri 392 193 408 209 ne
rect 408 193 452 209
tri 452 193 468 209 nw
rect 498 289 554 324
rect 498 255 510 289
rect 544 255 554 289
rect 498 221 554 255
tri 168 155 198 185 sw
tri 274 155 304 185 se
rect 304 163 362 187
tri 362 163 392 193 sw
tri 468 163 498 193 se
rect 498 187 510 221
rect 544 187 554 221
rect 498 163 554 187
rect 304 155 554 163
rect 112 151 554 155
rect 112 117 122 151
rect 156 117 316 151
rect 350 117 413 151
rect 447 117 510 151
rect 544 117 554 151
rect 112 101 554 117
rect 765 361 821 377
rect 765 327 775 361
rect 809 327 821 361
rect 765 289 821 327
rect 851 361 1011 377
rect 851 340 969 361
tri 851 324 867 340 ne
rect 867 327 969 340
rect 1003 327 1011 361
rect 867 324 1011 327
tri 927 294 957 324 ne
rect 765 255 775 289
rect 809 255 821 289
rect 765 221 821 255
rect 765 187 775 221
rect 809 187 821 221
tri 851 278 867 294 se
rect 867 278 911 294
tri 911 278 927 294 sw
rect 851 245 927 278
rect 851 211 871 245
rect 905 211 927 245
rect 851 209 927 211
tri 851 193 867 209 ne
rect 867 193 911 209
tri 911 193 927 209 nw
rect 957 289 1011 324
rect 957 255 969 289
rect 1003 255 1011 289
rect 957 221 1011 255
rect 765 163 821 187
tri 821 163 851 193 sw
tri 927 163 957 193 se
rect 957 187 969 221
rect 1003 187 1011 221
rect 957 163 1011 187
rect 765 151 1011 163
rect 765 117 775 151
rect 809 117 871 151
rect 905 117 969 151
rect 1003 117 1011 151
rect 765 101 1011 117
rect 1209 361 1265 377
rect 1209 327 1219 361
rect 1253 327 1265 361
rect 1209 289 1265 327
rect 1295 361 1455 377
rect 1295 340 1413 361
tri 1295 324 1311 340 ne
rect 1311 327 1413 340
rect 1447 327 1455 361
rect 1311 324 1455 327
tri 1371 294 1401 324 ne
rect 1209 255 1219 289
rect 1253 255 1265 289
rect 1209 221 1265 255
rect 1209 187 1219 221
rect 1253 187 1265 221
tri 1295 278 1311 294 se
rect 1311 278 1355 294
tri 1355 278 1371 294 sw
rect 1295 245 1371 278
rect 1295 211 1315 245
rect 1349 211 1371 245
rect 1295 209 1371 211
tri 1295 193 1311 209 ne
rect 1311 193 1355 209
tri 1355 193 1371 209 nw
rect 1401 289 1455 324
rect 1401 255 1413 289
rect 1447 255 1455 289
rect 1401 221 1455 255
rect 1209 163 1265 187
tri 1265 163 1295 193 sw
tri 1371 163 1401 193 se
rect 1401 187 1413 221
rect 1447 187 1455 221
rect 1401 163 1455 187
rect 1209 151 1455 163
rect 1209 117 1219 151
rect 1253 117 1315 151
rect 1349 117 1413 151
rect 1447 117 1455 151
rect 1209 101 1455 117
rect 1666 361 1722 377
rect 1666 327 1676 361
rect 1710 327 1722 361
rect 1666 289 1722 327
rect 1752 361 1916 377
rect 1752 332 1773 361
tri 1752 316 1768 332 ne
rect 1768 327 1773 332
rect 1807 327 1870 361
rect 1904 327 1916 361
rect 1768 316 1916 327
rect 1946 340 2108 377
tri 1946 324 1962 340 ne
rect 1962 324 2108 340
rect 1666 255 1676 289
rect 1710 255 1722 289
tri 1828 286 1858 316 ne
rect 1858 289 1916 316
tri 2022 294 2052 324 ne
rect 1666 221 1722 255
rect 1666 187 1676 221
rect 1710 187 1722 221
rect 1666 155 1722 187
tri 1752 270 1768 286 se
rect 1768 270 1812 286
tri 1812 270 1828 286 sw
rect 1752 236 1828 270
rect 1752 202 1773 236
rect 1807 202 1828 236
rect 1752 201 1828 202
tri 1752 185 1768 201 ne
rect 1768 185 1812 201
tri 1812 185 1828 201 nw
rect 1858 255 1870 289
rect 1904 255 1916 289
rect 1858 221 1916 255
rect 1858 187 1870 221
rect 1904 187 1916 221
tri 1946 278 1962 294 se
rect 1962 278 2006 294
tri 2006 278 2022 294 sw
rect 1946 245 2022 278
rect 1946 211 1967 245
rect 2001 211 2022 245
rect 1946 209 2022 211
tri 1946 193 1962 209 ne
rect 1962 193 2006 209
tri 2006 193 2022 209 nw
rect 2052 289 2108 324
rect 2052 255 2064 289
rect 2098 255 2108 289
rect 2052 221 2108 255
tri 1722 155 1752 185 sw
tri 1828 155 1858 185 se
rect 1858 163 1916 187
tri 1916 163 1946 193 sw
tri 2022 163 2052 193 se
rect 2052 187 2064 221
rect 2098 187 2108 221
rect 2052 163 2108 187
rect 1858 155 2108 163
rect 1666 151 2108 155
rect 1666 117 1676 151
rect 1710 117 1870 151
rect 1904 117 1967 151
rect 2001 117 2064 151
rect 2098 117 2108 151
rect 1666 101 2108 117
rect 2332 361 2388 377
rect 2332 327 2342 361
rect 2376 327 2388 361
rect 2332 289 2388 327
rect 2418 361 2582 377
rect 2418 332 2439 361
tri 2418 316 2434 332 ne
rect 2434 327 2439 332
rect 2473 327 2536 361
rect 2570 327 2582 361
rect 2434 316 2582 327
rect 2612 340 2774 377
tri 2612 324 2628 340 ne
rect 2628 324 2774 340
rect 2332 255 2342 289
rect 2376 255 2388 289
tri 2494 286 2524 316 ne
rect 2524 289 2582 316
tri 2688 294 2718 324 ne
rect 2332 221 2388 255
rect 2332 187 2342 221
rect 2376 187 2388 221
rect 2332 155 2388 187
tri 2418 270 2434 286 se
rect 2434 270 2478 286
tri 2478 270 2494 286 sw
rect 2418 236 2494 270
rect 2418 202 2439 236
rect 2473 202 2494 236
rect 2418 201 2494 202
tri 2418 185 2434 201 ne
rect 2434 185 2478 201
tri 2478 185 2494 201 nw
rect 2524 255 2536 289
rect 2570 255 2582 289
rect 2524 221 2582 255
rect 2524 187 2536 221
rect 2570 187 2582 221
tri 2612 278 2628 294 se
rect 2628 278 2672 294
tri 2672 278 2688 294 sw
rect 2612 245 2688 278
rect 2612 211 2633 245
rect 2667 211 2688 245
rect 2612 209 2688 211
tri 2612 193 2628 209 ne
rect 2628 193 2672 209
tri 2672 193 2688 209 nw
rect 2718 289 2774 324
rect 2718 255 2730 289
rect 2764 255 2774 289
rect 2718 221 2774 255
tri 2388 155 2418 185 sw
tri 2494 155 2524 185 se
rect 2524 163 2582 187
tri 2582 163 2612 193 sw
tri 2688 163 2718 193 se
rect 2718 187 2730 221
rect 2764 187 2774 221
rect 2718 163 2774 187
rect 2524 155 2774 163
rect 2332 151 2774 155
rect 2332 117 2342 151
rect 2376 117 2536 151
rect 2570 117 2633 151
rect 2667 117 2730 151
rect 2764 117 2774 151
rect 2332 101 2774 117
rect 2985 361 3145 377
rect 2985 327 2993 361
rect 3027 340 3145 361
rect 3027 327 3129 340
rect 2985 324 3129 327
tri 3129 324 3145 340 nw
rect 3175 361 3231 377
rect 3175 327 3187 361
rect 3221 327 3231 361
rect 2985 289 3039 324
tri 3039 294 3069 324 nw
rect 2985 255 2993 289
rect 3027 255 3039 289
rect 2985 221 3039 255
rect 2985 187 2993 221
rect 3027 187 3039 221
tri 3069 278 3085 294 se
rect 3085 278 3129 294
tri 3129 278 3145 294 sw
rect 3069 245 3145 278
rect 3069 211 3091 245
rect 3125 211 3145 245
rect 3069 209 3145 211
tri 3069 193 3085 209 ne
rect 3085 193 3129 209
tri 3129 193 3145 209 nw
rect 3175 289 3231 327
rect 3175 255 3187 289
rect 3221 255 3231 289
rect 3175 221 3231 255
rect 2985 163 3039 187
tri 3039 163 3069 193 sw
tri 3145 163 3175 193 se
rect 3175 187 3187 221
rect 3221 187 3231 221
rect 3175 163 3231 187
rect 2985 151 3231 163
rect 2985 117 2993 151
rect 3027 117 3091 151
rect 3125 117 3187 151
rect 3221 117 3231 151
rect 2985 101 3231 117
<< pdiff >>
rect 131 1412 187 1450
rect 131 1378 141 1412
rect 175 1378 187 1412
rect 131 1344 187 1378
rect 131 1310 141 1344
rect 175 1310 187 1344
rect 131 1276 187 1310
rect 131 1242 141 1276
rect 175 1242 187 1276
rect 131 1208 187 1242
rect 131 1174 141 1208
rect 175 1174 187 1208
rect 131 1139 187 1174
rect 131 1105 141 1139
rect 175 1105 187 1139
rect 131 1050 187 1105
rect 217 1412 275 1450
rect 217 1378 229 1412
rect 263 1378 275 1412
rect 217 1344 275 1378
rect 217 1310 229 1344
rect 263 1310 275 1344
rect 217 1276 275 1310
rect 217 1242 229 1276
rect 263 1242 275 1276
rect 217 1208 275 1242
rect 217 1174 229 1208
rect 263 1174 275 1208
rect 217 1139 275 1174
rect 217 1105 229 1139
rect 263 1105 275 1139
rect 217 1050 275 1105
rect 305 1412 363 1450
rect 305 1378 317 1412
rect 351 1378 363 1412
rect 305 1344 363 1378
rect 305 1310 317 1344
rect 351 1310 363 1344
rect 305 1276 363 1310
rect 305 1242 317 1276
rect 351 1242 363 1276
rect 305 1208 363 1242
rect 305 1174 317 1208
rect 351 1174 363 1208
rect 305 1050 363 1174
rect 393 1412 451 1450
rect 393 1378 405 1412
rect 439 1378 451 1412
rect 393 1344 451 1378
rect 393 1310 405 1344
rect 439 1310 451 1344
rect 393 1276 451 1310
rect 393 1242 405 1276
rect 439 1242 451 1276
rect 393 1208 451 1242
rect 393 1174 405 1208
rect 439 1174 451 1208
rect 393 1139 451 1174
rect 393 1105 405 1139
rect 439 1105 451 1139
rect 393 1050 451 1105
rect 481 1412 535 1450
rect 481 1378 493 1412
rect 527 1378 535 1412
rect 481 1344 535 1378
rect 481 1310 493 1344
rect 527 1310 535 1344
rect 481 1276 535 1310
rect 481 1242 493 1276
rect 527 1242 535 1276
rect 481 1208 535 1242
rect 481 1174 493 1208
rect 527 1174 535 1208
rect 481 1050 535 1174
rect 773 1412 829 1450
rect 773 1378 783 1412
rect 817 1378 829 1412
rect 773 1344 829 1378
rect 773 1310 783 1344
rect 817 1310 829 1344
rect 773 1276 829 1310
rect 773 1242 783 1276
rect 817 1242 829 1276
rect 773 1208 829 1242
rect 773 1174 783 1208
rect 817 1174 829 1208
rect 773 1139 829 1174
rect 773 1105 783 1139
rect 817 1105 829 1139
rect 773 1050 829 1105
rect 859 1412 917 1450
rect 859 1378 871 1412
rect 905 1378 917 1412
rect 859 1344 917 1378
rect 859 1310 871 1344
rect 905 1310 917 1344
rect 859 1276 917 1310
rect 859 1242 871 1276
rect 905 1242 917 1276
rect 859 1208 917 1242
rect 859 1174 871 1208
rect 905 1174 917 1208
rect 859 1139 917 1174
rect 859 1105 871 1139
rect 905 1105 917 1139
rect 859 1050 917 1105
rect 947 1412 1001 1450
rect 947 1378 959 1412
rect 993 1378 1001 1412
rect 947 1344 1001 1378
rect 947 1310 959 1344
rect 993 1310 1001 1344
rect 947 1276 1001 1310
rect 947 1242 959 1276
rect 993 1242 1001 1276
rect 947 1208 1001 1242
rect 947 1174 959 1208
rect 993 1174 1001 1208
rect 947 1139 1001 1174
rect 947 1105 959 1139
rect 993 1105 1001 1139
rect 947 1050 1001 1105
rect 1217 1412 1273 1450
rect 1217 1378 1227 1412
rect 1261 1378 1273 1412
rect 1217 1344 1273 1378
rect 1217 1310 1227 1344
rect 1261 1310 1273 1344
rect 1217 1276 1273 1310
rect 1217 1242 1227 1276
rect 1261 1242 1273 1276
rect 1217 1208 1273 1242
rect 1217 1174 1227 1208
rect 1261 1174 1273 1208
rect 1217 1139 1273 1174
rect 1217 1105 1227 1139
rect 1261 1105 1273 1139
rect 1217 1050 1273 1105
rect 1303 1412 1361 1450
rect 1303 1378 1315 1412
rect 1349 1378 1361 1412
rect 1303 1344 1361 1378
rect 1303 1310 1315 1344
rect 1349 1310 1361 1344
rect 1303 1276 1361 1310
rect 1303 1242 1315 1276
rect 1349 1242 1361 1276
rect 1303 1208 1361 1242
rect 1303 1174 1315 1208
rect 1349 1174 1361 1208
rect 1303 1139 1361 1174
rect 1303 1105 1315 1139
rect 1349 1105 1361 1139
rect 1303 1050 1361 1105
rect 1391 1412 1445 1450
rect 1391 1378 1403 1412
rect 1437 1378 1445 1412
rect 1391 1344 1445 1378
rect 1391 1310 1403 1344
rect 1437 1310 1445 1344
rect 1391 1276 1445 1310
rect 1391 1242 1403 1276
rect 1437 1242 1445 1276
rect 1391 1208 1445 1242
rect 1391 1174 1403 1208
rect 1437 1174 1445 1208
rect 1391 1139 1445 1174
rect 1391 1105 1403 1139
rect 1437 1105 1445 1139
rect 1391 1050 1445 1105
rect 1685 1411 1741 1451
rect 1685 1377 1695 1411
rect 1729 1377 1741 1411
rect 1685 1343 1741 1377
rect 1685 1309 1695 1343
rect 1729 1309 1741 1343
rect 1685 1275 1741 1309
rect 1685 1241 1695 1275
rect 1729 1241 1741 1275
rect 1685 1207 1741 1241
rect 1685 1173 1695 1207
rect 1729 1173 1741 1207
rect 1685 1139 1741 1173
rect 1685 1105 1695 1139
rect 1729 1105 1741 1139
rect 1685 1051 1741 1105
rect 1771 1343 1829 1451
rect 1771 1309 1783 1343
rect 1817 1309 1829 1343
rect 1771 1275 1829 1309
rect 1771 1241 1783 1275
rect 1817 1241 1829 1275
rect 1771 1207 1829 1241
rect 1771 1173 1783 1207
rect 1817 1173 1829 1207
rect 1771 1051 1829 1173
rect 1859 1411 1917 1451
rect 1859 1377 1871 1411
rect 1905 1377 1917 1411
rect 1859 1343 1917 1377
rect 1859 1309 1871 1343
rect 1905 1309 1917 1343
rect 1859 1275 1917 1309
rect 1859 1241 1871 1275
rect 1905 1241 1917 1275
rect 1859 1207 1917 1241
rect 1859 1173 1871 1207
rect 1905 1173 1917 1207
rect 1859 1139 1917 1173
rect 1859 1105 1871 1139
rect 1905 1105 1917 1139
rect 1859 1051 1917 1105
rect 1947 1343 2005 1451
rect 1947 1309 1959 1343
rect 1993 1309 2005 1343
rect 1947 1275 2005 1309
rect 1947 1241 1959 1275
rect 1993 1241 2005 1275
rect 1947 1207 2005 1241
rect 1947 1173 1959 1207
rect 1993 1173 2005 1207
rect 1947 1139 2005 1173
rect 1947 1105 1959 1139
rect 1993 1105 2005 1139
rect 1947 1051 2005 1105
rect 2035 1411 2089 1451
rect 2035 1377 2047 1411
rect 2081 1377 2089 1411
rect 2035 1343 2089 1377
rect 2035 1309 2047 1343
rect 2081 1309 2089 1343
rect 2035 1275 2089 1309
rect 2035 1241 2047 1275
rect 2081 1241 2089 1275
rect 2035 1207 2089 1241
rect 2035 1173 2047 1207
rect 2081 1173 2089 1207
rect 2035 1051 2089 1173
rect 2351 1411 2407 1451
rect 2351 1377 2361 1411
rect 2395 1377 2407 1411
rect 2351 1343 2407 1377
rect 2351 1309 2361 1343
rect 2395 1309 2407 1343
rect 2351 1275 2407 1309
rect 2351 1241 2361 1275
rect 2395 1241 2407 1275
rect 2351 1207 2407 1241
rect 2351 1173 2361 1207
rect 2395 1173 2407 1207
rect 2351 1139 2407 1173
rect 2351 1105 2361 1139
rect 2395 1105 2407 1139
rect 2351 1051 2407 1105
rect 2437 1343 2495 1451
rect 2437 1309 2449 1343
rect 2483 1309 2495 1343
rect 2437 1275 2495 1309
rect 2437 1241 2449 1275
rect 2483 1241 2495 1275
rect 2437 1207 2495 1241
rect 2437 1173 2449 1207
rect 2483 1173 2495 1207
rect 2437 1051 2495 1173
rect 2525 1411 2583 1451
rect 2525 1377 2537 1411
rect 2571 1377 2583 1411
rect 2525 1343 2583 1377
rect 2525 1309 2537 1343
rect 2571 1309 2583 1343
rect 2525 1275 2583 1309
rect 2525 1241 2537 1275
rect 2571 1241 2583 1275
rect 2525 1207 2583 1241
rect 2525 1173 2537 1207
rect 2571 1173 2583 1207
rect 2525 1139 2583 1173
rect 2525 1105 2537 1139
rect 2571 1105 2583 1139
rect 2525 1051 2583 1105
rect 2613 1343 2671 1451
rect 2613 1309 2625 1343
rect 2659 1309 2671 1343
rect 2613 1275 2671 1309
rect 2613 1241 2625 1275
rect 2659 1241 2671 1275
rect 2613 1207 2671 1241
rect 2613 1173 2625 1207
rect 2659 1173 2671 1207
rect 2613 1139 2671 1173
rect 2613 1105 2625 1139
rect 2659 1105 2671 1139
rect 2613 1051 2671 1105
rect 2701 1411 2755 1451
rect 2701 1377 2713 1411
rect 2747 1377 2755 1411
rect 2701 1343 2755 1377
rect 2701 1309 2713 1343
rect 2747 1309 2755 1343
rect 2701 1275 2755 1309
rect 2701 1241 2713 1275
rect 2747 1241 2755 1275
rect 2701 1207 2755 1241
rect 2701 1173 2713 1207
rect 2747 1173 2755 1207
rect 2701 1051 2755 1173
rect 2995 1412 3049 1450
rect 2995 1378 3003 1412
rect 3037 1378 3049 1412
rect 2995 1344 3049 1378
rect 2995 1310 3003 1344
rect 3037 1310 3049 1344
rect 2995 1276 3049 1310
rect 2995 1242 3003 1276
rect 3037 1242 3049 1276
rect 2995 1208 3049 1242
rect 2995 1174 3003 1208
rect 3037 1174 3049 1208
rect 2995 1139 3049 1174
rect 2995 1105 3003 1139
rect 3037 1105 3049 1139
rect 2995 1050 3049 1105
rect 3079 1412 3137 1450
rect 3079 1378 3091 1412
rect 3125 1378 3137 1412
rect 3079 1344 3137 1378
rect 3079 1310 3091 1344
rect 3125 1310 3137 1344
rect 3079 1276 3137 1310
rect 3079 1242 3091 1276
rect 3125 1242 3137 1276
rect 3079 1208 3137 1242
rect 3079 1174 3091 1208
rect 3125 1174 3137 1208
rect 3079 1139 3137 1174
rect 3079 1105 3091 1139
rect 3125 1105 3137 1139
rect 3079 1050 3137 1105
rect 3167 1412 3223 1450
rect 3167 1378 3179 1412
rect 3213 1378 3223 1412
rect 3167 1344 3223 1378
rect 3167 1310 3179 1344
rect 3213 1310 3223 1344
rect 3167 1276 3223 1310
rect 3167 1242 3179 1276
rect 3213 1242 3223 1276
rect 3167 1208 3223 1242
rect 3167 1174 3179 1208
rect 3213 1174 3223 1208
rect 3167 1139 3223 1174
rect 3167 1105 3179 1139
rect 3213 1105 3223 1139
rect 3167 1050 3223 1105
<< ndiffc >>
rect 122 327 156 361
rect 219 327 253 361
rect 316 327 350 361
rect 122 255 156 289
rect 122 187 156 221
rect 219 202 253 236
rect 316 255 350 289
rect 316 187 350 221
rect 413 211 447 245
rect 510 255 544 289
rect 510 187 544 221
rect 122 117 156 151
rect 316 117 350 151
rect 413 117 447 151
rect 510 117 544 151
rect 775 327 809 361
rect 969 327 1003 361
rect 775 255 809 289
rect 775 187 809 221
rect 871 211 905 245
rect 969 255 1003 289
rect 969 187 1003 221
rect 775 117 809 151
rect 871 117 905 151
rect 969 117 1003 151
rect 1219 327 1253 361
rect 1413 327 1447 361
rect 1219 255 1253 289
rect 1219 187 1253 221
rect 1315 211 1349 245
rect 1413 255 1447 289
rect 1413 187 1447 221
rect 1219 117 1253 151
rect 1315 117 1349 151
rect 1413 117 1447 151
rect 1676 327 1710 361
rect 1773 327 1807 361
rect 1870 327 1904 361
rect 1676 255 1710 289
rect 1676 187 1710 221
rect 1773 202 1807 236
rect 1870 255 1904 289
rect 1870 187 1904 221
rect 1967 211 2001 245
rect 2064 255 2098 289
rect 2064 187 2098 221
rect 1676 117 1710 151
rect 1870 117 1904 151
rect 1967 117 2001 151
rect 2064 117 2098 151
rect 2342 327 2376 361
rect 2439 327 2473 361
rect 2536 327 2570 361
rect 2342 255 2376 289
rect 2342 187 2376 221
rect 2439 202 2473 236
rect 2536 255 2570 289
rect 2536 187 2570 221
rect 2633 211 2667 245
rect 2730 255 2764 289
rect 2730 187 2764 221
rect 2342 117 2376 151
rect 2536 117 2570 151
rect 2633 117 2667 151
rect 2730 117 2764 151
rect 2993 327 3027 361
rect 3187 327 3221 361
rect 2993 255 3027 289
rect 2993 187 3027 221
rect 3091 211 3125 245
rect 3187 255 3221 289
rect 3187 187 3221 221
rect 2993 117 3027 151
rect 3091 117 3125 151
rect 3187 117 3221 151
<< pdiffc >>
rect 141 1378 175 1412
rect 141 1310 175 1344
rect 141 1242 175 1276
rect 141 1174 175 1208
rect 141 1105 175 1139
rect 229 1378 263 1412
rect 229 1310 263 1344
rect 229 1242 263 1276
rect 229 1174 263 1208
rect 229 1105 263 1139
rect 317 1378 351 1412
rect 317 1310 351 1344
rect 317 1242 351 1276
rect 317 1174 351 1208
rect 405 1378 439 1412
rect 405 1310 439 1344
rect 405 1242 439 1276
rect 405 1174 439 1208
rect 405 1105 439 1139
rect 493 1378 527 1412
rect 493 1310 527 1344
rect 493 1242 527 1276
rect 493 1174 527 1208
rect 783 1378 817 1412
rect 783 1310 817 1344
rect 783 1242 817 1276
rect 783 1174 817 1208
rect 783 1105 817 1139
rect 871 1378 905 1412
rect 871 1310 905 1344
rect 871 1242 905 1276
rect 871 1174 905 1208
rect 871 1105 905 1139
rect 959 1378 993 1412
rect 959 1310 993 1344
rect 959 1242 993 1276
rect 959 1174 993 1208
rect 959 1105 993 1139
rect 1227 1378 1261 1412
rect 1227 1310 1261 1344
rect 1227 1242 1261 1276
rect 1227 1174 1261 1208
rect 1227 1105 1261 1139
rect 1315 1378 1349 1412
rect 1315 1310 1349 1344
rect 1315 1242 1349 1276
rect 1315 1174 1349 1208
rect 1315 1105 1349 1139
rect 1403 1378 1437 1412
rect 1403 1310 1437 1344
rect 1403 1242 1437 1276
rect 1403 1174 1437 1208
rect 1403 1105 1437 1139
rect 1695 1377 1729 1411
rect 1695 1309 1729 1343
rect 1695 1241 1729 1275
rect 1695 1173 1729 1207
rect 1695 1105 1729 1139
rect 1783 1309 1817 1343
rect 1783 1241 1817 1275
rect 1783 1173 1817 1207
rect 1871 1377 1905 1411
rect 1871 1309 1905 1343
rect 1871 1241 1905 1275
rect 1871 1173 1905 1207
rect 1871 1105 1905 1139
rect 1959 1309 1993 1343
rect 1959 1241 1993 1275
rect 1959 1173 1993 1207
rect 1959 1105 1993 1139
rect 2047 1377 2081 1411
rect 2047 1309 2081 1343
rect 2047 1241 2081 1275
rect 2047 1173 2081 1207
rect 2361 1377 2395 1411
rect 2361 1309 2395 1343
rect 2361 1241 2395 1275
rect 2361 1173 2395 1207
rect 2361 1105 2395 1139
rect 2449 1309 2483 1343
rect 2449 1241 2483 1275
rect 2449 1173 2483 1207
rect 2537 1377 2571 1411
rect 2537 1309 2571 1343
rect 2537 1241 2571 1275
rect 2537 1173 2571 1207
rect 2537 1105 2571 1139
rect 2625 1309 2659 1343
rect 2625 1241 2659 1275
rect 2625 1173 2659 1207
rect 2625 1105 2659 1139
rect 2713 1377 2747 1411
rect 2713 1309 2747 1343
rect 2713 1241 2747 1275
rect 2713 1173 2747 1207
rect 3003 1378 3037 1412
rect 3003 1310 3037 1344
rect 3003 1242 3037 1276
rect 3003 1174 3037 1208
rect 3003 1105 3037 1139
rect 3091 1378 3125 1412
rect 3091 1310 3125 1344
rect 3091 1242 3125 1276
rect 3091 1174 3125 1208
rect 3091 1105 3125 1139
rect 3179 1378 3213 1412
rect 3179 1310 3213 1344
rect 3179 1242 3213 1276
rect 3179 1174 3213 1208
rect 3179 1105 3213 1139
<< psubdiff >>
rect -31 546 3361 572
rect -31 512 -17 546
rect 17 512 649 546
rect 683 512 1093 546
rect 1127 512 1537 546
rect 1571 512 2203 546
rect 2237 512 2869 546
rect 2903 512 3313 546
rect 3347 512 3361 546
rect -31 510 3361 512
rect -31 474 31 510
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect -31 368 -17 402
rect 17 368 31 402
rect 635 474 697 510
rect 635 440 649 474
rect 683 440 697 474
rect 635 402 697 440
rect 1079 474 1141 510
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect 635 368 649 402
rect 683 368 697 402
rect 1079 440 1093 474
rect 1127 440 1141 474
rect 1079 402 1141 440
rect 1523 474 1585 510
rect 635 330 697 368
rect 635 296 649 330
rect 683 296 697 330
rect 635 258 697 296
rect 635 224 649 258
rect 683 224 697 258
rect 635 186 697 224
rect 635 152 649 186
rect 683 152 697 186
rect 635 114 697 152
rect -31 47 31 80
rect 635 80 649 114
rect 683 80 697 114
rect 1079 368 1093 402
rect 1127 368 1141 402
rect 1523 440 1537 474
rect 1571 440 1585 474
rect 1523 402 1585 440
rect 1079 330 1141 368
rect 1079 296 1093 330
rect 1127 296 1141 330
rect 1079 258 1141 296
rect 1079 224 1093 258
rect 1127 224 1141 258
rect 1079 186 1141 224
rect 1079 152 1093 186
rect 1127 152 1141 186
rect 1079 114 1141 152
rect 635 47 697 80
rect 1079 80 1093 114
rect 1127 80 1141 114
rect 1523 368 1537 402
rect 1571 368 1585 402
rect 2189 474 2251 510
rect 2189 440 2203 474
rect 2237 440 2251 474
rect 2189 402 2251 440
rect 1523 330 1585 368
rect 1523 296 1537 330
rect 1571 296 1585 330
rect 1523 258 1585 296
rect 1523 224 1537 258
rect 1571 224 1585 258
rect 1523 186 1585 224
rect 1523 152 1537 186
rect 1571 152 1585 186
rect 1523 114 1585 152
rect 1079 47 1141 80
rect 1523 80 1537 114
rect 1571 80 1585 114
rect 2189 368 2203 402
rect 2237 368 2251 402
rect 2855 474 2917 510
rect 2855 440 2869 474
rect 2903 440 2917 474
rect 2855 402 2917 440
rect 2189 330 2251 368
rect 2189 296 2203 330
rect 2237 296 2251 330
rect 2189 258 2251 296
rect 2189 224 2203 258
rect 2237 224 2251 258
rect 2189 186 2251 224
rect 2189 152 2203 186
rect 2237 152 2251 186
rect 2189 114 2251 152
rect 1523 47 1585 80
rect 2189 80 2203 114
rect 2237 80 2251 114
rect 2855 368 2869 402
rect 2903 368 2917 402
rect 3299 474 3361 510
rect 3299 440 3313 474
rect 3347 440 3361 474
rect 3299 402 3361 440
rect 2855 330 2917 368
rect 2855 296 2869 330
rect 2903 296 2917 330
rect 2855 258 2917 296
rect 2855 224 2869 258
rect 2903 224 2917 258
rect 2855 186 2917 224
rect 2855 152 2869 186
rect 2903 152 2917 186
rect 2855 114 2917 152
rect 2189 47 2251 80
rect 2855 80 2869 114
rect 2903 80 2917 114
rect 3299 368 3313 402
rect 3347 368 3361 402
rect 3299 330 3361 368
rect 3299 296 3313 330
rect 3347 296 3361 330
rect 3299 258 3361 296
rect 3299 224 3313 258
rect 3347 224 3361 258
rect 3299 186 3361 224
rect 3299 152 3313 186
rect 3347 152 3361 186
rect 3299 114 3361 152
rect 2855 47 2917 80
rect 3299 80 3313 114
rect 3347 80 3361 114
rect 3299 47 3361 80
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 361 47
rect 395 13 433 47
rect 467 13 505 47
rect 539 13 577 47
rect 611 13 721 47
rect 755 13 793 47
rect 827 13 871 47
rect 905 13 949 47
rect 983 13 1021 47
rect 1055 13 1165 47
rect 1199 13 1237 47
rect 1271 13 1315 47
rect 1349 13 1393 47
rect 1427 13 1465 47
rect 1499 13 1609 47
rect 1643 13 1681 47
rect 1715 13 1753 47
rect 1787 13 1825 47
rect 1859 13 1915 47
rect 1949 13 1987 47
rect 2021 13 2059 47
rect 2093 13 2131 47
rect 2165 13 2275 47
rect 2309 13 2347 47
rect 2381 13 2419 47
rect 2453 13 2491 47
rect 2525 13 2581 47
rect 2615 13 2653 47
rect 2687 13 2725 47
rect 2759 13 2797 47
rect 2831 13 2941 47
rect 2975 13 3013 47
rect 3047 13 3091 47
rect 3125 13 3169 47
rect 3203 13 3241 47
rect 3275 13 3361 47
rect -31 11 31 13
rect 635 11 697 13
rect 1079 11 1141 13
rect 1523 11 1585 13
rect 2189 11 2251 13
rect 2855 11 2917 13
rect 3299 11 3361 13
<< nsubdiff >>
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 361 1539
rect 395 1505 433 1539
rect 467 1505 505 1539
rect 539 1505 577 1539
rect 611 1505 721 1539
rect 755 1505 793 1539
rect 827 1505 871 1539
rect 905 1505 949 1539
rect 983 1505 1021 1539
rect 1055 1505 1165 1539
rect 1199 1505 1237 1539
rect 1271 1505 1315 1539
rect 1349 1505 1393 1539
rect 1427 1505 1465 1539
rect 1499 1505 1609 1539
rect 1643 1505 1681 1539
rect 1715 1505 1753 1539
rect 1787 1505 1825 1539
rect 1859 1505 1915 1539
rect 1949 1505 1987 1539
rect 2021 1505 2059 1539
rect 2093 1505 2131 1539
rect 2165 1505 2275 1539
rect 2309 1505 2347 1539
rect 2381 1505 2419 1539
rect 2453 1505 2491 1539
rect 2525 1505 2581 1539
rect 2615 1505 2653 1539
rect 2687 1505 2725 1539
rect 2759 1505 2797 1539
rect 2831 1505 2941 1539
rect 2975 1505 3013 1539
rect 3047 1505 3091 1539
rect 3125 1505 3169 1539
rect 3203 1505 3241 1539
rect 3275 1505 3361 1539
rect -31 1470 31 1505
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect 635 1470 697 1505
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect -31 1038 31 1076
rect 635 1436 649 1470
rect 683 1436 697 1470
rect 1079 1470 1141 1505
rect 635 1398 697 1436
rect 635 1364 649 1398
rect 683 1364 697 1398
rect 635 1326 697 1364
rect 635 1292 649 1326
rect 683 1292 697 1326
rect 635 1254 697 1292
rect 635 1220 649 1254
rect 683 1220 697 1254
rect 635 1182 697 1220
rect 635 1148 649 1182
rect 683 1148 697 1182
rect 635 1110 697 1148
rect 635 1076 649 1110
rect 683 1076 697 1110
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect 635 1038 697 1076
rect 1079 1436 1093 1470
rect 1127 1436 1141 1470
rect 1523 1470 1585 1505
rect 1079 1398 1141 1436
rect 1079 1364 1093 1398
rect 1127 1364 1141 1398
rect 1079 1326 1141 1364
rect 1079 1292 1093 1326
rect 1127 1292 1141 1326
rect 1079 1254 1141 1292
rect 1079 1220 1093 1254
rect 1127 1220 1141 1254
rect 1079 1182 1141 1220
rect 1079 1148 1093 1182
rect 1127 1148 1141 1182
rect 1079 1110 1141 1148
rect 1079 1076 1093 1110
rect 1127 1076 1141 1110
rect 635 1004 649 1038
rect 683 1004 697 1038
rect 635 966 697 1004
rect -31 930 31 932
rect 635 932 649 966
rect 683 932 697 966
rect 1079 1038 1141 1076
rect 1523 1436 1537 1470
rect 1571 1436 1585 1470
rect 2189 1470 2251 1505
rect 1523 1398 1585 1436
rect 1523 1364 1537 1398
rect 1571 1364 1585 1398
rect 1523 1326 1585 1364
rect 1523 1292 1537 1326
rect 1571 1292 1585 1326
rect 1523 1254 1585 1292
rect 1523 1220 1537 1254
rect 1571 1220 1585 1254
rect 1523 1182 1585 1220
rect 1523 1148 1537 1182
rect 1571 1148 1585 1182
rect 1523 1110 1585 1148
rect 1523 1076 1537 1110
rect 1571 1076 1585 1110
rect 1079 1004 1093 1038
rect 1127 1004 1141 1038
rect 1079 966 1141 1004
rect 635 930 697 932
rect 1079 932 1093 966
rect 1127 932 1141 966
rect 1523 1038 1585 1076
rect 2189 1436 2203 1470
rect 2237 1436 2251 1470
rect 2855 1470 2917 1505
rect 2189 1398 2251 1436
rect 2189 1364 2203 1398
rect 2237 1364 2251 1398
rect 2189 1326 2251 1364
rect 2189 1292 2203 1326
rect 2237 1292 2251 1326
rect 2189 1254 2251 1292
rect 2189 1220 2203 1254
rect 2237 1220 2251 1254
rect 2189 1182 2251 1220
rect 2189 1148 2203 1182
rect 2237 1148 2251 1182
rect 2189 1110 2251 1148
rect 2189 1076 2203 1110
rect 2237 1076 2251 1110
rect 1523 1004 1537 1038
rect 1571 1004 1585 1038
rect 1523 966 1585 1004
rect 1079 930 1141 932
rect 1523 932 1537 966
rect 1571 932 1585 966
rect 2189 1038 2251 1076
rect 2855 1436 2869 1470
rect 2903 1436 2917 1470
rect 3299 1470 3361 1505
rect 2855 1398 2917 1436
rect 2855 1364 2869 1398
rect 2903 1364 2917 1398
rect 2855 1326 2917 1364
rect 2855 1292 2869 1326
rect 2903 1292 2917 1326
rect 2855 1254 2917 1292
rect 2855 1220 2869 1254
rect 2903 1220 2917 1254
rect 2855 1182 2917 1220
rect 2855 1148 2869 1182
rect 2903 1148 2917 1182
rect 2855 1110 2917 1148
rect 2855 1076 2869 1110
rect 2903 1076 2917 1110
rect 2189 1004 2203 1038
rect 2237 1004 2251 1038
rect 2189 966 2251 1004
rect 1523 930 1585 932
rect 2189 932 2203 966
rect 2237 932 2251 966
rect 2855 1038 2917 1076
rect 3299 1436 3313 1470
rect 3347 1436 3361 1470
rect 3299 1398 3361 1436
rect 3299 1364 3313 1398
rect 3347 1364 3361 1398
rect 3299 1326 3361 1364
rect 3299 1292 3313 1326
rect 3347 1292 3361 1326
rect 3299 1254 3361 1292
rect 3299 1220 3313 1254
rect 3347 1220 3361 1254
rect 3299 1182 3361 1220
rect 3299 1148 3313 1182
rect 3347 1148 3361 1182
rect 3299 1110 3361 1148
rect 3299 1076 3313 1110
rect 3347 1076 3361 1110
rect 2855 1004 2869 1038
rect 2903 1004 2917 1038
rect 2855 966 2917 1004
rect 3299 1038 3361 1076
rect 2189 930 2251 932
rect 2855 932 2869 966
rect 2903 932 2917 966
rect 3299 1004 3313 1038
rect 3347 1004 3361 1038
rect 3299 966 3361 1004
rect 2855 930 2917 932
rect 3299 932 3313 966
rect 3347 932 3361 966
rect 3299 930 3361 932
rect -31 868 3361 930
<< psubdiffcont >>
rect -17 512 17 546
rect 649 512 683 546
rect 1093 512 1127 546
rect 1537 512 1571 546
rect 2203 512 2237 546
rect 2869 512 2903 546
rect 3313 512 3347 546
rect -17 440 17 474
rect -17 368 17 402
rect 649 440 683 474
rect -17 296 17 330
rect -17 224 17 258
rect -17 152 17 186
rect -17 80 17 114
rect 649 368 683 402
rect 1093 440 1127 474
rect 649 296 683 330
rect 649 224 683 258
rect 649 152 683 186
rect 649 80 683 114
rect 1093 368 1127 402
rect 1537 440 1571 474
rect 1093 296 1127 330
rect 1093 224 1127 258
rect 1093 152 1127 186
rect 1093 80 1127 114
rect 1537 368 1571 402
rect 2203 440 2237 474
rect 1537 296 1571 330
rect 1537 224 1571 258
rect 1537 152 1571 186
rect 1537 80 1571 114
rect 2203 368 2237 402
rect 2869 440 2903 474
rect 2203 296 2237 330
rect 2203 224 2237 258
rect 2203 152 2237 186
rect 2203 80 2237 114
rect 2869 368 2903 402
rect 3313 440 3347 474
rect 2869 296 2903 330
rect 2869 224 2903 258
rect 2869 152 2903 186
rect 2869 80 2903 114
rect 3313 368 3347 402
rect 3313 296 3347 330
rect 3313 224 3347 258
rect 3313 152 3347 186
rect 3313 80 3347 114
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 361 13 395 47
rect 433 13 467 47
rect 505 13 539 47
rect 577 13 611 47
rect 721 13 755 47
rect 793 13 827 47
rect 871 13 905 47
rect 949 13 983 47
rect 1021 13 1055 47
rect 1165 13 1199 47
rect 1237 13 1271 47
rect 1315 13 1349 47
rect 1393 13 1427 47
rect 1465 13 1499 47
rect 1609 13 1643 47
rect 1681 13 1715 47
rect 1753 13 1787 47
rect 1825 13 1859 47
rect 1915 13 1949 47
rect 1987 13 2021 47
rect 2059 13 2093 47
rect 2131 13 2165 47
rect 2275 13 2309 47
rect 2347 13 2381 47
rect 2419 13 2453 47
rect 2491 13 2525 47
rect 2581 13 2615 47
rect 2653 13 2687 47
rect 2725 13 2759 47
rect 2797 13 2831 47
rect 2941 13 2975 47
rect 3013 13 3047 47
rect 3091 13 3125 47
rect 3169 13 3203 47
rect 3241 13 3275 47
<< nsubdiffcont >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 361 1505 395 1539
rect 433 1505 467 1539
rect 505 1505 539 1539
rect 577 1505 611 1539
rect 721 1505 755 1539
rect 793 1505 827 1539
rect 871 1505 905 1539
rect 949 1505 983 1539
rect 1021 1505 1055 1539
rect 1165 1505 1199 1539
rect 1237 1505 1271 1539
rect 1315 1505 1349 1539
rect 1393 1505 1427 1539
rect 1465 1505 1499 1539
rect 1609 1505 1643 1539
rect 1681 1505 1715 1539
rect 1753 1505 1787 1539
rect 1825 1505 1859 1539
rect 1915 1505 1949 1539
rect 1987 1505 2021 1539
rect 2059 1505 2093 1539
rect 2131 1505 2165 1539
rect 2275 1505 2309 1539
rect 2347 1505 2381 1539
rect 2419 1505 2453 1539
rect 2491 1505 2525 1539
rect 2581 1505 2615 1539
rect 2653 1505 2687 1539
rect 2725 1505 2759 1539
rect 2797 1505 2831 1539
rect 2941 1505 2975 1539
rect 3013 1505 3047 1539
rect 3091 1505 3125 1539
rect 3169 1505 3203 1539
rect 3241 1505 3275 1539
rect -17 1436 17 1470
rect -17 1364 17 1398
rect -17 1292 17 1326
rect -17 1220 17 1254
rect -17 1148 17 1182
rect -17 1076 17 1110
rect 649 1436 683 1470
rect 649 1364 683 1398
rect 649 1292 683 1326
rect 649 1220 683 1254
rect 649 1148 683 1182
rect 649 1076 683 1110
rect -17 1004 17 1038
rect -17 932 17 966
rect 1093 1436 1127 1470
rect 1093 1364 1127 1398
rect 1093 1292 1127 1326
rect 1093 1220 1127 1254
rect 1093 1148 1127 1182
rect 1093 1076 1127 1110
rect 649 1004 683 1038
rect 649 932 683 966
rect 1537 1436 1571 1470
rect 1537 1364 1571 1398
rect 1537 1292 1571 1326
rect 1537 1220 1571 1254
rect 1537 1148 1571 1182
rect 1537 1076 1571 1110
rect 1093 1004 1127 1038
rect 1093 932 1127 966
rect 2203 1436 2237 1470
rect 2203 1364 2237 1398
rect 2203 1292 2237 1326
rect 2203 1220 2237 1254
rect 2203 1148 2237 1182
rect 2203 1076 2237 1110
rect 1537 1004 1571 1038
rect 1537 932 1571 966
rect 2869 1436 2903 1470
rect 2869 1364 2903 1398
rect 2869 1292 2903 1326
rect 2869 1220 2903 1254
rect 2869 1148 2903 1182
rect 2869 1076 2903 1110
rect 2203 1004 2237 1038
rect 2203 932 2237 966
rect 3313 1436 3347 1470
rect 3313 1364 3347 1398
rect 3313 1292 3347 1326
rect 3313 1220 3347 1254
rect 3313 1148 3347 1182
rect 3313 1076 3347 1110
rect 2869 1004 2903 1038
rect 2869 932 2903 966
rect 3313 1004 3347 1038
rect 3313 932 3347 966
<< poly >>
rect 187 1450 217 1476
rect 275 1450 305 1476
rect 363 1450 393 1476
rect 451 1450 481 1476
rect 829 1450 859 1476
rect 917 1450 947 1476
rect 187 1019 217 1050
rect 275 1019 305 1050
rect 363 1019 393 1050
rect 451 1019 481 1050
rect 187 1003 305 1019
rect 187 989 205 1003
rect 195 969 205 989
rect 239 989 305 1003
rect 349 1003 481 1019
rect 239 969 249 989
rect 195 953 249 969
rect 349 969 359 1003
rect 393 989 481 1003
rect 1273 1450 1303 1476
rect 1361 1450 1391 1476
rect 829 1019 859 1050
rect 917 1019 947 1050
rect 393 969 403 989
rect 349 953 403 969
rect 787 1003 947 1019
rect 787 969 797 1003
rect 831 989 947 1003
rect 1741 1451 1771 1477
rect 1829 1451 1859 1477
rect 1917 1451 1947 1477
rect 2005 1451 2035 1477
rect 1273 1019 1303 1050
rect 1361 1019 1391 1050
rect 831 969 841 989
rect 787 953 841 969
rect 1231 1003 1391 1019
rect 1231 969 1241 1003
rect 1275 989 1391 1003
rect 2407 1451 2437 1477
rect 2495 1451 2525 1477
rect 2583 1451 2613 1477
rect 2671 1451 2701 1477
rect 1275 969 1285 989
rect 1231 953 1285 969
rect 1741 1020 1771 1051
rect 1829 1020 1859 1051
rect 1741 1004 1859 1020
rect 1741 990 1759 1004
rect 1749 970 1759 990
rect 1793 990 1859 1004
rect 1917 1020 1947 1051
rect 2005 1020 2035 1051
rect 1917 1004 2035 1020
rect 1917 990 1981 1004
rect 1793 970 1803 990
rect 1749 954 1803 970
rect 1971 970 1981 990
rect 2015 990 2035 1004
rect 3049 1450 3079 1476
rect 3137 1450 3167 1476
rect 2015 970 2025 990
rect 1971 954 2025 970
rect 2407 1020 2437 1051
rect 2495 1020 2525 1051
rect 2407 1004 2525 1020
rect 2407 990 2425 1004
rect 2415 970 2425 990
rect 2459 990 2525 1004
rect 2583 1020 2613 1051
rect 2671 1020 2701 1051
rect 2583 1004 2701 1020
rect 2583 990 2647 1004
rect 2459 970 2469 990
rect 2415 954 2469 970
rect 2637 970 2647 990
rect 2681 990 2701 1004
rect 2681 970 2691 990
rect 2637 954 2691 970
rect 3049 1019 3079 1050
rect 3137 1019 3167 1050
rect 3049 1003 3209 1019
rect 3049 989 3165 1003
rect 3155 969 3165 989
rect 3199 969 3209 1003
rect 3155 953 3209 969
rect 195 461 249 477
rect 195 441 205 461
rect 168 427 205 441
rect 239 427 249 461
rect 168 411 249 427
rect 343 461 397 477
rect 343 427 353 461
rect 387 427 397 461
rect 343 411 397 427
rect 168 377 198 411
rect 362 377 392 411
rect 787 461 841 477
rect 787 427 797 461
rect 831 441 841 461
rect 831 427 851 441
rect 787 411 851 427
rect 821 377 851 411
rect 1231 461 1285 477
rect 1231 427 1241 461
rect 1275 441 1285 461
rect 1275 427 1295 441
rect 1231 411 1295 427
rect 1265 377 1295 411
rect 1749 461 1803 477
rect 1749 441 1759 461
rect 1722 427 1759 441
rect 1793 427 1803 461
rect 1971 461 2025 477
rect 1971 441 1981 461
rect 1722 411 1803 427
rect 1916 427 1981 441
rect 2015 427 2025 461
rect 1916 411 2025 427
rect 2415 461 2469 477
rect 2415 441 2425 461
rect 1722 377 1752 411
rect 1916 377 1946 411
rect 2388 427 2425 441
rect 2459 427 2469 461
rect 2637 461 2691 477
rect 2637 441 2647 461
rect 2388 411 2469 427
rect 2582 427 2647 441
rect 2681 427 2691 461
rect 2582 411 2691 427
rect 3155 461 3209 477
rect 3155 441 3165 461
rect 2388 377 2418 411
rect 2582 377 2612 411
rect 3145 427 3165 441
rect 3199 427 3209 461
rect 3145 411 3209 427
rect 3145 377 3175 411
<< polycont >>
rect 205 969 239 1003
rect 359 969 393 1003
rect 797 969 831 1003
rect 1241 969 1275 1003
rect 1759 970 1793 1004
rect 1981 970 2015 1004
rect 2425 970 2459 1004
rect 2647 970 2681 1004
rect 3165 969 3199 1003
rect 205 427 239 461
rect 353 427 387 461
rect 797 427 831 461
rect 1241 427 1275 461
rect 1759 427 1793 461
rect 1981 427 2015 461
rect 2425 427 2459 461
rect 2647 427 2681 461
rect 3165 427 3199 461
<< locali >>
rect -31 1539 3361 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 361 1539
rect 395 1505 433 1539
rect 467 1505 505 1539
rect 539 1505 577 1539
rect 611 1505 721 1539
rect 755 1505 793 1539
rect 827 1505 871 1539
rect 905 1505 949 1539
rect 983 1505 1021 1539
rect 1055 1505 1165 1539
rect 1199 1505 1237 1539
rect 1271 1505 1315 1539
rect 1349 1505 1393 1539
rect 1427 1505 1465 1539
rect 1499 1505 1609 1539
rect 1643 1505 1681 1539
rect 1715 1505 1753 1539
rect 1787 1505 1825 1539
rect 1859 1505 1915 1539
rect 1949 1505 1987 1539
rect 2021 1505 2059 1539
rect 2093 1505 2131 1539
rect 2165 1505 2275 1539
rect 2309 1505 2347 1539
rect 2381 1505 2419 1539
rect 2453 1505 2491 1539
rect 2525 1505 2581 1539
rect 2615 1505 2653 1539
rect 2687 1505 2725 1539
rect 2759 1505 2797 1539
rect 2831 1505 2941 1539
rect 2975 1505 3013 1539
rect 3047 1505 3091 1539
rect 3125 1505 3169 1539
rect 3203 1505 3241 1539
rect 3275 1505 3361 1539
rect -31 1492 3361 1505
rect -31 1470 31 1492
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect -31 1038 31 1076
rect 141 1412 175 1492
rect 141 1344 175 1378
rect 141 1276 175 1310
rect 141 1208 175 1242
rect 141 1139 175 1174
rect 141 1073 175 1105
rect 229 1412 263 1450
rect 229 1344 263 1378
rect 229 1276 263 1310
rect 229 1208 263 1242
rect 229 1139 263 1174
rect 317 1412 351 1492
rect 317 1344 351 1378
rect 317 1276 351 1310
rect 317 1208 351 1242
rect 317 1157 351 1174
rect 405 1412 439 1450
rect 405 1344 439 1378
rect 405 1276 439 1310
rect 405 1208 439 1242
rect 229 1103 263 1105
rect 405 1139 439 1174
rect 493 1412 527 1492
rect 493 1344 527 1378
rect 493 1276 527 1310
rect 493 1208 527 1242
rect 493 1157 527 1174
rect 635 1470 697 1492
rect 635 1436 649 1470
rect 683 1436 697 1470
rect 635 1398 697 1436
rect 635 1364 649 1398
rect 683 1364 697 1398
rect 635 1326 697 1364
rect 635 1292 649 1326
rect 683 1292 697 1326
rect 635 1254 697 1292
rect 635 1220 649 1254
rect 683 1220 697 1254
rect 635 1182 697 1220
rect 405 1103 439 1105
rect 635 1148 649 1182
rect 683 1148 697 1182
rect 635 1110 697 1148
rect 229 1069 535 1103
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect -31 868 31 932
rect 205 1003 239 1019
rect 359 1003 393 1019
rect 205 905 239 969
rect -31 546 31 572
rect -31 512 -17 546
rect 17 512 31 546
rect -31 474 31 512
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect 205 461 239 871
rect 205 411 239 427
rect 353 969 359 988
rect 353 953 393 969
rect 353 757 387 953
rect 353 461 387 723
rect 353 411 387 427
rect 501 683 535 1069
rect 635 1076 649 1110
rect 683 1076 697 1110
rect 783 1412 817 1492
rect 783 1344 817 1378
rect 783 1276 817 1310
rect 783 1208 817 1242
rect 783 1139 817 1174
rect 783 1083 817 1105
rect 871 1412 905 1450
rect 871 1344 905 1378
rect 871 1276 905 1310
rect 871 1208 905 1242
rect 871 1139 905 1174
rect 635 1038 697 1076
rect 635 1004 649 1038
rect 683 1004 697 1038
rect 635 966 697 1004
rect 635 932 649 966
rect 683 932 697 966
rect 635 868 697 932
rect 797 1003 831 1019
rect -31 368 -17 402
rect 17 368 31 402
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect 122 361 156 377
rect 316 361 350 377
rect 501 376 535 649
rect 797 683 831 969
rect 871 979 905 1105
rect 959 1412 993 1492
rect 959 1344 993 1378
rect 959 1276 993 1310
rect 959 1208 993 1242
rect 959 1139 993 1174
rect 959 1083 993 1105
rect 1079 1470 1141 1492
rect 1079 1436 1093 1470
rect 1127 1436 1141 1470
rect 1079 1398 1141 1436
rect 1079 1364 1093 1398
rect 1127 1364 1141 1398
rect 1079 1326 1141 1364
rect 1079 1292 1093 1326
rect 1127 1292 1141 1326
rect 1079 1254 1141 1292
rect 1079 1220 1093 1254
rect 1127 1220 1141 1254
rect 1079 1182 1141 1220
rect 1079 1148 1093 1182
rect 1127 1148 1141 1182
rect 1079 1110 1141 1148
rect 1079 1076 1093 1110
rect 1127 1076 1141 1110
rect 1227 1412 1261 1492
rect 1227 1344 1261 1378
rect 1227 1276 1261 1310
rect 1227 1208 1261 1242
rect 1227 1139 1261 1174
rect 1227 1083 1261 1105
rect 1315 1412 1349 1450
rect 1315 1344 1349 1378
rect 1315 1276 1349 1310
rect 1315 1208 1349 1242
rect 1315 1139 1349 1174
rect 1079 1038 1141 1076
rect 1079 1004 1093 1038
rect 1127 1004 1141 1038
rect 871 945 979 979
rect 156 327 219 361
rect 253 327 316 361
rect 122 289 156 327
rect 122 221 156 255
rect 316 289 350 327
rect 122 151 156 187
rect 122 101 156 117
rect 219 236 253 252
rect -31 62 31 80
rect 219 62 253 202
rect 316 221 350 255
rect 413 342 535 376
rect 635 546 697 572
rect 635 512 649 546
rect 683 512 697 546
rect 635 474 697 512
rect 635 440 649 474
rect 683 440 697 474
rect 635 402 697 440
rect 797 461 831 649
rect 945 609 979 945
rect 1079 966 1141 1004
rect 1079 932 1093 966
rect 1127 932 1141 966
rect 1079 868 1141 932
rect 1241 1003 1275 1019
rect 1241 905 1275 969
rect 1315 979 1349 1105
rect 1403 1412 1437 1492
rect 1403 1344 1437 1378
rect 1403 1276 1437 1310
rect 1403 1208 1437 1242
rect 1403 1139 1437 1174
rect 1403 1083 1437 1105
rect 1523 1470 1585 1492
rect 1523 1436 1537 1470
rect 1571 1436 1585 1470
rect 1523 1398 1585 1436
rect 1523 1364 1537 1398
rect 1571 1364 1585 1398
rect 1523 1326 1585 1364
rect 1523 1292 1537 1326
rect 1571 1292 1585 1326
rect 1523 1254 1585 1292
rect 1523 1220 1537 1254
rect 1571 1220 1585 1254
rect 1523 1182 1585 1220
rect 1523 1148 1537 1182
rect 1571 1148 1585 1182
rect 1523 1110 1585 1148
rect 1523 1076 1537 1110
rect 1571 1076 1585 1110
rect 1523 1038 1585 1076
rect 1695 1411 1729 1427
rect 1695 1343 1729 1377
rect 1695 1275 1729 1309
rect 1695 1207 1729 1241
rect 1695 1139 1729 1173
rect 1783 1343 1817 1492
rect 2189 1470 2251 1492
rect 1783 1275 1817 1309
rect 1783 1207 1817 1241
rect 1783 1157 1817 1173
rect 1871 1411 2081 1445
rect 1871 1343 1905 1377
rect 1871 1275 1905 1309
rect 1871 1207 1905 1241
rect 1871 1139 1905 1173
rect 1695 1071 1905 1105
rect 1959 1343 1993 1359
rect 1959 1275 1993 1309
rect 1959 1207 1993 1241
rect 1959 1139 1993 1173
rect 2047 1343 2081 1377
rect 2047 1275 2081 1309
rect 2047 1207 2081 1241
rect 2047 1157 2081 1173
rect 2189 1436 2203 1470
rect 2237 1436 2251 1470
rect 2189 1398 2251 1436
rect 2189 1364 2203 1398
rect 2237 1364 2251 1398
rect 2189 1326 2251 1364
rect 2189 1292 2203 1326
rect 2237 1292 2251 1326
rect 2189 1254 2251 1292
rect 2189 1220 2203 1254
rect 2237 1220 2251 1254
rect 2189 1182 2251 1220
rect 2189 1148 2203 1182
rect 2237 1148 2251 1182
rect 2189 1110 2251 1148
rect 1959 1071 2089 1105
rect 1523 1004 1537 1038
rect 1571 1004 1585 1038
rect 1315 945 1423 979
rect 945 461 979 575
rect 797 411 831 427
rect 871 427 979 461
rect 1079 546 1141 572
rect 1079 512 1093 546
rect 1127 512 1141 546
rect 1079 474 1141 512
rect 1079 440 1093 474
rect 1127 440 1141 474
rect 635 368 649 402
rect 683 368 697 402
rect 413 245 447 342
rect 635 330 697 368
rect 413 195 447 211
rect 510 289 544 305
rect 510 221 544 255
rect 316 151 350 187
rect 510 151 544 187
rect 350 117 413 151
rect 447 117 510 151
rect 316 101 350 117
rect 510 101 544 117
rect 635 296 649 330
rect 683 296 697 330
rect 635 258 697 296
rect 635 224 649 258
rect 683 224 697 258
rect 635 186 697 224
rect 635 152 649 186
rect 683 152 697 186
rect 635 114 697 152
rect 635 80 649 114
rect 683 80 697 114
rect 635 62 697 80
rect 775 361 809 377
rect 775 289 809 327
rect 775 221 809 255
rect 871 245 905 427
rect 1079 402 1141 440
rect 1241 461 1275 871
rect 1389 683 1423 945
rect 1523 966 1585 1004
rect 1523 932 1537 966
rect 1571 932 1585 966
rect 1523 868 1585 932
rect 1759 1004 1793 1020
rect 1759 905 1793 970
rect 1981 1004 2015 1020
rect 1389 461 1423 649
rect 1241 411 1275 427
rect 1315 427 1423 461
rect 1523 546 1585 572
rect 1523 512 1537 546
rect 1571 512 1585 546
rect 1523 474 1585 512
rect 1523 440 1537 474
rect 1571 440 1585 474
rect 871 195 905 211
rect 969 361 1003 377
rect 969 289 1003 327
rect 969 221 1003 255
rect 775 151 809 187
rect 969 151 1003 187
rect 809 117 871 151
rect 905 117 969 151
rect 775 62 809 117
rect 872 62 906 117
rect 969 62 1003 117
rect 1079 368 1093 402
rect 1127 368 1141 402
rect 1079 330 1141 368
rect 1079 296 1093 330
rect 1127 296 1141 330
rect 1079 258 1141 296
rect 1079 224 1093 258
rect 1127 224 1141 258
rect 1079 186 1141 224
rect 1079 152 1093 186
rect 1127 152 1141 186
rect 1079 114 1141 152
rect 1079 80 1093 114
rect 1127 80 1141 114
rect 1079 62 1141 80
rect 1219 361 1253 377
rect 1219 289 1253 327
rect 1219 221 1253 255
rect 1315 245 1349 427
rect 1523 402 1585 440
rect 1759 461 1793 871
rect 1907 905 1941 921
rect 1907 757 1941 871
rect 1981 831 2015 970
rect 1981 781 2015 797
rect 1907 707 1941 723
rect 2055 757 2089 1071
rect 2189 1076 2203 1110
rect 2237 1076 2251 1110
rect 2189 1038 2251 1076
rect 2361 1411 2395 1427
rect 2361 1343 2395 1377
rect 2361 1275 2395 1309
rect 2361 1207 2395 1241
rect 2361 1139 2395 1173
rect 2449 1343 2483 1492
rect 2855 1470 2917 1492
rect 2449 1275 2483 1309
rect 2449 1207 2483 1241
rect 2449 1157 2483 1173
rect 2537 1411 2747 1445
rect 2537 1343 2571 1377
rect 2537 1275 2571 1309
rect 2537 1207 2571 1241
rect 2537 1139 2571 1173
rect 2361 1071 2571 1105
rect 2625 1343 2659 1359
rect 2625 1275 2659 1309
rect 2625 1207 2659 1241
rect 2625 1139 2659 1173
rect 2713 1343 2747 1377
rect 2713 1275 2747 1309
rect 2713 1207 2747 1241
rect 2713 1157 2747 1173
rect 2855 1436 2869 1470
rect 2903 1436 2917 1470
rect 2855 1398 2917 1436
rect 2855 1364 2869 1398
rect 2903 1364 2917 1398
rect 2855 1326 2917 1364
rect 2855 1292 2869 1326
rect 2903 1292 2917 1326
rect 2855 1254 2917 1292
rect 2855 1220 2869 1254
rect 2903 1220 2917 1254
rect 2855 1182 2917 1220
rect 2855 1148 2869 1182
rect 2903 1148 2917 1182
rect 2855 1110 2917 1148
rect 2625 1071 2755 1105
rect 2189 1004 2203 1038
rect 2237 1004 2251 1038
rect 2189 966 2251 1004
rect 2189 932 2203 966
rect 2237 932 2251 966
rect 2189 868 2251 932
rect 2425 1004 2459 1020
rect 2425 905 2459 970
rect 2425 855 2459 871
rect 2647 1004 2681 1020
rect 1759 411 1793 427
rect 1981 535 2015 551
rect 1981 461 2015 501
rect 1981 411 2015 427
rect 1315 195 1349 211
rect 1413 361 1447 377
rect 1413 289 1447 327
rect 1413 221 1447 255
rect 1219 151 1253 187
rect 1413 151 1447 187
rect 1253 117 1315 151
rect 1349 117 1413 151
rect 1219 62 1253 117
rect 1316 62 1350 117
rect 1413 62 1447 117
rect 1523 368 1537 402
rect 1571 368 1585 402
rect 1523 330 1585 368
rect 1523 296 1537 330
rect 1571 296 1585 330
rect 1523 258 1585 296
rect 1523 224 1537 258
rect 1571 224 1585 258
rect 1523 186 1585 224
rect 1523 152 1537 186
rect 1571 152 1585 186
rect 1523 114 1585 152
rect 1523 80 1537 114
rect 1571 80 1585 114
rect 1676 361 1710 377
rect 1870 361 1904 377
rect 2055 375 2089 723
rect 2647 683 2681 970
rect 2425 609 2459 625
rect 1710 327 1773 361
rect 1807 327 1870 361
rect 1676 289 1710 327
rect 1676 221 1710 255
rect 1870 289 1904 327
rect 1676 151 1710 187
rect 1676 101 1710 117
rect 1773 236 1807 252
rect 1523 62 1585 80
rect 1773 62 1807 202
rect 1870 221 1904 255
rect 1967 341 2089 375
rect 2189 546 2251 572
rect 2189 512 2203 546
rect 2237 512 2251 546
rect 2189 474 2251 512
rect 2189 440 2203 474
rect 2237 440 2251 474
rect 2189 402 2251 440
rect 2425 461 2459 575
rect 2425 411 2459 427
rect 2647 461 2681 649
rect 2647 411 2681 427
rect 2721 757 2755 1071
rect 2855 1076 2869 1110
rect 2903 1076 2917 1110
rect 3003 1412 3037 1492
rect 3003 1344 3037 1378
rect 3003 1276 3037 1310
rect 3003 1208 3037 1242
rect 3003 1139 3037 1174
rect 3003 1083 3037 1105
rect 3091 1412 3125 1450
rect 3091 1344 3125 1378
rect 3091 1276 3125 1310
rect 3091 1208 3125 1242
rect 3091 1139 3125 1174
rect 2855 1038 2917 1076
rect 2855 1004 2869 1038
rect 2903 1004 2917 1038
rect 2855 966 2917 1004
rect 3091 979 3125 1105
rect 3179 1412 3213 1492
rect 3179 1344 3213 1378
rect 3179 1276 3213 1310
rect 3179 1208 3213 1242
rect 3179 1139 3213 1174
rect 3179 1083 3213 1105
rect 3299 1470 3361 1492
rect 3299 1436 3313 1470
rect 3347 1436 3361 1470
rect 3299 1398 3361 1436
rect 3299 1364 3313 1398
rect 3347 1364 3361 1398
rect 3299 1326 3361 1364
rect 3299 1292 3313 1326
rect 3347 1292 3361 1326
rect 3299 1254 3361 1292
rect 3299 1220 3313 1254
rect 3347 1220 3361 1254
rect 3299 1182 3361 1220
rect 3299 1148 3313 1182
rect 3347 1148 3361 1182
rect 3299 1110 3361 1148
rect 3299 1076 3313 1110
rect 3347 1076 3361 1110
rect 3299 1038 3361 1076
rect 2855 932 2869 966
rect 2903 932 2917 966
rect 2855 868 2917 932
rect 3017 945 3125 979
rect 3165 1003 3199 1019
rect 2189 368 2203 402
rect 2237 368 2251 402
rect 1967 245 2001 341
rect 2189 330 2251 368
rect 1967 195 2001 211
rect 2064 289 2098 305
rect 2064 221 2098 255
rect 1870 151 1904 187
rect 2064 151 2098 187
rect 1904 117 1967 151
rect 2001 117 2064 151
rect 1870 101 1904 117
rect 2064 101 2098 117
rect 2189 296 2203 330
rect 2237 296 2251 330
rect 2189 258 2251 296
rect 2189 224 2203 258
rect 2237 224 2251 258
rect 2189 186 2251 224
rect 2189 152 2203 186
rect 2237 152 2251 186
rect 2189 114 2251 152
rect 2189 80 2203 114
rect 2237 80 2251 114
rect 2342 361 2376 377
rect 2536 361 2570 377
rect 2721 375 2755 723
rect 3017 831 3051 945
rect 3017 609 3051 797
rect 2376 327 2439 361
rect 2473 327 2536 361
rect 2342 289 2376 327
rect 2342 221 2376 255
rect 2536 289 2570 327
rect 2342 151 2376 187
rect 2342 101 2376 117
rect 2439 236 2473 252
rect 2189 62 2251 80
rect 2439 62 2473 202
rect 2536 221 2570 255
rect 2633 341 2755 375
rect 2855 546 2917 572
rect 2855 512 2869 546
rect 2903 512 2917 546
rect 2855 474 2917 512
rect 2855 440 2869 474
rect 2903 440 2917 474
rect 2855 402 2917 440
rect 3017 461 3051 575
rect 3165 905 3199 969
rect 3165 535 3199 871
rect 3299 1004 3313 1038
rect 3347 1004 3361 1038
rect 3299 966 3361 1004
rect 3299 932 3313 966
rect 3347 932 3361 966
rect 3299 868 3361 932
rect 3165 461 3199 501
rect 3017 427 3125 461
rect 2855 368 2869 402
rect 2903 368 2917 402
rect 2633 245 2667 341
rect 2855 330 2917 368
rect 2633 195 2667 211
rect 2730 289 2764 305
rect 2730 221 2764 255
rect 2536 151 2570 187
rect 2730 151 2764 187
rect 2570 117 2633 151
rect 2667 117 2730 151
rect 2536 101 2570 117
rect 2730 101 2764 117
rect 2855 296 2869 330
rect 2903 296 2917 330
rect 2855 258 2917 296
rect 2855 224 2869 258
rect 2903 224 2917 258
rect 2855 186 2917 224
rect 2855 152 2869 186
rect 2903 152 2917 186
rect 2855 114 2917 152
rect 2855 80 2869 114
rect 2903 80 2917 114
rect 2855 62 2917 80
rect 2993 361 3027 377
rect 2993 289 3027 327
rect 2993 221 3027 255
rect 3091 245 3125 427
rect 3165 411 3199 427
rect 3299 546 3361 572
rect 3299 512 3313 546
rect 3347 512 3361 546
rect 3299 474 3361 512
rect 3299 440 3313 474
rect 3347 440 3361 474
rect 3299 402 3361 440
rect 3091 195 3125 211
rect 3187 361 3221 377
rect 3187 289 3221 327
rect 3187 221 3221 255
rect 2993 151 3027 187
rect 3187 151 3221 187
rect 3027 117 3091 151
rect 3125 117 3187 151
rect 2993 62 3027 117
rect 3090 62 3124 117
rect 3187 62 3221 117
rect 3299 368 3313 402
rect 3347 368 3361 402
rect 3299 330 3361 368
rect 3299 296 3313 330
rect 3347 296 3361 330
rect 3299 258 3361 296
rect 3299 224 3313 258
rect 3347 224 3361 258
rect 3299 186 3361 224
rect 3299 152 3313 186
rect 3347 152 3361 186
rect 3299 114 3361 152
rect 3299 80 3313 114
rect 3347 80 3361 114
rect 3299 62 3361 80
rect -31 47 3361 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 361 47
rect 395 13 433 47
rect 467 13 505 47
rect 539 13 577 47
rect 611 13 721 47
rect 755 13 793 47
rect 827 13 871 47
rect 905 13 949 47
rect 983 13 1021 47
rect 1055 13 1165 47
rect 1199 13 1237 47
rect 1271 13 1315 47
rect 1349 13 1393 47
rect 1427 13 1465 47
rect 1499 13 1609 47
rect 1643 13 1681 47
rect 1715 13 1753 47
rect 1787 13 1825 47
rect 1859 13 1915 47
rect 1949 13 1987 47
rect 2021 13 2059 47
rect 2093 13 2131 47
rect 2165 13 2275 47
rect 2309 13 2347 47
rect 2381 13 2419 47
rect 2453 13 2491 47
rect 2525 13 2581 47
rect 2615 13 2653 47
rect 2687 13 2725 47
rect 2759 13 2797 47
rect 2831 13 2941 47
rect 2975 13 3013 47
rect 3047 13 3091 47
rect 3125 13 3169 47
rect 3203 13 3241 47
rect 3275 13 3361 47
rect -31 0 3361 13
<< viali >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 361 1505 395 1539
rect 433 1505 467 1539
rect 505 1505 539 1539
rect 577 1505 611 1539
rect 721 1505 755 1539
rect 793 1505 827 1539
rect 871 1505 905 1539
rect 949 1505 983 1539
rect 1021 1505 1055 1539
rect 1165 1505 1199 1539
rect 1237 1505 1271 1539
rect 1315 1505 1349 1539
rect 1393 1505 1427 1539
rect 1465 1505 1499 1539
rect 1609 1505 1643 1539
rect 1681 1505 1715 1539
rect 1753 1505 1787 1539
rect 1825 1505 1859 1539
rect 1915 1505 1949 1539
rect 1987 1505 2021 1539
rect 2059 1505 2093 1539
rect 2131 1505 2165 1539
rect 2275 1505 2309 1539
rect 2347 1505 2381 1539
rect 2419 1505 2453 1539
rect 2491 1505 2525 1539
rect 2581 1505 2615 1539
rect 2653 1505 2687 1539
rect 2725 1505 2759 1539
rect 2797 1505 2831 1539
rect 2941 1505 2975 1539
rect 3013 1505 3047 1539
rect 3091 1505 3125 1539
rect 3169 1505 3203 1539
rect 3241 1505 3275 1539
rect 205 871 239 905
rect 353 723 387 757
rect 501 649 535 683
rect 797 649 831 683
rect 1241 871 1275 905
rect 945 575 979 609
rect 1759 871 1793 905
rect 1389 649 1423 683
rect 1907 871 1941 905
rect 1981 797 2015 831
rect 1907 723 1941 757
rect 2425 871 2459 905
rect 2055 723 2089 757
rect 1981 501 2015 535
rect 2647 649 2681 683
rect 2425 575 2459 609
rect 2721 723 2755 757
rect 3017 797 3051 831
rect 3017 575 3051 609
rect 3165 871 3199 905
rect 3165 501 3199 535
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 361 13 395 47
rect 433 13 467 47
rect 505 13 539 47
rect 577 13 611 47
rect 721 13 755 47
rect 793 13 827 47
rect 871 13 905 47
rect 949 13 983 47
rect 1021 13 1055 47
rect 1165 13 1199 47
rect 1237 13 1271 47
rect 1315 13 1349 47
rect 1393 13 1427 47
rect 1465 13 1499 47
rect 1609 13 1643 47
rect 1681 13 1715 47
rect 1753 13 1787 47
rect 1825 13 1859 47
rect 1915 13 1949 47
rect 1987 13 2021 47
rect 2059 13 2093 47
rect 2131 13 2165 47
rect 2275 13 2309 47
rect 2347 13 2381 47
rect 2419 13 2453 47
rect 2491 13 2525 47
rect 2581 13 2615 47
rect 2653 13 2687 47
rect 2725 13 2759 47
rect 2797 13 2831 47
rect 2941 13 2975 47
rect 3013 13 3047 47
rect 3091 13 3125 47
rect 3169 13 3203 47
rect 3241 13 3275 47
<< metal1 >>
rect -31 1539 3361 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 361 1539
rect 395 1505 433 1539
rect 467 1505 505 1539
rect 539 1505 577 1539
rect 611 1505 721 1539
rect 755 1505 793 1539
rect 827 1505 871 1539
rect 905 1505 949 1539
rect 983 1505 1021 1539
rect 1055 1505 1165 1539
rect 1199 1505 1237 1539
rect 1271 1505 1315 1539
rect 1349 1505 1393 1539
rect 1427 1505 1465 1539
rect 1499 1505 1609 1539
rect 1643 1505 1681 1539
rect 1715 1505 1753 1539
rect 1787 1505 1825 1539
rect 1859 1505 1915 1539
rect 1949 1505 1987 1539
rect 2021 1505 2059 1539
rect 2093 1505 2131 1539
rect 2165 1505 2275 1539
rect 2309 1505 2347 1539
rect 2381 1505 2419 1539
rect 2453 1505 2491 1539
rect 2525 1505 2581 1539
rect 2615 1505 2653 1539
rect 2687 1505 2725 1539
rect 2759 1505 2797 1539
rect 2831 1505 2941 1539
rect 2975 1505 3013 1539
rect 3047 1505 3091 1539
rect 3125 1505 3169 1539
rect 3203 1505 3241 1539
rect 3275 1505 3361 1539
rect -31 1492 3361 1505
rect 199 905 245 911
rect 1235 905 1281 911
rect 1753 905 1799 911
rect 1901 905 1947 911
rect 2419 905 2465 911
rect 3159 905 3205 911
rect 193 871 205 905
rect 239 871 1241 905
rect 1275 871 1759 905
rect 1793 871 1805 905
rect 1895 871 1907 905
rect 1941 871 2425 905
rect 2459 871 3165 905
rect 3199 871 3211 905
rect 199 865 245 871
rect 1235 865 1281 871
rect 1753 865 1799 871
rect 1901 865 1947 871
rect 2419 865 2465 871
rect 3159 865 3205 871
rect 1975 831 2021 837
rect 3011 831 3057 837
rect 1969 797 1981 831
rect 2015 797 3017 831
rect 3051 797 3063 831
rect 1975 791 2021 797
rect 3011 791 3057 797
rect 347 757 393 763
rect 1901 757 1947 763
rect 2049 757 2095 763
rect 2715 757 2761 763
rect 341 723 353 757
rect 387 723 1907 757
rect 1941 723 1953 757
rect 2043 723 2055 757
rect 2089 723 2721 757
rect 2755 723 2767 757
rect 347 717 393 723
rect 1901 717 1947 723
rect 2049 717 2095 723
rect 2715 717 2761 723
rect 495 683 541 689
rect 791 683 837 689
rect 1383 683 1429 689
rect 2641 683 2687 689
rect 489 649 501 683
rect 535 649 797 683
rect 831 649 843 683
rect 1377 649 1389 683
rect 1423 649 2647 683
rect 2681 649 2693 683
rect 495 643 541 649
rect 791 643 837 649
rect 1383 643 1429 649
rect 2641 643 2687 649
rect 939 609 985 615
rect 2419 609 2465 615
rect 3011 609 3057 615
rect 909 575 945 609
rect 979 575 991 609
rect 2413 575 2425 609
rect 2459 575 3017 609
rect 3051 575 3063 609
rect 939 569 985 575
rect 2419 569 2465 575
rect 3011 569 3057 575
rect 1975 535 2021 541
rect 3159 535 3205 541
rect 1969 501 1981 535
rect 2015 501 3165 535
rect 3199 501 3211 535
rect 1975 495 2021 501
rect 3159 495 3205 501
rect -31 47 3361 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 361 47
rect 395 13 433 47
rect 467 13 505 47
rect 539 13 577 47
rect 611 13 721 47
rect 755 13 793 47
rect 827 13 871 47
rect 905 13 949 47
rect 983 13 1021 47
rect 1055 13 1165 47
rect 1199 13 1237 47
rect 1271 13 1315 47
rect 1349 13 1393 47
rect 1427 13 1465 47
rect 1499 13 1609 47
rect 1643 13 1681 47
rect 1715 13 1753 47
rect 1787 13 1825 47
rect 1859 13 1915 47
rect 1949 13 1987 47
rect 2021 13 2059 47
rect 2093 13 2131 47
rect 2165 13 2275 47
rect 2309 13 2347 47
rect 2381 13 2419 47
rect 2453 13 2491 47
rect 2525 13 2581 47
rect 2615 13 2653 47
rect 2687 13 2725 47
rect 2759 13 2797 47
rect 2831 13 2941 47
rect 2975 13 3013 47
rect 3047 13 3091 47
rect 3125 13 3169 47
rect 3203 13 3241 47
rect 3275 13 3361 47
rect -31 0 3361 13
<< labels >>
rlabel metal1 2721 723 2755 757 1 SUM
port 1 n
rlabel metal1 945 575 979 609 1 COUT
port 2 n
rlabel metal1 205 871 239 905 1 A
port 3 n
rlabel metal1 353 723 387 757 1 B
port 4 n
rlabel metal1 55 1505 89 1539 1 VDD
port 5 n
rlabel metal1 55 13 89 47 1 VSS
port 6 n
<< end >>
