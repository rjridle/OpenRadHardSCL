* SPICE3 file created from MUX2X1.ext - technology: sky130A

.subckt MUX2X1 Y A0 A1 S VDD GND
X0 GND S.t1 a_556_101.t0 GND sky130_fd_pr__nfet_01v8 ad=1.6781p pd=1.281u as=0p ps=0u w=0u l=0u
X1 VDD.t15 a_185_209.t3 a_1327_1050.t2 @d%��U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X2 a_185_209.t0 S.t0 VDD.t11 0#��U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X3 a_661_1050.t2 A0.t0 VDD.t9  ����U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X4 VDD.t21 A1.t0 a_1327_1050.t3 �!���U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X5 a_661_1050.t4 S.t3 VDD.t23  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X6 a_1327_1050.t1 a_185_209.t4 VDD.t13 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X7 VDD.t19 a_1327_1050.t6 Y.t3 �+|6� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X8 VDD.t27 S.t4 a_661_1050.t3  ,|6� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X9 VDD.t7 a_661_1050.t5 Y.t1 �+|6� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X10 a_1327_1050.t0 A1.t2 VDD.t3  ,|6� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X11 VDD.t25 S.t5 a_185_209.t2 �+|6� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X12 Y.t0 a_661_1050.t6 VDD.t1  ,|6� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X13 GND a_661_1050.t7 a_1888_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X14 GND a_185_209.t5 a_1222_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X15 Y.t2 a_1327_1050.t7 VDD.t17 �+|6� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X16 Y a_1327_1050.t5 a_1888_101.t0 GND sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=0p ps=0u w=0u l=0u
X17 VDD.t5 A0.t2 a_661_1050.t1  ,|6� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
C0 A0 S 0.27fF
C1 A1 VDD 0.33fF
C2 A0 VDD 0.32fF
C3 S VDD 0.70fF
C4 Y VDD 1.85fF
R0 a_185_209.n1 a_185_209.t3 480.392
R1 a_185_209.n1 a_185_209.t4 403.272
R2 a_185_209.n2 a_185_209.t5 329.345
R3 a_185_209.n5 a_185_209.n3 278.973
R4 a_185_209.n3 a_185_209.n0 271.281
R5 a_185_209.n2 a_185_209.n1 199.147
R6 a_185_209.n5 a_185_209.n4 15.218
R7 a_185_209.n0 a_185_209.t2 14.282
R8 a_185_209.n0 a_185_209.t0 14.282
R9 a_185_209.n3 a_185_209.n2 13.063
R10 a_185_209.n6 a_185_209.n5 12.014
R11 a_1327_1050.n3 a_1327_1050.t6 472.359
R12 a_1327_1050.n3 a_1327_1050.t7 384.527
R13 a_1327_1050.n4 a_1327_1050.t5 287.037
R14 a_1327_1050.n7 a_1327_1050.n5 284.244
R15 a_1327_1050.n4 a_1327_1050.n3 210.673
R16 a_1327_1050.n5 a_1327_1050.n2 187.858
R17 a_1327_1050.n2 a_1327_1050.n1 157.964
R18 a_1327_1050.n2 a_1327_1050.n0 91.706
R19 a_1327_1050.n7 a_1327_1050.n6 15.218
R20 a_1327_1050.n0 a_1327_1050.t3 14.282
R21 a_1327_1050.n0 a_1327_1050.t0 14.282
R22 a_1327_1050.n1 a_1327_1050.t2 14.282
R23 a_1327_1050.n1 a_1327_1050.t1 14.282
R24 a_1327_1050.n8 a_1327_1050.n7 12.014
R25 a_1327_1050.n5 a_1327_1050.n4 11.159
R26 VDD.n161 VDD.n150 144.705
R27 VDD.n79 VDD.n68 144.705
R28 VDD.n215 VDD.n208 144.705
R29 VDD.n201 VDD.t5 143.754
R30 VDD.n84 VDD.t21 143.754
R31 VDD.n26 VDD.t19 143.754
R32 VDD.n134 VDD.t11 135.17
R33 VDD.n141 VDD.t25 135.17
R34 VDD.n177 VDD.t23 135.17
R35 VDD.n104 VDD.t13 135.17
R36 VDD.n46 VDD.t1 135.17
R37 VDD.n192 VDD.n191 129.472
R38 VDD.n93 VDD.n92 129.472
R39 VDD.n35 VDD.n34 129.472
R40 VDD.n64 VDD.n63 92.5
R41 VDD.n62 VDD.n61 92.5
R42 VDD.n60 VDD.n59 92.5
R43 VDD.n58 VDD.n57 92.5
R44 VDD.n66 VDD.n65 92.5
R45 VDD.n228 VDD.n227 92.5
R46 VDD.n226 VDD.n225 92.5
R47 VDD.n224 VDD.n223 92.5
R48 VDD.n222 VDD.n221 92.5
R49 VDD.n230 VDD.n229 92.5
R50 VDD.n171 VDD.n170 92.5
R51 VDD.n169 VDD.n168 92.5
R52 VDD.n167 VDD.n166 92.5
R53 VDD.n165 VDD.n164 92.5
R54 VDD.n173 VDD.n172 92.5
R55 VDD.n120 VDD.n119 92.5
R56 VDD.n118 VDD.n117 92.5
R57 VDD.n116 VDD.n115 92.5
R58 VDD.n114 VDD.n113 92.5
R59 VDD.n122 VDD.n121 92.5
R60 VDD.n14 VDD.n1 92.5
R61 VDD.n5 VDD.n4 92.5
R62 VDD.n7 VDD.n6 92.5
R63 VDD.n9 VDD.n8 92.5
R64 VDD.n11 VDD.n10 92.5
R65 VDD.n13 VDD.n12 92.5
R66 VDD.n21 VDD.n20 92.059
R67 VDD.n78 VDD.n77 92.059
R68 VDD.n214 VDD.n213 92.059
R69 VDD.n160 VDD.n159 92.059
R70 VDD.n128 VDD.n127 92.059
R71 VDD.n20 VDD.n16 67.194
R72 VDD.n20 VDD.n17 67.194
R73 VDD.n20 VDD.n18 67.194
R74 VDD.n20 VDD.n19 67.194
R75 VDD.n112 VDD.n111 44.141
R76 VDD.n220 VDD.n219 44.141
R77 VDD.n5 VDD.n3 44.141
R78 VDD.n219 VDD.n217 44.107
R79 VDD.n111 VDD.n109 44.107
R80 VDD.n3 VDD.n2 44.107
R81 VDD.n142 �+|6� 43.472
R82 VDD.n132 0#��U 43.472
R83 VDD.n20 VDD.n15 41.052
R84 VDD.n72 VDD.n70 39.742
R85 VDD.n72 VDD.n71 39.742
R86 VDD.n74 VDD.n73 39.742
R87 VDD.n210 VDD.n209 39.742
R88 VDD.n124 VDD.n123 39.742
R89 VDD.n158 VDD.n155 39.742
R90 VDD.n158 VDD.n157 39.742
R91 VDD.n154 VDD.n153 39.742
R92 VDD.n219 VDD.n218 38
R93 VDD.n111 VDD.n110 38
R94 VDD.n217 VDD.n216 36.774
R95 VDD.n70 VDD.n69 36.774
R96 VDD.n157 VDD.n156 36.774
R97 VDD.n1 VDD.n0 30.923
R98 VDD.n77 VDD.n75 26.38
R99 VDD.n77 VDD.n74 26.38
R100 VDD.n77 VDD.n72 26.38
R101 VDD.n77 VDD.n76 26.38
R102 VDD.n213 VDD.n211 26.38
R103 VDD.n213 VDD.n210 26.38
R104 VDD.n213 VDD.n212 26.38
R105 VDD.n127 VDD.n125 26.38
R106 VDD.n127 VDD.n124 26.38
R107 VDD.n127 VDD.n126 26.38
R108 VDD.n159 VDD.n158 26.38
R109 VDD.n159 VDD.n154 26.38
R110 VDD.n159 VDD.n152 26.38
R111 VDD.n159 VDD.n151 26.38
R112 VDD.n130 VDD.n122 22.915
R113 VDD.n23 VDD.n14 22.915
R114 VDD.n29 �+|6� 20.457
R115 VDD.n87 �!���U 20.457
R116 VDD.n195  ,|6� 20.457
R117 VDD.n42  ,|6� 17.9
R118 VDD.n100 VDD.t12 17.9
R119 VDD.n182  ���U 17.9
R120 VDD.n122 VDD.n120 14.864
R121 VDD.n120 VDD.n118 14.864
R122 VDD.n118 VDD.n116 14.864
R123 VDD.n116 VDD.n114 14.864
R124 VDD.n114 VDD.n112 14.864
R125 VDD.n230 VDD.n228 14.864
R126 VDD.n228 VDD.n226 14.864
R127 VDD.n226 VDD.n224 14.864
R128 VDD.n224 VDD.n222 14.864
R129 VDD.n222 VDD.n220 14.864
R130 VDD.n66 VDD.n64 14.864
R131 VDD.n64 VDD.n62 14.864
R132 VDD.n62 VDD.n60 14.864
R133 VDD.n60 VDD.n58 14.864
R134 VDD.n58 VDD.n56 14.864
R135 VDD.n56 VDD.n55 14.864
R136 VDD.n173 VDD.n171 14.864
R137 VDD.n171 VDD.n169 14.864
R138 VDD.n169 VDD.n167 14.864
R139 VDD.n167 VDD.n165 14.864
R140 VDD.n165 VDD.n163 14.864
R141 VDD.n163 VDD.n162 14.864
R142 VDD.n14 VDD.n13 14.864
R143 VDD.n13 VDD.n11 14.864
R144 VDD.n11 VDD.n9 14.864
R145 VDD.n9 VDD.n7 14.864
R146 VDD.n7 VDD.n5 14.864
R147 VDD.n80 VDD.n67 14.864
R148 VDD.n232 VDD.n231 14.864
R149 VDD.n175 VDD.n174 14.864
R150 VDD.n191 VDD.t9 14.282
R151 VDD.n191 VDD.t27 14.282
R152 VDD.n92 VDD.t3 14.282
R153 VDD.n92 VDD.t15 14.282
R154 VDD.n34 VDD.t17 14.282
R155 VDD.n34 VDD.t7 14.282
R156 VDD.n36 VDD.n35 9.083
R157 VDD.n94 VDD.n93 9.083
R158 VDD.n193 VDD.n192 9.083
R159 VDD.n23 VDD.n22 8.855
R160 VDD.n22 VDD.n21 8.855
R161 VDD.n27 VDD.n25 8.855
R162 VDD.n25 VDD.n24 8.855
R163 VDD.n31 VDD.n30 8.855
R164 VDD.n30 VDD.n29 8.855
R165 VDD.n36 VDD.n33 8.855
R166 VDD.n33 �+|6� 8.855
R167 VDD.n40 VDD.n39 8.855
R168 VDD.n39 VDD.n38 8.855
R169 VDD.n44 VDD.n43 8.855
R170 VDD.n43 VDD.n42 8.855
R171 VDD.n49 VDD.n48 8.855
R172 VDD.n48 VDD.n47 8.855
R173 VDD.n53 VDD.n52 8.855
R174 VDD.n52 VDD.n51 8.855
R175 VDD.n80 VDD.n79 8.855
R176 VDD.n79 VDD.n78 8.855
R177 VDD.n85 VDD.n83 8.855
R178 VDD.n83 VDD.n82 8.855
R179 VDD.n89 VDD.n88 8.855
R180 VDD.n88 VDD.n87 8.855
R181 VDD.n94 VDD.n91 8.855
R182 VDD.n91  ,|6� 8.855
R183 VDD.n98 VDD.n97 8.855
R184 VDD.n97 VDD.n96 8.855
R185 VDD.n102 VDD.n101 8.855
R186 VDD.n101 VDD.n100 8.855
R187 VDD.n107 VDD.n106 8.855
R188 VDD.n106 VDD.n105 8.855
R189 VDD.n232 VDD.n215 8.855
R190 VDD.n215 VDD.n214 8.855
R191 VDD.n206 VDD.n205 8.855
R192 VDD.n205 VDD.n204 8.855
R193 VDD.n202 VDD.n200 8.855
R194 VDD.n200 VDD.n199 8.855
R195 VDD.n197 VDD.n196 8.855
R196 VDD.n196 VDD.n195 8.855
R197 VDD.n193 VDD.n190 8.855
R198 VDD.n190  ����U 8.855
R199 VDD.n188 VDD.n187 8.855
R200 VDD.n187 VDD.n186 8.855
R201 VDD.n184 VDD.n183 8.855
R202 VDD.n183 VDD.n182 8.855
R203 VDD.n180 VDD.n179 8.855
R204 VDD.n179 VDD.n178 8.855
R205 VDD.n175 VDD.n161 8.855
R206 VDD.n161 VDD.n160 8.855
R207 VDD.n148 VDD.n147 8.855
R208 VDD.n147 VDD.n146 8.855
R209 VDD.n144 VDD.n143 8.855
R210 VDD.n143 VDD.n142 8.855
R211 VDD.n139 VDD.n138 8.855
R212 VDD.n138 VDD.n137 8.855
R213 VDD.n135 VDD.n133 8.855
R214 VDD.n133 VDD.n132 8.855
R215 VDD.n130 VDD.n129 8.855
R216 VDD.n129 VDD.n128 8.855
R217 VDD.n231 VDD.n230 8.051
R218 VDD.n67 VDD.n66 8.051
R219 VDD.n174 VDD.n173 8.051
R220 VDD.n32 VDD.n31 4.65
R221 VDD.n37 VDD.n36 4.65
R222 VDD.n41 VDD.n40 4.65
R223 VDD.n45 VDD.n44 4.65
R224 VDD.n50 VDD.n49 4.65
R225 VDD.n54 VDD.n53 4.65
R226 VDD.n81 VDD.n80 4.65
R227 VDD.n86 VDD.n85 4.65
R228 VDD.n90 VDD.n89 4.65
R229 VDD.n95 VDD.n94 4.65
R230 VDD.n99 VDD.n98 4.65
R231 VDD.n103 VDD.n102 4.65
R232 VDD.n108 VDD.n107 4.65
R233 VDD.n233 VDD.n232 4.65
R234 VDD.n207 VDD.n206 4.65
R235 VDD.n203 VDD.n202 4.65
R236 VDD.n198 VDD.n197 4.65
R237 VDD.n194 VDD.n193 4.65
R238 VDD.n189 VDD.n188 4.65
R239 VDD.n185 VDD.n184 4.65
R240 VDD.n181 VDD.n180 4.65
R241 VDD.n176 VDD.n175 4.65
R242 VDD.n149 VDD.n148 4.65
R243 VDD.n145 VDD.n144 4.65
R244 VDD.n140 VDD.n139 4.65
R245 VDD.n136 VDD.n135 4.65
R246 VDD.n131 VDD.n130 4.65
R247 VDD.n28 VDD.n23 2.933
R248 VDD.n49 VDD.n46 2.89
R249 VDD.n107 VDD.n104 2.89
R250 VDD.n180 VDD.n177 2.89
R251 VDD.n28 VDD.n27 2.844
R252 VDD.n38 �+|6� 2.557
R253 VDD.n96 @d%��U 2.557
R254 VDD.n186  ,|6� 2.557
R255 VDD.n27 VDD.n26 2.477
R256 VDD.n85 VDD.n84 2.477
R257 VDD.n202 VDD.n201 2.477
R258 VDD.n144 VDD.n141 2.064
R259 VDD.n135 VDD.n134 2.064
R260 VDD.n32 VDD.n28 1.063
R261 VDD.n81 VDD.n54 0.29
R262 VDD.n233 VDD.n207 0.29
R263 VDD.n176 VDD.n149 0.29
R264 VDD.n131 VDD 0.207
R265 VDD.n41 VDD.n37 0.181
R266 VDD.n99 VDD.n95 0.181
R267 VDD.n194 VDD.n189 0.181
R268 VDD.n145 VDD.n140 0.157
R269 VDD.n140 VDD.n136 0.157
R270 VDD.n37 VDD.n32 0.145
R271 VDD.n45 VDD.n41 0.145
R272 VDD.n50 VDD.n45 0.145
R273 VDD.n54 VDD.n50 0.145
R274 VDD.n86 VDD.n81 0.145
R275 VDD.n90 VDD.n86 0.145
R276 VDD.n95 VDD.n90 0.145
R277 VDD.n103 VDD.n99 0.145
R278 VDD.n108 VDD.n103 0.145
R279 VDD.n207 VDD.n203 0.145
R280 VDD.n203 VDD.n198 0.145
R281 VDD.n198 VDD.n194 0.145
R282 VDD.n189 VDD.n185 0.145
R283 VDD.n185 VDD.n181 0.145
R284 VDD.n181 VDD.n176 0.145
R285 VDD.n149 VDD.n145 0.145
R286 VDD.n136 VDD.n131 0.145
R287 VDD VDD.n233 0.078
R288 VDD VDD.n108 0.066
R289 S.n2 S.t5 512.525
R290 S.n0 S.t4 480.392
R291 S.n0 S.t3 403.272
R292 S.n2 S.t0 371.139
R293 S.n1 S.t1 301.486
R294 S.n3 S.n2 275.206
R295 S.n3 S.t2 254.993
R296 S.n1 S.n0 227.006
R297 S.n4 S.n1 6.509
R298 S.n4 S.n3 4.65
R299 S.n4 S 0.046
R300 a_1888_101.t0 a_1888_101.n6 93.333
R301 a_1888_101.n5 a_1888_101.n4 51.907
R302 a_1888_101.n5 a_1888_101.n3 51.594
R303 a_1888_101.n2 a_1888_101.n0 41.528
R304 a_1888_101.t0 a_1888_101.n5 38.864
R305 a_1888_101.t0 a_1888_101.n7 8.137
R306 a_1888_101.n2 a_1888_101.n1 3.644
R307 a_1888_101.t0 a_1888_101.n2 1.093
R308 Y.n4 Y.n3 299.461
R309 Y.n4 Y.n2 187.858
R310 Y.n2 Y.n1 157.964
R311 Y.n2 Y.n0 91.706
R312 Y.n0 Y.t3 14.282
R313 Y.n0 Y.t2 14.282
R314 Y.n1 Y.t1 14.282
R315 Y.n1 Y.t0 14.282
R316 Y.n5 Y.n4 4.65
R317 Y.n5 Y 0.046
R318 GND.n84 GND.n83 237.558
R319 GND.n28 GND.n27 237.558
R320 GND.n117 GND.n116 237.558
R321 GND.n25 GND.n24 210.82
R322 GND.n86 GND.n85 210.82
R323 GND.n119 GND.n118 210.82
R324 GND.n14 GND.n13 172.612
R325 GND.n47 GND.n46 151.605
R326 GND.n97 GND.n96 151.605
R327 GND.n64 GND.n63 37.582
R328 GND.t4 GND.n61 32.601
R329 GND.n46 GND.n45 28.421
R330 GND.n96 GND.n95 28.421
R331 GND.n46 GND.n44 25.263
R332 GND.n96 GND.n94 25.263
R333 GND.n44 GND.n43 24.383
R334 GND.n94 GND.n93 24.383
R335 GND.n61 GND.n60 21.734
R336 GND.n76 GND.n75 20.705
R337 GND.n70 GND.n69 20.705
R338 GND.n65 GND.n64 20.705
R339 GND.n75 GND.n74 19.952
R340 GND.n26 GND.n25 18.953
R341 GND.n87 GND.n86 18.953
R342 GND.n120 GND.n119 18.953
R343 GND.n63 GND.t4 15.644
R344 GND.n29 GND.n26 14.864
R345 GND.n121 GND.n120 14.864
R346 GND.n88 GND.n87 14.864
R347 GND.n63 GND.n62 13.541
R348 GND.n66 GND.n57 9.154
R349 GND.n72 GND.n71 9.154
R350 GND.n78 GND.n77 9.154
R351 GND.n81 GND.n80 9.154
R352 GND.n88 GND.n84 9.154
R353 GND.n91 GND.n90 9.154
R354 GND.n99 GND.n98 9.154
R355 GND.n102 GND.n101 9.154
R356 GND.n105 GND.n104 9.154
R357 GND.n108 GND.n107 9.154
R358 GND.n111 GND.n110 9.154
R359 GND.n114 GND.n113 9.154
R360 GND.n121 GND.n117 9.154
R361 GND.n52 GND.n51 9.154
R362 GND.n49 GND.n48 9.154
R363 GND.n41 GND.n40 9.154
R364 GND.n38 GND.n37 9.154
R365 GND.n35 GND.n34 9.154
R366 GND.n32 GND.n31 9.154
R367 GND.n29 GND.n28 9.154
R368 GND.n22 GND.n21 9.154
R369 GND.n19 GND.n18 9.154
R370 GND.n16 GND.n15 9.154
R371 GND.n11 GND.n10 9.154
R372 GND.n8 GND.n7 9.154
R373 GND.n5 GND.n4 9.154
R374 GND.n2 GND.n1 9.154
R375 GND.n56 GND.n55 4.65
R376 GND.n6 GND.n5 4.65
R377 GND.n9 GND.n8 4.65
R378 GND.n12 GND.n11 4.65
R379 GND.n17 GND.n16 4.65
R380 GND.n20 GND.n19 4.65
R381 GND.n23 GND.n22 4.65
R382 GND.n30 GND.n29 4.65
R383 GND.n33 GND.n32 4.65
R384 GND.n36 GND.n35 4.65
R385 GND.n39 GND.n38 4.65
R386 GND.n42 GND.n41 4.65
R387 GND.n50 GND.n49 4.65
R388 GND.n53 GND.n52 4.65
R389 GND.n122 GND.n121 4.65
R390 GND.n115 GND.n114 4.65
R391 GND.n112 GND.n111 4.65
R392 GND.n109 GND.n108 4.65
R393 GND.n106 GND.n105 4.65
R394 GND.n103 GND.n102 4.65
R395 GND.n100 GND.n99 4.65
R396 GND.n92 GND.n91 4.65
R397 GND.n89 GND.n88 4.65
R398 GND.n82 GND.n81 4.65
R399 GND.n79 GND.n78 4.65
R400 GND.n73 GND.n72 4.65
R401 GND.n67 GND.n66 4.65
R402 GND.n59 GND.n58 4.504
R403 GND.n16 GND.n14 4.129
R404 GND.n49 GND.n47 4.129
R405 GND.n99 GND.n97 4.129
R406 GND.n78 GND.n76 4.129
R407 GND.n66 GND.n65 3.716
R408 GND.n3 GND.n0 3.407
R409 GND.n3 GND.n2 2.844
R410 GND.t4 GND.n59 2.452
R411 GND.n6 GND.n3 1.063
R412 GND.n55 GND.n54 0.474
R413 GND.n69 GND.n68 0.376
R414 GND.n30 GND.n23 0.29
R415 GND.n122 GND.n115 0.29
R416 GND.n89 GND.n82 0.29
R417 GND.n56 GND 0.207
R418 GND.n72 GND.n70 0.206
R419 GND.n12 GND.n9 0.181
R420 GND.n42 GND.n39 0.181
R421 GND.n106 GND.n103 0.181
R422 GND.n79 GND.n73 0.157
R423 GND.n73 GND.n67 0.157
R424 GND.n9 GND.n6 0.145
R425 GND.n17 GND.n12 0.145
R426 GND.n20 GND.n17 0.145
R427 GND.n23 GND.n20 0.145
R428 GND.n33 GND.n30 0.145
R429 GND.n36 GND.n33 0.145
R430 GND.n39 GND.n36 0.145
R431 GND.n50 GND.n42 0.145
R432 GND.n53 GND.n50 0.145
R433 GND.n115 GND.n112 0.145
R434 GND.n112 GND.n109 0.145
R435 GND.n109 GND.n106 0.145
R436 GND.n103 GND.n100 0.145
R437 GND.n100 GND.n92 0.145
R438 GND.n92 GND.n89 0.145
R439 GND.n82 GND.n79 0.145
R440 GND.n67 GND.n56 0.145
R441 GND GND.n122 0.078
R442 GND GND.n53 0.066
R443 A0.n0 A0.t2 472.359
R444 A0.n0 A0.t0 384.527
R445 A0.n1 A0.t1 314.896
R446 A0.n1 A0.n0 182.814
R447 A0.n2 A0.n1 4.65
R448 A0.n2 A0 0.046
R449 a_661_1050.n0 a_661_1050.t5 480.392
R450 a_661_1050.n0 a_661_1050.t6 403.272
R451 a_661_1050.n1 a_661_1050.t7 301.486
R452 a_661_1050.n6 a_661_1050.n5 249.863
R453 a_661_1050.n1 a_661_1050.n0 227.006
R454 a_661_1050.n8 a_661_1050.n6 215.717
R455 a_661_1050.n8 a_661_1050.n7 157.964
R456 a_661_1050.n9 a_661_1050.n8 91.705
R457 a_661_1050.n5 a_661_1050.n4 30
R458 a_661_1050.n3 a_661_1050.n2 24.383
R459 a_661_1050.n5 a_661_1050.n3 23.684
R460 a_661_1050.n7 a_661_1050.t3 14.282
R461 a_661_1050.n7 a_661_1050.t4 14.282
R462 a_661_1050.n9 a_661_1050.t1 14.282
R463 a_661_1050.t2 a_661_1050.n9 14.282
R464 a_661_1050.n6 a_661_1050.n1 13.063
R465 a_556_101.n3 a_556_101.n1 42.788
R466 a_556_101.t0 a_556_101.n0 8.137
R467 a_556_101.n3 a_556_101.n2 4.665
R468 a_556_101.t0 a_556_101.n3 0.06
R469 A1.n0 A1.t0 472.359
R470 A1.n0 A1.t2 384.527
R471 A1.n1 A1.t1 342.755
R472 A1.n1 A1.n0 154.955
R473 A1.n2 A1.n1 4.65
R474 A1.n2 A1 0.046
R475 a_1222_101.n11 a_1222_101.n10 68.43
R476 a_1222_101.n3 a_1222_101.n2 62.817
R477 a_1222_101.n7 a_1222_101.n6 38.626
R478 a_1222_101.n6 a_1222_101.n5 35.955
R479 a_1222_101.n3 a_1222_101.n1 26.202
R480 a_1222_101.t0 a_1222_101.n3 19.737
R481 a_1222_101.t1 a_1222_101.n8 8.137
R482 a_1222_101.t0 a_1222_101.n4 7.273
R483 a_1222_101.t0 a_1222_101.n0 6.109
R484 a_1222_101.t1 a_1222_101.n7 4.864
R485 a_1222_101.t0 a_1222_101.n12 2.074
R486 a_1222_101.n12 a_1222_101.t1 0.937
R487 a_1222_101.t1 a_1222_101.n11 0.763
R488 a_1222_101.n11 a_1222_101.n9 0.185
C5 S GND 0.86fF
C6 VDD GND 4.01fF
C7 a_1222_101.n0 GND 0.02fF
C8 a_1222_101.n1 GND 0.09fF
C9 a_1222_101.n2 GND 0.08fF
C10 a_1222_101.n3 GND 0.03fF
C11 a_1222_101.n4 GND 0.01fF
C12 a_1222_101.n5 GND 0.04fF
C13 a_1222_101.n6 GND 0.04fF
C14 a_1222_101.n7 GND 0.02fF
C15 a_1222_101.n8 GND 0.05fF
C16 a_1222_101.n9 GND 0.15fF
C17 a_1222_101.n10 GND 0.08fF
C18 a_1222_101.n11 GND 0.08fF
C19 a_1222_101.t1 GND 0.23fF
C20 a_1222_101.n12 GND 0.01fF
C21 a_556_101.n0 GND 0.05fF
C22 a_556_101.n1 GND 0.12fF
C23 a_556_101.n2 GND 0.04fF
C24 a_556_101.n3 GND 0.17fF
C25 a_661_1050.n0 GND 0.37fF
C26 a_661_1050.n1 GND 0.83fF
C27 a_661_1050.n2 GND 0.04fF
C28 a_661_1050.n3 GND 0.05fF
C29 a_661_1050.n4 GND 0.03fF
C30 a_661_1050.n5 GND 0.16fF
C31 a_661_1050.n6 GND 0.90fF
C32 a_661_1050.n7 GND 0.47fF
C33 a_661_1050.n8 GND 0.61fF
C34 a_661_1050.n9 GND 0.37fF
C35 Y.n0 GND 0.34fF
C36 Y.n1 GND 0.43fF
C37 Y.n2 GND 0.53fF
C38 Y.n3 GND 0.27fF
C39 Y.n4 GND 0.45fF
C40 Y.n5 GND 0.01fF
C41 a_1888_101.n0 GND 0.08fF
C42 a_1888_101.n1 GND 0.02fF
C43 a_1888_101.n2 GND 0.02fF
C44 a_1888_101.n3 GND 0.09fF
C45 a_1888_101.n4 GND 0.07fF
C46 a_1888_101.n5 GND 0.04fF
C47 a_1888_101.n6 GND 0.02fF
C48 a_1888_101.n7 GND 0.05fF
C49 S.n0 GND 0.28fF
C50 S.n1 GND 0.36fF
C51 S.n2 GND 0.28fF
C52 S.t2 GND 0.36fF
C53 S.n3 GND 0.32fF
C54 S.n4 GND 0.29fF
C55 VDD.n1 GND 0.03fF
C56 VDD.n2 GND 0.11fF
C57 VDD.n3 GND 0.02fF
C58 VDD.n4 GND 0.02fF
C59 VDD.n5 GND 0.05fF
C60 VDD.n6 GND 0.02fF
C61 VDD.n7 GND 0.02fF
C62 VDD.n8 GND 0.02fF
C63 VDD.n9 GND 0.02fF
C64 VDD.n10 GND 0.02fF
C65 VDD.n11 GND 0.02fF
C66 VDD.n12 GND 0.02fF
C67 VDD.n13 GND 0.02fF
C68 VDD.n14 GND 0.03fF
C69 VDD.n15 GND 0.01fF
C70 VDD.n20 GND 0.36fF
C71 VDD.n21 GND 0.21fF
C72 VDD.n22 GND 0.02fF
C73 VDD.n23 GND 0.03fF
C74 VDD.n24 GND 0.19fF
C75 VDD.n25 GND 0.01fF
C76 VDD.n26 GND 0.05fF
C77 VDD.n27 GND 0.01fF
C78 VDD.n28 GND 0.01fF
C79 VDD.n29 GND 0.13fF
C80 VDD.n30 GND 0.01fF
C81 VDD.n31 GND 0.02fF
C82 VDD.n32 GND 0.06fF
C83 VDD.n33 GND 0.01fF
C84 VDD.n34 GND 0.06fF
C85 VDD.n35 GND 0.04fF
C86 VDD.n36 GND 0.01fF
C87 VDD.n37 GND 0.02fF
C88 VDD.n38 GND 0.11fF
C89 VDD.n39 GND 0.01fF
C90 VDD.n40 GND 0.01fF
C91 VDD.n41 GND 0.02fF
C92 VDD.n42 GND 0.13fF
C93 VDD.n43 GND 0.01fF
C94 VDD.n44 GND 0.02fF
C95 VDD.n45 GND 0.02fF
C96 VDD.n46 GND 0.05fF
C97 VDD.n47 GND 0.19fF
C98 VDD.n48 GND 0.01fF
C99 VDD.n49 GND 0.01fF
C100 VDD.n50 GND 0.02fF
C101 VDD.n51 GND 0.21fF
C102 VDD.n52 GND 0.01fF
C103 VDD.n53 GND 0.02fF
C104 VDD.n54 GND 0.03fF
C105 VDD.n55 GND 0.04fF
C106 VDD.n56 GND 0.02fF
C107 VDD.n57 GND 0.02fF
C108 VDD.n58 GND 0.02fF
C109 VDD.n59 GND 0.02fF
C110 VDD.n60 GND 0.02fF
C111 VDD.n61 GND 0.02fF
C112 VDD.n62 GND 0.02fF
C113 VDD.n63 GND 0.02fF
C114 VDD.n64 GND 0.02fF
C115 VDD.n65 GND 0.02fF
C116 VDD.n66 GND 0.01fF
C117 VDD.n67 GND 0.02fF
C118 VDD.n68 GND 0.02fF
C119 VDD.n69 GND 0.17fF
C120 VDD.n70 GND 0.02fF
C121 VDD.n71 GND 0.02fF
C122 VDD.n73 GND 0.02fF
C123 VDD.n77 GND 0.21fF
C124 VDD.n78 GND 0.21fF
C125 VDD.n79 GND 0.01fF
C126 VDD.n80 GND 0.02fF
C127 VDD.n81 GND 0.03fF
C128 VDD.n82 GND 0.19fF
C129 VDD.n83 GND 0.01fF
C130 VDD.n84 GND 0.05fF
C131 VDD.n85 GND 0.01fF
C132 VDD.n86 GND 0.02fF
C133 VDD.n87 GND 0.13fF
C134 VDD.n88 GND 0.01fF
C135 VDD.n89 GND 0.02fF
C136 VDD.n90 GND 0.02fF
C137 VDD.n91 GND 0.01fF
C138 VDD.n92 GND 0.06fF
C139 VDD.n93 GND 0.04fF
C140 VDD.n94 GND 0.01fF
C141 VDD.n95 GND 0.02fF
C142 VDD.n96 GND 0.11fF
C143 VDD.n97 GND 0.01fF
C144 VDD.n98 GND 0.01fF
C145 VDD.n99 GND 0.02fF
C146 VDD.n100 GND 0.13fF
C147 VDD.n101 GND 0.01fF
C148 VDD.n102 GND 0.02fF
C149 VDD.n103 GND 0.02fF
C150 VDD.n104 GND 0.05fF
C151 VDD.n105 GND 0.19fF
C152 VDD.n106 GND 0.01fF
C153 VDD.n107 GND 0.01fF
C154 VDD.n108 GND 0.01fF
C155 VDD.n109 GND 0.08fF
C156 VDD.n110 GND 0.02fF
C157 VDD.n111 GND 0.01fF
C158 VDD.n112 GND 0.05fF
C159 VDD.n113 GND 0.02fF
C160 VDD.n114 GND 0.02fF
C161 VDD.n115 GND 0.02fF
C162 VDD.n116 GND 0.02fF
C163 VDD.n117 GND 0.02fF
C164 VDD.n118 GND 0.02fF
C165 VDD.n119 GND 0.02fF
C166 VDD.n120 GND 0.02fF
C167 VDD.n121 GND 0.03fF
C168 VDD.n122 GND 0.03fF
C169 VDD.n123 GND 0.02fF
C170 VDD.n127 GND 0.36fF
C171 VDD.n128 GND 0.21fF
C172 VDD.n129 GND 0.02fF
C173 VDD.n130 GND 0.02fF
C174 VDD.n131 GND 0.02fF
C175 VDD.n132 GND 0.16fF
C176 VDD.n133 GND 0.01fF
C177 VDD.n134 GND 0.05fF
C178 VDD.n135 GND 0.01fF
C179 VDD.n136 GND 0.02fF
C180 VDD.n