magic
tech sky130
magscale 1 2
timestamp 1645050501
<< locali >>
rect 17 -17 49 17
<< viali >>
rect -17 -17 17 17
<< metal1 >>
rect -17 23 17 29
rect -23 17 23 23
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -23 23 -17
rect -17 -53 17 -23
<< end >>
