magic
tech sky130A
magscale 1 2
timestamp 1648490770
<< nwell >>
rect 55 1505 89 1539
<< psubdiffcont >>
rect 55 13 89 47
<< nsubdiffcont >>
rect 55 1505 89 1539
<< viali >>
rect 55 1505 89 1539
rect 55 13 89 47
<< metal1 >>
rect 4235 945 15915 979
rect 427 797 13414 831
rect 17817 797 17851 831
rect 15411 723 16694 757
rect 1604 649 14368 683
rect 9451 501 15707 535
rect 1353 427 11782 461
use dffrnqx1_pcell  dffrnqx1_pcell_0 pcells
timestamp 1648484181
transform 1 0 0 0 1 0
box -84 0 5264 1575
use dffrnqx1_pcell  dffrnqx1_pcell_1
timestamp 1648484181
transform 1 0 5180 0 1 0
box -84 0 5264 1575
use li1_M1_contact  li1_M1_contact_14 pcells
timestamp 1648061256
transform -1 0 4218 0 -1 962
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform -1 0 5032 0 -1 962
box -53 -33 29 33
use dffrnqx1_pcell  dffrnqx1_pcell_2
timestamp 1648484181
transform 1 0 10360 0 1 0
box -84 0 5264 1575
use li1_M1_contact  li1_M1_contact_13
timestamp 1648061256
transform 1 0 10212 0 1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform -1 0 9398 0 -1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_6
timestamp 1648061256
transform 1 0 15910 0 -1 962
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_15
timestamp 1648061256
transform -1 0 15392 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_12
timestamp 1648061256
transform 1 0 16724 0 -1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_16
timestamp 1648061256
transform -1 0 17834 0 -1 814
box -53 -33 29 33
use voter3x1_pcell  voter3x1_pcell_0 pcells
timestamp 1648490579
transform 1 0 15540 0 1 0
box -84 0 2526 1575
<< labels >>
rlabel metal1 17817 797 17851 831 1 Q
port 1 n
rlabel metal1 1389 427 1423 461 1 D
port 2 n
rlabel metal1 427 797 461 831 1 CLK
port 3 n
rlabel metal1 1611 649 1645 683 1 RN
port 4 n
rlabel metal1 72 1522 72 1522 1 VDD
port 5 n
rlabel metal1 72 30 72 30 1 VSS
port 6 n
<< end >>
