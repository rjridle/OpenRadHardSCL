magic
tech sky130A
magscale 1 2
timestamp 1645649939
<< nmos >>
rect 19 210 49 272
rect 19 180 125 210
tri 125 180 155 210 sw
rect 19 80 49 180
tri 49 164 65 180 nw
tri 109 164 125 180 ne
tri 49 80 65 96 sw
tri 109 80 125 96 se
rect 125 80 155 180
tri 19 50 49 80 ne
rect 49 50 125 80
tri 125 50 155 80 nw
<< ndiff >>
rect -37 256 19 272
rect -37 222 -27 256
rect 7 222 19 256
rect -37 185 19 222
rect 49 256 211 272
rect 49 222 65 256
rect 99 222 167 256
rect 201 222 211 256
rect 49 210 211 222
rect -37 151 -27 185
rect 7 151 19 185
tri 125 180 155 210 ne
rect 155 185 211 210
rect -37 117 19 151
rect -37 83 -27 117
rect 7 83 19 117
rect -37 50 19 83
tri 49 164 65 180 se
rect 65 164 109 180
tri 109 164 125 180 sw
rect 49 140 125 164
rect 49 106 70 140
rect 104 106 125 140
rect 49 96 125 106
tri 49 80 65 96 ne
rect 65 80 109 96
tri 109 80 125 96 nw
rect 155 151 167 185
rect 201 151 211 185
rect 155 117 211 151
rect 155 83 167 117
rect 201 83 211 117
tri 19 50 49 80 sw
tri 125 50 155 80 se
rect 155 50 211 83
rect -37 46 211 50
rect -37 12 -27 46
rect 7 12 167 46
rect 201 12 211 46
rect -37 -4 211 12
<< ndiffc >>
rect -27 222 7 256
rect 65 222 99 256
rect 167 222 201 256
rect -27 151 7 185
rect -27 83 7 117
rect 70 106 104 140
rect 167 151 201 185
rect 167 83 201 117
rect -27 12 7 46
rect 167 12 201 46
<< poly >>
rect 19 272 49 298
<< locali >>
rect -27 256 7 272
rect 167 256 201 272
rect 7 222 65 256
rect 99 222 167 256
rect -27 185 7 222
rect 167 185 201 222
rect -27 117 7 151
rect 70 140 104 156
rect 70 90 104 106
rect 167 117 201 151
rect -27 46 7 83
rect -27 -4 7 12
rect 167 46 201 83
rect 167 -4 201 12
<< end >>
