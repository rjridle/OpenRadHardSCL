* SPICE3 file created from VOTER3X1.ext - technology: sky130A

.subckt VOTER3X1 Y A B C VDD GND
X0 Y.t2 a_392_209.t7 VDD.t18  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X1 GND B.t1 a_778_101.t0 GND sky130_fd_pr__nfet_01v8 ad=1.6781p pd=1.281u as=0p ps=0u w=0u l=0u
X2 GND B.t2 a_112_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X3 GND C.t1 a_1444_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X4 a_392_209.t0 A.t0 a_881_1051.t7 �a�u�U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X5 VDD.t1 B.t0 a_217_1051.t3 |u�U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X6 VDD.t16 a_392_209.t8 Y.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X7 a_881_1051.t4 C.t0 a_217_1051.t1 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X8 VDD.t8 A.t1 a_217_1051.t7  �x�7 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X9 a_881_1051.t0 B.t3 a_217_1051.t5 ��x�7 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X10 a_881_1051.t3 C.t2 a_392_209.t5  �x�7 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X11 Y a_392_209.t9 GND.t0 GND sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=0p ps=0u w=0u l=0u
X12 a_217_1051.t2 B.t4 VDD.t3 ��x�7 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X13 a_217_1051.t4 B.t5 a_881_1051.t2  �x�7 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X14 a_217_1051.t6 A.t4 VDD.t11 ��x�7 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X15 a_881_1051.t6 A.t5 a_392_209.t1  �x�7 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X16 a_217_1051.t0 C.t4 a_881_1051.t1 ��x�7 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X17 a_392_209.t6 C.t5 a_881_1051.t5  �x�7 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
C0 VDD A 1.95fF
C1 B VDD 1.14fF
C2 A C 0.26fF
C3 B C 0.15fF
C4 B A 0.96fF
C5 VDD Y 1.06fF
C6 VDD C 0.73fF
R0 a_392_209.n3 a_392_209.t8 512.525
R1 a_392_209.n3 a_392_209.t7 371.139
R2 a_392_209.n4 a_392_209.t9 338.57
R3 a_392_209.n13 a_392_209.n5 227.387
R4 a_392_209.n4 a_392_209.n3 191.629
R5 a_392_209.n2 a_392_209.n1 165.613
R6 a_392_209.n5 a_392_209.n2 132.893
R7 a_392_209.n12 a_392_209.n11 128.294
R8 a_392_209.n12 a_392_209.n8 126.225
R9 a_392_209.n15 a_392_209.n13 112.91
R10 a_392_209.n2 a_392_209.n0 99.355
R11 a_392_209.n8 a_392_209.n7 22.578
R12 a_392_209.n11 a_392_209.n10 22.578
R13 a_392_209.n15 a_392_209.n14 15.001
R14 a_392_209.n0 a_392_209.t1 14.282
R15 a_392_209.n0 a_392_209.t0 14.282
R16 a_392_209.n1 a_392_209.t5 14.282
R17 a_392_209.n1 a_392_209.t6 14.282
R18 a_392_209.n16 a_392_209.n15 12.632
R19 a_392_209.n5 a_392_209.n4 10.343
R20 a_392_209.n8 a_392_209.n6 8.58
R21 a_392_209.n11 a_392_209.n9 8.58
R22 a_392_209.n13 a_392_209.n12 7.053
R23 VDD.n119 VDD.n112 144.705
R24 VDD.n200 VDD.n189 144.705
R25 VDD.n66 VDD.n55 144.705
R26 VDD.n145 VDD.t3 135.539
R27 VDD.n167 VDD.t8 135.539
R28 VDD.n35 VDD.t18 135.17
R29 VDD.n24 VDD.t16 135.17
R30 VDD.n159 VDD.n158 129.849
R31 VDD.n51 VDD.n50 92.5
R32 VDD.n49 VDD.n48 92.5
R33 VDD.n47 VDD.n46 92.5
R34 VDD.n45 VDD.n44 92.5
R35 VDD.n53 VDD.n52 92.5
R36 VDD.n108 VDD.n107 92.5
R37 VDD.n106 VDD.n105 92.5
R38 VDD.n104 VDD.n103 92.5
R39 VDD.n102 VDD.n101 92.5
R40 VDD.n110 VDD.n109 92.5
R41 VDD.n185 VDD.n184 92.5
R42 VDD.n183 VDD.n182 92.5
R43 VDD.n181 VDD.n180 92.5
R44 VDD.n179 VDD.n178 92.5
R45 VDD.n187 VDD.n186 92.5
R46 VDD.n133 VDD.n132 92.5
R47 VDD.n131 VDD.n130 92.5
R48 VDD.n129 VDD.n128 92.5
R49 VDD.n127 VDD.n126 92.5
R50 VDD.n135 VDD.n134 92.5
R51 VDD.n14 VDD.n1 92.5
R52 VDD.n5 VDD.n4 92.5
R53 VDD.n7 VDD.n6 92.5
R54 VDD.n9 VDD.n8 92.5
R55 VDD.n11 VDD.n10 92.5
R56 VDD.n13 VDD.n12 92.5
R57 VDD.n21 VDD.n20 92.059
R58 VDD.n65 VDD.n64 92.059
R59 VDD.n118 VDD.n117 92.059
R60 VDD.n199 VDD.n198 92.059
R61 VDD.n141 VDD.n140 92.059
R62 VDD.n20 VDD.n16 67.194
R63 VDD.n20 VDD.n17 67.194
R64 VDD.n20 VDD.n18 67.194
R65 VDD.n20 VDD.n19 67.194
R66 VDD.n125 VDD.n124 44.141
R67 VDD.n100 VDD.n99 44.141
R68 VDD.n5 VDD.n3 44.141
R69 VDD.n99 VDD.n97 44.107
R70 VDD.n124 VDD.n122 44.107
R71 VDD.n3 VDD.n2 44.107
R72 VDD.n25  43.472
R73 VDD.n33  43.472
R74 VDD.n20 VDD.n15 41.052
R75 VDD.n59 VDD.n57 39.742
R76 VDD.n59 VDD.n58 39.742
R77 VDD.n61 VDD.n60 39.742
R78 VDD.n114 VDD.n113 39.742
R79 VDD.n137 VDD.n136 39.742
R80 VDD.n197 VDD.n194 39.742
R81 VDD.n197 VDD.n196 39.742
R82 VDD.n193 VDD.n192 39.742
R83 VDD.n99 VDD.n98 38
R84 VDD.n124 VDD.n123 38
R85 VDD.n97 VDD.n96 36.774
R86 VDD.n57 VDD.n56 36.774
R87 VDD.n196 VDD.n195 36.774
R88 VDD.n1 VDD.n0 30.923
R89 VDD.n64 VDD.n62 26.38
R90 VDD.n64 VDD.n61 26.38
R91 VDD.n64 VDD.n59 26.38
R92 VDD.n64 VDD.n63 26.38
R93 VDD.n117 VDD.n115 26.38
R94 VDD.n117 VDD.n114 26.38
R95 VDD.n117 VDD.n116 26.38
R96 VDD.n140 VDD.n138 26.38
R97 VDD.n140 VDD.n137 26.38
R98 VDD.n140 VDD.n139 26.38
R99 VDD.n198 VDD.n197 26.38
R100 VDD.n198 VDD.n193 26.38
R101 VDD.n198 VDD.n191 26.38
R102 VDD.n198 VDD.n190 26.38
R103 VDD.n143 VDD.n135 22.915
R104 VDD.n23 VDD.n14 22.915
R105 VDD.n73  �x�7 20.457
R106 VDD.n207 ��x�7 20.457
R107 VDD.n163  �x�7 20.457
R108 VDD.n84  �x�7 17.9
R109 VDD.n218 ��x�7 17.9
R110 VDD.n150 ��x�7 17.9
R111 VDD.n135 VDD.n133 14.864
R112 VDD.n133 VDD.n131 14.864
R113 VDD.n131 VDD.n129 14.864
R114 VDD.n129 VDD.n127 14.864
R115 VDD.n127 VDD.n125 14.864
R116 VDD.n110 VDD.n108 14.864
R117 VDD.n108 VDD.n106 14.864
R118 VDD.n106 VDD.n104 14.864
R119 VDD.n104 VDD.n102 14.864
R120 VDD.n102 VDD.n100 14.864
R121 VDD.n53 VDD.n51 14.864
R122 VDD.n51 VDD.n49 14.864
R123 VDD.n49 VDD.n47 14.864
R124 VDD.n47 VDD.n45 14.864
R125 VDD.n45 VDD.n43 14.864
R126 VDD.n43 VDD.n42 14.864
R127 VDD.n187 VDD.n185 14.864
R128 VDD.n185 VDD.n183 14.864
R129 VDD.n183 VDD.n181 14.864
R130 VDD.n181 VDD.n179 14.864
R131 VDD.n179 VDD.n177 14.864
R132 VDD.n177 VDD.n176 14.864
R133 VDD.n14 VDD.n13 14.864
R134 VDD.n13 VDD.n11 14.864
R135 VDD.n11 VDD.n9 14.864
R136 VDD.n9 VDD.n7 14.864
R137 VDD.n7 VDD.n5 14.864
R138 VDD.n67 VDD.n54 14.864
R139 VDD.n120 VDD.n111 14.864
R140 VDD.n201 VDD.n188 14.864
R141 VDD.n158 VDD.t11 14.282
R142 VDD.n158 VDD.t1 14.282
R143 VDD.n161 VDD.n159 9.083
R144 VDD.n23 VDD.n22 8.855
R145 VDD.n22 VDD.n21 8.855
R146 VDD.n27 VDD.n26 8.855
R147 VDD.n26 VDD.n25 8.855
R148 VDD.n31 VDD.n30 8.855
R149 VDD.n30 VDD.n29 8.855
R150 VDD.n36 VDD.n34 8.855
R151 VDD.n34 VDD.n33 8.855
R152 VDD.n40 VDD.n39 8.855
R153 VDD.n39 VDD.n38 8.855
R154 VDD.n67 VDD.n66 8.855
R155 VDD.n66 VDD.n65 8.855
R156 VDD.n71 VDD.n70 8.855
R157 VDD.n70 VDD.n69 8.855
R158 VDD.n75 VDD.n74 8.855
R159 VDD.n74 VDD.n73 8.855
R160 VDD.n78 VDD.n77 8.855
R161 VDD.n77 �a�u�U 8.855
R162 VDD.n82 VDD.n81 8.855
R163 VDD.n81 VDD.n80 8.855
R164 VDD.n86 VDD.n85 8.855
R165 VDD.n85 VDD.n84 8.855
R166 VDD.n90 VDD.n89 8.855
R167 VDD.n89 VDD.n88 8.855
R168 VDD.n94 VDD.n93 8.855
R169 VDD.n93 VDD.n92 8.855
R170 VDD.n120 VDD.n119 8.855
R171 VDD.n119 VDD.n118 8.855
R172 VDD.n224 VDD.n223 8.855
R173 VDD.n223 VDD.n222 8.855
R174 VDD.n220 VDD.n219 8.855
R175 VDD.n219 VDD.n218 8.855
R176 VDD.n216 VDD.n215 8.855
R177 VDD.n215 VDD.n214 8.855
R178 VDD.n212 VDD.n211 8.855
R179 VDD.n211  �x�7 8.855
R180 VDD.n209 VDD.n208 8.855
R181 VDD.n208 VDD.n207 8.855
R182 VDD.n205 VDD.n204 8.855
R183 VDD.n204 VDD.n203 8.855
R184 VDD.n201 VDD.n200 8.855
R185 VDD.n200 VDD.n199 8.855
R186 VDD.n174 VDD.n173 8.855
R187 VDD.n173 VDD.n172 8.855
R188 VDD.n170 VDD.n169 8.855
R189 VDD.n169 VDD.n168 8.855
R190 VDD.n165 VDD.n164 8.855
R191 VDD.n164 VDD.n163 8.855
R192 VDD.n161 VDD.n160 8.855
R193 VDD.n160 ��x�7 8.855
R194 VDD.n156 VDD.n155 8.855
R195 VDD.n155 VDD.n154 8.855
R196 VDD.n152 VDD.n151 8.855
R197 VDD.n151 VDD.n150 8.855
R198 VDD.n148 VDD.n147 8.855
R199 VDD.n147 VDD.n146 8.855
R200 VDD.n143 VDD.n142 8.855
R201 VDD.n142 VDD.n141 8.855
R202 VDD.n111 VDD.n110 8.051
R203 VDD.n54 VDD.n53 8.051
R204 VDD.n188 VDD.n187 8.051
R205 VDD.n28 VDD.n23 4.795
R206 VDD.n28 VDD.n27 4.65
R207 VDD.n32 VDD.n31 4.65
R208 VDD.n37 VDD.n36 4.65
R209 VDD.n41 VDD.n40 4.65
R210 VDD.n68 VDD.n67 4.65
R211 VDD.n72 VDD.n71 4.65
R212 VDD.n76 VDD.n75 4.65
R213 VDD.n79 VDD.n78 4.65
R214 VDD.n83 VDD.n82 4.65
R215 VDD.n87 VDD.n86 4.65
R216 VDD.n91 VDD.n90 4.65
R217 VDD.n95 VDD.n94 4.65
R218 VDD.n121 VDD.n120 4.65
R219 VDD.n225 VDD.n224 4.65
R220 VDD.n221 VDD.n220 4.65
R221 VDD.n217 VDD.n216 4.65
R222 VDD.n213 VDD.n212 4.65
R223 VDD.n210 VDD.n209 4.65
R224 VDD.n206 VDD.n205 4.65
R225 VDD.n202 VDD.n201 4.65
R226 VDD.n175 VDD.n174 4.65
R227 VDD.n171 VDD.n170 4.65
R228 VDD.n166 VDD.n165 4.65
R229 VDD.n162 VDD.n161 4.65
R230 VDD.n157 VDD.n156 4.65
R231 VDD.n153 VDD.n152 4.65
R232 VDD.n149 VDD.n148 4.65
R233 VDD.n144 VDD.n143 4.65
R234 VDD.n148 VDD.n145 2.89
R235 VDD.n80  �x�7 2.557
R236 VDD.n214 VDD.t14 2.557
R237 VDD.n154 |u�U 2.557
R238 VDD.n170 VDD.n167 2.477
R239 VDD.n27 VDD.n24 2.064
R240 VDD.n36 VDD.n35 2.064
R241 VDD.n68 VDD.n41 0.29
R242 VDD.n121 VDD.n95 0.29
R243 VDD.n202 VDD.n175 0.29
R244 VDD.n144 VDD 0.207
R245 VDD.n83 VDD.n79 0.181
R246 VDD.n217 VDD.n213 0.181
R247 VDD.n162 VDD.n157 0.181
R248 VDD.n32 VDD.n28 0.157
R249 VDD.n37 VDD.n32 0.157
R250 VDD.n41 VDD.n37 0.145
R251 VDD.n72 VDD.n68 0.145
R252 VDD.n76 VDD.n72 0.145
R253 VDD.n79 VDD.n76 0.145
R254 VDD.n87 VDD.n83 0.145
R255 VDD.n91 VDD.n87 0.145
R256 VDD.n95 VDD.n91 0.145
R257 VDD.n225 VDD.n221 0.145
R258 VDD.n221 VDD.n217 0.145
R259 VDD.n213 VDD.n210 0.145
R260 VDD.n210 VDD.n206 0.145
R261 VDD.n206 VDD.n202 0.145
R262 VDD.n175 VDD.n171 0.145
R263 VDD.n171 VDD.n166 0.145
R264 VDD.n166 VDD.n162 0.145
R265 VDD.n157 VDD.n153 0.145
R266 VDD.n153 VDD.n149 0.145
R267 VDD.n149 VDD.n144 0.145
R268 VDD VDD.n121 0.078
R269 VDD VDD.n225 0.066
R270 Y.n5 Y.n4 328.545
R271 Y.n5 Y.n0 215.188
R272 Y.n4 Y.n3 30
R273 Y.n2 Y.n1 24.383
R274 Y.n4 Y.n2 23.684
R275 Y.n0 Y.t1 14.282
R276 Y.n0 Y.t2 14.282
R277 Y.n6 Y.n5 4.65
R278 Y.n6 Y 0.046
R279 A.n0 A.t5 475.572
R280 A.n2 A.t1 469.145
R281 A.n2 A.t4 384.527
R282 A.n0 A.t0 384.527
R283 A.n3 A.t3 370.613
R284 A.n1 A.t2 370.613
R285 A.n1 A.n0 128.028
R286 A.n3 A.n2 126.97
R287 A.n4 A.n1 9.501
R288 A.n4 A.n3 4.65
R289 A.n4 A 0.046
R290 a_881_1051.t6 a_881_1051.n5 179.898
R291 a_881_1051.n3 a_881_1051.n2 165.613
R292 a_881_1051.n3 a_881_1051.n1 142.653
R293 a_881_1051.n5 a_881_1051.n4 106.183
R294 a_881_1051.n5 a_881_1051.n0 99.355
R295 a_881_1051.n4 a_881_1051.n3 82.665
R296 a_881_1051.n4 a_881_1051.t5 73.712
R297 a_881_1051.n1 a_881_1051.t1 14.282
R298 a_881_1051.n1 a_881_1051.t4 14.282
R299 a_881_1051.n2 a_881_1051.t2 14.282
R300 a_881_1051.n2 a_881_1051.t0 14.282
R301 a_881_1051.n0 a_881_1051.t7 14.282
R302 a_881_1051.n0 a_881_1051.t3 14.282
R303 B.n2 B.t0 512.525
R304 B.n0 B.t5 477.179
R305 B.n1 B.t1 440.954
R306 B.n3 B.t2 434.527
R307 B.n0 B.t3 406.485
R308 B.n2 B.t4 371.139
R309 B.n3 B.n2 77.972
R310 B.n1 B.n0 21.4
R311 B.n4 B.n1 4.754
R312 B.n4 B.n3 2.079
R313 B.n4 B 0.046
R314 a_217_1051.n2 a_217_1051.t0 179.895
R315 a_217_1051.n5 a_217_1051.n4 157.021
R316 a_217_1051.n4 a_217_1051.n0 124.955
R317 a_217_1051.n3 a_217_1051.n2 106.183
R318 a_217_1051.n2 a_217_1051.n1 99.355
R319 a_217_1051.n4 a_217_1051.n3 82.65
R320 a_217_1051.n3 a_217_1051.t5 73.712
R321 a_217_1051.n0 a_217_1051.t7 14.282
R322 a_217_1051.n0 a_217_1051.t6 14.282
R323 a_217_1051.n1 a_217_1051.t1 14.282
R324 a_217_1051.n1 a_217_1051.t4 14.282
R325 a_217_1051.t3 a_217_1051.n5 14.282
R326 a_217_1051.n5 a_217_1051.t2 14.282
R327 C.n2 C.t0 512.525
R328 C.n0 C.t2 512.525
R329 C.n2 C.t4 371.139
R330 C.n0 C.t5 371.139
R331 C.n3 C.n2 343.521
R332 C.n1 C.n0 343.521
R333 C.n1 C.t1 172.106
R334 C.n3 C.t3 165.68
R335 C.n4 C.n1 5.693
R336 C.n4 C.n3 4.65
R337 C.n4 C 0.046
R338 a_778_101.t0 a_778_101.n0 93.333
R339 a_778_101.n3 a_778_101.n1 79.053
R340 a_778_101.n3 a_778_101.n2 2.109
R341 a_778_101.t0 a_778_101.n3 0.195
R342 GND.n32 GND.n31 237.558
R343 GND.n65 GND.n64 237.558
R344 GND.n98 GND.n97 237.558
R345 GND.n29 GND.n28 210.82
R346 GND.n62 GND.n61 210.82
R347 GND.n100 GND.n99 210.82
R348 GND.n108 GND.n107 172.612
R349 GND.n78 GND.n77 151.605
R350 GND.n51 GND.n50 151.605
R351 GND.n20 GND.n19 37.582
R352 GND.t0 GND.n17 32.601
R353 GND.n77 GND.n76 28.421
R354 GND.n50 GND.n49 28.421
R355 GND.n77 GND.n75 25.263
R356 GND.n50 GND.n48 25.263
R357 GND.n75 GND.n74 24.383
R358 GND.n48 GND.n47 24.383
R359 GND.n17 GND.n16 21.734
R360 GND.n4 GND.n3 20.705
R361 GND.n10 GND.n9 20.705
R362 GND.n21 GND.n20 20.705
R363 GND.n3 GND.n2 19.952
R364 GND.n30 GND.n29 18.953
R365 GND.n63 GND.n62 18.953
R366 GND.n101 GND.n100 18.953
R367 GND.n19 GND.t0 15.644
R368 GND.n33 GND.n30 14.864
R369 GND.n66 GND.n63 14.864
R370 GND.n102 GND.n101 14.864
R371 GND.n19 GND.n18 13.541
R372 GND.n72 GND.n71 9.154
R373 GND.n80 GND.n79 9.154
R374 GND.n83 GND.n82 9.154
R375 GND.n86 GND.n85 9.154
R376 GND.n89 GND.n88 9.154
R377 GND.n92 GND.n91 9.154
R378 GND.n95 GND.n94 9.154
R379 GND.n102 GND.n98 9.154
R380 GND.n105 GND.n104 9.154
R381 GND.n110 GND.n109 9.154
R382 GND.n113 GND.n112 9.154
R383 GND.n116 GND.n115 9.154
R384 GND.n6 GND.n5 9.154
R385 GND.n12 GND.n11 9.154
R386 GND.n23 GND.n22 9.154
R387 GND.n26 GND.n25 9.154
R388 GND.n33 GND.n32 9.154
R389 GND.n36 GND.n35 9.154
R390 GND.n39 GND.n38 9.154
R391 GND.n42 GND.n41 9.154
R392 GND.n45 GND.n44 9.154
R393 GND.n53 GND.n52 9.154
R394 GND.n56 GND.n55 9.154
R395 GND.n59 GND.n58 9.154
R396 GND.n66 GND.n65 9.154
R397 GND.n122 GND.n121 9.154
R398 GND.n119 GND.n118 9.154
R399 GND.n7 GND.n1 4.795
R400 GND.n70 GND.n69 4.65
R401 GND.n117 GND.n116 4.65
R402 GND.n114 GND.n113 4.65
R403 GND.n111 GND.n110 4.65
R404 GND.n106 GND.n105 4.65
R405 GND.n103 GND.n102 4.65
R406 GND.n96 GND.n95 4.65
R407 GND.n93 GND.n92 4.65
R408 GND.n90 GND.n89 4.65
R409 GND.n87 GND.n86 4.65
R410 GND.n84 GND.n83 4.65
R411 GND.n81 GND.n80 4.65
R412 GND.n73 GND.n72 4.65
R413 GND.n7 GND.n6 4.65
R414 GND.n13 GND.n12 4.65
R415 GND.n24 GND.n23 4.65
R416 GND.n27 GND.n26 4.65
R417 GND.n34 GND.n33 4.65
R418 GND.n37 GND.n36 4.65
R419 GND.n40 GND.n39 4.65
R420 GND.n43 GND.n42 4.65
R421 GND.n46 GND.n45 4.65
R422 GND.n54 GND.n53 4.65
R423 GND.n57 GND.n56 4.65
R424 GND.n60 GND.n59 4.65
R425 GND.n67 GND.n66 4.65
R426 GND.n123 GND.n122 4.65
R427 GND.n120 GND.n119 4.65
R428 GND.n15 GND.n14 4.504
R429 GND.n6 GND.n4 4.129
R430 GND.n53 GND.n51 4.129
R431 GND.n110 GND.n108 4.129
R432 GND.n80 GND.n78 4.129
R433 GND.n23 GND.n21 3.716
R434 GND.t0 GND.n15 2.452
R435 GND.n1 GND.n0 0.475
R436 GND.n69 GND.n68 0.474
R437 GND.n9 GND.n8 0.376
R438 GND.n34 GND.n27 0.29
R439 GND.n67 GND.n60 0.29
R440 GND.n103 GND.n96 0.29
R441 GND.n70 GND 0.207
R442 GND.n12 GND.n10 0.206
R443 GND.n46 GND.n43 0.181
R444 GND.n117 GND.n114 0.181
R445 GND.n87 GND.n84 0.181
R446 GND.n13 GND.n7 0.157
R447 GND.n24 GND.n13 0.157
R448 GND.n27 GND.n24 0.145
R449 GND.n37 GND.n34 0.145
R450 GND.n40 GND.n37 0.145
R451 GND.n43 GND.n40 0.145
R452 GND.n54 GND.n46 0.145
R453 GND.n57 GND.n54 0.145
R454 GND.n60 GND.n57 0.145
R455 GND.n123 GND.n120 0.145
R456 GND.n120 GND.n117 0.145
R457 GND.n114 GND.n111 0.145
R458 GND.n111 GND.n106 0.145
R459 GND.n106 GND.n103 0.145
R460 GND.n96 GND.n93 0.145
R461 GND.n93 GND.n90 0.145
R462 GND.n90 GND.n87 0.145
R463 GND.n84 GND.n81 0.145
R464 GND.n81 GND.n73 0.145
R465 GND.n73 GND.n70 0.145
R466 GND GND.n67 0.078
R467 GND GND.n123 0.066
R468 a_112_101.n3 a_112_101.n2 62.817
R469 a_112_101.n11 a_112_101.n10 46.054
R470 a_112_101.n7 a_112_101.n6 38.626
R471 a_112_101.n6 a_112_101.n5 35.955
R472 a_112_101.n12 a_112_101.n11 27.923
R473 a_112_101.n3 a_112_101.n1 26.202
R474 a_112_101.t0 a_112_101.n3 19.737
R475 a_112_101.t0 a_112_101.n4 7.273
R476 a_112_101.n9 a_112_101.n8 6.883
R477 a_112_101.t0 a_112_101.n0 6.109
R478 a_112_101.t1 a_112_101.n7 4.864
R479 a_112_101.t0 a_112_101.n13 2.074
R480 a_112_101.t1 a_112_101.n9 1.179
R481 a_112_101.t1 a_112_101.n12 0.958
R482 a_112_101.n13 a_112_101.t1 0.937
R483 a_1444_101.n3 a_1444_101.n1 42.788
R484 a_1444_101.t0 a_1444_101.n0 8.137
R485 a_1444_101.n3 a_1444_101.n2 4.665
R486 a_1444_101.t0 a_1444_101.n3 0.06
C7 VDD GND 4.85fF
C8 a_1444_101.n0 GND 0.06fF
C9 a_1444_101.n1 GND 0.13fF
C10 a_1444_101.n2 GND 0.04fF
C11 a_1444_101.n3 GND 0.19fF
C12 a_112_101.n0 GND 0.02fF
C13 a_112_101.n1 GND 0.08fF
C14 a_112_101.n2 GND 0.07fF
C15 a_112_101.n3 GND 0.03fF
C16 a_112_101.n4 GND 0.01fF
C17 a_112_101.n5 GND 0.03fF
C18 a_112_101.n6 GND 0.04fF
C19 a_112_101.n7 GND 0.02fF
C20 a_112_101.n8 GND 0.04fF
C21 a_112_101.n9 GND 0.07fF
C22 a_112_101.n10 GND 0.04fF
C23 a_112_101.n11 GND 0.11fF
C24 a_112_101.n12 GND 0.14fF
C25 a_112_101.t1 GND 0.15fF
C26 a_112_101.n13 GND 0.01fF
C27 a_778_101.n0 GND 0.02fF
C28 a_778_101.n1 GND 0.13fF
C29 a_778_101.n2 GND 0.13fF
C30 a_778_101.n3 GND 0.15fF
C31 a_217_1051.n0 GND 0.36fF
C32 a_217_1051.n1 GND 0.32fF
C33 a_217_1051.n2 GND 0.52fF
C34 a_217_1051.n3 GND 0.30fF
C35 a_217_1051.n4 GND 0.79fF
C36 a_217_1051.n5 GND 0.42fF
C37 a_881_1051.n0 GND 0.29fF
C38 a_881_1051.n1 GND 0.28fF
C39 a_881_1051.n2 GND 0.37fF
C40 a_881_1051.n3 GND 0.70fF
C41 a_881_1051.n4 GND 0.27fF
C42 a_881_1051.n5 GND 0.45fF
C43 Y.n0 GND 0.58fF
C44 Y.n1 GND 0.04fF
C45 Y.n2 GND 0.05fF
C46 Y.n3 GND 0.03fF
C47 Y.n4 GND 0.25fF
C48 Y.n5 GND 0.64fF
C49 Y.n6 GND 0.01fF
C50 VDD.n1 GND 0.03fF
C51 VDD.n2 GND 0.10fF
C52 VDD.n3 GND 0.03fF
C53 VDD.n4 GND 0.02fF
C54 VDD.n5 GND 0.06fF
C55 VDD.n6 GND 0.02fF
C56 VDD.n7 GND 0.02fF
C57 VDD.n8 GND 0.02fF
C58 VDD.n9 GND 0.02fF
C59 VDD.n10 GND 0.02fF
C60 VDD.n11 GND 0.02fF
C61 VDD.n12 GND 0.02fF
C62 VDD.n13 GND 0.02fF
C63 VDD.n14 GND 0.04fF
C64 VDD.n15 GND 0.01fF
C65 VDD.n20 GND 0.47fF
C66 VDD.n21 GND 0.28fF
C67 VDD.n22 GND 0.02fF
C68 VDD.n23 GND 0.03fF
C69 VDD.n24 GND 0.06fF
C70 VDD.n25 GND 0.21fF
C71 VDD.n26 GND 0.01fF
C72 VDD.n27 GND 0.01fF
C73 VDD.n28 GND 0.07fF
C74 VDD.n29 GND 0.17fF
C75 VDD.n30 GND 0.01fF
C76 VDD.n31 GND 0.03fF
C77 VDD.n32 GND 0.03fF
C78 VDD.n33 GND 0.21fF
C79 VDD.n34 GND 0.01fF
C80 VDD.n35 GND 0.06fF
C81 VDD.n36 GND 0.01fF
C82 VDD.n37 GND 0.02fF
C83 VDD.n38 GND 0.28fF
C84 VDD.n39 GND 0.01fF
C85 VDD.n40 GND 0.02fF
C86 VDD.n41 GND 0.04fF
C87 VDD.n42 GND 0.06fF
C88 VDD.n43 GND 0.02fF
C89 VDD.n44 GND 0.02fF
C90 VDD.n45 GND 0.02fF
C91 VDD.n46 GND 0.02fF
C92 VDD.n47 GND 0.02fF
C93 VDD.n48 GND 0.02fF
C94 VDD.n49 GND 0.02fF
C95 VDD.n50 GND 0.02fF
C96 VDD.n51 GND 0.02fF
C97 VDD.n52 GND 0.02fF
C98 VDD.n53 GND 0.02fF
C99 VDD.n54 GND 0.03fF
C100 VDD.n55 GND 0.02fF
C101 VDD.n56 GND 0.19fF
C102 VDD.n57 GND 0.02fF
C103 VDD.n58 GND 0.02fF
C104 VDD.n60 GND 0.02fF
C105 VDD.n64 GND 0.28fF
C106 VDD.n65 GND 0.28fF
C107 VDD.n66 GND 0.01fF
C108 VDD.n67 GND 0.02fF
C109 VDD.n68 GND 0.04fF
C110 VDD.n69 GND 0.25fF
C111 VDD.n70 GND 0.01fF
C112 VDD.n71 GND 0.02fF
C113 VDD.n72 GND 0.02fF
C114 VDD.n73 GND 0.17fF
C115 VDD.n74 GND 0.01fF
C116 VDD.n75 GND 0.02fF
C117 VDD.n76 GND 0.02fF
C118 VDD.n77 GND 0.01fF
C119 VDD.n78 GND 0.03fF
C120 VDD.n79 GND 0.03fF
C121 VDD.n80 GND 0.14fF
C122 VDD.n81 GND 0.01fF
C123 VDD.n82 GND 0.03fF
C124 VDD.n83 GND 0.03fF
C125 VDD.n84 GND 0.17fF
C126 VDD.n85 GND 0.01fF
C127 VDD.n86 GND 0.02fF
C128 VDD.n87 GND 0.02fF
C129 VDD.n88 GND 0.25fF
C130 VDD.n89 GND 0.01fF
C131 VDD.n90 GND 0.02fF
C132 VDD.n91 GND 0.02fF
C133 VDD.n92 GND 0.28fF
C134 VDD.n93 GND 0.01fF
C135 VDD.n94 GND 0.02fF
C136 VDD.n95 GND 0.04fF
C137 VDD.n96 GND 0.22fF
C138 VDD.n97 GND 0.02fF
C139 VDD.n98 GND 0.02fF
C140 VDD.n99 GND 0.02fF
C141 VDD.n100 GND 0.06fF
C142 VDD.n101 GND 0.02fF
C143 VDD.n102 GND 0.02fF
C144 VDD.n103 GND 0.02fF
C145 VDD.n104 GND 0.02fF
C146 VDD.n105 GND 0.02fF
C147 VDD.n106 GND 0.02fF
C148 VDD.n107 GND 0.02fF
C149 VDD.n108 GND 0.02fF
C150 VDD.n109 GND 0.02fF
C151 VDD.n110 GND 0.02fF
C152 VDD.n111 GND 0.03fF
C153 VDD.n112 GND 0.02fF
C154 VDD.n113 GND 0.02fF
C155 VDD.n117 GND 0.28fF
C156 VDD.n118 GND 0.28fF
C157 VDD.n119 GND 0.01fF
C158 VDD.n120 GND 0.02fF
C159 VDD.n121 GND 0.03fF
C160 VDD.n122 GND 0.14fF
C161 VDD.n123 GND 0.02fF
C162 VDD.n124 GND 0.02fF
C163 VDD.n125 GND 0.06fF
C164 VDD.n126 GND 0.02fF
C165 VDD.n127 GND 0.02fF
C166 VDD.n128 GND 0.02fF
C167 VDD.n129 GND 0.02fF
C168 VDD.n130 GND 0.02fF
C169 VDD.n131 GND 0.02fF
C170 VDD.n132 GND 0.02fF
C171 VDD.n133 GND 0.02fF
C172 VDD.n134 GND 0.03fF
C173 VDD.n135 GND 0.04fF
C174 VDD.n136 GND 0.02fF
C175 VDD.n140 GND 0.47fF
C176 VDD.n141 GND 0.28fF
C177 VDD.n142 GND 0.02fF
C178 VDD.n143 GND 0.03fF
C179 VDD.n144 GND 0.03fF
C180 VDD.n145 GND 0.07fF
C181 VDD.n146 GND 0.25fF
C182 VDD.n147 GND 0.01fF
C183 VDD.n148 GND 0.01fF
C184 VDD.n149 GND 0.02fF
C185 VDD.n150 GND 0.17fF
C186 VDD.n151 GND 0.01fF
C187 VDD.n152 GND 0.02fF
C188 VDD.n153 GND