** sch_path: /home/rjridle/OpenRadHardSCL/lib/xschem/schematics/NAND2X2.sch
.subckt NAND2X2 A B YN
*.PININFO A:I B:I YN:O
M1 YN A VDD VDD pmos w=2u l=0.15u m=1
M2 YN B VDD VDD pmos w=2u l=0.15u m=1
M4 YN A net1 GND nmos w=3u l=0.15u m=1
M5 net1 B GND GND nmos w=3u l=0.15u m=1
M3 YN A VDD VDD pmos w=2u l=0.15u m=1
M6 YN B VDD VDD pmos w=2u l=0.15u m=1
.ends
.GLOBAL GND
.GLOBAL VDD
.end
