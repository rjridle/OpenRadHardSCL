# Standard Cell LEF generated in Magic




MACRO AND2X1
  CLASS BLOCK ;
  FOREIGN AND2X1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 6.390 BY 7.950 ;
  PIN Y
    ANTENNADIFFAREA 0.771900 ;
    PORT
      LAYER li1 ;
        RECT 4.355 4.895 4.525 7.250 ;
        RECT 4.355 4.725 4.895 4.895 ;
        RECT 4.725 2.305 4.895 4.725 ;
        RECT 4.355 2.135 4.895 2.305 ;
        RECT 4.355 0.975 4.525 2.135 ;
      LAYER mcon ;
        RECT 4.725 3.245 4.895 3.415 ;
      LAYER met1 ;
        RECT 4.695 3.415 4.925 3.445 ;
        RECT 4.665 3.245 5.075 3.415 ;
        RECT 4.695 3.215 4.925 3.245 ;
    END
  END Y
  PIN A
    ANTENNAGATEAREA 1.033250 ;
    PORT
      LAYER li1 ;
        RECT 1.025 2.055 1.195 5.095 ;
      LAYER mcon ;
        RECT 1.025 3.985 1.195 4.155 ;
      LAYER met1 ;
        RECT 0.995 4.155 1.225 4.185 ;
        RECT 0.845 3.985 1.255 4.155 ;
        RECT 0.995 3.955 1.225 3.985 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 1.027250 ;
    PORT
      LAYER li1 ;
        RECT 1.795 4.940 1.965 5.095 ;
        RECT 1.765 4.765 1.965 4.940 ;
        RECT 1.765 2.055 1.935 4.765 ;
      LAYER mcon ;
        RECT 1.765 3.615 1.935 3.785 ;
      LAYER met1 ;
        RECT 1.735 3.785 1.965 3.815 ;
        RECT 1.585 3.615 1.995 3.785 ;
        RECT 1.735 3.585 1.965 3.615 ;
    END
  END B
  PIN VDD
    ANTENNADIFFAREA 8.266550 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 5.970 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 5.705 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 0.705 5.365 0.875 7.460 ;
        RECT 1.585 5.785 1.755 7.460 ;
        RECT 2.465 5.785 2.635 7.460 ;
        RECT 3.175 4.340 3.485 7.460 ;
        RECT 3.915 5.415 4.085 7.460 ;
        RECT 4.795 5.415 4.965 7.460 ;
        RECT 5.395 4.340 5.705 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 0.995 7.525 1.165 7.695 ;
        RECT 1.355 7.525 1.525 7.695 ;
        RECT 1.805 7.525 1.975 7.695 ;
        RECT 2.165 7.525 2.335 7.695 ;
        RECT 2.525 7.525 2.695 7.695 ;
        RECT 2.885 7.525 3.055 7.695 ;
        RECT 3.605 7.525 3.775 7.695 ;
        RECT 3.965 7.525 4.135 7.695 ;
        RECT 4.355 7.525 4.525 7.695 ;
        RECT 4.745 7.525 4.915 7.695 ;
        RECT 5.105 7.525 5.275 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 5.705 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 6.344700 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 5.835 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 3.045 -0.075 3.615 -0.065 ;
        RECT 5.265 -0.075 5.835 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 1.095 0.310 1.265 1.260 ;
        RECT 3.175 0.310 3.485 2.860 ;
        RECT 3.875 0.755 4.045 1.885 ;
        RECT 4.845 0.755 5.015 1.885 ;
        RECT 3.875 0.585 5.015 0.755 ;
        RECT 3.875 0.310 4.045 0.585 ;
        RECT 4.360 0.310 4.530 0.585 ;
        RECT 4.845 0.310 5.015 0.585 ;
        RECT 5.395 0.310 5.705 2.860 ;
        RECT -0.155 0.000 5.705 0.310 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 0.995 0.065 1.165 0.235 ;
        RECT 1.355 0.065 1.525 0.235 ;
        RECT 1.805 0.065 1.975 0.235 ;
        RECT 2.165 0.065 2.335 0.235 ;
        RECT 2.525 0.065 2.695 0.235 ;
        RECT 2.885 0.065 3.055 0.235 ;
        RECT 3.605 0.065 3.775 0.235 ;
        RECT 3.965 0.065 4.135 0.235 ;
        RECT 4.355 0.065 4.525 0.235 ;
        RECT 4.745 0.065 4.915 0.235 ;
        RECT 5.105 0.065 5.275 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 5.705 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 1.145 5.515 1.315 7.250 ;
        RECT 2.025 5.515 2.195 7.250 ;
        RECT 1.145 5.345 2.675 5.515 ;
        RECT 0.610 1.805 0.780 1.885 ;
        RECT 1.580 1.805 1.750 1.885 ;
        RECT 2.505 1.880 2.675 5.345 ;
        RECT 3.985 2.055 4.155 5.095 ;
        RECT 0.610 1.635 1.750 1.805 ;
        RECT 0.610 0.505 0.780 1.635 ;
        RECT 1.580 0.755 1.750 1.635 ;
        RECT 2.065 1.710 2.675 1.880 ;
        RECT 2.065 0.975 2.235 1.710 ;
        RECT 2.550 0.755 2.720 1.525 ;
        RECT 1.580 0.585 2.720 0.755 ;
        RECT 1.580 0.505 1.750 0.585 ;
        RECT 2.550 0.505 2.720 0.585 ;
      LAYER mcon ;
        RECT 2.505 3.245 2.675 3.415 ;
        RECT 3.985 3.245 4.155 3.415 ;
      LAYER met1 ;
        RECT 2.475 3.415 2.705 3.445 ;
        RECT 3.955 3.415 4.185 3.445 ;
        RECT 2.445 3.245 4.215 3.415 ;
        RECT 2.475 3.215 2.705 3.245 ;
        RECT 3.955 3.215 4.185 3.245 ;
  END
END AND2X1






MACRO AND3X1
  CLASS BLOCK ;
  FOREIGN AND3X1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 7.870 BY 7.950 ;
  PIN Y
    ANTENNADIFFAREA 0.771900 ;
    PORT
      LAYER li1 ;
        RECT 5.835 4.895 6.005 7.250 ;
        RECT 5.835 4.725 6.375 4.895 ;
        RECT 6.205 2.305 6.375 4.725 ;
        RECT 5.835 2.135 6.375 2.305 ;
        RECT 5.835 0.975 6.005 2.135 ;
      LAYER mcon ;
        RECT 6.205 3.245 6.375 3.415 ;
      LAYER met1 ;
        RECT 6.175 3.415 6.405 3.445 ;
        RECT 6.145 3.245 6.555 3.415 ;
        RECT 6.175 3.215 6.405 3.245 ;
    END
  END Y
  PIN A
    ANTENNAGATEAREA 1.033250 ;
    PORT
      LAYER li1 ;
        RECT 1.025 2.055 1.195 5.095 ;
      LAYER mcon ;
        RECT 1.025 3.985 1.195 4.155 ;
      LAYER met1 ;
        RECT 0.995 4.155 1.225 4.185 ;
        RECT 0.845 3.985 1.255 4.155 ;
        RECT 0.995 3.955 1.225 3.985 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 1.014850 ;
    PORT
      LAYER li1 ;
        RECT 2.135 2.055 2.305 5.095 ;
      LAYER mcon ;
        RECT 2.135 3.615 2.305 3.785 ;
      LAYER met1 ;
        RECT 2.105 3.785 2.335 3.815 ;
        RECT 1.955 3.615 2.365 3.785 ;
        RECT 2.105 3.585 2.335 3.615 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA 1.027250 ;
    PORT
      LAYER li1 ;
        RECT 3.245 2.055 3.415 5.095 ;
      LAYER mcon ;
        RECT 3.245 3.245 3.415 3.415 ;
      LAYER met1 ;
        RECT 3.215 3.415 3.445 3.445 ;
        RECT 3.065 3.245 3.475 3.415 ;
        RECT 3.215 3.215 3.445 3.245 ;
    END
  END C
  PIN VDD
    ANTENNADIFFAREA 9.556950 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 7.450 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 7.185 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 1.005 5.445 1.175 7.460 ;
        RECT 1.885 5.785 2.055 7.460 ;
        RECT 2.765 5.785 2.935 7.460 ;
        RECT 3.645 5.785 3.815 7.460 ;
        RECT 4.655 4.340 4.965 7.460 ;
        RECT 5.395 5.415 5.565 7.460 ;
        RECT 6.275 5.415 6.445 7.460 ;
        RECT 6.875 4.340 7.185 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 0.995 7.525 1.165 7.695 ;
        RECT 1.355 7.525 1.525 7.695 ;
        RECT 1.715 7.525 1.885 7.695 ;
        RECT 2.075 7.525 2.245 7.695 ;
        RECT 2.565 7.525 2.735 7.695 ;
        RECT 2.925 7.525 3.095 7.695 ;
        RECT 3.285 7.525 3.455 7.695 ;
        RECT 3.645 7.525 3.815 7.695 ;
        RECT 4.005 7.525 4.175 7.695 ;
        RECT 4.365 7.525 4.535 7.695 ;
        RECT 5.085 7.525 5.255 7.695 ;
        RECT 5.445 7.525 5.615 7.695 ;
        RECT 5.835 7.525 6.005 7.695 ;
        RECT 6.225 7.525 6.395 7.695 ;
        RECT 6.585 7.525 6.755 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 7.185 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 7.055100 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 7.315 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 4.525 -0.075 5.095 -0.065 ;
        RECT 6.745 -0.075 7.315 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 0.990 0.310 1.160 1.270 ;
        RECT 4.655 0.310 4.965 2.860 ;
        RECT 5.355 0.755 5.525 1.885 ;
        RECT 6.325 0.755 6.495 1.885 ;
        RECT 5.355 0.585 6.495 0.755 ;
        RECT 5.355 0.310 5.525 0.585 ;
        RECT 5.840 0.310 6.010 0.585 ;
        RECT 6.325 0.310 6.495 0.585 ;
        RECT 6.875 0.310 7.185 2.860 ;
        RECT -0.155 0.000 7.185 0.310 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 0.995 0.065 1.165 0.235 ;
        RECT 1.355 0.065 1.525 0.235 ;
        RECT 1.715 0.065 1.885 0.235 ;
        RECT 2.075 0.065 2.245 0.235 ;
        RECT 2.565 0.065 2.735 0.235 ;
        RECT 2.925 0.065 3.095 0.235 ;
        RECT 3.285 0.065 3.455 0.235 ;
        RECT 3.645 0.065 3.815 0.235 ;
        RECT 4.005 0.065 4.175 0.235 ;
        RECT 4.365 0.065 4.535 0.235 ;
        RECT 5.085 0.065 5.255 0.235 ;
        RECT 5.445 0.065 5.615 0.235 ;
        RECT 5.835 0.065 6.005 0.235 ;
        RECT 6.225 0.065 6.395 0.235 ;
        RECT 6.585 0.065 6.755 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 7.185 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 1.445 5.470 1.615 7.250 ;
        RECT 2.325 5.470 2.495 7.250 ;
        RECT 3.205 5.470 3.375 7.250 ;
        RECT 1.445 5.300 4.155 5.470 ;
        RECT 0.505 1.815 0.675 1.895 ;
        RECT 1.475 1.815 1.645 1.895 ;
        RECT 2.445 1.815 2.615 1.895 ;
        RECT 0.505 1.645 2.615 1.815 ;
        RECT 0.505 0.515 0.675 1.645 ;
        RECT 1.475 0.765 1.645 1.645 ;
        RECT 2.445 1.565 2.615 1.645 ;
        RECT 1.965 1.220 2.135 1.300 ;
        RECT 3.015 1.220 3.185 1.895 ;
        RECT 3.985 1.890 4.155 5.300 ;
        RECT 5.465 2.055 5.635 5.095 ;
        RECT 1.965 1.050 3.185 1.220 ;
        RECT 1.965 0.970 2.135 1.050 ;
        RECT 2.445 0.765 2.615 0.845 ;
        RECT 1.475 0.595 2.615 0.765 ;
        RECT 1.475 0.515 1.645 0.595 ;
        RECT 2.445 0.515 2.615 0.595 ;
        RECT 3.015 0.765 3.185 1.050 ;
        RECT 3.500 1.720 4.155 1.890 ;
        RECT 3.500 0.985 3.670 1.720 ;
        RECT 3.985 0.765 4.155 1.535 ;
        RECT 3.015 0.595 4.155 0.765 ;
        RECT 3.015 0.515 3.185 0.595 ;
        RECT 3.985 0.515 4.155 0.595 ;
      LAYER mcon ;
        RECT 3.985 3.245 4.155 3.415 ;
        RECT 5.465 3.245 5.635 3.415 ;
      LAYER met1 ;
        RECT 3.955 3.415 4.185 3.445 ;
        RECT 5.435 3.415 5.665 3.445 ;
        RECT 3.925 3.245 5.695 3.415 ;
        RECT 3.955 3.215 4.185 3.245 ;
        RECT 5.435 3.215 5.665 3.245 ;
  END
END AND3X1






MACRO AO3X1
  CLASS BLOCK ;
  FOREIGN AO3X1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 9.720 BY 7.950 ;
  PIN A
    ANTENNAGATEAREA 1.033250 ;
    PORT
      LAYER li1 ;
        RECT 1.025 2.055 1.195 5.095 ;
      LAYER mcon ;
        RECT 1.025 2.875 1.195 3.045 ;
      LAYER met1 ;
        RECT 0.995 3.045 1.225 3.075 ;
        RECT 0.845 2.875 1.255 3.045 ;
        RECT 0.995 2.845 1.225 2.875 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 1.027250 ;
    PORT
      LAYER li1 ;
        RECT 1.795 4.940 1.965 5.095 ;
        RECT 1.765 4.765 1.965 4.940 ;
        RECT 1.765 2.055 1.935 4.765 ;
      LAYER mcon ;
        RECT 1.765 3.245 1.935 3.415 ;
      LAYER met1 ;
        RECT 1.735 3.415 1.965 3.445 ;
        RECT 1.585 3.245 1.995 3.415 ;
        RECT 1.735 3.215 1.965 3.245 ;
    END
  END B
  PIN VDD
    ANTENNADIFFAREA 11.336200 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 9.300 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 9.035 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 0.705 5.365 0.875 7.460 ;
        RECT 1.585 5.785 1.755 7.460 ;
        RECT 2.465 5.785 2.635 7.460 ;
        RECT 3.175 4.340 3.485 7.460 ;
        RECT 4.475 5.785 4.645 7.460 ;
        RECT 6.505 4.340 6.815 7.460 ;
        RECT 7.245 5.415 7.415 7.460 ;
        RECT 8.125 5.415 8.295 7.460 ;
        RECT 8.725 4.340 9.035 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 0.995 7.525 1.165 7.695 ;
        RECT 1.355 7.525 1.525 7.695 ;
        RECT 1.805 7.525 1.975 7.695 ;
        RECT 2.165 7.525 2.335 7.695 ;
        RECT 2.525 7.525 2.695 7.695 ;
        RECT 2.885 7.525 3.055 7.695 ;
        RECT 3.605 7.525 3.775 7.695 ;
        RECT 3.965 7.525 4.135 7.695 ;
        RECT 4.325 7.525 4.495 7.695 ;
        RECT 4.685 7.525 4.855 7.695 ;
        RECT 5.135 7.525 5.305 7.695 ;
        RECT 5.495 7.525 5.665 7.695 ;
        RECT 5.855 7.525 6.025 7.695 ;
        RECT 6.215 7.525 6.385 7.695 ;
        RECT 6.935 7.525 7.105 7.695 ;
        RECT 7.295 7.525 7.465 7.695 ;
        RECT 7.685 7.525 7.855 7.695 ;
        RECT 8.075 7.525 8.245 7.695 ;
        RECT 8.435 7.525 8.605 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 9.035 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 10.674350 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 9.165 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 3.045 -0.075 3.615 -0.065 ;
        RECT 6.375 -0.075 6.945 -0.065 ;
        RECT 8.595 -0.075 9.165 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 1.095 0.310 1.265 1.260 ;
        RECT 3.175 0.310 3.485 2.860 ;
        RECT 3.940 0.755 4.110 1.885 ;
        RECT 4.910 0.755 5.080 1.530 ;
        RECT 5.880 0.755 6.050 1.530 ;
        RECT 3.940 0.585 6.050 0.755 ;
        RECT 3.940 0.310 4.110 0.585 ;
        RECT 4.425 0.310 4.595 0.585 ;
        RECT 4.910 0.310 5.080 0.585 ;
        RECT 5.395 0.310 5.565 0.585 ;
        RECT 5.880 0.310 6.050 0.585 ;
        RECT 6.505 0.310 6.815 2.860 ;
        RECT 7.205 0.755 7.375 1.885 ;
        RECT 8.175 0.755 8.345 1.885 ;
        RECT 7.205 0.585 8.345 0.755 ;
        RECT 7.205 0.310 7.375 0.585 ;
        RECT 7.690 0.310 7.860 0.585 ;
        RECT 8.175 0.310 8.345 0.585 ;
        RECT 8.725 0.310 9.035 2.860 ;
        RECT -0.155 0.000 9.035 0.310 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 0.995 0.065 1.165 0.235 ;
        RECT 1.355 0.065 1.525 0.235 ;
        RECT 1.805 0.065 1.975 0.235 ;
        RECT 2.165 0.065 2.335 0.235 ;
        RECT 2.525 0.065 2.695 0.235 ;
        RECT 2.885 0.065 3.055 0.235 ;
        RECT 3.605 0.065 3.775 0.235 ;
        RECT 3.965 0.065 4.135 0.235 ;
        RECT 4.325 0.065 4.495 0.235 ;
        RECT 4.685 0.065 4.855 0.235 ;
        RECT 5.135 0.065 5.305 0.235 ;
        RECT 5.495 0.065 5.665 0.235 ;
        RECT 5.855 0.065 6.025 0.235 ;
        RECT 6.215 0.065 6.385 0.235 ;
        RECT 6.935 0.065 7.105 0.235 ;
        RECT 7.295 0.065 7.465 0.235 ;
        RECT 7.685 0.065 7.855 0.235 ;
        RECT 8.075 0.065 8.245 0.235 ;
        RECT 8.435 0.065 8.605 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 9.035 0.310 ;
    END
  END VSS
  PIN C
    ANTENNAGATEAREA 1.026450 ;
    PORT
      LAYER li1 ;
        RECT 5.130 4.940 5.300 5.100 ;
        RECT 5.095 4.770 5.300 4.940 ;
        RECT 5.095 2.055 5.265 4.770 ;
      LAYER mcon ;
        RECT 5.095 3.615 5.265 3.785 ;
      LAYER met1 ;
        RECT 5.065 3.785 5.295 3.815 ;
        RECT 4.915 3.615 5.325 3.785 ;
        RECT 5.065 3.585 5.295 3.615 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA 0.771900 ;
    PORT
      LAYER li1 ;
        RECT 7.685 4.895 7.855 7.250 ;
        RECT 7.685 4.725 8.225 4.895 ;
        RECT 8.055 2.305 8.225 4.725 ;
        RECT 7.685 2.135 8.225 2.305 ;
        RECT 7.685 0.975 7.855 2.135 ;
      LAYER mcon ;
        RECT 8.055 3.985 8.225 4.155 ;
      LAYER met1 ;
        RECT 8.025 4.155 8.255 4.185 ;
        RECT 7.995 3.985 8.405 4.155 ;
        RECT 8.025 3.955 8.255 3.985 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 1.145 5.515 1.315 7.250 ;
        RECT 2.025 5.515 2.195 7.250 ;
        RECT 4.035 5.525 4.205 7.255 ;
        RECT 4.915 7.055 5.965 7.225 ;
        RECT 4.915 5.525 5.085 7.055 ;
        RECT 1.145 5.345 2.675 5.515 ;
        RECT 4.035 5.355 5.085 5.525 ;
        RECT 5.355 5.525 5.525 6.795 ;
        RECT 5.795 5.785 5.965 7.055 ;
        RECT 5.355 5.355 6.005 5.525 ;
        RECT 0.610 1.805 0.780 1.885 ;
        RECT 1.580 1.805 1.750 1.885 ;
        RECT 2.505 1.880 2.675 5.345 ;
        RECT 4.200 4.940 4.370 5.100 ;
        RECT 4.200 4.770 4.525 4.940 ;
        RECT 4.355 2.055 4.525 4.770 ;
        RECT 5.835 1.880 6.005 5.355 ;
        RECT 7.315 2.055 7.485 5.095 ;
        RECT 0.610 1.635 1.750 1.805 ;
        RECT 0.610 0.505 0.780 1.635 ;
        RECT 1.580 0.755 1.750 1.635 ;
        RECT 2.065 1.710 2.675 1.880 ;
        RECT 4.425 1.710 6.005 1.880 ;
        RECT 2.065 0.975 2.235 1.710 ;
        RECT 2.550 0.755 2.720 1.525 ;
        RECT 4.425 0.975 4.595 1.710 ;
        RECT 5.395 0.975 5.565 1.710 ;
        RECT 1.580 0.585 2.720 0.755 ;
        RECT 1.580 0.505 1.750 0.585 ;
        RECT 2.550 0.505 2.720 0.585 ;
      LAYER mcon ;
        RECT 2.505 2.505 2.675 2.675 ;
        RECT 4.355 2.505 4.525 2.675 ;
        RECT 5.835 2.505 6.005 2.675 ;
        RECT 7.315 2.505 7.485 2.675 ;
      LAYER met1 ;
        RECT 2.475 2.675 2.705 2.705 ;
        RECT 4.325 2.675 4.555 2.705 ;
        RECT 5.805 2.675 6.035 2.705 ;
        RECT 7.285 2.675 7.515 2.705 ;
        RECT 2.445 2.505 4.585 2.675 ;
        RECT 5.775 2.505 7.545 2.675 ;
        RECT 2.475 2.475 2.705 2.505 ;
        RECT 4.325 2.475 4.555 2.505 ;
        RECT 5.805 2.475 6.035 2.505 ;
        RECT 7.285 2.475 7.515 2.505 ;
  END
END AO3X1






MACRO AOA4X1
  CLASS BLOCK ;
  FOREIGN AOA4X1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 13.050 BY 7.950 ;
  PIN Y
    ANTENNADIFFAREA 0.771900 ;
    PORT
      LAYER li1 ;
        RECT 11.015 4.895 11.185 7.250 ;
        RECT 11.015 4.725 11.555 4.895 ;
        RECT 11.385 2.305 11.555 4.725 ;
        RECT 11.015 2.135 11.555 2.305 ;
        RECT 11.015 0.975 11.185 2.135 ;
      LAYER mcon ;
        RECT 11.385 2.875 11.555 3.045 ;
      LAYER met1 ;
        RECT 11.355 3.045 11.585 3.075 ;
        RECT 11.325 2.875 11.735 3.045 ;
        RECT 11.355 2.845 11.585 2.875 ;
    END
  END Y
  PIN A
    ANTENNAGATEAREA 1.033250 ;
    PORT
      LAYER li1 ;
        RECT 1.025 2.055 1.195 5.095 ;
      LAYER mcon ;
        RECT 1.025 2.875 1.195 3.045 ;
      LAYER met1 ;
        RECT 0.995 3.045 1.225 3.075 ;
        RECT 0.845 2.875 1.255 3.045 ;
        RECT 0.995 2.845 1.225 2.875 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 1.027250 ;
    PORT
      LAYER li1 ;
        RECT 1.795 4.940 1.965 5.095 ;
        RECT 1.765 4.765 1.965 4.940 ;
        RECT 1.765 2.055 1.935 4.765 ;
      LAYER mcon ;
        RECT 1.765 3.245 1.935 3.415 ;
      LAYER met1 ;
        RECT 1.735 3.415 1.965 3.445 ;
        RECT 1.585 3.245 1.995 3.415 ;
        RECT 1.735 3.215 1.965 3.245 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA 1.026450 ;
    PORT
      LAYER li1 ;
        RECT 5.130 4.940 5.300 5.100 ;
        RECT 5.095 4.770 5.300 4.940 ;
        RECT 5.095 2.055 5.265 4.770 ;
      LAYER mcon ;
        RECT 5.095 3.615 5.265 3.785 ;
      LAYER met1 ;
        RECT 5.065 3.785 5.295 3.815 ;
        RECT 4.915 3.615 5.325 3.785 ;
        RECT 5.065 3.585 5.295 3.615 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA 1.027250 ;
    PORT
      LAYER li1 ;
        RECT 8.455 4.940 8.625 5.095 ;
        RECT 8.425 4.765 8.625 4.940 ;
        RECT 8.425 2.055 8.595 4.765 ;
      LAYER mcon ;
        RECT 8.425 3.985 8.595 4.155 ;
      LAYER met1 ;
        RECT 8.395 4.155 8.625 4.185 ;
        RECT 8.245 3.985 8.655 4.155 ;
        RECT 8.395 3.955 8.625 3.985 ;
    END
  END D
  PIN VDD
    ANTENNADIFFAREA 15.505850 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 12.630 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 12.365 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 0.705 5.365 0.875 7.460 ;
        RECT 1.585 5.785 1.755 7.460 ;
        RECT 2.465 5.785 2.635 7.460 ;
        RECT 3.175 4.340 3.485 7.460 ;
        RECT 4.475 5.785 4.645 7.460 ;
        RECT 6.505 4.340 6.815 7.460 ;
        RECT 7.365 5.365 7.535 7.460 ;
        RECT 8.245 5.785 8.415 7.460 ;
        RECT 9.125 5.785 9.295 7.460 ;
        RECT 9.835 4.340 10.145 7.460 ;
        RECT 10.575 5.415 10.745 7.460 ;
        RECT 11.455 5.415 11.625 7.460 ;
        RECT 12.055 4.340 12.365 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 0.995 7.525 1.165 7.695 ;
        RECT 1.355 7.525 1.525 7.695 ;
        RECT 1.805 7.525 1.975 7.695 ;
        RECT 2.165 7.525 2.335 7.695 ;
        RECT 2.525 7.525 2.695 7.695 ;
        RECT 2.885 7.525 3.055 7.695 ;
        RECT 3.605 7.525 3.775 7.695 ;
        RECT 3.965 7.525 4.135 7.695 ;
        RECT 4.325 7.525 4.495 7.695 ;
        RECT 4.685 7.525 4.855 7.695 ;
        RECT 5.135 7.525 5.305 7.695 ;
        RECT 5.495 7.525 5.665 7.695 ;
        RECT 5.855 7.525 6.025 7.695 ;
        RECT 6.215 7.525 6.385 7.695 ;
        RECT 6.935 7.525 7.105 7.695 ;
        RECT 7.295 7.525 7.465 7.695 ;
        RECT 7.655 7.525 7.825 7.695 ;
        RECT 8.015 7.525 8.185 7.695 ;
        RECT 8.465 7.525 8.635 7.695 ;
        RECT 8.825 7.525 8.995 7.695 ;
        RECT 9.185 7.525 9.355 7.695 ;
        RECT 9.545 7.525 9.715 7.695 ;
        RECT 10.265 7.525 10.435 7.695 ;
        RECT 10.625 7.525 10.795 7.695 ;
        RECT 11.015 7.525 11.185 7.695 ;
        RECT 11.405 7.525 11.575 7.695 ;
        RECT 11.765 7.525 11.935 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 12.365 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 13.185400 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 12.495 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 3.045 -0.075 3.615 -0.065 ;
        RECT 6.375 -0.075 6.945 -0.065 ;
        RECT 9.705 -0.075 10.275 -0.065 ;
        RECT 11.925 -0.075 12.495 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 1.095 0.310 1.265 1.260 ;
        RECT 3.175 0.310 3.485 2.860 ;
        RECT 3.940 0.755 4.110 1.885 ;
        RECT 4.910 0.755 5.080 1.530 ;
        RECT 5.880 0.755 6.050 1.530 ;
        RECT 3.940 0.585 6.050 0.755 ;
        RECT 3.940 0.310 4.110 0.585 ;
        RECT 4.425 0.310 4.595 0.585 ;
        RECT 4.910 0.310 5.080 0.585 ;
        RECT 5.395 0.310 5.565 0.585 ;
        RECT 5.880 0.310 6.050 0.585 ;
        RECT 6.505 0.310 6.815 2.860 ;
        RECT 7.755 0.310 7.925 1.260 ;
        RECT 9.835 0.310 10.145 2.860 ;
        RECT 10.535 0.755 10.705 1.885 ;
        RECT 11.505 0.755 11.675 1.885 ;
        RECT 10.535 0.585 11.675 0.755 ;
        RECT 10.535 0.310 10.705 0.585 ;
        RECT 11.020 0.310 11.190 0.585 ;
        RECT 11.505 0.310 11.675 0.585 ;
        RECT 12.055 0.310 12.365 2.860 ;
        RECT -0.155 0.000 12.365 0.310 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 0.995 0.065 1.165 0.235 ;
        RECT 1.355 0.065 1.525 0.235 ;
        RECT 1.805 0.065 1.975 0.235 ;
        RECT 2.165 0.065 2.335 0.235 ;
        RECT 2.525 0.065 2.695 0.235 ;
        RECT 2.885 0.065 3.055 0.235 ;
        RECT 3.605 0.065 3.775 0.235 ;
        RECT 3.965 0.065 4.135 0.235 ;
        RECT 4.325 0.065 4.495 0.235 ;
        RECT 4.685 0.065 4.855 0.235 ;
        RECT 5.135 0.065 5.305 0.235 ;
        RECT 5.495 0.065 5.665 0.235 ;
        RECT 5.855 0.065 6.025 0.235 ;
        RECT 6.215 0.065 6.385 0.235 ;
        RECT 6.935 0.065 7.105 0.235 ;
        RECT 7.295 0.065 7.465 0.235 ;
        RECT 7.655 0.065 7.825 0.235 ;
        RECT 8.015 0.065 8.185 0.235 ;
        RECT 8.465 0.065 8.635 0.235 ;
        RECT 8.825 0.065 8.995 0.235 ;
        RECT 9.185 0.065 9.355 0.235 ;
        RECT 9.545 0.065 9.715 0.235 ;
        RECT 10.265 0.065 10.435 0.235 ;
        RECT 10.625 0.065 10.795 0.235 ;
        RECT 11.015 0.065 11.185 0.235 ;
        RECT 11.405 0.065 11.575 0.235 ;
        RECT 11.765 0.065 11.935 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 12.365 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 1.145 5.515 1.315 7.250 ;
        RECT 2.025 5.515 2.195 7.250 ;
        RECT 4.035 5.525 4.205 7.255 ;
        RECT 4.915 7.055 5.965 7.225 ;
        RECT 4.915 5.525 5.085 7.055 ;
        RECT 1.145 5.345 2.675 5.515 ;
        RECT 4.035 5.355 5.085 5.525 ;
        RECT 5.355 5.525 5.525 6.795 ;
        RECT 5.795 5.785 5.965 7.055 ;
        RECT 5.355 5.355 6.005 5.525 ;
        RECT 0.610 1.805 0.780 1.885 ;
        RECT 1.580 1.805 1.750 1.885 ;
        RECT 2.505 1.880 2.675 5.345 ;
        RECT 4.200 4.940 4.370 5.100 ;
        RECT 4.200 4.770 4.525 4.940 ;
        RECT 4.355 2.055 4.525 4.770 ;
        RECT 5.835 1.880 6.005 5.355 ;
        RECT 7.805 5.515 7.975 7.250 ;
        RECT 8.685 5.515 8.855 7.250 ;
        RECT 7.805 5.345 9.335 5.515 ;
        RECT 7.685 2.055 7.855 5.095 ;
        RECT 0.610 1.635 1.750 1.805 ;
        RECT 0.610 0.505 0.780 1.635 ;
        RECT 1.580 0.755 1.750 1.635 ;
        RECT 2.065 1.710 2.675 1.880 ;
        RECT 4.425 1.710 6.005 1.880 ;
        RECT 7.270 1.805 7.440 1.885 ;
        RECT 8.240 1.805 8.410 1.885 ;
        RECT 9.165 1.880 9.335 5.345 ;
        RECT 10.645 2.055 10.815 5.095 ;
        RECT 2.065 0.975 2.235 1.710 ;
        RECT 2.550 0.755 2.720 1.525 ;
        RECT 4.425 0.975 4.595 1.710 ;
        RECT 5.395 0.975 5.565 1.710 ;
        RECT 7.270 1.635 8.410 1.805 ;
        RECT 1.580 0.585 2.720 0.755 ;
        RECT 1.580 0.505 1.750 0.585 ;
        RECT 2.550 0.505 2.720 0.585 ;
        RECT 7.270 0.505 7.440 1.635 ;
        RECT 8.240 0.755 8.410 1.635 ;
        RECT 8.725 1.710 9.335 1.880 ;
        RECT 8.725 0.975 8.895 1.710 ;
        RECT 9.210 0.755 9.380 1.525 ;
        RECT 8.240 0.585 9.380 0.755 ;
        RECT 8.240 0.505 8.410 0.585 ;
        RECT 9.210 0.505 9.380 0.585 ;
      LAYER mcon ;
        RECT 2.505 2.505 2.675 2.675 ;
        RECT 4.355 2.505 4.525 2.675 ;
        RECT 5.835 2.505 6.005 2.675 ;
        RECT 7.685 2.505 7.855 2.675 ;
        RECT 9.165 2.505 9.335 2.675 ;
        RECT 10.645 2.505 10.815 2.675 ;
      LAYER met1 ;
        RECT 2.475 2.675 2.705 2.705 ;
        RECT 4.325 2.675 4.555 2.705 ;
        RECT 5.805 2.675 6.035 2.705 ;
        RECT 7.655 2.675 7.885 2.705 ;
        RECT 9.135 2.675 9.365 2.705 ;
        RECT 10.615 2.675 10.845 2.705 ;
        RECT 2.445 2.505 4.585 2.675 ;
        RECT 5.775 2.505 7.915 2.675 ;
        RECT 9.105 2.505 10.875 2.675 ;
        RECT 2.475 2.475 2.705 2.505 ;
        RECT 4.325 2.475 4.555 2.505 ;
        RECT 5.805 2.475 6.035 2.505 ;
        RECT 7.655 2.475 7.885 2.505 ;
        RECT 9.135 2.475 9.365 2.505 ;
        RECT 10.615 2.475 10.845 2.505 ;
  END
END AOA4X1






MACRO AOAI4X1
  CLASS BLOCK ;
  FOREIGN AOAI4X1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 10.830 BY 7.950 ;
  PIN YN
    ANTENNADIFFAREA 1.351900 ;
    PORT
      LAYER li1 ;
        RECT 7.805 5.515 7.975 7.250 ;
        RECT 8.685 5.515 8.855 7.250 ;
        RECT 7.805 5.345 9.335 5.515 ;
        RECT 9.165 1.880 9.335 5.345 ;
        RECT 8.725 1.710 9.335 1.880 ;
        RECT 8.725 0.975 8.895 1.710 ;
      LAYER mcon ;
        RECT 9.165 2.875 9.335 3.045 ;
      LAYER met1 ;
        RECT 9.135 3.045 9.365 3.075 ;
        RECT 9.105 2.875 9.515 3.045 ;
        RECT 9.135 2.845 9.365 2.875 ;
    END
  END YN
  PIN A
    ANTENNAGATEAREA 1.033250 ;
    PORT
      LAYER li1 ;
        RECT 1.025 2.055 1.195 5.095 ;
      LAYER mcon ;
        RECT 1.025 2.875 1.195 3.045 ;
      LAYER met1 ;
        RECT 0.995 3.045 1.225 3.075 ;
        RECT 0.845 2.875 1.255 3.045 ;
        RECT 0.995 2.845 1.225 2.875 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 1.027250 ;
    PORT
      LAYER li1 ;
        RECT 1.795 4.940 1.965 5.095 ;
        RECT 1.765 4.765 1.965 4.940 ;
        RECT 1.765 2.055 1.935 4.765 ;
      LAYER mcon ;
        RECT 1.765 3.245 1.935 3.415 ;
      LAYER met1 ;
        RECT 1.735 3.415 1.965 3.445 ;
        RECT 1.585 3.245 1.995 3.415 ;
        RECT 1.735 3.215 1.965 3.245 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA 1.026450 ;
    PORT
      LAYER li1 ;
        RECT 5.130 4.940 5.300 5.100 ;
        RECT 5.095 4.770 5.300 4.940 ;
        RECT 5.095 2.055 5.265 4.770 ;
      LAYER mcon ;
        RECT 5.095 3.615 5.265 3.785 ;
      LAYER met1 ;
        RECT 5.065 3.785 5.295 3.815 ;
        RECT 4.915 3.615 5.325 3.785 ;
        RECT 5.065 3.585 5.295 3.615 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA 1.027250 ;
    PORT
      LAYER li1 ;
        RECT 8.455 4.940 8.625 5.095 ;
        RECT 8.425 4.765 8.625 4.940 ;
        RECT 8.425 2.055 8.595 4.765 ;
      LAYER mcon ;
        RECT 8.425 3.985 8.595 4.155 ;
      LAYER met1 ;
        RECT 8.395 4.155 8.625 4.185 ;
        RECT 8.245 3.985 8.655 4.155 ;
        RECT 8.395 3.955 8.625 3.985 ;
    END
  END D
  PIN VDD
    ANTENNADIFFAREA 12.448999 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 10.410 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 10.145 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 0.705 5.365 0.875 7.460 ;
        RECT 1.585 5.785 1.755 7.460 ;
        RECT 2.465 5.785 2.635 7.460 ;
        RECT 3.175 4.340 3.485 7.460 ;
        RECT 4.475 5.785 4.645 7.460 ;
        RECT 6.505 4.340 6.815 7.460 ;
        RECT 7.365 5.365 7.535 7.460 ;
        RECT 8.245 5.785 8.415 7.460 ;
        RECT 9.125 5.785 9.295 7.460 ;
        RECT 9.835 4.340 10.145 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 0.995 7.525 1.165 7.695 ;
        RECT 1.355 7.525 1.525 7.695 ;
        RECT 1.805 7.525 1.975 7.695 ;
        RECT 2.165 7.525 2.335 7.695 ;
        RECT 2.525 7.525 2.695 7.695 ;
        RECT 2.885 7.525 3.055 7.695 ;
        RECT 3.605 7.525 3.775 7.695 ;
        RECT 3.965 7.525 4.135 7.695 ;
        RECT 4.325 7.525 4.495 7.695 ;
        RECT 4.685 7.525 4.855 7.695 ;
        RECT 5.135 7.525 5.305 7.695 ;
        RECT 5.495 7.525 5.665 7.695 ;
        RECT 5.855 7.525 6.025 7.695 ;
        RECT 6.215 7.525 6.385 7.695 ;
        RECT 6.935 7.525 7.105 7.695 ;
        RECT 7.295 7.525 7.465 7.695 ;
        RECT 7.655 7.525 7.825 7.695 ;
        RECT 8.015 7.525 8.185 7.695 ;
        RECT 8.465 7.525 8.635 7.695 ;
        RECT 8.825 7.525 8.995 7.695 ;
        RECT 9.185 7.525 9.355 7.695 ;
        RECT 9.545 7.525 9.715 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 10.145 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 10.221300 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 10.275 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 3.045 -0.075 3.615 -0.065 ;
        RECT 6.375 -0.075 6.945 -0.065 ;
        RECT 9.705 -0.075 10.275 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 1.095 0.310 1.265 1.260 ;
        RECT 3.175 0.310 3.485 2.860 ;
        RECT 3.940 0.755 4.110 1.885 ;
        RECT 4.910 0.755 5.080 1.530 ;
        RECT 5.880 0.755 6.050 1.530 ;
        RECT 3.940 0.585 6.050 0.755 ;
        RECT 3.940 0.310 4.110 0.585 ;
        RECT 4.425 0.310 4.595 0.585 ;
        RECT 4.910 0.310 5.080 0.585 ;
        RECT 5.395 0.310 5.565 0.585 ;
        RECT 5.880 0.310 6.050 0.585 ;
        RECT 6.505 0.310 6.815 2.860 ;
        RECT 7.755 0.310 7.925 1.260 ;
        RECT 9.835 0.310 10.145 2.860 ;
        RECT -0.155 0.000 10.145 0.310 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 0.995 0.065 1.165 0.235 ;
        RECT 1.355 0.065 1.525 0.235 ;
        RECT 1.805 0.065 1.975 0.235 ;
        RECT 2.165 0.065 2.335 0.235 ;
        RECT 2.525 0.065 2.695 0.235 ;
        RECT 2.885 0.065 3.055 0.235 ;
        RECT 3.605 0.065 3.775 0.235 ;
        RECT 3.965 0.065 4.135 0.235 ;
        RECT 4.325 0.065 4.495 0.235 ;
        RECT 4.685 0.065 4.855 0.235 ;
        RECT 5.135 0.065 5.305 0.235 ;
        RECT 5.495 0.065 5.665 0.235 ;
        RECT 5.855 0.065 6.025 0.235 ;
        RECT 6.215 0.065 6.385 0.235 ;
        RECT 6.935 0.065 7.105 0.235 ;
        RECT 7.295 0.065 7.465 0.235 ;
        RECT 7.655 0.065 7.825 0.235 ;
        RECT 8.015 0.065 8.185 0.235 ;
        RECT 8.465 0.065 8.635 0.235 ;
        RECT 8.825 0.065 8.995 0.235 ;
        RECT 9.185 0.065 9.355 0.235 ;
        RECT 9.545 0.065 9.715 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 10.145 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 1.145 5.515 1.315 7.250 ;
        RECT 2.025 5.515 2.195 7.250 ;
        RECT 4.035 5.525 4.205 7.255 ;
        RECT 4.915 7.055 5.965 7.225 ;
        RECT 4.915 5.525 5.085 7.055 ;
        RECT 1.145 5.345 2.675 5.515 ;
        RECT 4.035 5.355 5.085 5.525 ;
        RECT 5.355 5.525 5.525 6.795 ;
        RECT 5.795 5.785 5.965 7.055 ;
        RECT 5.355 5.355 6.005 5.525 ;
        RECT 0.610 1.805 0.780 1.885 ;
        RECT 1.580 1.805 1.750 1.885 ;
        RECT 2.505 1.880 2.675 5.345 ;
        RECT 4.200 4.940 4.370 5.100 ;
        RECT 4.200 4.770 4.525 4.940 ;
        RECT 4.355 2.055 4.525 4.770 ;
        RECT 5.835 1.880 6.005 5.355 ;
        RECT 7.685 2.055 7.855 5.095 ;
        RECT 0.610 1.635 1.750 1.805 ;
        RECT 0.610 0.505 0.780 1.635 ;
        RECT 1.580 0.755 1.750 1.635 ;
        RECT 2.065 1.710 2.675 1.880 ;
        RECT 4.425 1.710 6.005 1.880 ;
        RECT 7.270 1.805 7.440 1.885 ;
        RECT 8.240 1.805 8.410 1.885 ;
        RECT 2.065 0.975 2.235 1.710 ;
        RECT 2.550 0.755 2.720 1.525 ;
        RECT 4.425 0.975 4.595 1.710 ;
        RECT 5.395 0.975 5.565 1.710 ;
        RECT 7.270 1.635 8.410 1.805 ;
        RECT 1.580 0.585 2.720 0.755 ;
        RECT 1.580 0.505 1.750 0.585 ;
        RECT 2.550 0.505 2.720 0.585 ;
        RECT 7.270 0.505 7.440 1.635 ;
        RECT 8.240 0.755 8.410 1.635 ;
        RECT 9.210 0.755 9.380 1.525 ;
        RECT 8.240 0.585 9.380 0.755 ;
        RECT 8.240 0.505 8.410 0.585 ;
        RECT 9.210 0.505 9.380 0.585 ;
      LAYER mcon ;
        RECT 2.505 2.505 2.675 2.675 ;
        RECT 4.355 2.505 4.525 2.675 ;
        RECT 5.835 2.505 6.005 2.675 ;
        RECT 7.685 2.505 7.855 2.675 ;
      LAYER met1 ;
        RECT 2.475 2.675 2.705 2.705 ;
        RECT 4.325 2.675 4.555 2.705 ;
        RECT 5.805 2.675 6.035 2.705 ;
        RECT 7.655 2.675 7.885 2.705 ;
        RECT 2.445 2.505 4.585 2.675 ;
        RECT 5.775 2.505 7.915 2.675 ;
        RECT 2.475 2.475 2.705 2.505 ;
        RECT 4.325 2.475 4.555 2.505 ;
        RECT 5.805 2.475 6.035 2.505 ;
        RECT 7.655 2.475 7.885 2.505 ;
  END
END AOAI4X1






MACRO AOI3X1
  CLASS BLOCK ;
  FOREIGN AOI3X1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 7.500 BY 7.950 ;
  PIN YN
    ANTENNADIFFAREA 0.963050 ;
    PORT
      LAYER li1 ;
        RECT 5.355 5.525 5.525 6.795 ;
        RECT 5.355 5.355 6.005 5.525 ;
        RECT 5.835 1.880 6.005 5.355 ;
        RECT 4.425 1.710 6.005 1.880 ;
        RECT 4.425 0.975 4.595 1.710 ;
        RECT 5.395 0.975 5.565 1.710 ;
      LAYER mcon ;
        RECT 5.835 3.985 6.005 4.155 ;
      LAYER met1 ;
        RECT 5.805 4.155 6.035 4.185 ;
        RECT 5.775 3.985 6.185 4.155 ;
        RECT 5.805 3.955 6.035 3.985 ;
    END
  END YN
  PIN A
    ANTENNAGATEAREA 1.033250 ;
    PORT
      LAYER li1 ;
        RECT 1.025 2.055 1.195 5.095 ;
      LAYER mcon ;
        RECT 1.025 2.875 1.195 3.045 ;
      LAYER met1 ;
        RECT 0.995 3.045 1.225 3.075 ;
        RECT 0.845 2.875 1.255 3.045 ;
        RECT 0.995 2.845 1.225 2.875 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 1.027250 ;
    PORT
      LAYER li1 ;
        RECT 1.795 4.940 1.965 5.095 ;
        RECT 1.765 4.765 1.965 4.940 ;
        RECT 1.765 2.055 1.935 4.765 ;
      LAYER mcon ;
        RECT 1.765 3.245 1.935 3.415 ;
      LAYER met1 ;
        RECT 1.735 3.415 1.965 3.445 ;
        RECT 1.585 3.245 1.995 3.415 ;
        RECT 1.735 3.215 1.965 3.245 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA 1.026450 ;
    PORT
      LAYER li1 ;
        RECT 5.130 4.940 5.300 5.100 ;
        RECT 5.095 4.770 5.300 4.940 ;
        RECT 5.095 2.055 5.265 4.770 ;
      LAYER mcon ;
        RECT 5.095 3.615 5.265 3.785 ;
      LAYER met1 ;
        RECT 5.065 3.785 5.295 3.815 ;
        RECT 4.915 3.615 5.325 3.785 ;
        RECT 5.065 3.585 5.295 3.615 ;
    END
  END C
  PIN VDD
    ANTENNADIFFAREA 8.279349 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 7.080 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 6.815 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 0.705 5.365 0.875 7.460 ;
        RECT 1.585 5.785 1.755 7.460 ;
        RECT 2.465 5.785 2.635 7.460 ;
        RECT 3.175 4.340 3.485 7.460 ;
        RECT 4.475 5.785 4.645 7.460 ;
        RECT 6.505 4.340 6.815 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 0.995 7.525 1.165 7.695 ;
        RECT 1.355 7.525 1.525 7.695 ;
        RECT 1.805 7.525 1.975 7.695 ;
        RECT 2.165 7.525 2.335 7.695 ;
        RECT 2.525 7.525 2.695 7.695 ;
        RECT 2.885 7.525 3.055 7.695 ;
        RECT 3.605 7.525 3.775 7.695 ;
        RECT 3.965 7.525 4.135 7.695 ;
        RECT 4.325 7.525 4.495 7.695 ;
        RECT 4.685 7.525 4.855 7.695 ;
        RECT 5.135 7.525 5.305 7.695 ;
        RECT 5.495 7.525 5.665 7.695 ;
        RECT 5.855 7.525 6.025 7.695 ;
        RECT 6.215 7.525 6.385 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 6.815 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 7.710250 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 6.945 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 3.045 -0.075 3.615 -0.065 ;
        RECT 6.375 -0.075 6.945 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 1.095 0.310 1.265 1.260 ;
        RECT 3.175 0.310 3.485 2.860 ;
        RECT 3.940 0.755 4.110 1.885 ;
        RECT 4.910 0.755 5.080 1.530 ;
        RECT 5.880 0.755 6.050 1.530 ;
        RECT 3.940 0.585 6.050 0.755 ;
        RECT 3.940 0.310 4.110 0.585 ;
        RECT 4.425 0.310 4.595 0.585 ;
        RECT 4.910 0.310 5.080 0.585 ;
        RECT 5.395 0.310 5.565 0.585 ;
        RECT 5.880 0.310 6.050 0.585 ;
        RECT 6.505 0.310 6.815 2.860 ;
        RECT -0.155 0.000 6.815 0.310 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 0.995 0.065 1.165 0.235 ;
        RECT 1.355 0.065 1.525 0.235 ;
        RECT 1.805 0.065 1.975 0.235 ;
        RECT 2.165 0.065 2.335 0.235 ;
        RECT 2.525 0.065 2.695 0.235 ;
        RECT 2.885 0.065 3.055 0.235 ;
        RECT 3.605 0.065 3.775 0.235 ;
        RECT 3.965 0.065 4.135 0.235 ;
        RECT 4.325 0.065 4.495 0.235 ;
        RECT 4.685 0.065 4.855 0.235 ;
        RECT 5.135 0.065 5.305 0.235 ;
        RECT 5.495 0.065 5.665 0.235 ;
        RECT 5.855 0.065 6.025 0.235 ;
        RECT 6.215 0.065 6.385 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 6.815 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 1.145 5.515 1.315 7.250 ;
        RECT 2.025 5.515 2.195 7.250 ;
        RECT 4.035 5.525 4.205 7.255 ;
        RECT 4.915 7.055 5.965 7.225 ;
        RECT 4.915 5.525 5.085 7.055 ;
        RECT 5.795 5.785 5.965 7.055 ;
        RECT 1.145 5.345 2.675 5.515 ;
        RECT 4.035 5.355 5.085 5.525 ;
        RECT 0.610 1.805 0.780 1.885 ;
        RECT 1.580 1.805 1.750 1.885 ;
        RECT 2.505 1.880 2.675 5.345 ;
        RECT 4.200 4.940 4.370 5.100 ;
        RECT 4.200 4.770 4.525 4.940 ;
        RECT 4.355 2.055 4.525 4.770 ;
        RECT 0.610 1.635 1.750 1.805 ;
        RECT 0.610 0.505 0.780 1.635 ;
        RECT 1.580 0.755 1.750 1.635 ;
        RECT 2.065 1.710 2.675 1.880 ;
        RECT 2.065 0.975 2.235 1.710 ;
        RECT 2.550 0.755 2.720 1.525 ;
        RECT 1.580 0.585 2.720 0.755 ;
        RECT 1.580 0.505 1.750 0.585 ;
        RECT 2.550 0.505 2.720 0.585 ;
      LAYER mcon ;
        RECT 2.505 2.505 2.675 2.675 ;
        RECT 4.355 2.505 4.525 2.675 ;
      LAYER met1 ;
        RECT 2.475 2.675 2.705 2.705 ;
        RECT 4.325 2.675 4.555 2.705 ;
        RECT 2.445 2.505 4.585 2.675 ;
        RECT 2.475 2.475 2.705 2.505 ;
        RECT 4.325 2.475 4.555 2.505 ;
  END
END AOI3X1






MACRO BUFX1
  CLASS BLOCK ;
  FOREIGN BUFX1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 5.280 BY 7.950 ;
  PIN Y
    ANTENNADIFFAREA 0.771900 ;
    PORT
      LAYER li1 ;
        RECT 3.245 4.895 3.415 7.250 ;
        RECT 3.245 4.725 3.785 4.895 ;
        RECT 3.615 2.305 3.785 4.725 ;
        RECT 3.245 2.135 3.785 2.305 ;
        RECT 3.245 0.975 3.415 2.135 ;
      LAYER mcon ;
        RECT 3.615 3.245 3.785 3.415 ;
      LAYER met1 ;
        RECT 3.585 3.415 3.815 3.445 ;
        RECT 3.555 3.245 3.965 3.415 ;
        RECT 3.585 3.215 3.815 3.245 ;
    END
  END Y
  PIN A
    ANTENNAGATEAREA 1.027250 ;
    PORT
      LAYER li1 ;
        RECT 0.655 2.055 0.825 5.095 ;
      LAYER mcon ;
        RECT 0.655 3.245 0.825 3.415 ;
      LAYER met1 ;
        RECT 0.625 3.415 0.855 3.445 ;
        RECT 0.475 3.245 0.885 3.415 ;
        RECT 0.625 3.215 0.855 3.245 ;
    END
  END A
  PIN VDD
    ANTENNADIFFAREA 7.153750 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 4.860 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 4.595 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 0.585 5.415 0.755 7.460 ;
        RECT 1.465 5.415 1.635 7.460 ;
        RECT 2.065 4.340 2.375 7.460 ;
        RECT 2.805 5.415 2.975 7.460 ;
        RECT 3.685 5.415 3.855 7.460 ;
        RECT 4.285 4.340 4.595 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 1.025 7.525 1.195 7.695 ;
        RECT 1.415 7.525 1.585 7.695 ;
        RECT 1.775 7.525 1.945 7.695 ;
        RECT 2.495 7.525 2.665 7.695 ;
        RECT 2.855 7.525 3.025 7.695 ;
        RECT 3.245 7.525 3.415 7.695 ;
        RECT 3.635 7.525 3.805 7.695 ;
        RECT 3.995 7.525 4.165 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 4.595 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 6.797750 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 4.725 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 1.935 -0.075 2.505 -0.065 ;
        RECT 4.155 -0.075 4.725 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 0.545 0.755 0.715 1.885 ;
        RECT 1.515 0.755 1.685 1.885 ;
        RECT 0.545 0.585 1.685 0.755 ;
        RECT 0.545 0.310 0.715 0.585 ;
        RECT 1.030 0.310 1.200 0.585 ;
        RECT 1.515 0.310 1.685 0.585 ;
        RECT 2.065 0.310 2.375 2.860 ;
        RECT 2.765 0.755 2.935 1.885 ;
        RECT 3.735 0.755 3.905 1.885 ;
        RECT 2.765 0.585 3.905 0.755 ;
        RECT 2.765 0.310 2.935 0.585 ;
        RECT 3.250 0.310 3.420 0.585 ;
        RECT 3.735 0.310 3.905 0.585 ;
        RECT 4.285 0.310 4.595 2.860 ;
        RECT -0.155 0.000 4.595 0.310 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 1.025 0.065 1.195 0.235 ;
        RECT 1.415 0.065 1.585 0.235 ;
        RECT 1.775 0.065 1.945 0.235 ;
        RECT 2.495 0.065 2.665 0.235 ;
        RECT 2.855 0.065 3.025 0.235 ;
        RECT 3.245 0.065 3.415 0.235 ;
        RECT 3.635 0.065 3.805 0.235 ;
        RECT 3.995 0.065 4.165 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 4.595 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 1.025 4.895 1.195 7.250 ;
        RECT 1.025 4.725 1.565 4.895 ;
        RECT 1.395 2.305 1.565 4.725 ;
        RECT 1.025 2.135 1.565 2.305 ;
        RECT 1.025 0.975 1.195 2.135 ;
        RECT 2.875 2.055 3.045 5.095 ;
      LAYER mcon ;
        RECT 1.395 2.505 1.565 2.675 ;
        RECT 2.875 2.505 3.045 2.675 ;
      LAYER met1 ;
        RECT 1.365 2.675 1.595 2.705 ;
        RECT 2.845 2.675 3.075 2.705 ;
        RECT 1.335 2.505 3.105 2.675 ;
        RECT 1.365 2.475 1.595 2.505 ;
        RECT 2.845 2.475 3.075 2.505 ;
  END
END BUFX1






MACRO DFFQNX1
  CLASS BLOCK ;
  FOREIGN DFFQNX1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 22.300 BY 7.950 ;
  PIN QN
    ANTENNAGATEAREA 1.033250 ;
    ANTENNADIFFAREA 1.351900 ;
    PORT
      LAYER li1 ;
        RECT 15.945 5.515 16.115 7.250 ;
        RECT 16.825 5.515 16.995 7.250 ;
        RECT 15.945 5.345 17.475 5.515 ;
        RECT 17.305 1.880 17.475 5.345 ;
        RECT 19.155 2.055 19.325 5.095 ;
        RECT 16.865 1.710 17.475 1.880 ;
        RECT 16.865 0.975 17.035 1.710 ;
      LAYER mcon ;
        RECT 17.305 3.615 17.475 3.785 ;
        RECT 19.155 3.615 19.325 3.785 ;
      LAYER met1 ;
        RECT 17.275 3.785 17.505 3.815 ;
        RECT 19.125 3.785 19.355 3.815 ;
        RECT 17.245 3.615 19.385 3.785 ;
        RECT 17.275 3.585 17.505 3.615 ;
        RECT 19.125 3.585 19.355 3.615 ;
    END
  END QN
  PIN D
    ANTENNAGATEAREA 1.027250 ;
    PORT
      LAYER li1 ;
        RECT 6.605 4.940 6.775 5.095 ;
        RECT 6.575 4.765 6.775 4.940 ;
        RECT 6.575 2.055 6.745 4.765 ;
      LAYER mcon ;
        RECT 6.575 3.245 6.745 3.415 ;
        RECT 6.575 2.135 6.745 2.305 ;
      LAYER met1 ;
        RECT 6.545 3.415 6.775 3.445 ;
        RECT 6.395 3.245 6.805 3.415 ;
        RECT 6.545 3.215 6.775 3.245 ;
        RECT 6.545 2.305 6.775 2.335 ;
        RECT 6.395 2.135 6.805 2.305 ;
        RECT 6.545 2.105 6.775 2.135 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 2.042100 ;
    PORT
      LAYER li1 ;
        RECT 2.135 2.055 2.305 5.095 ;
        RECT 13.265 4.975 13.435 5.095 ;
        RECT 13.235 4.765 13.435 4.975 ;
        RECT 13.235 2.055 13.405 4.765 ;
      LAYER mcon ;
        RECT 2.135 4.725 2.305 4.895 ;
        RECT 13.235 4.725 13.405 4.895 ;
      LAYER met1 ;
        RECT 2.105 4.895 2.335 4.925 ;
        RECT 13.205 4.895 13.435 4.925 ;
        RECT 2.075 4.725 13.465 4.895 ;
        RECT 2.105 4.695 2.335 4.725 ;
        RECT 13.205 4.695 13.435 4.725 ;
    END
  END CLK
  PIN VDD
    ANTENNADIFFAREA 27.348349 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 21.880 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 21.615 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 1.005 5.445 1.175 7.460 ;
        RECT 1.885 5.785 2.055 7.460 ;
        RECT 2.765 5.785 2.935 7.460 ;
        RECT 3.645 5.785 3.815 7.460 ;
        RECT 4.655 4.340 4.965 7.460 ;
        RECT 5.515 5.365 5.685 7.460 ;
        RECT 6.395 5.785 6.565 7.460 ;
        RECT 7.275 5.785 7.445 7.460 ;
        RECT 7.985 4.340 8.295 7.460 ;
        RECT 8.845 5.365 9.015 7.460 ;
        RECT 9.725 5.785 9.895 7.460 ;
        RECT 10.605 5.785 10.775 7.460 ;
        RECT 11.315 4.340 11.625 7.460 ;
        RECT 12.175 5.365 12.345 7.460 ;
        RECT 13.055 5.785 13.225 7.460 ;
        RECT 13.935 5.785 14.105 7.460 ;
        RECT 14.645 4.340 14.955 7.460 ;
        RECT 15.505 5.365 15.675 7.460 ;
        RECT 16.385 5.785 16.555 7.460 ;
        RECT 17.265 5.785 17.435 7.460 ;
        RECT 17.975 4.340 18.285 7.460 ;
        RECT 18.835 5.365 19.005 7.460 ;
        RECT 19.715 5.785 19.885 7.460 ;
        RECT 20.595 5.785 20.765 7.460 ;
        RECT 21.305 4.340 21.615 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 0.995 7.525 1.165 7.695 ;
        RECT 1.355 7.525 1.525 7.695 ;
        RECT 1.715 7.525 1.885 7.695 ;
        RECT 2.075 7.525 2.245 7.695 ;
        RECT 2.565 7.525 2.735 7.695 ;
        RECT 2.925 7.525 3.095 7.695 ;
        RECT 3.285 7.525 3.455 7.695 ;
        RECT 3.645 7.525 3.815 7.695 ;
        RECT 4.005 7.525 4.175 7.695 ;
        RECT 4.365 7.525 4.535 7.695 ;
        RECT 5.085 7.525 5.255 7.695 ;
        RECT 5.445 7.525 5.615 7.695 ;
        RECT 5.805 7.525 5.975 7.695 ;
        RECT 6.165 7.525 6.335 7.695 ;
        RECT 6.615 7.525 6.785 7.695 ;
        RECT 6.975 7.525 7.145 7.695 ;
        RECT 7.335 7.525 7.505 7.695 ;
        RECT 7.695 7.525 7.865 7.695 ;
        RECT 8.415 7.525 8.585 7.695 ;
        RECT 8.775 7.525 8.945 7.695 ;
        RECT 9.135 7.525 9.305 7.695 ;
        RECT 9.495 7.525 9.665 7.695 ;
        RECT 9.945 7.525 10.115 7.695 ;
        RECT 10.305 7.525 10.475 7.695 ;
        RECT 10.665 7.525 10.835 7.695 ;
        RECT 11.025 7.525 11.195 7.695 ;
        RECT 11.745 7.525 11.915 7.695 ;
        RECT 12.105 7.525 12.275 7.695 ;
        RECT 12.465 7.525 12.635 7.695 ;
        RECT 12.825 7.525 12.995 7.695 ;
        RECT 13.275 7.525 13.445 7.695 ;
        RECT 13.635 7.525 13.805 7.695 ;
        RECT 13.995 7.525 14.165 7.695 ;
        RECT 14.355 7.525 14.525 7.695 ;
        RECT 15.075 7.525 15.245 7.695 ;
        RECT 15.435 7.525 15.605 7.695 ;
        RECT 15.795 7.525 15.965 7.695 ;
        RECT 16.155 7.525 16.325 7.695 ;
        RECT 16.605 7.525 16.775 7.695 ;
        RECT 16.965 7.525 17.135 7.695 ;
        RECT 17.325 7.525 17.495 7.695 ;
        RECT 17.685 7.525 17.855 7.695 ;
        RECT 18.405 7.525 18.575 7.695 ;
        RECT 18.765 7.525 18.935 7.695 ;
        RECT 19.125 7.525 19.295 7.695 ;
        RECT 19.485 7.525 19.655 7.695 ;
        RECT 19.935 7.525 20.105 7.695 ;
        RECT 20.295 7.525 20.465 7.695 ;
        RECT 20.655 7.525 20.825 7.695 ;
        RECT 21.015 7.525 21.185 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 21.615 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 16.646250 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 21.745 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 4.525 -0.075 5.095 -0.065 ;
        RECT 7.855 -0.075 8.425 -0.065 ;
        RECT 11.185 -0.075 11.755 -0.065 ;
        RECT 14.515 -0.075 15.085 -0.065 ;
        RECT 17.845 -0.075 18.415 -0.065 ;
        RECT 21.175 -0.075 21.745 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 0.990 0.310 1.160 1.270 ;
        RECT 4.655 0.310 4.965 2.860 ;
        RECT 5.905 0.310 6.075 1.260 ;
        RECT 7.985 0.310 8.295 2.860 ;
        RECT 9.235 0.310 9.405 1.260 ;
        RECT 11.315 0.310 11.625 2.860 ;
        RECT 12.565 0.310 12.735 1.260 ;
        RECT 14.645 0.310 14.955 2.860 ;
        RECT 15.895 0.310 16.065 1.260 ;
        RECT 17.975 0.310 18.285 2.860 ;
        RECT 19.225 0.310 19.395 1.260 ;
        RECT 21.305 0.310 21.615 2.860 ;
        RECT -0.155 0.000 21.615 0.310 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 0.995 0.065 1.165 0.235 ;
        RECT 1.355 0.065 1.525 0.235 ;
        RECT 1.715 0.065 1.885 0.235 ;
        RECT 2.075 0.065 2.245 0.235 ;
        RECT 2.565 0.065 2.735 0.235 ;
        RECT 2.925 0.065 3.095 0.235 ;
        RECT 3.285 0.065 3.455 0.235 ;
        RECT 3.645 0.065 3.815 0.235 ;
        RECT 4.005 0.065 4.175 0.235 ;
        RECT 4.365 0.065 4.535 0.235 ;
        RECT 5.085 0.065 5.255 0.235 ;
        RECT 5.445 0.065 5.615 0.235 ;
        RECT 5.805 0.065 5.975 0.235 ;
        RECT 6.165 0.065 6.335 0.235 ;
        RECT 6.615 0.065 6.785 0.235 ;
        RECT 6.975 0.065 7.145 0.235 ;
        RECT 7.335 0.065 7.505 0.235 ;
        RECT 7.695 0.065 7.865 0.235 ;
        RECT 8.415 0.065 8.585 0.235 ;
        RECT 8.775 0.065 8.945 0.235 ;
        RECT 9.135 0.065 9.305 0.235 ;
        RECT 9.495 0.065 9.665 0.235 ;
        RECT 9.945 0.065 10.115 0.235 ;
        RECT 10.305 0.065 10.475 0.235 ;
        RECT 10.665 0.065 10.835 0.235 ;
        RECT 11.025 0.065 11.195 0.235 ;
        RECT 11.745 0.065 11.915 0.235 ;
        RECT 12.105 0.065 12.275 0.235 ;
        RECT 12.465 0.065 12.635 0.235 ;
        RECT 12.825 0.065 12.995 0.235 ;
        RECT 13.275 0.065 13.445 0.235 ;
        RECT 13.635 0.065 13.805 0.235 ;
        RECT 13.995 0.065 14.165 0.235 ;
        RECT 14.355 0.065 14.525 0.235 ;
        RECT 15.075 0.065 15.245 0.235 ;
        RECT 15.435 0.065 15.605 0.235 ;
        RECT 15.795 0.065 15.965 0.235 ;
        RECT 16.155 0.065 16.325 0.235 ;
        RECT 16.605 0.065 16.775 0.235 ;
        RECT 16.965 0.065 17.135 0.235 ;
        RECT 17.325 0.065 17.495 0.235 ;
        RECT 17.685 0.065 17.855 0.235 ;
        RECT 18.405 0.065 18.575 0.235 ;
        RECT 18.765 0.065 18.935 0.235 ;
        RECT 19.125 0.065 19.295 0.235 ;
        RECT 19.485 0.065 19.655 0.235 ;
        RECT 19.935 0.065 20.105 0.235 ;
        RECT 20.295 0.065 20.465 0.235 ;
        RECT 20.655 0.065 20.825 0.235 ;
        RECT 21.015 0.065 21.185 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 21.615 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 1.445 5.470 1.615 7.250 ;
        RECT 2.325 5.470 2.495 7.250 ;
        RECT 3.205 5.470 3.375 7.250 ;
        RECT 5.955 5.515 6.125 7.250 ;
        RECT 6.835 5.515 7.005 7.250 ;
        RECT 9.285 5.515 9.455 7.250 ;
        RECT 10.165 5.515 10.335 7.250 ;
        RECT 12.615 5.515 12.785 7.250 ;
        RECT 13.495 5.515 13.665 7.250 ;
        RECT 19.275 5.515 19.445 7.250 ;
        RECT 20.155 5.515 20.325 7.250 ;
        RECT 1.445 5.300 4.155 5.470 ;
        RECT 5.955 5.345 7.485 5.515 ;
        RECT 9.285 5.345 10.815 5.515 ;
        RECT 12.615 5.345 14.145 5.515 ;
        RECT 19.275 5.345 20.805 5.515 ;
        RECT 1.025 2.055 1.195 5.095 ;
        RECT 3.245 2.055 3.415 5.095 ;
        RECT 0.505 1.815 0.675 1.895 ;
        RECT 1.475 1.815 1.645 1.895 ;
        RECT 2.445 1.815 2.615 1.895 ;
        RECT 0.505 1.645 2.615 1.815 ;
        RECT 0.505 0.515 0.675 1.645 ;
        RECT 1.475 0.765 1.645 1.645 ;
        RECT 2.445 1.565 2.615 1.645 ;
        RECT 1.965 1.220 2.135 1.300 ;
        RECT 3.015 1.220 3.185 1.895 ;
        RECT 3.985 1.890 4.155 5.300 ;
        RECT 5.835 2.055 6.005 5.095 ;
        RECT 1.965 1.050 3.185 1.220 ;
        RECT 1.965 0.970 2.135 1.050 ;
        RECT 2.445 0.765 2.615 0.845 ;
        RECT 1.475 0.595 2.615 0.765 ;
        RECT 1.475 0.515 1.645 0.595 ;
        RECT 2.445 0.515 2.615 0.595 ;
        RECT 3.015 0.765 3.185 1.050 ;
        RECT 3.500 1.720 4.155 1.890 ;
        RECT 5.420 1.805 5.590 1.885 ;
        RECT 6.390 1.805 6.560 1.885 ;
        RECT 7.315 1.880 7.485 5.345 ;
        RECT 9.165 2.055 9.335 5.095 ;
        RECT 9.935 4.940 10.105 5.095 ;
        RECT 9.905 4.765 10.105 4.940 ;
        RECT 9.905 2.055 10.075 4.765 ;
        RECT 3.500 0.985 3.670 1.720 ;
        RECT 5.420 1.635 6.560 1.805 ;
        RECT 3.985 0.765 4.155 1.535 ;
        RECT 3.015 0.595 4.155 0.765 ;
        RECT 3.015 0.515 3.185 0.595 ;
        RECT 3.985 0.515 4.155 0.595 ;
        RECT 5.420 0.505 5.590 1.635 ;
        RECT 6.390 0.755 6.560 1.635 ;
        RECT 6.875 1.710 7.485 1.880 ;
        RECT 8.750 1.805 8.920 1.885 ;
        RECT 9.720 1.805 9.890 1.885 ;
        RECT 10.645 1.880 10.815 5.345 ;
        RECT 12.495 2.055 12.665 5.095 ;
        RECT 6.875 0.975 7.045 1.710 ;
        RECT 8.750 1.635 9.890 1.805 ;
        RECT 7.360 0.755 7.530 1.525 ;
        RECT 6.390 0.585 7.530 0.755 ;
        RECT 6.390 0.505 6.560 0.585 ;
        RECT 7.360 0.505 7.530 0.585 ;
        RECT 8.750 0.505 8.920 1.635 ;
        RECT 9.720 0.755 9.890 1.635 ;
        RECT 10.205 1.710 10.815 1.880 ;
        RECT 12.080 1.805 12.250 1.885 ;
        RECT 13.050 1.805 13.220 1.885 ;
        RECT 13.975 1.880 14.145 5.345 ;
        RECT 15.825 2.055 15.995 5.095 ;
        RECT 16.595 4.940 16.765 5.095 ;
        RECT 19.925 4.940 20.095 5.095 ;
        RECT 16.565 4.765 16.765 4.940 ;
        RECT 19.895 4.765 20.095 4.940 ;
        RECT 16.565 2.055 16.735 4.765 ;
        RECT 19.895 2.055 20.065 4.765 ;
        RECT 10.205 0.975 10.375 1.710 ;
        RECT 12.080 1.635 13.220 1.805 ;
        RECT 10.690 0.755 10.860 1.525 ;
        RECT 9.720 0.585 10.860 0.755 ;
        RECT 9.720 0.505 9.890 0.585 ;
        RECT 10.690 0.505 10.860 0.585 ;
        RECT 12.080 0.505 12.250 1.635 ;
        RECT 13.050 0.755 13.220 1.635 ;
        RECT 13.535 1.710 14.145 1.880 ;
        RECT 15.410 1.805 15.580 1.885 ;
        RECT 16.380 1.805 16.550 1.885 ;
        RECT 13.535 0.975 13.705 1.710 ;
        RECT 15.410 1.635 16.550 1.805 ;
        RECT 14.020 0.755 14.190 1.525 ;
        RECT 13.050 0.585 14.190 0.755 ;
        RECT 13.050 0.505 13.220 0.585 ;
        RECT 14.020 0.505 14.190 0.585 ;
        RECT 15.410 0.505 15.580 1.635 ;
        RECT 16.380 0.755 16.550 1.635 ;
        RECT 18.740 1.805 18.910 1.885 ;
        RECT 19.710 1.805 19.880 1.885 ;
        RECT 20.635 1.880 20.805 5.345 ;
        RECT 18.740 1.635 19.880 1.805 ;
        RECT 17.350 0.755 17.520 1.525 ;
        RECT 16.380 0.585 17.520 0.755 ;
        RECT 16.380 0.505 16.550 0.585 ;
        RECT 17.350 0.505 17.520 0.585 ;
        RECT 18.740 0.505 18.910 1.635 ;
        RECT 19.710 0.755 19.880 1.635 ;
        RECT 20.195 1.710 20.805 1.880 ;
        RECT 20.195 0.975 20.365 1.710 ;
        RECT 20.680 0.755 20.850 1.525 ;
        RECT 19.710 0.585 20.850 0.755 ;
        RECT 19.710 0.505 19.880 0.585 ;
        RECT 20.680 0.505 20.850 0.585 ;
      LAYER mcon ;
        RECT 1.025 4.355 1.195 4.525 ;
        RECT 3.245 3.615 3.415 3.785 ;
        RECT 3.985 3.985 4.155 4.155 ;
        RECT 5.835 3.985 6.005 4.155 ;
        RECT 7.315 3.615 7.485 3.785 ;
        RECT 9.165 3.615 9.335 3.785 ;
        RECT 9.905 4.355 10.075 4.525 ;
        RECT 10.645 3.615 10.815 3.785 ;
        RECT 12.495 3.615 12.665 3.785 ;
        RECT 13.975 4.355 14.145 4.525 ;
        RECT 15.825 3.985 15.995 4.155 ;
        RECT 16.565 3.985 16.735 4.155 ;
        RECT 19.895 4.355 20.065 4.525 ;
        RECT 20.635 3.985 20.805 4.155 ;
      LAYER met1 ;
        RECT 0.995 4.525 1.225 4.555 ;
        RECT 9.875 4.525 10.105 4.555 ;
        RECT 13.945 4.525 14.175 4.555 ;
        RECT 19.865 4.525 20.095 4.555 ;
        RECT 0.965 4.355 20.125 4.525 ;
        RECT 0.995 4.325 1.225 4.355 ;
        RECT 9.875 4.325 10.105 4.355 ;
        RECT 13.945 4.325 14.175 4.355 ;
        RECT 19.865 4.325 20.095 4.355 ;
        RECT 3.955 4.155 4.185 4.185 ;
        RECT 5.805 4.155 6.035 4.185 ;
        RECT 15.795 4.155 16.025 4.185 ;
        RECT 16.535 4.155 16.765 4.185 ;
        RECT 20.605 4.155 20.835 4.185 ;
        RECT 3.925 3.985 16.055 4.155 ;
        RECT 16.505 3.985 20.865 4.155 ;
        RECT 3.955 3.955 4.185 3.985 ;
        RECT 5.805 3.955 6.035 3.985 ;
        RECT 15.795 3.955 16.025 3.985 ;
        RECT 16.535 3.955 16.765 3.985 ;
        RECT 20.605 3.955 20.835 3.985 ;
        RECT 3.215 3.785 3.445 3.815 ;
        RECT 7.285 3.785 7.515 3.815 ;
        RECT 9.135 3.785 9.365 3.815 ;
        RECT 10.615 3.785 10.845 3.815 ;
        RECT 12.465 3.785 12.695 3.815 ;
        RECT 3.185 3.615 9.395 3.785 ;
        RECT 10.585 3.615 12.725 3.785 ;
        RECT 3.215 3.585 3.445 3.615 ;
        RECT 7.285 3.585 7.515 3.615 ;
        RECT 9.135 3.585 9.365 3.615 ;
        RECT 10.615 3.585 10.845 3.615 ;
        RECT 12.465 3.585 12.695 3.615 ;
  END
END DFFQNX1






MACRO DFFQX1
  CLASS BLOCK ;
  FOREIGN DFFQX1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 22.300 BY 7.950 ;
  PIN Q
    ANTENNAGATEAREA 1.027250 ;
    ANTENNADIFFAREA 1.351900 ;
    PORT
      LAYER li1 ;
        RECT 19.275 5.515 19.445 7.250 ;
        RECT 20.155 5.515 20.325 7.250 ;
        RECT 19.275 5.345 20.805 5.515 ;
        RECT 16.595 4.940 16.765 5.095 ;
        RECT 16.565 4.765 16.765 4.940 ;
        RECT 16.565 2.055 16.735 4.765 ;
        RECT 20.635 1.880 20.805 5.345 ;
        RECT 20.195 1.710 20.805 1.880 ;
        RECT 20.195 0.975 20.365 1.710 ;
      LAYER mcon ;
        RECT 16.565 3.985 16.735 4.155 ;
        RECT 20.635 3.985 20.805 4.155 ;
      LAYER met1 ;
        RECT 16.535 4.155 16.765 4.185 ;
        RECT 20.605 4.155 20.835 4.185 ;
        RECT 16.505 3.985 20.865 4.155 ;
        RECT 16.535 3.955 16.765 3.985 ;
        RECT 20.605 3.955 20.835 3.985 ;
    END
  END Q
  PIN D
    ANTENNAGATEAREA 1.027250 ;
    PORT
      LAYER li1 ;
        RECT 6.605 4.940 6.775 5.095 ;
        RECT 6.575 4.765 6.775 4.940 ;
        RECT 6.575 2.055 6.745 4.765 ;
      LAYER mcon ;
        RECT 6.575 3.245 6.745 3.415 ;
        RECT 6.575 2.135 6.745 2.305 ;
      LAYER met1 ;
        RECT 6.545 3.415 6.775 3.445 ;
        RECT 6.395 3.245 6.805 3.415 ;
        RECT 6.545 3.215 6.775 3.245 ;
        RECT 6.545 2.305 6.775 2.335 ;
        RECT 6.395 2.135 6.805 2.305 ;
        RECT 6.545 2.105 6.775 2.135 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 2.042100 ;
    PORT
      LAYER li1 ;
        RECT 2.135 2.055 2.305 5.095 ;
        RECT 13.265 4.975 13.435 5.095 ;
        RECT 13.235 4.765 13.435 4.975 ;
        RECT 13.235 2.055 13.405 4.765 ;
      LAYER mcon ;
        RECT 2.135 4.725 2.305 4.895 ;
        RECT 13.235 4.725 13.405 4.895 ;
      LAYER met1 ;
        RECT 2.105 4.895 2.335 4.925 ;
        RECT 13.205 4.895 13.435 4.925 ;
        RECT 2.075 4.725 13.465 4.895 ;
        RECT 2.105 4.695 2.335 4.725 ;
        RECT 13.205 4.695 13.435 4.725 ;
    END
  END CLK
  PIN VDD
    ANTENNADIFFAREA 27.348349 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 21.880 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 21.615 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 1.005 5.445 1.175 7.460 ;
        RECT 1.885 5.785 2.055 7.460 ;
        RECT 2.765 5.785 2.935 7.460 ;
        RECT 3.645 5.785 3.815 7.460 ;
        RECT 4.655 4.340 4.965 7.460 ;
        RECT 5.515 5.365 5.685 7.460 ;
        RECT 6.395 5.785 6.565 7.460 ;
        RECT 7.275 5.785 7.445 7.460 ;
        RECT 7.985 4.340 8.295 7.460 ;
        RECT 8.845 5.365 9.015 7.460 ;
        RECT 9.725 5.785 9.895 7.460 ;
        RECT 10.605 5.785 10.775 7.460 ;
        RECT 11.315 4.340 11.625 7.460 ;
        RECT 12.175 5.365 12.345 7.460 ;
        RECT 13.055 5.785 13.225 7.460 ;
        RECT 13.935 5.785 14.105 7.460 ;
        RECT 14.645 4.340 14.955 7.460 ;
        RECT 15.505 5.365 15.675 7.460 ;
        RECT 16.385 5.785 16.555 7.460 ;
        RECT 17.265 5.785 17.435 7.460 ;
        RECT 17.975 4.340 18.285 7.460 ;
        RECT 18.835 5.365 19.005 7.460 ;
        RECT 19.715 5.785 19.885 7.460 ;
        RECT 20.595 5.785 20.765 7.460 ;
        RECT 21.305 4.340 21.615 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 0.995 7.525 1.165 7.695 ;
        RECT 1.355 7.525 1.525 7.695 ;
        RECT 1.715 7.525 1.885 7.695 ;
        RECT 2.075 7.525 2.245 7.695 ;
        RECT 2.565 7.525 2.735 7.695 ;
        RECT 2.925 7.525 3.095 7.695 ;
        RECT 3.285 7.525 3.455 7.695 ;
        RECT 3.645 7.525 3.815 7.695 ;
        RECT 4.005 7.525 4.175 7.695 ;
        RECT 4.365 7.525 4.535 7.695 ;
        RECT 5.085 7.525 5.255 7.695 ;
        RECT 5.445 7.525 5.615 7.695 ;
        RECT 5.805 7.525 5.975 7.695 ;
        RECT 6.165 7.525 6.335 7.695 ;
        RECT 6.615 7.525 6.785 7.695 ;
        RECT 6.975 7.525 7.145 7.695 ;
        RECT 7.335 7.525 7.505 7.695 ;
        RECT 7.695 7.525 7.865 7.695 ;
        RECT 8.415 7.525 8.585 7.695 ;
        RECT 8.775 7.525 8.945 7.695 ;
        RECT 9.135 7.525 9.305 7.695 ;
        RECT 9.495 7.525 9.665 7.695 ;
        RECT 9.945 7.525 10.115 7.695 ;
        RECT 10.305 7.525 10.475 7.695 ;
        RECT 10.665 7.525 10.835 7.695 ;
        RECT 11.025 7.525 11.195 7.695 ;
        RECT 11.745 7.525 11.915 7.695 ;
        RECT 12.105 7.525 12.275 7.695 ;
        RECT 12.465 7.525 12.635 7.695 ;
        RECT 12.825 7.525 12.995 7.695 ;
        RECT 13.275 7.525 13.445 7.695 ;
        RECT 13.635 7.525 13.805 7.695 ;
        RECT 13.995 7.525 14.165 7.695 ;
        RECT 14.355 7.525 14.525 7.695 ;
        RECT 15.075 7.525 15.245 7.695 ;
        RECT 15.435 7.525 15.605 7.695 ;
        RECT 15.795 7.525 15.965 7.695 ;
        RECT 16.155 7.525 16.325 7.695 ;
        RECT 16.605 7.525 16.775 7.695 ;
        RECT 16.965 7.525 17.135 7.695 ;
        RECT 17.325 7.525 17.495 7.695 ;
        RECT 17.685 7.525 17.855 7.695 ;
        RECT 18.405 7.525 18.575 7.695 ;
        RECT 18.765 7.525 18.935 7.695 ;
        RECT 19.125 7.525 19.295 7.695 ;
        RECT 19.485 7.525 19.655 7.695 ;
        RECT 19.935 7.525 20.105 7.695 ;
        RECT 20.295 7.525 20.465 7.695 ;
        RECT 20.655 7.525 20.825 7.695 ;
        RECT 21.015 7.525 21.185 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 21.615 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 16.646250 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 21.745 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 4.525 -0.075 5.095 -0.065 ;
        RECT 7.855 -0.075 8.425 -0.065 ;
        RECT 11.185 -0.075 11.755 -0.065 ;
        RECT 14.515 -0.075 15.085 -0.065 ;
        RECT 17.845 -0.075 18.415 -0.065 ;
        RECT 21.175 -0.075 21.745 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 0.990 0.310 1.160 1.270 ;
        RECT 4.655 0.310 4.965 2.860 ;
        RECT 5.905 0.310 6.075 1.260 ;
        RECT 7.985 0.310 8.295 2.860 ;
        RECT 9.235 0.310 9.405 1.260 ;
        RECT 11.315 0.310 11.625 2.860 ;
        RECT 12.565 0.310 12.735 1.260 ;
        RECT 14.645 0.310 14.955 2.860 ;
        RECT 15.895 0.310 16.065 1.260 ;
        RECT 17.975 0.310 18.285 2.860 ;
        RECT 19.225 0.310 19.395 1.260 ;
        RECT 21.305 0.310 21.615 2.860 ;
        RECT -0.155 0.000 21.615 0.310 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 0.995 0.065 1.165 0.235 ;
        RECT 1.355 0.065 1.525 0.235 ;
        RECT 1.715 0.065 1.885 0.235 ;
        RECT 2.075 0.065 2.245 0.235 ;
        RECT 2.565 0.065 2.735 0.235 ;
        RECT 2.925 0.065 3.095 0.235 ;
        RECT 3.285 0.065 3.455 0.235 ;
        RECT 3.645 0.065 3.815 0.235 ;
        RECT 4.005 0.065 4.175 0.235 ;
        RECT 4.365 0.065 4.535 0.235 ;
        RECT 5.085 0.065 5.255 0.235 ;
        RECT 5.445 0.065 5.615 0.235 ;
        RECT 5.805 0.065 5.975 0.235 ;
        RECT 6.165 0.065 6.335 0.235 ;
        RECT 6.615 0.065 6.785 0.235 ;
        RECT 6.975 0.065 7.145 0.235 ;
        RECT 7.335 0.065 7.505 0.235 ;
        RECT 7.695 0.065 7.865 0.235 ;
        RECT 8.415 0.065 8.585 0.235 ;
        RECT 8.775 0.065 8.945 0.235 ;
        RECT 9.135 0.065 9.305 0.235 ;
        RECT 9.495 0.065 9.665 0.235 ;
        RECT 9.945 0.065 10.115 0.235 ;
        RECT 10.305 0.065 10.475 0.235 ;
        RECT 10.665 0.065 10.835 0.235 ;
        RECT 11.025 0.065 11.195 0.235 ;
        RECT 11.745 0.065 11.915 0.235 ;
        RECT 12.105 0.065 12.275 0.235 ;
        RECT 12.465 0.065 12.635 0.235 ;
        RECT 12.825 0.065 12.995 0.235 ;
        RECT 13.275 0.065 13.445 0.235 ;
        RECT 13.635 0.065 13.805 0.235 ;
        RECT 13.995 0.065 14.165 0.235 ;
        RECT 14.355 0.065 14.525 0.235 ;
        RECT 15.075 0.065 15.245 0.235 ;
        RECT 15.435 0.065 15.605 0.235 ;
        RECT 15.795 0.065 15.965 0.235 ;
        RECT 16.155 0.065 16.325 0.235 ;
        RECT 16.605 0.065 16.775 0.235 ;
        RECT 16.965 0.065 17.135 0.235 ;
        RECT 17.325 0.065 17.495 0.235 ;
        RECT 17.685 0.065 17.855 0.235 ;
        RECT 18.405 0.065 18.575 0.235 ;
        RECT 18.765 0.065 18.935 0.235 ;
        RECT 19.125 0.065 19.295 0.235 ;
        RECT 19.485 0.065 19.655 0.235 ;
        RECT 19.935 0.065 20.105 0.235 ;
        RECT 20.295 0.065 20.465 0.235 ;
        RECT 20.655 0.065 20.825 0.235 ;
        RECT 21.015 0.065 21.185 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 21.615 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 1.445 5.470 1.615 7.250 ;
        RECT 2.325 5.470 2.495 7.250 ;
        RECT 3.205 5.470 3.375 7.250 ;
        RECT 5.955 5.515 6.125 7.250 ;
        RECT 6.835 5.515 7.005 7.250 ;
        RECT 9.285 5.515 9.455 7.250 ;
        RECT 10.165 5.515 10.335 7.250 ;
        RECT 12.615 5.515 12.785 7.250 ;
        RECT 13.495 5.515 13.665 7.250 ;
        RECT 15.945 5.515 16.115 7.250 ;
        RECT 16.825 5.515 16.995 7.250 ;
        RECT 1.445 5.300 4.155 5.470 ;
        RECT 5.955 5.345 7.485 5.515 ;
        RECT 9.285 5.345 10.815 5.515 ;
        RECT 12.615 5.345 14.145 5.515 ;
        RECT 15.945 5.345 17.475 5.515 ;
        RECT 1.025 2.055 1.195 5.095 ;
        RECT 3.245 2.055 3.415 5.095 ;
        RECT 0.505 1.815 0.675 1.895 ;
        RECT 1.475 1.815 1.645 1.895 ;
        RECT 2.445 1.815 2.615 1.895 ;
        RECT 0.505 1.645 2.615 1.815 ;
        RECT 0.505 0.515 0.675 1.645 ;
        RECT 1.475 0.765 1.645 1.645 ;
        RECT 2.445 1.565 2.615 1.645 ;
        RECT 1.965 1.220 2.135 1.300 ;
        RECT 3.015 1.220 3.185 1.895 ;
        RECT 3.985 1.890 4.155 5.300 ;
        RECT 5.835 2.055 6.005 5.095 ;
        RECT 1.965 1.050 3.185 1.220 ;
        RECT 1.965 0.970 2.135 1.050 ;
        RECT 2.445 0.765 2.615 0.845 ;
        RECT 1.475 0.595 2.615 0.765 ;
        RECT 1.475 0.515 1.645 0.595 ;
        RECT 2.445 0.515 2.615 0.595 ;
        RECT 3.015 0.765 3.185 1.050 ;
        RECT 3.500 1.720 4.155 1.890 ;
        RECT 5.420 1.805 5.590 1.885 ;
        RECT 6.390 1.805 6.560 1.885 ;
        RECT 7.315 1.880 7.485 5.345 ;
        RECT 9.165 2.055 9.335 5.095 ;
        RECT 9.935 4.940 10.105 5.095 ;
        RECT 9.905 4.765 10.105 4.940 ;
        RECT 9.905 2.055 10.075 4.765 ;
        RECT 3.500 0.985 3.670 1.720 ;
        RECT 5.420 1.635 6.560 1.805 ;
        RECT 3.985 0.765 4.155 1.535 ;
        RECT 3.015 0.595 4.155 0.765 ;
        RECT 3.015 0.515 3.185 0.595 ;
        RECT 3.985 0.515 4.155 0.595 ;
        RECT 5.420 0.505 5.590 1.635 ;
        RECT 6.390 0.755 6.560 1.635 ;
        RECT 6.875 1.710 7.485 1.880 ;
        RECT 8.750 1.805 8.920 1.885 ;
        RECT 9.720 1.805 9.890 1.885 ;
        RECT 10.645 1.880 10.815 5.345 ;
        RECT 12.495 2.055 12.665 5.095 ;
        RECT 6.875 0.975 7.045 1.710 ;
        RECT 8.750 1.635 9.890 1.805 ;
        RECT 7.360 0.755 7.530 1.525 ;
        RECT 6.390 0.585 7.530 0.755 ;
        RECT 6.390 0.505 6.560 0.585 ;
        RECT 7.360 0.505 7.530 0.585 ;
        RECT 8.750 0.505 8.920 1.635 ;
        RECT 9.720 0.755 9.890 1.635 ;
        RECT 10.205 1.710 10.815 1.880 ;
        RECT 12.080 1.805 12.250 1.885 ;
        RECT 13.050 1.805 13.220 1.885 ;
        RECT 13.975 1.880 14.145 5.345 ;
        RECT 15.825 2.055 15.995 5.095 ;
        RECT 10.205 0.975 10.375 1.710 ;
        RECT 12.080 1.635 13.220 1.805 ;
        RECT 10.690 0.755 10.860 1.525 ;
        RECT 9.720 0.585 10.860 0.755 ;
        RECT 9.720 0.505 9.890 0.585 ;
        RECT 10.690 0.505 10.860 0.585 ;
        RECT 12.080 0.505 12.250 1.635 ;
        RECT 13.050 0.755 13.220 1.635 ;
        RECT 13.535 1.710 14.145 1.880 ;
        RECT 15.410 1.805 15.580 1.885 ;
        RECT 16.380 1.805 16.550 1.885 ;
        RECT 17.305 1.880 17.475 5.345 ;
        RECT 19.155 2.055 19.325 5.095 ;
        RECT 19.925 4.940 20.095 5.095 ;
        RECT 19.895 4.765 20.095 4.940 ;
        RECT 19.895 2.055 20.065 4.765 ;
        RECT 13.535 0.975 13.705 1.710 ;
        RECT 15.410 1.635 16.550 1.805 ;
        RECT 14.020 0.755 14.190 1.525 ;
        RECT 13.050 0.585 14.190 0.755 ;
        RECT 13.050 0.505 13.220 0.585 ;
        RECT 14.020 0.505 14.190 0.585 ;
        RECT 15.410 0.505 15.580 1.635 ;
        RECT 16.380 0.755 16.550 1.635 ;
        RECT 16.865 1.710 17.475 1.880 ;
        RECT 18.740 1.805 18.910 1.885 ;
        RECT 19.710 1.805 19.880 1.885 ;
        RECT 16.865 0.975 17.035 1.710 ;
        RECT 18.740 1.635 19.880 1.805 ;
        RECT 17.350 0.755 17.520 1.525 ;
        RECT 16.380 0.585 17.520 0.755 ;
        RECT 16.380 0.505 16.550 0.585 ;
        RECT 17.350 0.505 17.520 0.585 ;
        RECT 18.740 0.505 18.910 1.635 ;
        RECT 19.710 0.755 19.880 1.635 ;
        RECT 20.680 0.755 20.850 1.525 ;
        RECT 19.710 0.585 20.850 0.755 ;
        RECT 19.710 0.505 19.880 0.585 ;
        RECT 20.680 0.505 20.850 0.585 ;
      LAYER mcon ;
        RECT 1.025 4.355 1.195 4.525 ;
        RECT 3.245 3.615 3.415 3.785 ;
        RECT 3.985 3.985 4.155 4.155 ;
        RECT 5.835 3.985 6.005 4.155 ;
        RECT 7.315 3.615 7.485 3.785 ;
        RECT 9.165 3.615 9.335 3.785 ;
        RECT 9.905 4.355 10.075 4.525 ;
        RECT 10.645 3.615 10.815 3.785 ;
        RECT 12.495 3.615 12.665 3.785 ;
        RECT 13.975 4.355 14.145 4.525 ;
        RECT 15.825 3.985 15.995 4.155 ;
        RECT 17.305 3.615 17.475 3.785 ;
        RECT 19.155 3.615 19.325 3.785 ;
        RECT 19.895 4.355 20.065 4.525 ;
      LAYER met1 ;
        RECT 0.995 4.525 1.225 4.555 ;
        RECT 9.875 4.525 10.105 4.555 ;
        RECT 13.945 4.525 14.175 4.555 ;
        RECT 19.865 4.525 20.095 4.555 ;
        RECT 0.965 4.355 20.125 4.525 ;
        RECT 0.995 4.325 1.225 4.355 ;
        RECT 9.875 4.325 10.105 4.355 ;
        RECT 13.945 4.325 14.175 4.355 ;
        RECT 19.865 4.325 20.095 4.355 ;
        RECT 3.955 4.155 4.185 4.185 ;
        RECT 5.805 4.155 6.035 4.185 ;
        RECT 15.795 4.155 16.025 4.185 ;
        RECT 3.925 3.985 16.055 4.155 ;
        RECT 3.955 3.955 4.185 3.985 ;
        RECT 5.805 3.955 6.035 3.985 ;
        RECT 15.795 3.955 16.025 3.985 ;
        RECT 3.215 3.785 3.445 3.815 ;
        RECT 7.285 3.785 7.515 3.815 ;
        RECT 9.135 3.785 9.365 3.815 ;
        RECT 10.615 3.785 10.845 3.815 ;
        RECT 12.465 3.785 12.695 3.815 ;
        RECT 17.275 3.785 17.505 3.815 ;
        RECT 19.125 3.785 19.355 3.815 ;
        RECT 3.185 3.615 9.395 3.785 ;
        RECT 10.585 3.615 12.725 3.785 ;
        RECT 17.245 3.615 19.385 3.785 ;
        RECT 3.215 3.585 3.445 3.615 ;
        RECT 7.285 3.585 7.515 3.615 ;
        RECT 9.135 3.585 9.365 3.615 ;
        RECT 10.615 3.585 10.845 3.615 ;
        RECT 12.465 3.585 12.695 3.615 ;
        RECT 17.275 3.585 17.505 3.615 ;
        RECT 19.125 3.585 19.355 3.615 ;
  END
END DFFQX1






MACRO DFFRNQNX1
  CLASS BLOCK ;
  FOREIGN DFFRNQNX1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 26.740 BY 7.950 ;
  PIN QN
    ANTENNAGATEAREA 1.033250 ;
    ANTENNADIFFAREA 1.931900 ;
    PORT
      LAYER li1 ;
        RECT 19.205 5.470 19.375 7.250 ;
        RECT 20.085 5.470 20.255 7.250 ;
        RECT 20.965 5.470 21.135 7.250 ;
        RECT 19.205 5.300 21.915 5.470 ;
        RECT 21.745 1.890 21.915 5.300 ;
        RECT 23.595 2.055 23.765 5.095 ;
        RECT 21.260 1.720 21.915 1.890 ;
        RECT 21.260 0.985 21.430 1.720 ;
      LAYER mcon ;
        RECT 21.745 3.615 21.915 3.785 ;
        RECT 23.595 3.615 23.765 3.785 ;
      LAYER met1 ;
        RECT 21.715 3.785 21.945 3.815 ;
        RECT 23.565 3.785 23.795 3.815 ;
        RECT 21.685 3.615 23.825 3.785 ;
        RECT 21.715 3.585 21.945 3.615 ;
        RECT 23.565 3.585 23.795 3.615 ;
    END
  END QN
  PIN D
    ANTENNAGATEAREA 1.014850 ;
    PORT
      LAYER li1 ;
        RECT 6.945 2.055 7.115 5.095 ;
      LAYER mcon ;
        RECT 6.945 3.245 7.115 3.415 ;
      LAYER met1 ;
        RECT 6.915 3.415 7.145 3.445 ;
        RECT 6.765 3.245 7.175 3.415 ;
        RECT 6.915 3.215 7.145 3.245 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 2.029700 ;
    PORT
      LAYER li1 ;
        RECT 2.135 2.055 2.305 5.095 ;
        RECT 15.085 2.055 15.255 5.095 ;
      LAYER mcon ;
        RECT 2.135 4.725 2.305 4.895 ;
        RECT 15.085 4.725 15.255 4.895 ;
      LAYER met1 ;
        RECT 2.105 4.895 2.335 4.925 ;
        RECT 15.055 4.895 15.285 4.925 ;
        RECT 2.075 4.725 15.315 4.895 ;
        RECT 2.105 4.695 2.335 4.725 ;
        RECT 15.055 4.695 15.285 4.725 ;
    END
  END CLK
  PIN RN
    ANTENNAGATEAREA 3.069350 ;
    PORT
      LAYER li1 ;
        RECT 8.055 2.055 8.225 5.095 ;
        RECT 16.195 2.055 16.365 5.095 ;
        RECT 19.895 2.055 20.065 5.095 ;
      LAYER mcon ;
        RECT 8.055 2.505 8.225 2.675 ;
        RECT 16.195 2.505 16.365 2.675 ;
        RECT 19.895 2.505 20.065 2.675 ;
      LAYER met1 ;
        RECT 8.025 2.675 8.255 2.705 ;
        RECT 16.165 2.675 16.395 2.705 ;
        RECT 19.865 2.675 20.095 2.705 ;
        RECT 7.995 2.505 20.125 2.675 ;
        RECT 8.025 2.475 8.255 2.505 ;
        RECT 16.165 2.475 16.395 2.505 ;
        RECT 19.865 2.475 20.095 2.505 ;
    END
  END RN
  PIN VDD
    ANTENNADIFFAREA 31.219549 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 26.320 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 26.055 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 1.005 5.445 1.175 7.460 ;
        RECT 1.885 5.785 2.055 7.460 ;
        RECT 2.765 5.785 2.935 7.460 ;
        RECT 3.645 5.785 3.815 7.460 ;
        RECT 4.655 4.340 4.965 7.460 ;
        RECT 5.815 5.445 5.985 7.460 ;
        RECT 6.695 5.785 6.865 7.460 ;
        RECT 7.575 5.785 7.745 7.460 ;
        RECT 8.455 5.785 8.625 7.460 ;
        RECT 9.465 4.340 9.775 7.460 ;
        RECT 10.325 5.365 10.495 7.460 ;
        RECT 11.205 5.785 11.375 7.460 ;
        RECT 12.085 5.785 12.255 7.460 ;
        RECT 12.795 4.340 13.105 7.460 ;
        RECT 13.955 5.445 14.125 7.460 ;
        RECT 14.835 5.785 15.005 7.460 ;
        RECT 15.715 5.785 15.885 7.460 ;
        RECT 16.595 5.785 16.765 7.460 ;
        RECT 17.605 4.340 17.915 7.460 ;
        RECT 18.765 5.445 18.935 7.460 ;
        RECT 19.645 5.785 19.815 7.460 ;
        RECT 20.525 5.785 20.695 7.460 ;
        RECT 21.405 5.785 21.575 7.460 ;
        RECT 22.415 4.340 22.725 7.460 ;
        RECT 23.275 5.365 23.445 7.460 ;
        RECT 24.155 5.785 24.325 7.460 ;
        RECT 25.035 5.785 25.205 7.460 ;
        RECT 25.745 4.340 26.055 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 0.995 7.525 1.165 7.695 ;
        RECT 1.355 7.525 1.525 7.695 ;
        RECT 1.715 7.525 1.885 7.695 ;
        RECT 2.075 7.525 2.245 7.695 ;
        RECT 2.565 7.525 2.735 7.695 ;
        RECT 2.925 7.525 3.095 7.695 ;
        RECT 3.285 7.525 3.455 7.695 ;
        RECT 3.645 7.525 3.815 7.695 ;
        RECT 4.005 7.525 4.175 7.695 ;
        RECT 4.365 7.525 4.535 7.695 ;
        RECT 5.085 7.525 5.255 7.695 ;
        RECT 5.445 7.525 5.615 7.695 ;
        RECT 5.805 7.525 5.975 7.695 ;
        RECT 6.165 7.525 6.335 7.695 ;
        RECT 6.525 7.525 6.695 7.695 ;
        RECT 6.885 7.525 7.055 7.695 ;
        RECT 7.375 7.525 7.545 7.695 ;
        RECT 7.735 7.525 7.905 7.695 ;
        RECT 8.095 7.525 8.265 7.695 ;
        RECT 8.455 7.525 8.625 7.695 ;
        RECT 8.815 7.525 8.985 7.695 ;
        RECT 9.175 7.525 9.345 7.695 ;
        RECT 9.895 7.525 10.065 7.695 ;
        RECT 10.255 7.525 10.425 7.695 ;
        RECT 10.615 7.525 10.785 7.695 ;
        RECT 10.975 7.525 11.145 7.695 ;
        RECT 11.425 7.525 11.595 7.695 ;
        RECT 11.785 7.525 11.955 7.695 ;
        RECT 12.145 7.525 12.315 7.695 ;
        RECT 12.505 7.525 12.675 7.695 ;
        RECT 13.225 7.525 13.395 7.695 ;
        RECT 13.585 7.525 13.755 7.695 ;
        RECT 13.945 7.525 14.115 7.695 ;
        RECT 14.305 7.525 14.475 7.695 ;
        RECT 14.665 7.525 14.835 7.695 ;
        RECT 15.025 7.525 15.195 7.695 ;
        RECT 15.515 7.525 15.685 7.695 ;
        RECT 15.875 7.525 16.045 7.695 ;
        RECT 16.235 7.525 16.405 7.695 ;
        RECT 16.595 7.525 16.765 7.695 ;
        RECT 16.955 7.525 17.125 7.695 ;
        RECT 17.315 7.525 17.485 7.695 ;
        RECT 18.035 7.525 18.205 7.695 ;
        RECT 18.395 7.525 18.565 7.695 ;
        RECT 18.755 7.525 18.925 7.695 ;
        RECT 19.115 7.525 19.285 7.695 ;
        RECT 19.475 7.525 19.645 7.695 ;
        RECT 19.835 7.525 20.005 7.695 ;
        RECT 20.325 7.525 20.495 7.695 ;
        RECT 20.685 7.525 20.855 7.695 ;
        RECT 21.045 7.525 21.215 7.695 ;
        RECT 21.405 7.525 21.575 7.695 ;
        RECT 21.765 7.525 21.935 7.695 ;
        RECT 22.125 7.525 22.295 7.695 ;
        RECT 22.845 7.525 23.015 7.695 ;
        RECT 23.205 7.525 23.375 7.695 ;
        RECT 23.565 7.525 23.735 7.695 ;
        RECT 23.925 7.525 24.095 7.695 ;
        RECT 24.375 7.525 24.545 7.695 ;
        RECT 24.735 7.525 24.905 7.695 ;
        RECT 25.095 7.525 25.265 7.695 ;
        RECT 25.455 7.525 25.625 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 26.055 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 18.777449 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 26.185 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 4.525 -0.075 5.095 -0.065 ;
        RECT 9.335 -0.075 9.905 -0.065 ;
        RECT 12.665 -0.075 13.235 -0.065 ;
        RECT 17.475 -0.075 18.045 -0.065 ;
        RECT 22.285 -0.075 22.855 -0.065 ;
        RECT 25.615 -0.075 26.185 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 0.990 0.310 1.160 1.270 ;
        RECT 4.655 0.310 4.965 2.860 ;
        RECT 5.800 0.310 5.970 1.270 ;
        RECT 9.465 0.310 9.775 2.860 ;
        RECT 10.715 0.310 10.885 1.260 ;
        RECT 12.795 0.310 13.105 2.860 ;
        RECT 13.940 0.310 14.110 1.270 ;
        RECT 17.605 0.310 17.915 2.860 ;
        RECT 18.750 0.310 18.920 1.270 ;
        RECT 22.415 0.310 22.725 2.860 ;
        RECT 23.665 0.310 23.835 1.260 ;
        RECT 25.745 0.310 26.055 2.860 ;
        RECT -0.155 0.000 26.055 0.310 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 0.995 0.065 1.165 0.235 ;
        RECT 1.355 0.065 1.525 0.235 ;
        RECT 1.715 0.065 1.885 0.235 ;
        RECT 2.075 0.065 2.245 0.235 ;
        RECT 2.565 0.065 2.735 0.235 ;
        RECT 2.925 0.065 3.095 0.235 ;
        RECT 3.285 0.065 3.455 0.235 ;
        RECT 3.645 0.065 3.815 0.235 ;
        RECT 4.005 0.065 4.175 0.235 ;
        RECT 4.365 0.065 4.535 0.235 ;
        RECT 5.085 0.065 5.255 0.235 ;
        RECT 5.445 0.065 5.615 0.235 ;
        RECT 5.805 0.065 5.975 0.235 ;
        RECT 6.165 0.065 6.335 0.235 ;
        RECT 6.525 0.065 6.695 0.235 ;
        RECT 6.885 0.065 7.055 0.235 ;
        RECT 7.375 0.065 7.545 0.235 ;
        RECT 7.735 0.065 7.905 0.235 ;
        RECT 8.095 0.065 8.265 0.235 ;
        RECT 8.455 0.065 8.625 0.235 ;
        RECT 8.815 0.065 8.985 0.235 ;
        RECT 9.175 0.065 9.345 0.235 ;
        RECT 9.895 0.065 10.065 0.235 ;
        RECT 10.255 0.065 10.425 0.235 ;
        RECT 10.615 0.065 10.785 0.235 ;
        RECT 10.975 0.065 11.145 0.235 ;
        RECT 11.425 0.065 11.595 0.235 ;
        RECT 11.785 0.065 11.955 0.235 ;
        RECT 12.145 0.065 12.315 0.235 ;
        RECT 12.505 0.065 12.675 0.235 ;
        RECT 13.225 0.065 13.395 0.235 ;
        RECT 13.585 0.065 13.755 0.235 ;
        RECT 13.945 0.065 14.115 0.235 ;
        RECT 14.305 0.065 14.475 0.235 ;
        RECT 14.665 0.065 14.835 0.235 ;
        RECT 15.025 0.065 15.195 0.235 ;
        RECT 15.515 0.065 15.685 0.235 ;
        RECT 15.875 0.065 16.045 0.235 ;
        RECT 16.235 0.065 16.405 0.235 ;
        RECT 16.595 0.065 16.765 0.235 ;
        RECT 16.955 0.065 17.125 0.235 ;
        RECT 17.315 0.065 17.485 0.235 ;
        RECT 18.035 0.065 18.205 0.235 ;
        RECT 18.395 0.065 18.565 0.235 ;
        RECT 18.755 0.065 18.925 0.235 ;
        RECT 19.115 0.065 19.285 0.235 ;
        RECT 19.475 0.065 19.645 0.235 ;
        RECT 19.835 0.065 20.005 0.235 ;
        RECT 20.325 0.065 20.495 0.235 ;
        RECT 20.685 0.065 20.855 0.235 ;
        RECT 21.045 0.065 21.215 0.235 ;
        RECT 21.405 0.065 21.575 0.235 ;
        RECT 21.765 0.065 21.935 0.235 ;
        RECT 22.125 0.065 22.295 0.235 ;
        RECT 22.845 0.065 23.015 0.235 ;
        RECT 23.205 0.065 23.375 0.235 ;
        RECT 23.565 0.065 23.735 0.235 ;
        RECT 23.925 0.065 24.095 0.235 ;
        RECT 24.375 0.065 24.545 0.235 ;
        RECT 24.735 0.065 24.905 0.235 ;
        RECT 25.095 0.065 25.265 0.235 ;
        RECT 25.455 0.065 25.625 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 26.055 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 1.445 5.470 1.615 7.250 ;
        RECT 2.325 5.470 2.495 7.250 ;
        RECT 3.205 5.470 3.375 7.250 ;
        RECT 6.255 5.470 6.425 7.250 ;
        RECT 7.135 5.470 7.305 7.250 ;
        RECT 8.015 5.470 8.185 7.250 ;
        RECT 10.765 5.515 10.935 7.250 ;
        RECT 11.645 5.515 11.815 7.250 ;
        RECT 1.445 5.300 4.155 5.470 ;
        RECT 6.255 5.300 8.965 5.470 ;
        RECT 10.765 5.345 12.295 5.515 ;
        RECT 1.025 2.055 1.195 5.095 ;
        RECT 3.245 2.055 3.415 5.095 ;
        RECT 0.505 1.815 0.675 1.895 ;
        RECT 1.475 1.815 1.645 1.895 ;
        RECT 2.445 1.815 2.615 1.895 ;
        RECT 0.505 1.645 2.615 1.815 ;
        RECT 0.505 0.515 0.675 1.645 ;
        RECT 1.475 0.765 1.645 1.645 ;
        RECT 2.445 1.565 2.615 1.645 ;
        RECT 1.965 1.220 2.135 1.300 ;
        RECT 3.015 1.220 3.185 1.895 ;
        RECT 3.985 1.890 4.155 5.300 ;
        RECT 5.835 2.055 6.005 5.095 ;
        RECT 1.965 1.050 3.185 1.220 ;
        RECT 1.965 0.970 2.135 1.050 ;
        RECT 2.445 0.765 2.615 0.845 ;
        RECT 1.475 0.595 2.615 0.765 ;
        RECT 1.475 0.515 1.645 0.595 ;
        RECT 2.445 0.515 2.615 0.595 ;
        RECT 3.015 0.765 3.185 1.050 ;
        RECT 3.500 1.720 4.155 1.890 ;
        RECT 5.315 1.815 5.485 1.895 ;
        RECT 6.285 1.815 6.455 1.895 ;
        RECT 7.255 1.815 7.425 1.895 ;
        RECT 3.500 0.985 3.670 1.720 ;
        RECT 5.315 1.645 7.425 1.815 ;
        RECT 3.985 0.765 4.155 1.535 ;
        RECT 3.015 0.595 4.155 0.765 ;
        RECT 3.015 0.515 3.185 0.595 ;
        RECT 3.985 0.515 4.155 0.595 ;
        RECT 5.315 0.515 5.485 1.645 ;
        RECT 6.285 0.765 6.455 1.645 ;
        RECT 7.255 1.565 7.425 1.645 ;
        RECT 6.775 1.220 6.945 1.300 ;
        RECT 7.825 1.220 7.995 1.895 ;
        RECT 8.795 1.890 8.965 5.300 ;
        RECT 10.645 2.055 10.815 5.095 ;
        RECT 11.415 4.940 11.585 5.095 ;
        RECT 11.385 4.765 11.585 4.940 ;
        RECT 11.385 2.055 11.555 4.765 ;
        RECT 6.775 1.050 7.995 1.220 ;
        RECT 6.775 0.970 6.945 1.050 ;
        RECT 7.255 0.765 7.425 0.845 ;
        RECT 6.285 0.595 7.425 0.765 ;
        RECT 6.285 0.515 6.455 0.595 ;
        RECT 7.255 0.515 7.425 0.595 ;
        RECT 7.825 0.765 7.995 1.050 ;
        RECT 8.310 1.720 8.965 1.890 ;
        RECT 10.230 1.805 10.400 1.885 ;
        RECT 11.200 1.805 11.370 1.885 ;
        RECT 12.125 1.880 12.295 5.345 ;
        RECT 14.395 5.470 14.565 7.250 ;
        RECT 15.275 5.470 15.445 7.250 ;
        RECT 16.155 5.470 16.325 7.250 ;
        RECT 23.715 5.515 23.885 7.250 ;
        RECT 24.595 5.515 24.765 7.250 ;
        RECT 14.395 5.300 17.105 5.470 ;
        RECT 23.715 5.345 25.245 5.515 ;
        RECT 13.975 2.055 14.145 5.095 ;
        RECT 8.310 0.985 8.480 1.720 ;
        RECT 10.230 1.635 11.370 1.805 ;
        RECT 8.795 0.765 8.965 1.535 ;
        RECT 7.825 0.595 8.965 0.765 ;
        RECT 7.825 0.515 7.995 0.595 ;
        RECT 8.795 0.515 8.965 0.595 ;
        RECT 10.230 0.505 10.400 1.635 ;
        RECT 11.200 0.755 11.370 1.635 ;
        RECT 11.685 1.710 12.295 1.880 ;
        RECT 13.455 1.815 13.625 1.895 ;
        RECT 14.425 1.815 14.595 1.895 ;
        RECT 15.395 1.815 15.565 1.895 ;
        RECT 11.685 0.975 11.855 1.710 ;
        RECT 13.455 1.645 15.565 1.815 ;
        RECT 12.170 0.755 12.340 1.525 ;
        RECT 11.200 0.585 12.340 0.755 ;
        RECT 11.200 0.505 11.370 0.585 ;
        RECT 12.170 0.505 12.340 0.585 ;
        RECT 13.455 0.515 13.625 1.645 ;
        RECT 14.425 0.765 14.595 1.645 ;
        RECT 15.395 1.565 15.565 1.645 ;
        RECT 14.915 1.220 15.085 1.300 ;
        RECT 15.965 1.220 16.135 1.895 ;
        RECT 16.935 1.890 17.105 5.300 ;
        RECT 18.785 2.055 18.955 5.095 ;
        RECT 21.005 2.055 21.175 5.095 ;
        RECT 24.365 4.940 24.535 5.095 ;
        RECT 24.335 4.765 24.535 4.940 ;
        RECT 24.335 2.055 24.505 4.765 ;
        RECT 14.915 1.050 16.135 1.220 ;
        RECT 14.915 0.970 15.085 1.050 ;
        RECT 15.395 0.765 15.565 0.845 ;
        RECT 14.425 0.595 15.565 0.765 ;
        RECT 14.425 0.515 14.595 0.595 ;
        RECT 15.395 0.515 15.565 0.595 ;
        RECT 15.965 0.765 16.135 1.050 ;
        RECT 16.450 1.720 17.105 1.890 ;
        RECT 18.265 1.815 18.435 1.895 ;
        RECT 19.235 1.815 19.405 1.895 ;
        RECT 20.205 1.815 20.375 1.895 ;
        RECT 16.450 0.985 16.620 1.720 ;
        RECT 18.265 1.645 20.375 1.815 ;
        RECT 16.935 0.765 17.105 1.535 ;
        RECT 15.965 0.595 17.105 0.765 ;
        RECT 15.965 0.515 16.135 0.595 ;
        RECT 16.935 0.515 17.105 0.595 ;
        RECT 18.265 0.515 18.435 1.645 ;
        RECT 19.235 0.765 19.405 1.645 ;
        RECT 20.205 1.565 20.375 1.645 ;
        RECT 19.725 1.220 19.895 1.300 ;
        RECT 20.775 1.220 20.945 1.895 ;
        RECT 23.180 1.805 23.350 1.885 ;
        RECT 24.150 1.805 24.320 1.885 ;
        RECT 25.075 1.880 25.245 5.345 ;
        RECT 23.180 1.635 24.320 1.805 ;
        RECT 19.725 1.050 20.945 1.220 ;
        RECT 19.725 0.970 19.895 1.050 ;
        RECT 20.205 0.765 20.375 0.845 ;
        RECT 19.235 0.595 20.375 0.765 ;
        RECT 19.235 0.515 19.405 0.595 ;
        RECT 20.205 0.515 20.375 0.595 ;
        RECT 20.775 0.765 20.945 1.050 ;
        RECT 21.745 0.765 21.915 1.535 ;
        RECT 20.775 0.595 21.915 0.765 ;
        RECT 20.775 0.515 20.945 0.595 ;
        RECT 21.745 0.515 21.915 0.595 ;
        RECT 23.180 0.505 23.350 1.635 ;
        RECT 24.150 0.755 24.320 1.635 ;
        RECT 24.635 1.710 25.245 1.880 ;
        RECT 24.635 0.975 24.805 1.710 ;
        RECT 25.120 0.755 25.290 1.525 ;
        RECT 24.150 0.585 25.290 0.755 ;
        RECT 24.150 0.505 24.320 0.585 ;
        RECT 25.120 0.505 25.290 0.585 ;
      LAYER mcon ;
        RECT 1.025 4.355 1.195 4.525 ;
        RECT 3.245 3.615 3.415 3.785 ;
        RECT 3.985 3.985 4.155 4.155 ;
        RECT 5.835 3.985 6.005 4.155 ;
        RECT 8.795 3.615 8.965 3.785 ;
        RECT 10.645 3.615 10.815 3.785 ;
        RECT 11.385 4.355 11.555 4.525 ;
        RECT 12.125 3.615 12.295 3.785 ;
        RECT 13.975 3.615 14.145 3.785 ;
        RECT 16.935 4.355 17.105 4.525 ;
        RECT 18.785 3.985 18.955 4.155 ;
        RECT 21.005 3.985 21.175 4.155 ;
        RECT 24.335 4.355 24.505 4.525 ;
        RECT 25.075 3.985 25.245 4.155 ;
      LAYER met1 ;
        RECT 0.995 4.525 1.225 4.555 ;
        RECT 11.355 4.525 11.585 4.555 ;
        RECT 16.905 4.525 17.135 4.555 ;
        RECT 24.305 4.525 24.535 4.555 ;
        RECT 0.965 4.355 24.565 4.525 ;
        RECT 0.995 4.325 1.225 4.355 ;
        RECT 11.355 4.325 11.585 4.355 ;
        RECT 16.905 4.325 17.135 4.355 ;
        RECT 24.305 4.325 24.535 4.355 ;
        RECT 3.955 4.155 4.185 4.185 ;
        RECT 5.805 4.155 6.035 4.185 ;
        RECT 18.755 4.155 18.985 4.185 ;
        RECT 20.975 4.155 21.205 4.185 ;
        RECT 25.045 4.155 25.275 4.185 ;
        RECT 3.925 3.985 19.015 4.155 ;
        RECT 20.945 3.985 25.305 4.155 ;
        RECT 3.955 3.955 4.185 3.985 ;
        RECT 5.805 3.955 6.035 3.985 ;
        RECT 18.755 3.955 18.985 3.985 ;
        RECT 20.975 3.955 21.205 3.985 ;
        RECT 25.045 3.955 25.275 3.985 ;
        RECT 3.215 3.785 3.445 3.815 ;
        RECT 8.765 3.785 8.995 3.815 ;
        RECT 10.615 3.785 10.845 3.815 ;
        RECT 12.095 3.785 12.325 3.815 ;
        RECT 13.945 3.785 14.175 3.815 ;
        RECT 3.185 3.615 10.875 3.785 ;
        RECT 12.065 3.615 14.205 3.785 ;
        RECT 3.215 3.585 3.445 3.615 ;
        RECT 8.765 3.585 8.995 3.615 ;
        RECT 10.615 3.585 10.845 3.615 ;
        RECT 12.095 3.585 12.325 3.615 ;
        RECT 13.945 3.585 14.175 3.615 ;
  END
END DFFRNQNX1






MACRO DFFRNQX1
  CLASS BLOCK ;
  FOREIGN DFFRNQX1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 26.740 BY 7.950 ;
  PIN Q
    ANTENNAGATEAREA 1.027250 ;
    ANTENNADIFFAREA 1.351900 ;
    PORT
      LAYER li1 ;
        RECT 23.715 5.515 23.885 7.250 ;
        RECT 24.595 5.515 24.765 7.250 ;
        RECT 23.715 5.345 25.245 5.515 ;
        RECT 21.005 2.055 21.175 5.095 ;
        RECT 25.075 1.880 25.245 5.345 ;
        RECT 24.635 1.710 25.245 1.880 ;
        RECT 24.635 0.975 24.805 1.710 ;
      LAYER mcon ;
        RECT 21.005 3.985 21.175 4.155 ;
        RECT 25.075 3.985 25.245 4.155 ;
      LAYER met1 ;
        RECT 20.975 4.155 21.205 4.185 ;
        RECT 25.045 4.155 25.275 4.185 ;
        RECT 20.945 3.985 25.305 4.155 ;
        RECT 20.975 3.955 21.205 3.985 ;
        RECT 25.045 3.955 25.275 3.985 ;
    END
  END Q
  PIN D
    ANTENNAGATEAREA 1.014850 ;
    PORT
      LAYER li1 ;
        RECT 6.945 2.055 7.115 5.095 ;
      LAYER mcon ;
        RECT 6.945 3.245 7.115 3.415 ;
      LAYER met1 ;
        RECT 6.915 3.415 7.145 3.445 ;
        RECT 6.765 3.245 7.175 3.415 ;
        RECT 6.915 3.215 7.145 3.245 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 2.029700 ;
    PORT
      LAYER li1 ;
        RECT 2.135 2.055 2.305 5.095 ;
        RECT 15.085 2.055 15.255 5.095 ;
      LAYER mcon ;
        RECT 2.135 4.725 2.305 4.895 ;
        RECT 15.085 4.725 15.255 4.895 ;
      LAYER met1 ;
        RECT 2.105 4.895 2.335 4.925 ;
        RECT 15.055 4.895 15.285 4.925 ;
        RECT 2.075 4.725 15.315 4.895 ;
        RECT 2.105 4.695 2.335 4.725 ;
        RECT 15.055 4.695 15.285 4.725 ;
    END
  END CLK
  PIN RN
    ANTENNAGATEAREA 3.069350 ;
    PORT
      LAYER li1 ;
        RECT 8.055 2.055 8.225 5.095 ;
        RECT 16.195 2.055 16.365 5.095 ;
        RECT 19.895 2.055 20.065 5.095 ;
      LAYER mcon ;
        RECT 8.055 2.505 8.225 2.675 ;
        RECT 16.195 2.505 16.365 2.675 ;
        RECT 19.895 2.505 20.065 2.675 ;
      LAYER met1 ;
        RECT 8.025 2.675 8.255 2.705 ;
        RECT 16.165 2.675 16.395 2.705 ;
        RECT 19.865 2.675 20.095 2.705 ;
        RECT 7.995 2.505 20.125 2.675 ;
        RECT 8.025 2.475 8.255 2.505 ;
        RECT 16.165 2.475 16.395 2.505 ;
        RECT 19.865 2.475 20.095 2.505 ;
    END
  END RN
  PIN VDD
    ANTENNADIFFAREA 31.219549 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 26.320 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 26.055 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 1.005 5.445 1.175 7.460 ;
        RECT 1.885 5.785 2.055 7.460 ;
        RECT 2.765 5.785 2.935 7.460 ;
        RECT 3.645 5.785 3.815 7.460 ;
        RECT 4.655 4.340 4.965 7.460 ;
        RECT 5.815 5.445 5.985 7.460 ;
        RECT 6.695 5.785 6.865 7.460 ;
        RECT 7.575 5.785 7.745 7.460 ;
        RECT 8.455 5.785 8.625 7.460 ;
        RECT 9.465 4.340 9.775 7.460 ;
        RECT 10.325 5.365 10.495 7.460 ;
        RECT 11.205 5.785 11.375 7.460 ;
        RECT 12.085 5.785 12.255 7.460 ;
        RECT 12.795 4.340 13.105 7.460 ;
        RECT 13.955 5.445 14.125 7.460 ;
        RECT 14.835 5.785 15.005 7.460 ;
        RECT 15.715 5.785 15.885 7.460 ;
        RECT 16.595 5.785 16.765 7.460 ;
        RECT 17.605 4.340 17.915 7.460 ;
        RECT 18.765 5.445 18.935 7.460 ;
        RECT 19.645 5.785 19.815 7.460 ;
        RECT 20.525 5.785 20.695 7.460 ;
        RECT 21.405 5.785 21.575 7.460 ;
        RECT 22.415 4.340 22.725 7.460 ;
        RECT 23.275 5.365 23.445 7.460 ;
        RECT 24.155 5.785 24.325 7.460 ;
        RECT 25.035 5.785 25.205 7.460 ;
        RECT 25.745 4.340 26.055 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 0.995 7.525 1.165 7.695 ;
        RECT 1.355 7.525 1.525 7.695 ;
        RECT 1.715 7.525 1.885 7.695 ;
        RECT 2.075 7.525 2.245 7.695 ;
        RECT 2.565 7.525 2.735 7.695 ;
        RECT 2.925 7.525 3.095 7.695 ;
        RECT 3.285 7.525 3.455 7.695 ;
        RECT 3.645 7.525 3.815 7.695 ;
        RECT 4.005 7.525 4.175 7.695 ;
        RECT 4.365 7.525 4.535 7.695 ;
        RECT 5.085 7.525 5.255 7.695 ;
        RECT 5.445 7.525 5.615 7.695 ;
        RECT 5.805 7.525 5.975 7.695 ;
        RECT 6.165 7.525 6.335 7.695 ;
        RECT 6.525 7.525 6.695 7.695 ;
        RECT 6.885 7.525 7.055 7.695 ;
        RECT 7.375 7.525 7.545 7.695 ;
        RECT 7.735 7.525 7.905 7.695 ;
        RECT 8.095 7.525 8.265 7.695 ;
        RECT 8.455 7.525 8.625 7.695 ;
        RECT 8.815 7.525 8.985 7.695 ;
        RECT 9.175 7.525 9.345 7.695 ;
        RECT 9.895 7.525 10.065 7.695 ;
        RECT 10.255 7.525 10.425 7.695 ;
        RECT 10.615 7.525 10.785 7.695 ;
        RECT 10.975 7.525 11.145 7.695 ;
        RECT 11.425 7.525 11.595 7.695 ;
        RECT 11.785 7.525 11.955 7.695 ;
        RECT 12.145 7.525 12.315 7.695 ;
        RECT 12.505 7.525 12.675 7.695 ;
        RECT 13.225 7.525 13.395 7.695 ;
        RECT 13.585 7.525 13.755 7.695 ;
        RECT 13.945 7.525 14.115 7.695 ;
        RECT 14.305 7.525 14.475 7.695 ;
        RECT 14.665 7.525 14.835 7.695 ;
        RECT 15.025 7.525 15.195 7.695 ;
        RECT 15.515 7.525 15.685 7.695 ;
        RECT 15.875 7.525 16.045 7.695 ;
        RECT 16.235 7.525 16.405 7.695 ;
        RECT 16.595 7.525 16.765 7.695 ;
        RECT 16.955 7.525 17.125 7.695 ;
        RECT 17.315 7.525 17.485 7.695 ;
        RECT 18.035 7.525 18.205 7.695 ;
        RECT 18.395 7.525 18.565 7.695 ;
        RECT 18.755 7.525 18.925 7.695 ;
        RECT 19.115 7.525 19.285 7.695 ;
        RECT 19.475 7.525 19.645 7.695 ;
        RECT 19.835 7.525 20.005 7.695 ;
        RECT 20.325 7.525 20.495 7.695 ;
        RECT 20.685 7.525 20.855 7.695 ;
        RECT 21.045 7.525 21.215 7.695 ;
        RECT 21.405 7.525 21.575 7.695 ;
        RECT 21.765 7.525 21.935 7.695 ;
        RECT 22.125 7.525 22.295 7.695 ;
        RECT 22.845 7.525 23.015 7.695 ;
        RECT 23.205 7.525 23.375 7.695 ;
        RECT 23.565 7.525 23.735 7.695 ;
        RECT 23.925 7.525 24.095 7.695 ;
        RECT 24.375 7.525 24.545 7.695 ;
        RECT 24.735 7.525 24.905 7.695 ;
        RECT 25.095 7.525 25.265 7.695 ;
        RECT 25.455 7.525 25.625 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 26.055 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 18.777449 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 26.185 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 4.525 -0.075 5.095 -0.065 ;
        RECT 9.335 -0.075 9.905 -0.065 ;
        RECT 12.665 -0.075 13.235 -0.065 ;
        RECT 17.475 -0.075 18.045 -0.065 ;
        RECT 22.285 -0.075 22.855 -0.065 ;
        RECT 25.615 -0.075 26.185 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 0.990 0.310 1.160 1.270 ;
        RECT 4.655 0.310 4.965 2.860 ;
        RECT 5.800 0.310 5.970 1.270 ;
        RECT 9.465 0.310 9.775 2.860 ;
        RECT 10.715 0.310 10.885 1.260 ;
        RECT 12.795 0.310 13.105 2.860 ;
        RECT 13.940 0.310 14.110 1.270 ;
        RECT 17.605 0.310 17.915 2.860 ;
        RECT 18.750 0.310 18.920 1.270 ;
        RECT 22.415 0.310 22.725 2.860 ;
        RECT 23.665 0.310 23.835 1.260 ;
        RECT 25.745 0.310 26.055 2.860 ;
        RECT -0.155 0.000 26.055 0.310 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 0.995 0.065 1.165 0.235 ;
        RECT 1.355 0.065 1.525 0.235 ;
        RECT 1.715 0.065 1.885 0.235 ;
        RECT 2.075 0.065 2.245 0.235 ;
        RECT 2.565 0.065 2.735 0.235 ;
        RECT 2.925 0.065 3.095 0.235 ;
        RECT 3.285 0.065 3.455 0.235 ;
        RECT 3.645 0.065 3.815 0.235 ;
        RECT 4.005 0.065 4.175 0.235 ;
        RECT 4.365 0.065 4.535 0.235 ;
        RECT 5.085 0.065 5.255 0.235 ;
        RECT 5.445 0.065 5.615 0.235 ;
        RECT 5.805 0.065 5.975 0.235 ;
        RECT 6.165 0.065 6.335 0.235 ;
        RECT 6.525 0.065 6.695 0.235 ;
        RECT 6.885 0.065 7.055 0.235 ;
        RECT 7.375 0.065 7.545 0.235 ;
        RECT 7.735 0.065 7.905 0.235 ;
        RECT 8.095 0.065 8.265 0.235 ;
        RECT 8.455 0.065 8.625 0.235 ;
        RECT 8.815 0.065 8.985 0.235 ;
        RECT 9.175 0.065 9.345 0.235 ;
        RECT 9.895 0.065 10.065 0.235 ;
        RECT 10.255 0.065 10.425 0.235 ;
        RECT 10.615 0.065 10.785 0.235 ;
        RECT 10.975 0.065 11.145 0.235 ;
        RECT 11.425 0.065 11.595 0.235 ;
        RECT 11.785 0.065 11.955 0.235 ;
        RECT 12.145 0.065 12.315 0.235 ;
        RECT 12.505 0.065 12.675 0.235 ;
        RECT 13.225 0.065 13.395 0.235 ;
        RECT 13.585 0.065 13.755 0.235 ;
        RECT 13.945 0.065 14.115 0.235 ;
        RECT 14.305 0.065 14.475 0.235 ;
        RECT 14.665 0.065 14.835 0.235 ;
        RECT 15.025 0.065 15.195 0.235 ;
        RECT 15.515 0.065 15.685 0.235 ;
        RECT 15.875 0.065 16.045 0.235 ;
        RECT 16.235 0.065 16.405 0.235 ;
        RECT 16.595 0.065 16.765 0.235 ;
        RECT 16.955 0.065 17.125 0.235 ;
        RECT 17.315 0.065 17.485 0.235 ;
        RECT 18.035 0.065 18.205 0.235 ;
        RECT 18.395 0.065 18.565 0.235 ;
        RECT 18.755 0.065 18.925 0.235 ;
        RECT 19.115 0.065 19.285 0.235 ;
        RECT 19.475 0.065 19.645 0.235 ;
        RECT 19.835 0.065 20.005 0.235 ;
        RECT 20.325 0.065 20.495 0.235 ;
        RECT 20.685 0.065 20.855 0.235 ;
        RECT 21.045 0.065 21.215 0.235 ;
        RECT 21.405 0.065 21.575 0.235 ;
        RECT 21.765 0.065 21.935 0.235 ;
        RECT 22.125 0.065 22.295 0.235 ;
        RECT 22.845 0.065 23.015 0.235 ;
        RECT 23.205 0.065 23.375 0.235 ;
        RECT 23.565 0.065 23.735 0.235 ;
        RECT 23.925 0.065 24.095 0.235 ;
        RECT 24.375 0.065 24.545 0.235 ;
        RECT 24.735 0.065 24.905 0.235 ;
        RECT 25.095 0.065 25.265 0.235 ;
        RECT 25.455 0.065 25.625 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 26.055 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 1.445 5.470 1.615 7.250 ;
        RECT 2.325 5.470 2.495 7.250 ;
        RECT 3.205 5.470 3.375 7.250 ;
        RECT 6.255 5.470 6.425 7.250 ;
        RECT 7.135 5.470 7.305 7.250 ;
        RECT 8.015 5.470 8.185 7.250 ;
        RECT 10.765 5.515 10.935 7.250 ;
        RECT 11.645 5.515 11.815 7.250 ;
        RECT 1.445 5.300 4.155 5.470 ;
        RECT 6.255 5.300 8.965 5.470 ;
        RECT 10.765 5.345 12.295 5.515 ;
        RECT 1.025 2.055 1.195 5.095 ;
        RECT 3.245 2.055 3.415 5.095 ;
        RECT 0.505 1.815 0.675 1.895 ;
        RECT 1.475 1.815 1.645 1.895 ;
        RECT 2.445 1.815 2.615 1.895 ;
        RECT 0.505 1.645 2.615 1.815 ;
        RECT 0.505 0.515 0.675 1.645 ;
        RECT 1.475 0.765 1.645 1.645 ;
        RECT 2.445 1.565 2.615 1.645 ;
        RECT 1.965 1.220 2.135 1.300 ;
        RECT 3.015 1.220 3.185 1.895 ;
        RECT 3.985 1.890 4.155 5.300 ;
        RECT 5.835 2.055 6.005 5.095 ;
        RECT 1.965 1.050 3.185 1.220 ;
        RECT 1.965 0.970 2.135 1.050 ;
        RECT 2.445 0.765 2.615 0.845 ;
        RECT 1.475 0.595 2.615 0.765 ;
        RECT 1.475 0.515 1.645 0.595 ;
        RECT 2.445 0.515 2.615 0.595 ;
        RECT 3.015 0.765 3.185 1.050 ;
        RECT 3.500 1.720 4.155 1.890 ;
        RECT 5.315 1.815 5.485 1.895 ;
        RECT 6.285 1.815 6.455 1.895 ;
        RECT 7.255 1.815 7.425 1.895 ;
        RECT 3.500 0.985 3.670 1.720 ;
        RECT 5.315 1.645 7.425 1.815 ;
        RECT 3.985 0.765 4.155 1.535 ;
        RECT 3.015 0.595 4.155 0.765 ;
        RECT 3.015 0.515 3.185 0.595 ;
        RECT 3.985 0.515 4.155 0.595 ;
        RECT 5.315 0.515 5.485 1.645 ;
        RECT 6.285 0.765 6.455 1.645 ;
        RECT 7.255 1.565 7.425 1.645 ;
        RECT 6.775 1.220 6.945 1.300 ;
        RECT 7.825 1.220 7.995 1.895 ;
        RECT 8.795 1.890 8.965 5.300 ;
        RECT 10.645 2.055 10.815 5.095 ;
        RECT 11.415 4.940 11.585 5.095 ;
        RECT 11.385 4.765 11.585 4.940 ;
        RECT 11.385 2.055 11.555 4.765 ;
        RECT 6.775 1.050 7.995 1.220 ;
        RECT 6.775 0.970 6.945 1.050 ;
        RECT 7.255 0.765 7.425 0.845 ;
        RECT 6.285 0.595 7.425 0.765 ;
        RECT 6.285 0.515 6.455 0.595 ;
        RECT 7.255 0.515 7.425 0.595 ;
        RECT 7.825 0.765 7.995 1.050 ;
        RECT 8.310 1.720 8.965 1.890 ;
        RECT 10.230 1.805 10.400 1.885 ;
        RECT 11.200 1.805 11.370 1.885 ;
        RECT 12.125 1.880 12.295 5.345 ;
        RECT 14.395 5.470 14.565 7.250 ;
        RECT 15.275 5.470 15.445 7.250 ;
        RECT 16.155 5.470 16.325 7.250 ;
        RECT 19.205 5.470 19.375 7.250 ;
        RECT 20.085 5.470 20.255 7.250 ;
        RECT 20.965 5.470 21.135 7.250 ;
        RECT 14.395 5.300 17.105 5.470 ;
        RECT 19.205 5.300 21.915 5.470 ;
        RECT 13.975 2.055 14.145 5.095 ;
        RECT 8.310 0.985 8.480 1.720 ;
        RECT 10.230 1.635 11.370 1.805 ;
        RECT 8.795 0.765 8.965 1.535 ;
        RECT 7.825 0.595 8.965 0.765 ;
        RECT 7.825 0.515 7.995 0.595 ;
        RECT 8.795 0.515 8.965 0.595 ;
        RECT 10.230 0.505 10.400 1.635 ;
        RECT 11.200 0.755 11.370 1.635 ;
        RECT 11.685 1.710 12.295 1.880 ;
        RECT 13.455 1.815 13.625 1.895 ;
        RECT 14.425 1.815 14.595 1.895 ;
        RECT 15.395 1.815 15.565 1.895 ;
        RECT 11.685 0.975 11.855 1.710 ;
        RECT 13.455 1.645 15.565 1.815 ;
        RECT 12.170 0.755 12.340 1.525 ;
        RECT 11.200 0.585 12.340 0.755 ;
        RECT 11.200 0.505 11.370 0.585 ;
        RECT 12.170 0.505 12.340 0.585 ;
        RECT 13.455 0.515 13.625 1.645 ;
        RECT 14.425 0.765 14.595 1.645 ;
        RECT 15.395 1.565 15.565 1.645 ;
        RECT 14.915 1.220 15.085 1.300 ;
        RECT 15.965 1.220 16.135 1.895 ;
        RECT 16.935 1.890 17.105 5.300 ;
        RECT 18.785 2.055 18.955 5.095 ;
        RECT 14.915 1.050 16.135 1.220 ;
        RECT 14.915 0.970 15.085 1.050 ;
        RECT 15.395 0.765 15.565 0.845 ;
        RECT 14.425 0.595 15.565 0.765 ;
        RECT 14.425 0.515 14.595 0.595 ;
        RECT 15.395 0.515 15.565 0.595 ;
        RECT 15.965 0.765 16.135 1.050 ;
        RECT 16.450 1.720 17.105 1.890 ;
        RECT 18.265 1.815 18.435 1.895 ;
        RECT 19.235 1.815 19.405 1.895 ;
        RECT 20.205 1.815 20.375 1.895 ;
        RECT 16.450 0.985 16.620 1.720 ;
        RECT 18.265 1.645 20.375 1.815 ;
        RECT 16.935 0.765 17.105 1.535 ;
        RECT 15.965 0.595 17.105 0.765 ;
        RECT 15.965 0.515 16.135 0.595 ;
        RECT 16.935 0.515 17.105 0.595 ;
        RECT 18.265 0.515 18.435 1.645 ;
        RECT 19.235 0.765 19.405 1.645 ;
        RECT 20.205 1.565 20.375 1.645 ;
        RECT 19.725 1.220 19.895 1.300 ;
        RECT 20.775 1.220 20.945 1.895 ;
        RECT 21.745 1.890 21.915 5.300 ;
        RECT 23.595 2.055 23.765 5.095 ;
        RECT 24.365 4.940 24.535 5.095 ;
        RECT 24.335 4.765 24.535 4.940 ;
        RECT 24.335 2.055 24.505 4.765 ;
        RECT 19.725 1.050 20.945 1.220 ;
        RECT 19.725 0.970 19.895 1.050 ;
        RECT 20.205 0.765 20.375 0.845 ;
        RECT 19.235 0.595 20.375 0.765 ;
        RECT 19.235 0.515 19.405 0.595 ;
        RECT 20.205 0.515 20.375 0.595 ;
        RECT 20.775 0.765 20.945 1.050 ;
        RECT 21.260 1.720 21.915 1.890 ;
        RECT 23.180 1.805 23.350 1.885 ;
        RECT 24.150 1.805 24.320 1.885 ;
        RECT 21.260 0.985 21.430 1.720 ;
        RECT 23.180 1.635 24.320 1.805 ;
        RECT 21.745 0.765 21.915 1.535 ;
        RECT 20.775 0.595 21.915 0.765 ;
        RECT 20.775 0.515 20.945 0.595 ;
        RECT 21.745 0.515 21.915 0.595 ;
        RECT 23.180 0.505 23.350 1.635 ;
        RECT 24.150 0.755 24.320 1.635 ;
        RECT 25.120 0.755 25.290 1.525 ;
        RECT 24.150 0.585 25.290 0.755 ;
        RECT 24.150 0.505 24.320 0.585 ;
        RECT 25.120 0.505 25.290 0.585 ;
      LAYER mcon ;
        RECT 1.025 4.355 1.195 4.525 ;
        RECT 3.245 3.615 3.415 3.785 ;
        RECT 3.985 3.985 4.155 4.155 ;
        RECT 5.835 3.985 6.005 4.155 ;
        RECT 8.795 3.615 8.965 3.785 ;
        RECT 10.645 3.615 10.815 3.785 ;
        RECT 11.385 4.355 11.555 4.525 ;
        RECT 12.125 3.615 12.295 3.785 ;
        RECT 13.975 3.615 14.145 3.785 ;
        RECT 16.935 4.355 17.105 4.525 ;
        RECT 18.785 3.985 18.955 4.155 ;
        RECT 21.745 3.615 21.915 3.785 ;
        RECT 23.595 3.615 23.765 3.785 ;
        RECT 24.335 4.355 24.505 4.525 ;
      LAYER met1 ;
        RECT 0.995 4.525 1.225 4.555 ;
        RECT 11.355 4.525 11.585 4.555 ;
        RECT 16.905 4.525 17.135 4.555 ;
        RECT 24.305 4.525 24.535 4.555 ;
        RECT 0.965 4.355 24.565 4.525 ;
        RECT 0.995 4.325 1.225 4.355 ;
        RECT 11.355 4.325 11.585 4.355 ;
        RECT 16.905 4.325 17.135 4.355 ;
        RECT 24.305 4.325 24.535 4.355 ;
        RECT 3.955 4.155 4.185 4.185 ;
        RECT 5.805 4.155 6.035 4.185 ;
        RECT 18.755 4.155 18.985 4.185 ;
        RECT 3.925 3.985 19.015 4.155 ;
        RECT 3.955 3.955 4.185 3.985 ;
        RECT 5.805 3.955 6.035 3.985 ;
        RECT 18.755 3.955 18.985 3.985 ;
        RECT 3.215 3.785 3.445 3.815 ;
        RECT 8.765 3.785 8.995 3.815 ;
        RECT 10.615 3.785 10.845 3.815 ;
        RECT 12.095 3.785 12.325 3.815 ;
        RECT 13.945 3.785 14.175 3.815 ;
        RECT 21.715 3.785 21.945 3.815 ;
        RECT 23.565 3.785 23.795 3.815 ;
        RECT 3.185 3.615 10.875 3.785 ;
        RECT 12.065 3.615 14.205 3.785 ;
        RECT 21.685 3.615 23.825 3.785 ;
        RECT 3.215 3.585 3.445 3.615 ;
        RECT 8.765 3.585 8.995 3.615 ;
        RECT 10.615 3.585 10.845 3.615 ;
        RECT 12.095 3.585 12.325 3.615 ;
        RECT 13.945 3.585 14.175 3.615 ;
        RECT 21.715 3.585 21.945 3.615 ;
        RECT 23.565 3.585 23.795 3.615 ;
  END
END DFFRNQX1






MACRO DFFRNX1
  CLASS BLOCK ;
  FOREIGN DFFRNX1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 26.740 BY 7.950 ;
  PIN Q
    ANTENNAGATEAREA 1.027250 ;
    ANTENNADIFFAREA 1.351900 ;
    PORT
      LAYER li1 ;
        RECT 23.715 5.515 23.885 7.250 ;
        RECT 24.595 5.515 24.765 7.250 ;
        RECT 23.715 5.345 25.245 5.515 ;
        RECT 21.005 2.055 21.175 5.095 ;
        RECT 25.075 1.880 25.245 5.345 ;
        RECT 24.635 1.710 25.245 1.880 ;
        RECT 24.635 0.975 24.805 1.710 ;
      LAYER mcon ;
        RECT 21.005 3.985 21.175 4.155 ;
        RECT 25.075 3.985 25.245 4.155 ;
      LAYER met1 ;
        RECT 20.975 4.155 21.205 4.185 ;
        RECT 25.045 4.155 25.275 4.185 ;
        RECT 20.945 3.985 25.305 4.155 ;
        RECT 20.975 3.955 21.205 3.985 ;
        RECT 25.045 3.955 25.275 3.985 ;
    END
  END Q
  PIN QN
    ANTENNAGATEAREA 1.033250 ;
    ANTENNADIFFAREA 1.931900 ;
    PORT
      LAYER li1 ;
        RECT 19.205 5.470 19.375 7.250 ;
        RECT 20.085 5.470 20.255 7.250 ;
        RECT 20.965 5.470 21.135 7.250 ;
        RECT 19.205 5.300 21.915 5.470 ;
        RECT 21.745 1.890 21.915 5.300 ;
        RECT 23.595 2.055 23.765 5.095 ;
        RECT 21.260 1.720 21.915 1.890 ;
        RECT 21.260 0.985 21.430 1.720 ;
      LAYER mcon ;
        RECT 21.745 3.615 21.915 3.785 ;
        RECT 23.595 3.615 23.765 3.785 ;
      LAYER met1 ;
        RECT 21.715 3.785 21.945 3.815 ;
        RECT 23.565 3.785 23.795 3.815 ;
        RECT 21.685 3.615 23.825 3.785 ;
        RECT 21.715 3.585 21.945 3.615 ;
        RECT 23.565 3.585 23.795 3.615 ;
    END
  END QN
  PIN D
    ANTENNAGATEAREA 1.014850 ;
    PORT
      LAYER li1 ;
        RECT 6.945 2.055 7.115 5.095 ;
      LAYER mcon ;
        RECT 6.945 3.245 7.115 3.415 ;
      LAYER met1 ;
        RECT 6.915 3.415 7.145 3.445 ;
        RECT 6.765 3.245 7.175 3.415 ;
        RECT 6.915 3.215 7.145 3.245 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 2.029700 ;
    PORT
      LAYER li1 ;
        RECT 2.135 2.055 2.305 5.095 ;
        RECT 15.085 2.055 15.255 5.095 ;
      LAYER mcon ;
        RECT 2.135 4.725 2.305 4.895 ;
        RECT 15.085 4.725 15.255 4.895 ;
      LAYER met1 ;
        RECT 2.105 4.895 2.335 4.925 ;
        RECT 15.055 4.895 15.285 4.925 ;
        RECT 2.075 4.725 15.315 4.895 ;
        RECT 2.105 4.695 2.335 4.725 ;
        RECT 15.055 4.695 15.285 4.725 ;
    END
  END CLK
  PIN RN
    ANTENNAGATEAREA 3.069350 ;
    PORT
      LAYER li1 ;
        RECT 8.055 2.055 8.225 5.095 ;
        RECT 16.195 2.055 16.365 5.095 ;
        RECT 19.895 2.055 20.065 5.095 ;
      LAYER mcon ;
        RECT 8.055 2.505 8.225 2.675 ;
        RECT 16.195 2.505 16.365 2.675 ;
        RECT 19.895 2.505 20.065 2.675 ;
      LAYER met1 ;
        RECT 8.025 2.675 8.255 2.705 ;
        RECT 16.165 2.675 16.395 2.705 ;
        RECT 19.865 2.675 20.095 2.705 ;
        RECT 7.995 2.505 20.125 2.675 ;
        RECT 8.025 2.475 8.255 2.505 ;
        RECT 16.165 2.475 16.395 2.505 ;
        RECT 19.865 2.475 20.095 2.505 ;
    END
  END RN
  PIN VDD
    ANTENNADIFFAREA 31.219549 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 26.320 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 26.055 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 1.005 5.445 1.175 7.460 ;
        RECT 1.885 5.785 2.055 7.460 ;
        RECT 2.765 5.785 2.935 7.460 ;
        RECT 3.645 5.785 3.815 7.460 ;
        RECT 4.655 4.340 4.965 7.460 ;
        RECT 5.815 5.445 5.985 7.460 ;
        RECT 6.695 5.785 6.865 7.460 ;
        RECT 7.575 5.785 7.745 7.460 ;
        RECT 8.455 5.785 8.625 7.460 ;
        RECT 9.465 4.340 9.775 7.460 ;
        RECT 10.325 5.365 10.495 7.460 ;
        RECT 11.205 5.785 11.375 7.460 ;
        RECT 12.085 5.785 12.255 7.460 ;
        RECT 12.795 4.340 13.105 7.460 ;
        RECT 13.955 5.445 14.125 7.460 ;
        RECT 14.835 5.785 15.005 7.460 ;
        RECT 15.715 5.785 15.885 7.460 ;
        RECT 16.595 5.785 16.765 7.460 ;
        RECT 17.605 4.340 17.915 7.460 ;
        RECT 18.765 5.445 18.935 7.460 ;
        RECT 19.645 5.785 19.815 7.460 ;
        RECT 20.525 5.785 20.695 7.460 ;
        RECT 21.405 5.785 21.575 7.460 ;
        RECT 22.415 4.340 22.725 7.460 ;
        RECT 23.275 5.365 23.445 7.460 ;
        RECT 24.155 5.785 24.325 7.460 ;
        RECT 25.035 5.785 25.205 7.460 ;
        RECT 25.745 4.340 26.055 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 0.995 7.525 1.165 7.695 ;
        RECT 1.355 7.525 1.525 7.695 ;
        RECT 1.715 7.525 1.885 7.695 ;
        RECT 2.075 7.525 2.245 7.695 ;
        RECT 2.565 7.525 2.735 7.695 ;
        RECT 2.925 7.525 3.095 7.695 ;
        RECT 3.285 7.525 3.455 7.695 ;
        RECT 3.645 7.525 3.815 7.695 ;
        RECT 4.005 7.525 4.175 7.695 ;
        RECT 4.365 7.525 4.535 7.695 ;
        RECT 5.085 7.525 5.255 7.695 ;
        RECT 5.445 7.525 5.615 7.695 ;
        RECT 5.805 7.525 5.975 7.695 ;
        RECT 6.165 7.525 6.335 7.695 ;
        RECT 6.525 7.525 6.695 7.695 ;
        RECT 6.885 7.525 7.055 7.695 ;
        RECT 7.375 7.525 7.545 7.695 ;
        RECT 7.735 7.525 7.905 7.695 ;
        RECT 8.095 7.525 8.265 7.695 ;
        RECT 8.455 7.525 8.625 7.695 ;
        RECT 8.815 7.525 8.985 7.695 ;
        RECT 9.175 7.525 9.345 7.695 ;
        RECT 9.895 7.525 10.065 7.695 ;
        RECT 10.255 7.525 10.425 7.695 ;
        RECT 10.615 7.525 10.785 7.695 ;
        RECT 10.975 7.525 11.145 7.695 ;
        RECT 11.425 7.525 11.595 7.695 ;
        RECT 11.785 7.525 11.955 7.695 ;
        RECT 12.145 7.525 12.315 7.695 ;
        RECT 12.505 7.525 12.675 7.695 ;
        RECT 13.225 7.525 13.395 7.695 ;
        RECT 13.585 7.525 13.755 7.695 ;
        RECT 13.945 7.525 14.115 7.695 ;
        RECT 14.305 7.525 14.475 7.695 ;
        RECT 14.665 7.525 14.835 7.695 ;
        RECT 15.025 7.525 15.195 7.695 ;
        RECT 15.515 7.525 15.685 7.695 ;
        RECT 15.875 7.525 16.045 7.695 ;
        RECT 16.235 7.525 16.405 7.695 ;
        RECT 16.595 7.525 16.765 7.695 ;
        RECT 16.955 7.525 17.125 7.695 ;
        RECT 17.315 7.525 17.485 7.695 ;
        RECT 18.035 7.525 18.205 7.695 ;
        RECT 18.395 7.525 18.565 7.695 ;
        RECT 18.755 7.525 18.925 7.695 ;
        RECT 19.115 7.525 19.285 7.695 ;
        RECT 19.475 7.525 19.645 7.695 ;
        RECT 19.835 7.525 20.005 7.695 ;
        RECT 20.325 7.525 20.495 7.695 ;
        RECT 20.685 7.525 20.855 7.695 ;
        RECT 21.045 7.525 21.215 7.695 ;
        RECT 21.405 7.525 21.575 7.695 ;
        RECT 21.765 7.525 21.935 7.695 ;
        RECT 22.125 7.525 22.295 7.695 ;
        RECT 22.845 7.525 23.015 7.695 ;
        RECT 23.205 7.525 23.375 7.695 ;
        RECT 23.565 7.525 23.735 7.695 ;
        RECT 23.925 7.525 24.095 7.695 ;
        RECT 24.375 7.525 24.545 7.695 ;
        RECT 24.735 7.525 24.905 7.695 ;
        RECT 25.095 7.525 25.265 7.695 ;
        RECT 25.455 7.525 25.625 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 26.055 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 18.777449 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 26.185 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 4.525 -0.075 5.095 -0.065 ;
        RECT 9.335 -0.075 9.905 -0.065 ;
        RECT 12.665 -0.075 13.235 -0.065 ;
        RECT 17.475 -0.075 18.045 -0.065 ;
        RECT 22.285 -0.075 22.855 -0.065 ;
        RECT 25.615 -0.075 26.185 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 0.990 0.310 1.160 1.270 ;
        RECT 4.655 0.310 4.965 2.860 ;
        RECT 5.800 0.310 5.970 1.270 ;
        RECT 9.465 0.310 9.775 2.860 ;
        RECT 10.715 0.310 10.885 1.260 ;
        RECT 12.795 0.310 13.105 2.860 ;
        RECT 13.940 0.310 14.110 1.270 ;
        RECT 17.605 0.310 17.915 2.860 ;
        RECT 18.750 0.310 18.920 1.270 ;
        RECT 22.415 0.310 22.725 2.860 ;
        RECT 23.665 0.310 23.835 1.260 ;
        RECT 25.745 0.310 26.055 2.860 ;
        RECT -0.155 0.000 26.055 0.310 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 0.995 0.065 1.165 0.235 ;
        RECT 1.355 0.065 1.525 0.235 ;
        RECT 1.715 0.065 1.885 0.235 ;
        RECT 2.075 0.065 2.245 0.235 ;
        RECT 2.565 0.065 2.735 0.235 ;
        RECT 2.925 0.065 3.095 0.235 ;
        RECT 3.285 0.065 3.455 0.235 ;
        RECT 3.645 0.065 3.815 0.235 ;
        RECT 4.005 0.065 4.175 0.235 ;
        RECT 4.365 0.065 4.535 0.235 ;
        RECT 5.085 0.065 5.255 0.235 ;
        RECT 5.445 0.065 5.615 0.235 ;
        RECT 5.805 0.065 5.975 0.235 ;
        RECT 6.165 0.065 6.335 0.235 ;
        RECT 6.525 0.065 6.695 0.235 ;
        RECT 6.885 0.065 7.055 0.235 ;
        RECT 7.375 0.065 7.545 0.235 ;
        RECT 7.735 0.065 7.905 0.235 ;
        RECT 8.095 0.065 8.265 0.235 ;
        RECT 8.455 0.065 8.625 0.235 ;
        RECT 8.815 0.065 8.985 0.235 ;
        RECT 9.175 0.065 9.345 0.235 ;
        RECT 9.895 0.065 10.065 0.235 ;
        RECT 10.255 0.065 10.425 0.235 ;
        RECT 10.615 0.065 10.785 0.235 ;
        RECT 10.975 0.065 11.145 0.235 ;
        RECT 11.425 0.065 11.595 0.235 ;
        RECT 11.785 0.065 11.955 0.235 ;
        RECT 12.145 0.065 12.315 0.235 ;
        RECT 12.505 0.065 12.675 0.235 ;
        RECT 13.225 0.065 13.395 0.235 ;
        RECT 13.585 0.065 13.755 0.235 ;
        RECT 13.945 0.065 14.115 0.235 ;
        RECT 14.305 0.065 14.475 0.235 ;
        RECT 14.665 0.065 14.835 0.235 ;
        RECT 15.025 0.065 15.195 0.235 ;
        RECT 15.515 0.065 15.685 0.235 ;
        RECT 15.875 0.065 16.045 0.235 ;
        RECT 16.235 0.065 16.405 0.235 ;
        RECT 16.595 0.065 16.765 0.235 ;
        RECT 16.955 0.065 17.125 0.235 ;
        RECT 17.315 0.065 17.485 0.235 ;
        RECT 18.035 0.065 18.205 0.235 ;
        RECT 18.395 0.065 18.565 0.235 ;
        RECT 18.755 0.065 18.925 0.235 ;
        RECT 19.115 0.065 19.285 0.235 ;
        RECT 19.475 0.065 19.645 0.235 ;
        RECT 19.835 0.065 20.005 0.235 ;
        RECT 20.325 0.065 20.495 0.235 ;
        RECT 20.685 0.065 20.855 0.235 ;
        RECT 21.045 0.065 21.215 0.235 ;
        RECT 21.405 0.065 21.575 0.235 ;
        RECT 21.765 0.065 21.935 0.235 ;
        RECT 22.125 0.065 22.295 0.235 ;
        RECT 22.845 0.065 23.015 0.235 ;
        RECT 23.205 0.065 23.375 0.235 ;
        RECT 23.565 0.065 23.735 0.235 ;
        RECT 23.925 0.065 24.095 0.235 ;
        RECT 24.375 0.065 24.545 0.235 ;
        RECT 24.735 0.065 24.905 0.235 ;
        RECT 25.095 0.065 25.265 0.235 ;
        RECT 25.455 0.065 25.625 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 26.055 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 1.445 5.470 1.615 7.250 ;
        RECT 2.325 5.470 2.495 7.250 ;
        RECT 3.205 5.470 3.375 7.250 ;
        RECT 6.255 5.470 6.425 7.250 ;
        RECT 7.135 5.470 7.305 7.250 ;
        RECT 8.015 5.470 8.185 7.250 ;
        RECT 10.765 5.515 10.935 7.250 ;
        RECT 11.645 5.515 11.815 7.250 ;
        RECT 1.445 5.300 4.155 5.470 ;
        RECT 6.255 5.300 8.965 5.470 ;
        RECT 10.765 5.345 12.295 5.515 ;
        RECT 1.025 2.055 1.195 5.095 ;
        RECT 3.245 2.055 3.415 5.095 ;
        RECT 0.505 1.815 0.675 1.895 ;
        RECT 1.475 1.815 1.645 1.895 ;
        RECT 2.445 1.815 2.615 1.895 ;
        RECT 0.505 1.645 2.615 1.815 ;
        RECT 0.505 0.515 0.675 1.645 ;
        RECT 1.475 0.765 1.645 1.645 ;
        RECT 2.445 1.565 2.615 1.645 ;
        RECT 1.965 1.220 2.135 1.300 ;
        RECT 3.015 1.220 3.185 1.895 ;
        RECT 3.985 1.890 4.155 5.300 ;
        RECT 5.835 2.055 6.005 5.095 ;
        RECT 1.965 1.050 3.185 1.220 ;
        RECT 1.965 0.970 2.135 1.050 ;
        RECT 2.445 0.765 2.615 0.845 ;
        RECT 1.475 0.595 2.615 0.765 ;
        RECT 1.475 0.515 1.645 0.595 ;
        RECT 2.445 0.515 2.615 0.595 ;
        RECT 3.015 0.765 3.185 1.050 ;
        RECT 3.500 1.720 4.155 1.890 ;
        RECT 5.315 1.815 5.485 1.895 ;
        RECT 6.285 1.815 6.455 1.895 ;
        RECT 7.255 1.815 7.425 1.895 ;
        RECT 3.500 0.985 3.670 1.720 ;
        RECT 5.315 1.645 7.425 1.815 ;
        RECT 3.985 0.765 4.155 1.535 ;
        RECT 3.015 0.595 4.155 0.765 ;
        RECT 3.015 0.515 3.185 0.595 ;
        RECT 3.985 0.515 4.155 0.595 ;
        RECT 5.315 0.515 5.485 1.645 ;
        RECT 6.285 0.765 6.455 1.645 ;
        RECT 7.255 1.565 7.425 1.645 ;
        RECT 6.775 1.220 6.945 1.300 ;
        RECT 7.825 1.220 7.995 1.895 ;
        RECT 8.795 1.890 8.965 5.300 ;
        RECT 10.645 2.055 10.815 5.095 ;
        RECT 11.415 4.940 11.585 5.095 ;
        RECT 11.385 4.765 11.585 4.940 ;
        RECT 11.385 2.055 11.555 4.765 ;
        RECT 6.775 1.050 7.995 1.220 ;
        RECT 6.775 0.970 6.945 1.050 ;
        RECT 7.255 0.765 7.425 0.845 ;
        RECT 6.285 0.595 7.425 0.765 ;
        RECT 6.285 0.515 6.455 0.595 ;
        RECT 7.255 0.515 7.425 0.595 ;
        RECT 7.825 0.765 7.995 1.050 ;
        RECT 8.310 1.720 8.965 1.890 ;
        RECT 10.230 1.805 10.400 1.885 ;
        RECT 11.200 1.805 11.370 1.885 ;
        RECT 12.125 1.880 12.295 5.345 ;
        RECT 14.395 5.470 14.565 7.250 ;
        RECT 15.275 5.470 15.445 7.250 ;
        RECT 16.155 5.470 16.325 7.250 ;
        RECT 14.395 5.300 17.105 5.470 ;
        RECT 13.975 2.055 14.145 5.095 ;
        RECT 8.310 0.985 8.480 1.720 ;
        RECT 10.230 1.635 11.370 1.805 ;
        RECT 8.795 0.765 8.965 1.535 ;
        RECT 7.825 0.595 8.965 0.765 ;
        RECT 7.825 0.515 7.995 0.595 ;
        RECT 8.795 0.515 8.965 0.595 ;
        RECT 10.230 0.505 10.400 1.635 ;
        RECT 11.200 0.755 11.370 1.635 ;
        RECT 11.685 1.710 12.295 1.880 ;
        RECT 13.455 1.815 13.625 1.895 ;
        RECT 14.425 1.815 14.595 1.895 ;
        RECT 15.395 1.815 15.565 1.895 ;
        RECT 11.685 0.975 11.855 1.710 ;
        RECT 13.455 1.645 15.565 1.815 ;
        RECT 12.170 0.755 12.340 1.525 ;
        RECT 11.200 0.585 12.340 0.755 ;
        RECT 11.200 0.505 11.370 0.585 ;
        RECT 12.170 0.505 12.340 0.585 ;
        RECT 13.455 0.515 13.625 1.645 ;
        RECT 14.425 0.765 14.595 1.645 ;
        RECT 15.395 1.565 15.565 1.645 ;
        RECT 14.915 1.220 15.085 1.300 ;
        RECT 15.965 1.220 16.135 1.895 ;
        RECT 16.935 1.890 17.105 5.300 ;
        RECT 18.785 2.055 18.955 5.095 ;
        RECT 24.365 4.940 24.535 5.095 ;
        RECT 24.335 4.765 24.535 4.940 ;
        RECT 24.335 2.055 24.505 4.765 ;
        RECT 14.915 1.050 16.135 1.220 ;
        RECT 14.915 0.970 15.085 1.050 ;
        RECT 15.395 0.765 15.565 0.845 ;
        RECT 14.425 0.595 15.565 0.765 ;
        RECT 14.425 0.515 14.595 0.595 ;
        RECT 15.395 0.515 15.565 0.595 ;
        RECT 15.965 0.765 16.135 1.050 ;
        RECT 16.450 1.720 17.105 1.890 ;
        RECT 18.265 1.815 18.435 1.895 ;
        RECT 19.235 1.815 19.405 1.895 ;
        RECT 20.205 1.815 20.375 1.895 ;
        RECT 16.450 0.985 16.620 1.720 ;
        RECT 18.265 1.645 20.375 1.815 ;
        RECT 16.935 0.765 17.105 1.535 ;
        RECT 15.965 0.595 17.105 0.765 ;
        RECT 15.965 0.515 16.135 0.595 ;
        RECT 16.935 0.515 17.105 0.595 ;
        RECT 18.265 0.515 18.435 1.645 ;
        RECT 19.235 0.765 19.405 1.645 ;
        RECT 20.205 1.565 20.375 1.645 ;
        RECT 19.725 1.220 19.895 1.300 ;
        RECT 20.775 1.220 20.945 1.895 ;
        RECT 23.180 1.805 23.350 1.885 ;
        RECT 24.150 1.805 24.320 1.885 ;
        RECT 23.180 1.635 24.320 1.805 ;
        RECT 19.725 1.050 20.945 1.220 ;
        RECT 19.725 0.970 19.895 1.050 ;
        RECT 20.205 0.765 20.375 0.845 ;
        RECT 19.235 0.595 20.375 0.765 ;
        RECT 19.235 0.515 19.405 0.595 ;
        RECT 20.205 0.515 20.375 0.595 ;
        RECT 20.775 0.765 20.945 1.050 ;
        RECT 21.745 0.765 21.915 1.535 ;
        RECT 20.775 0.595 21.915 0.765 ;
        RECT 20.775 0.515 20.945 0.595 ;
        RECT 21.745 0.515 21.915 0.595 ;
        RECT 23.180 0.505 23.350 1.635 ;
        RECT 24.150 0.755 24.320 1.635 ;
        RECT 25.120 0.755 25.290 1.525 ;
        RECT 24.150 0.585 25.290 0.755 ;
        RECT 24.150 0.505 24.320 0.585 ;
        RECT 25.120 0.505 25.290 0.585 ;
      LAYER mcon ;
        RECT 1.025 4.355 1.195 4.525 ;
        RECT 3.245 3.615 3.415 3.785 ;
        RECT 3.985 3.985 4.155 4.155 ;
        RECT 5.835 3.985 6.005 4.155 ;
        RECT 8.795 3.615 8.965 3.785 ;
        RECT 10.645 3.615 10.815 3.785 ;
        RECT 11.385 4.355 11.555 4.525 ;
        RECT 12.125 3.615 12.295 3.785 ;
        RECT 13.975 3.615 14.145 3.785 ;
        RECT 16.935 4.355 17.105 4.525 ;
        RECT 18.785 3.985 18.955 4.155 ;
        RECT 24.335 4.355 24.505 4.525 ;
      LAYER met1 ;
        RECT 0.995 4.525 1.225 4.555 ;
        RECT 11.355 4.525 11.585 4.555 ;
        RECT 16.905 4.525 17.135 4.555 ;
        RECT 24.305 4.525 24.535 4.555 ;
        RECT 0.965 4.355 24.565 4.525 ;
        RECT 0.995 4.325 1.225 4.355 ;
        RECT 11.355 4.325 11.585 4.355 ;
        RECT 16.905 4.325 17.135 4.355 ;
        RECT 24.305 4.325 24.535 4.355 ;
        RECT 3.955 4.155 4.185 4.185 ;
        RECT 5.805 4.155 6.035 4.185 ;
        RECT 18.755 4.155 18.985 4.185 ;
        RECT 3.925 3.985 19.015 4.155 ;
        RECT 3.955 3.955 4.185 3.985 ;
        RECT 5.805 3.955 6.035 3.985 ;
        RECT 18.755 3.955 18.985 3.985 ;
        RECT 3.215 3.785 3.445 3.815 ;
        RECT 8.765 3.785 8.995 3.815 ;
        RECT 10.615 3.785 10.845 3.815 ;
        RECT 12.095 3.785 12.325 3.815 ;
        RECT 13.945 3.785 14.175 3.815 ;
        RECT 3.185 3.615 10.875 3.785 ;
        RECT 12.065 3.615 14.205 3.785 ;
        RECT 3.215 3.585 3.445 3.615 ;
        RECT 8.765 3.585 8.995 3.615 ;
        RECT 10.615 3.585 10.845 3.615 ;
        RECT 12.095 3.585 12.325 3.615 ;
        RECT 13.945 3.585 14.175 3.615 ;
  END
END DFFRNX1






MACRO DFFSNQNX1
  CLASS BLOCK ;
  FOREIGN DFFSNQNX1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 25.260 BY 7.950 ;
  PIN QN
    ANTENNAGATEAREA 1.033250 ;
    ANTENNADIFFAREA 1.351900 ;
    PORT
      LAYER li1 ;
        RECT 17.425 5.515 17.595 7.250 ;
        RECT 18.305 5.515 18.475 7.250 ;
        RECT 17.425 5.345 18.955 5.515 ;
        RECT 18.785 1.880 18.955 5.345 ;
        RECT 20.635 2.055 20.805 5.095 ;
        RECT 18.345 1.710 18.955 1.880 ;
        RECT 18.345 0.975 18.515 1.710 ;
      LAYER mcon ;
        RECT 18.785 3.245 18.955 3.415 ;
        RECT 20.635 3.245 20.805 3.415 ;
      LAYER met1 ;
        RECT 18.755 3.415 18.985 3.445 ;
        RECT 20.605 3.415 20.835 3.445 ;
        RECT 18.725 3.245 20.865 3.415 ;
        RECT 18.755 3.215 18.985 3.245 ;
        RECT 20.605 3.215 20.835 3.245 ;
    END
  END QN
  PIN D
    ANTENNAGATEAREA 1.033250 ;
    PORT
      LAYER li1 ;
        RECT 1.025 2.055 1.195 5.095 ;
      LAYER mcon ;
        RECT 1.025 3.985 1.195 4.155 ;
      LAYER met1 ;
        RECT 0.995 4.155 1.225 4.185 ;
        RECT 0.845 3.985 1.255 4.155 ;
        RECT 0.995 3.955 1.225 3.985 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 2.042100 ;
    PORT
      LAYER li1 ;
        RECT 5.465 2.055 5.635 5.095 ;
        RECT 14.745 4.975 14.915 5.095 ;
        RECT 14.715 4.765 14.915 4.975 ;
        RECT 14.715 2.055 14.885 4.765 ;
      LAYER mcon ;
        RECT 5.465 4.725 5.635 4.895 ;
        RECT 14.715 4.725 14.885 4.895 ;
      LAYER met1 ;
        RECT 5.435 4.895 5.665 4.925 ;
        RECT 14.685 4.895 14.915 4.925 ;
        RECT 5.405 4.725 14.945 4.895 ;
        RECT 5.435 4.695 5.665 4.725 ;
        RECT 14.685 4.695 14.915 4.725 ;
    END
  END CLK
  PIN SN
    ANTENNAGATEAREA 2.029700 ;
    PORT
      LAYER li1 ;
        RECT 10.275 2.055 10.445 5.095 ;
        RECT 21.745 2.055 21.915 5.095 ;
      LAYER mcon ;
        RECT 10.275 2.505 10.445 2.675 ;
        RECT 21.745 2.505 21.915 2.675 ;
      LAYER met1 ;
        RECT 10.245 2.675 10.475 2.705 ;
        RECT 21.715 2.675 21.945 2.705 ;
        RECT 10.215 2.505 21.975 2.675 ;
        RECT 10.245 2.475 10.475 2.505 ;
        RECT 21.715 2.475 21.945 2.505 ;
    END
  END SN
  PIN VDD
    ANTENNADIFFAREA 29.929150 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 24.840 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 24.575 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 0.705 5.365 0.875 7.460 ;
        RECT 1.585 5.785 1.755 7.460 ;
        RECT 2.465 5.785 2.635 7.460 ;
        RECT 3.175 4.340 3.485 7.460 ;
        RECT 4.335 5.445 4.505 7.460 ;
        RECT 5.215 5.785 5.385 7.460 ;
        RECT 6.095 5.785 6.265 7.460 ;
        RECT 6.975 5.785 7.145 7.460 ;
        RECT 7.985 4.340 8.295 7.460 ;
        RECT 9.145 5.445 9.315 7.460 ;
        RECT 10.025 5.785 10.195 7.460 ;
        RECT 10.905 5.785 11.075 7.460 ;
        RECT 11.785 5.785 11.955 7.460 ;
        RECT 12.795 4.340 13.105 7.460 ;
        RECT 13.655 5.365 13.825 7.460 ;
        RECT 14.535 5.785 14.705 7.460 ;
        RECT 15.415 5.785 15.585 7.460 ;
        RECT 16.125 4.340 16.435 7.460 ;
        RECT 16.985 5.365 17.155 7.460 ;
        RECT 17.865 5.785 18.035 7.460 ;
        RECT 18.745 5.785 18.915 7.460 ;
        RECT 19.455 4.340 19.765 7.460 ;
        RECT 20.615 5.445 20.785 7.460 ;
        RECT 21.495 5.785 21.665 7.460 ;
        RECT 22.375 5.785 22.545 7.460 ;
        RECT 23.255 5.785 23.425 7.460 ;
        RECT 24.265 4.340 24.575 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 0.995 7.525 1.165 7.695 ;
        RECT 1.355 7.525 1.525 7.695 ;
        RECT 1.805 7.525 1.975 7.695 ;
        RECT 2.165 7.525 2.335 7.695 ;
        RECT 2.525 7.525 2.695 7.695 ;
        RECT 2.885 7.525 3.055 7.695 ;
        RECT 3.605 7.525 3.775 7.695 ;
        RECT 3.965 7.525 4.135 7.695 ;
        RECT 4.325 7.525 4.495 7.695 ;
        RECT 4.685 7.525 4.855 7.695 ;
        RECT 5.045 7.525 5.215 7.695 ;
        RECT 5.405 7.525 5.575 7.695 ;
        RECT 5.895 7.525 6.065 7.695 ;
        RECT 6.255 7.525 6.425 7.695 ;
        RECT 6.615 7.525 6.785 7.695 ;
        RECT 6.975 7.525 7.145 7.695 ;
        RECT 7.335 7.525 7.505 7.695 ;
        RECT 7.695 7.525 7.865 7.695 ;
        RECT 8.415 7.525 8.585 7.695 ;
        RECT 8.775 7.525 8.945 7.695 ;
        RECT 9.135 7.525 9.305 7.695 ;
        RECT 9.495 7.525 9.665 7.695 ;
        RECT 9.855 7.525 10.025 7.695 ;
        RECT 10.215 7.525 10.385 7.695 ;
        RECT 10.705 7.525 10.875 7.695 ;
        RECT 11.065 7.525 11.235 7.695 ;
        RECT 11.425 7.525 11.595 7.695 ;
        RECT 11.785 7.525 11.955 7.695 ;
        RECT 12.145 7.525 12.315 7.695 ;
        RECT 12.505 7.525 12.675 7.695 ;
        RECT 13.225 7.525 13.395 7.695 ;
        RECT 13.585 7.525 13.755 7.695 ;
        RECT 13.945 7.525 14.115 7.695 ;
        RECT 14.305 7.525 14.475 7.695 ;
        RECT 14.755 7.525 14.925 7.695 ;
        RECT 15.115 7.525 15.285 7.695 ;
        RECT 15.475 7.525 15.645 7.695 ;
        RECT 15.835 7.525 16.005 7.695 ;
        RECT 16.555 7.525 16.725 7.695 ;
        RECT 16.915 7.525 17.085 7.695 ;
        RECT 17.275 7.525 17.445 7.695 ;
        RECT 17.635 7.525 17.805 7.695 ;
        RECT 18.085 7.525 18.255 7.695 ;
        RECT 18.445 7.525 18.615 7.695 ;
        RECT 18.805 7.525 18.975 7.695 ;
        RECT 19.165 7.525 19.335 7.695 ;
        RECT 19.885 7.525 20.055 7.695 ;
        RECT 20.245 7.525 20.415 7.695 ;
        RECT 20.605 7.525 20.775 7.695 ;
        RECT 20.965 7.525 21.135 7.695 ;
        RECT 21.325 7.525 21.495 7.695 ;
        RECT 21.685 7.525 21.855 7.695 ;
        RECT 22.175 7.525 22.345 7.695 ;
        RECT 22.535 7.525 22.705 7.695 ;
        RECT 22.895 7.525 23.065 7.695 ;
        RECT 23.255 7.525 23.425 7.695 ;
        RECT 23.615 7.525 23.785 7.695 ;
        RECT 23.975 7.525 24.145 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 24.575 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 18.067049 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 24.705 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 3.045 -0.075 3.615 -0.065 ;
        RECT 7.855 -0.075 8.425 -0.065 ;
        RECT 12.665 -0.075 13.235 -0.065 ;
        RECT 15.995 -0.075 16.565 -0.065 ;
        RECT 19.325 -0.075 19.895 -0.065 ;
        RECT 24.135 -0.075 24.705 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 1.095 0.310 1.265 1.260 ;
        RECT 3.175 0.310 3.485 2.860 ;
        RECT 4.320 0.310 4.490 1.270 ;
        RECT 7.985 0.310 8.295 2.860 ;
        RECT 9.130 0.310 9.300 1.270 ;
        RECT 12.795 0.310 13.105 2.860 ;
        RECT 14.045 0.310 14.215 1.260 ;
        RECT 16.125 0.310 16.435 2.860 ;
        RECT 17.375 0.310 17.545 1.260 ;
        RECT 19.455 0.310 19.765 2.860 ;
        RECT 20.600 0.310 20.770 1.270 ;
        RECT 24.265 0.310 24.575 2.860 ;
        RECT -0.155 0.000 24.575 0.310 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 0.995 0.065 1.165 0.235 ;
        RECT 1.355 0.065 1.525 0.235 ;
        RECT 1.805 0.065 1.975 0.235 ;
        RECT 2.165 0.065 2.335 0.235 ;
        RECT 2.525 0.065 2.695 0.235 ;
        RECT 2.885 0.065 3.055 0.235 ;
        RECT 3.605 0.065 3.775 0.235 ;
        RECT 3.965 0.065 4.135 0.235 ;
        RECT 4.325 0.065 4.495 0.235 ;
        RECT 4.685 0.065 4.855 0.235 ;
        RECT 5.045 0.065 5.215 0.235 ;
        RECT 5.405 0.065 5.575 0.235 ;
        RECT 5.895 0.065 6.065 0.235 ;
        RECT 6.255 0.065 6.425 0.235 ;
        RECT 6.615 0.065 6.785 0.235 ;
        RECT 6.975 0.065 7.145 0.235 ;
        RECT 7.335 0.065 7.505 0.235 ;
        RECT 7.695 0.065 7.865 0.235 ;
        RECT 8.415 0.065 8.585 0.235 ;
        RECT 8.775 0.065 8.945 0.235 ;
        RECT 9.135 0.065 9.305 0.235 ;
        RECT 9.495 0.065 9.665 0.235 ;
        RECT 9.855 0.065 10.025 0.235 ;
        RECT 10.215 0.065 10.385 0.235 ;
        RECT 10.705 0.065 10.875 0.235 ;
        RECT 11.065 0.065 11.235 0.235 ;
        RECT 11.425 0.065 11.595 0.235 ;
        RECT 11.785 0.065 11.955 0.235 ;
        RECT 12.145 0.065 12.315 0.235 ;
        RECT 12.505 0.065 12.675 0.235 ;
        RECT 13.225 0.065 13.395 0.235 ;
        RECT 13.585 0.065 13.755 0.235 ;
        RECT 13.945 0.065 14.115 0.235 ;
        RECT 14.305 0.065 14.475 0.235 ;
        RECT 14.755 0.065 14.925 0.235 ;
        RECT 15.115 0.065 15.285 0.235 ;
        RECT 15.475 0.065 15.645 0.235 ;
        RECT 15.835 0.065 16.005 0.235 ;
        RECT 16.555 0.065 16.725 0.235 ;
        RECT 16.915 0.065 17.085 0.235 ;
        RECT 17.275 0.065 17.445 0.235 ;
        RECT 17.635 0.065 17.805 0.235 ;
        RECT 18.085 0.065 18.255 0.235 ;
        RECT 18.445 0.065 18.615 0.235 ;
        RECT 18.805 0.065 18.975 0.235 ;
        RECT 19.165 0.065 19.335 0.235 ;
        RECT 19.885 0.065 20.055 0.235 ;
        RECT 20.245 0.065 20.415 0.235 ;
        RECT 20.605 0.065 20.775 0.235 ;
        RECT 20.965 0.065 21.135 0.235 ;
        RECT 21.325 0.065 21.495 0.235 ;
        RECT 21.685 0.065 21.855 0.235 ;
        RECT 22.175 0.065 22.345 0.235 ;
        RECT 22.535 0.065 22.705 0.235 ;
        RECT 22.895 0.065 23.065 0.235 ;
        RECT 23.255 0.065 23.425 0.235 ;
        RECT 23.615 0.065 23.785 0.235 ;
        RECT 23.975 0.065 24.145 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 24.575 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 1.145 5.515 1.315 7.250 ;
        RECT 2.025 5.515 2.195 7.250 ;
        RECT 1.145 5.345 2.675 5.515 ;
        RECT 1.795 4.940 1.965 5.095 ;
        RECT 1.765 4.765 1.965 4.940 ;
        RECT 1.765 2.055 1.935 4.765 ;
        RECT 0.610 1.805 0.780 1.885 ;
        RECT 1.580 1.805 1.750 1.885 ;
        RECT 2.505 1.880 2.675 5.345 ;
        RECT 4.775 5.470 4.945 7.250 ;
        RECT 5.655 5.470 5.825 7.250 ;
        RECT 6.535 5.470 6.705 7.250 ;
        RECT 9.585 5.470 9.755 7.250 ;
        RECT 10.465 5.470 10.635 7.250 ;
        RECT 11.345 5.470 11.515 7.250 ;
        RECT 14.095 5.515 14.265 7.250 ;
        RECT 14.975 5.515 15.145 7.250 ;
        RECT 4.775 5.300 7.485 5.470 ;
        RECT 9.585 5.300 12.295 5.470 ;
        RECT 14.095 5.345 15.625 5.515 ;
        RECT 4.355 2.055 4.525 5.095 ;
        RECT 6.575 2.055 6.745 5.095 ;
        RECT 7.315 4.605 7.485 5.300 ;
        RECT 7.310 4.275 7.485 4.605 ;
        RECT 0.610 1.635 1.750 1.805 ;
        RECT 0.610 0.505 0.780 1.635 ;
        RECT 1.580 0.755 1.750 1.635 ;
        RECT 2.065 1.710 2.675 1.880 ;
        RECT 3.835 1.815 4.005 1.895 ;
        RECT 4.805 1.815 4.975 1.895 ;
        RECT 5.775 1.815 5.945 1.895 ;
        RECT 2.065 0.975 2.235 1.710 ;
        RECT 3.835 1.645 5.945 1.815 ;
        RECT 2.550 0.755 2.720 1.525 ;
        RECT 1.580 0.585 2.720 0.755 ;
        RECT 1.580 0.505 1.750 0.585 ;
        RECT 2.550 0.505 2.720 0.585 ;
        RECT 3.835 0.515 4.005 1.645 ;
        RECT 4.805 0.765 4.975 1.645 ;
        RECT 5.775 1.565 5.945 1.645 ;
        RECT 5.295 1.220 5.465 1.300 ;
        RECT 6.345 1.220 6.515 1.895 ;
        RECT 7.315 1.890 7.485 4.275 ;
        RECT 9.165 2.055 9.335 5.095 ;
        RECT 11.385 2.055 11.555 5.095 ;
        RECT 5.295 1.050 6.515 1.220 ;
        RECT 5.295 0.970 5.465 1.050 ;
        RECT 5.775 0.765 5.945 0.845 ;
        RECT 4.805 0.595 5.945 0.765 ;
        RECT 4.805 0.515 4.975 0.595 ;
        RECT 5.775 0.515 5.945 0.595 ;
        RECT 6.345 0.765 6.515 1.050 ;
        RECT 6.830 1.720 7.485 1.890 ;
        RECT 8.645 1.815 8.815 1.895 ;
        RECT 9.615 1.815 9.785 1.895 ;
        RECT 10.585 1.815 10.755 1.895 ;
        RECT 6.830 0.985 7.000 1.720 ;
        RECT 8.645 1.645 10.755 1.815 ;
        RECT 7.315 0.765 7.485 1.535 ;
        RECT 6.345 0.595 7.485 0.765 ;
        RECT 6.345 0.515 6.515 0.595 ;
        RECT 7.315 0.515 7.485 0.595 ;
        RECT 8.645 0.515 8.815 1.645 ;
        RECT 9.615 0.765 9.785 1.645 ;
        RECT 10.585 1.565 10.755 1.645 ;
        RECT 10.105 1.220 10.275 1.300 ;
        RECT 11.155 1.220 11.325 1.895 ;
        RECT 12.125 1.890 12.295 5.300 ;
        RECT 13.975 2.055 14.145 5.095 ;
        RECT 10.105 1.050 11.325 1.220 ;
        RECT 10.105 0.970 10.275 1.050 ;
        RECT 10.585 0.765 10.755 0.845 ;
        RECT 9.615 0.595 10.755 0.765 ;
        RECT 9.615 0.515 9.785 0.595 ;
        RECT 10.585 0.515 10.755 0.595 ;
        RECT 11.155 0.765 11.325 1.050 ;
        RECT 11.640 1.720 12.295 1.890 ;
        RECT 13.560 1.805 13.730 1.885 ;
        RECT 14.530 1.805 14.700 1.885 ;
        RECT 15.455 1.880 15.625 5.345 ;
        RECT 21.055 5.470 21.225 7.250 ;
        RECT 21.935 5.470 22.105 7.250 ;
        RECT 22.815 5.470 22.985 7.250 ;
        RECT 21.055 5.300 23.765 5.470 ;
        RECT 17.305 2.055 17.475 5.095 ;
        RECT 18.075 4.940 18.245 5.095 ;
        RECT 18.045 4.765 18.245 4.940 ;
        RECT 18.045 2.055 18.215 4.765 ;
        RECT 22.855 2.055 23.025 5.095 ;
        RECT 11.640 0.985 11.810 1.720 ;
        RECT 13.560 1.635 14.700 1.805 ;
        RECT 12.125 0.765 12.295 1.535 ;
        RECT 11.155 0.595 12.295 0.765 ;
        RECT 11.155 0.515 11.325 0.595 ;
        RECT 12.125 0.515 12.295 0.595 ;
        RECT 13.560 0.505 13.730 1.635 ;
        RECT 14.530 0.755 14.700 1.635 ;
        RECT 15.015 1.710 15.625 1.880 ;
        RECT 16.890 1.805 17.060 1.885 ;
        RECT 17.860 1.805 18.030 1.885 ;
        RECT 15.015 0.975 15.185 1.710 ;
        RECT 16.890 1.635 18.030 1.805 ;
        RECT 15.500 0.755 15.670 1.525 ;
        RECT 14.530 0.585 15.670 0.755 ;
        RECT 14.530 0.505 14.700 0.585 ;
        RECT 15.500 0.505 15.670 0.585 ;
        RECT 16.890 0.505 17.060 1.635 ;
        RECT 17.860 0.755 18.030 1.635 ;
        RECT 20.115 1.815 20.285 1.895 ;
        RECT 21.085 1.815 21.255 1.895 ;
        RECT 22.055 1.815 22.225 1.895 ;
        RECT 20.115 1.645 22.225 1.815 ;
        RECT 18.830 0.755 19.000 1.525 ;
        RECT 17.860 0.585 19.000 0.755 ;
        RECT 17.860 0.505 18.030 0.585 ;
        RECT 18.830 0.505 19.000 0.585 ;
        RECT 20.115 0.515 20.285 1.645 ;
        RECT 21.085 0.765 21.255 1.645 ;
        RECT 22.055 1.565 22.225 1.645 ;
        RECT 21.575 1.220 21.745 1.300 ;
        RECT 22.625 1.220 22.795 1.895 ;
        RECT 23.595 1.890 23.765 5.300 ;
        RECT 21.575 1.050 22.795 1.220 ;
        RECT 21.575 0.970 21.745 1.050 ;
        RECT 22.055 0.765 22.225 0.845 ;
        RECT 21.085 0.595 22.225 0.765 ;
        RECT 21.085 0.515 21.255 0.595 ;
        RECT 22.055 0.515 22.225 0.595 ;
        RECT 22.625 0.765 22.795 1.050 ;
        RECT 23.110 1.720 23.765 1.890 ;
        RECT 23.110 0.985 23.280 1.720 ;
        RECT 23.595 0.765 23.765 1.535 ;
        RECT 22.625 0.595 23.765 0.765 ;
        RECT 22.625 0.515 22.795 0.595 ;
        RECT 23.595 0.515 23.765 0.595 ;
      LAYER mcon ;
        RECT 1.765 4.355 1.935 4.525 ;
        RECT 2.505 2.875 2.675 3.045 ;
        RECT 4.355 2.870 4.525 3.040 ;
        RECT 7.310 4.355 7.480 4.525 ;
        RECT 6.575 3.985 6.745 4.155 ;
        RECT 9.165 2.875 9.335 3.045 ;
        RECT 11.385 3.985 11.555 4.155 ;
        RECT 12.125 2.875 12.295 3.045 ;
        RECT 13.975 2.875 14.145 3.045 ;
        RECT 15.455 3.985 15.625 4.155 ;
        RECT 17.305 4.355 17.475 4.525 ;
        RECT 18.045 3.615 18.215 3.785 ;
        RECT 22.855 3.985 23.025 4.155 ;
        RECT 23.595 3.615 23.765 3.785 ;
      LAYER met1 ;
        RECT 1.735 4.525 1.965 4.555 ;
        RECT 7.280 4.525 7.510 4.555 ;
        RECT 17.275 4.525 17.505 4.555 ;
        RECT 1.705 4.355 17.535 4.525 ;
        RECT 1.735 4.325 1.965 4.355 ;
        RECT 7.280 4.325 7.510 4.355 ;
        RECT 17.275 4.325 17.505 4.355 ;
        RECT 6.545 4.155 6.775 4.185 ;
        RECT 11.355 4.155 11.585 4.185 ;
        RECT 15.425 4.155 15.655 4.185 ;
        RECT 22.825 4.155 23.055 4.185 ;
        RECT 6.515 3.985 23.085 4.155 ;
        RECT 6.545 3.955 6.775 3.985 ;
        RECT 11.355 3.955 11.585 3.985 ;
        RECT 15.425 3.955 15.655 3.985 ;
        RECT 22.825 3.955 23.055 3.985 ;
        RECT 18.015 3.785 18.245 3.815 ;
        RECT 23.565 3.785 23.795 3.815 ;
        RECT 17.985 3.615 23.825 3.785 ;
        RECT 18.015 3.585 18.245 3.615 ;
        RECT 23.565 3.585 23.795 3.615 ;
        RECT 2.475 3.045 2.705 3.075 ;
        RECT 4.325 3.045 4.555 3.070 ;
        RECT 9.135 3.045 9.365 3.075 ;
        RECT 12.095 3.045 12.325 3.075 ;
        RECT 13.945 3.045 14.175 3.075 ;
        RECT 2.445 2.875 9.395 3.045 ;
        RECT 12.065 2.875 14.205 3.045 ;
        RECT 2.475 2.845 2.705 2.875 ;
        RECT 4.295 2.870 4.705 2.875 ;
        RECT 4.325 2.840 4.555 2.870 ;
        RECT 9.135 2.845 9.365 2.875 ;
        RECT 12.095 2.845 12.325 2.875 ;
        RECT 13.945 2.845 14.175 2.875 ;
  END
END DFFSNQNX1






MACRO DFFSNQX1
  CLASS BLOCK ;
  FOREIGN DFFSNQX1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 25.260 BY 7.950 ;
  PIN Q
    ANTENNAGATEAREA 1.027250 ;
    ANTENNADIFFAREA 1.931900 ;
    PORT
      LAYER li1 ;
        RECT 21.055 5.470 21.225 7.250 ;
        RECT 21.935 5.470 22.105 7.250 ;
        RECT 22.815 5.470 22.985 7.250 ;
        RECT 21.055 5.300 23.765 5.470 ;
        RECT 18.075 4.940 18.245 5.095 ;
        RECT 18.045 4.765 18.245 4.940 ;
        RECT 18.045 2.055 18.215 4.765 ;
        RECT 23.595 1.890 23.765 5.300 ;
        RECT 23.110 1.720 23.765 1.890 ;
        RECT 23.110 0.985 23.280 1.720 ;
      LAYER mcon ;
        RECT 18.045 3.615 18.215 3.785 ;
        RECT 23.595 3.615 23.765 3.785 ;
      LAYER met1 ;
        RECT 18.015 3.785 18.245 3.815 ;
        RECT 23.565 3.785 23.795 3.815 ;
        RECT 17.985 3.615 23.825 3.785 ;
        RECT 18.015 3.585 18.245 3.615 ;
        RECT 23.565 3.585 23.795 3.615 ;
    END
  END Q
  PIN D
    ANTENNAGATEAREA 1.033250 ;
    PORT
      LAYER li1 ;
        RECT 1.025 2.055 1.195 5.095 ;
      LAYER mcon ;
        RECT 1.025 3.985 1.195 4.155 ;
      LAYER met1 ;
        RECT 0.995 4.155 1.225 4.185 ;
        RECT 0.845 3.985 1.255 4.155 ;
        RECT 0.995 3.955 1.225 3.985 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 2.042100 ;
    PORT
      LAYER li1 ;
        RECT 5.465 2.055 5.635 5.095 ;
        RECT 14.745 4.975 14.915 5.095 ;
        RECT 14.715 4.765 14.915 4.975 ;
        RECT 14.715 2.055 14.885 4.765 ;
      LAYER mcon ;
        RECT 5.465 4.725 5.635 4.895 ;
        RECT 14.715 4.725 14.885 4.895 ;
      LAYER met1 ;
        RECT 5.435 4.895 5.665 4.925 ;
        RECT 14.685 4.895 14.915 4.925 ;
        RECT 5.405 4.725 14.945 4.895 ;
        RECT 5.435 4.695 5.665 4.725 ;
        RECT 14.685 4.695 14.915 4.725 ;
    END
  END CLK
  PIN SN
    ANTENNAGATEAREA 2.029700 ;
    PORT
      LAYER li1 ;
        RECT 10.275 2.055 10.445 5.095 ;
        RECT 21.745 2.055 21.915 5.095 ;
      LAYER mcon ;
        RECT 10.275 2.505 10.445 2.675 ;
        RECT 21.745 2.505 21.915 2.675 ;
      LAYER met1 ;
        RECT 10.245 2.675 10.475 2.705 ;
        RECT 21.715 2.675 21.945 2.705 ;
        RECT 10.215 2.505 21.975 2.675 ;
        RECT 10.245 2.475 10.475 2.505 ;
        RECT 21.715 2.475 21.945 2.505 ;
    END
  END SN
  PIN VDD
    ANTENNADIFFAREA 29.929150 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 24.840 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 24.575 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 0.705 5.365 0.875 7.460 ;
        RECT 1.585 5.785 1.755 7.460 ;
        RECT 2.465 5.785 2.635 7.460 ;
        RECT 3.175 4.340 3.485 7.460 ;
        RECT 4.335 5.445 4.505 7.460 ;
        RECT 5.215 5.785 5.385 7.460 ;
        RECT 6.095 5.785 6.265 7.460 ;
        RECT 6.975 5.785 7.145 7.460 ;
        RECT 7.985 4.340 8.295 7.460 ;
        RECT 9.145 5.445 9.315 7.460 ;
        RECT 10.025 5.785 10.195 7.460 ;
        RECT 10.905 5.785 11.075 7.460 ;
        RECT 11.785 5.785 11.955 7.460 ;
        RECT 12.795 4.340 13.105 7.460 ;
        RECT 13.655 5.365 13.825 7.460 ;
        RECT 14.535 5.785 14.705 7.460 ;
        RECT 15.415 5.785 15.585 7.460 ;
        RECT 16.125 4.340 16.435 7.460 ;
        RECT 16.985 5.365 17.155 7.460 ;
        RECT 17.865 5.785 18.035 7.460 ;
        RECT 18.745 5.785 18.915 7.460 ;
        RECT 19.455 4.340 19.765 7.460 ;
        RECT 20.615 5.445 20.785 7.460 ;
        RECT 21.495 5.785 21.665 7.460 ;
        RECT 22.375 5.785 22.545 7.460 ;
        RECT 23.255 5.785 23.425 7.460 ;
        RECT 24.265 4.340 24.575 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 0.995 7.525 1.165 7.695 ;
        RECT 1.355 7.525 1.525 7.695 ;
        RECT 1.805 7.525 1.975 7.695 ;
        RECT 2.165 7.525 2.335 7.695 ;
        RECT 2.525 7.525 2.695 7.695 ;
        RECT 2.885 7.525 3.055 7.695 ;
        RECT 3.605 7.525 3.775 7.695 ;
        RECT 3.965 7.525 4.135 7.695 ;
        RECT 4.325 7.525 4.495 7.695 ;
        RECT 4.685 7.525 4.855 7.695 ;
        RECT 5.045 7.525 5.215 7.695 ;
        RECT 5.405 7.525 5.575 7.695 ;
        RECT 5.895 7.525 6.065 7.695 ;
        RECT 6.255 7.525 6.425 7.695 ;
        RECT 6.615 7.525 6.785 7.695 ;
        RECT 6.975 7.525 7.145 7.695 ;
        RECT 7.335 7.525 7.505 7.695 ;
        RECT 7.695 7.525 7.865 7.695 ;
        RECT 8.415 7.525 8.585 7.695 ;
        RECT 8.775 7.525 8.945 7.695 ;
        RECT 9.135 7.525 9.305 7.695 ;
        RECT 9.495 7.525 9.665 7.695 ;
        RECT 9.855 7.525 10.025 7.695 ;
        RECT 10.215 7.525 10.385 7.695 ;
        RECT 10.705 7.525 10.875 7.695 ;
        RECT 11.065 7.525 11.235 7.695 ;
        RECT 11.425 7.525 11.595 7.695 ;
        RECT 11.785 7.525 11.955 7.695 ;
        RECT 12.145 7.525 12.315 7.695 ;
        RECT 12.505 7.525 12.675 7.695 ;
        RECT 13.225 7.525 13.395 7.695 ;
        RECT 13.585 7.525 13.755 7.695 ;
        RECT 13.945 7.525 14.115 7.695 ;
        RECT 14.305 7.525 14.475 7.695 ;
        RECT 14.755 7.525 14.925 7.695 ;
        RECT 15.115 7.525 15.285 7.695 ;
        RECT 15.475 7.525 15.645 7.695 ;
        RECT 15.835 7.525 16.005 7.695 ;
        RECT 16.555 7.525 16.725 7.695 ;
        RECT 16.915 7.525 17.085 7.695 ;
        RECT 17.275 7.525 17.445 7.695 ;
        RECT 17.635 7.525 17.805 7.695 ;
        RECT 18.085 7.525 18.255 7.695 ;
        RECT 18.445 7.525 18.615 7.695 ;
        RECT 18.805 7.525 18.975 7.695 ;
        RECT 19.165 7.525 19.335 7.695 ;
        RECT 19.885 7.525 20.055 7.695 ;
        RECT 20.245 7.525 20.415 7.695 ;
        RECT 20.605 7.525 20.775 7.695 ;
        RECT 20.965 7.525 21.135 7.695 ;
        RECT 21.325 7.525 21.495 7.695 ;
        RECT 21.685 7.525 21.855 7.695 ;
        RECT 22.175 7.525 22.345 7.695 ;
        RECT 22.535 7.525 22.705 7.695 ;
        RECT 22.895 7.525 23.065 7.695 ;
        RECT 23.255 7.525 23.425 7.695 ;
        RECT 23.615 7.525 23.785 7.695 ;
        RECT 23.975 7.525 24.145 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 24.575 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 18.067049 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 24.705 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 3.045 -0.075 3.615 -0.065 ;
        RECT 7.855 -0.075 8.425 -0.065 ;
        RECT 12.665 -0.075 13.235 -0.065 ;
        RECT 15.995 -0.075 16.565 -0.065 ;
        RECT 19.325 -0.075 19.895 -0.065 ;
        RECT 24.135 -0.075 24.705 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 1.095 0.310 1.265 1.260 ;
        RECT 3.175 0.310 3.485 2.860 ;
        RECT 4.320 0.310 4.490 1.270 ;
        RECT 7.985 0.310 8.295 2.860 ;
        RECT 9.130 0.310 9.300 1.270 ;
        RECT 12.795 0.310 13.105 2.860 ;
        RECT 14.045 0.310 14.215 1.260 ;
        RECT 16.125 0.310 16.435 2.860 ;
        RECT 17.375 0.310 17.545 1.260 ;
        RECT 19.455 0.310 19.765 2.860 ;
        RECT 20.600 0.310 20.770 1.270 ;
        RECT 24.265 0.310 24.575 2.860 ;
        RECT -0.155 0.000 24.575 0.310 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 0.995 0.065 1.165 0.235 ;
        RECT 1.355 0.065 1.525 0.235 ;
        RECT 1.805 0.065 1.975 0.235 ;
        RECT 2.165 0.065 2.335 0.235 ;
        RECT 2.525 0.065 2.695 0.235 ;
        RECT 2.885 0.065 3.055 0.235 ;
        RECT 3.605 0.065 3.775 0.235 ;
        RECT 3.965 0.065 4.135 0.235 ;
        RECT 4.325 0.065 4.495 0.235 ;
        RECT 4.685 0.065 4.855 0.235 ;
        RECT 5.045 0.065 5.215 0.235 ;
        RECT 5.405 0.065 5.575 0.235 ;
        RECT 5.895 0.065 6.065 0.235 ;
        RECT 6.255 0.065 6.425 0.235 ;
        RECT 6.615 0.065 6.785 0.235 ;
        RECT 6.975 0.065 7.145 0.235 ;
        RECT 7.335 0.065 7.505 0.235 ;
        RECT 7.695 0.065 7.865 0.235 ;
        RECT 8.415 0.065 8.585 0.235 ;
        RECT 8.775 0.065 8.945 0.235 ;
        RECT 9.135 0.065 9.305 0.235 ;
        RECT 9.495 0.065 9.665 0.235 ;
        RECT 9.855 0.065 10.025 0.235 ;
        RECT 10.215 0.065 10.385 0.235 ;
        RECT 10.705 0.065 10.875 0.235 ;
        RECT 11.065 0.065 11.235 0.235 ;
        RECT 11.425 0.065 11.595 0.235 ;
        RECT 11.785 0.065 11.955 0.235 ;
        RECT 12.145 0.065 12.315 0.235 ;
        RECT 12.505 0.065 12.675 0.235 ;
        RECT 13.225 0.065 13.395 0.235 ;
        RECT 13.585 0.065 13.755 0.235 ;
        RECT 13.945 0.065 14.115 0.235 ;
        RECT 14.305 0.065 14.475 0.235 ;
        RECT 14.755 0.065 14.925 0.235 ;
        RECT 15.115 0.065 15.285 0.235 ;
        RECT 15.475 0.065 15.645 0.235 ;
        RECT 15.835 0.065 16.005 0.235 ;
        RECT 16.555 0.065 16.725 0.235 ;
        RECT 16.915 0.065 17.085 0.235 ;
        RECT 17.275 0.065 17.445 0.235 ;
        RECT 17.635 0.065 17.805 0.235 ;
        RECT 18.085 0.065 18.255 0.235 ;
        RECT 18.445 0.065 18.615 0.235 ;
        RECT 18.805 0.065 18.975 0.235 ;
        RECT 19.165 0.065 19.335 0.235 ;
        RECT 19.885 0.065 20.055 0.235 ;
        RECT 20.245 0.065 20.415 0.235 ;
        RECT 20.605 0.065 20.775 0.235 ;
        RECT 20.965 0.065 21.135 0.235 ;
        RECT 21.325 0.065 21.495 0.235 ;
        RECT 21.685 0.065 21.855 0.235 ;
        RECT 22.175 0.065 22.345 0.235 ;
        RECT 22.535 0.065 22.705 0.235 ;
        RECT 22.895 0.065 23.065 0.235 ;
        RECT 23.255 0.065 23.425 0.235 ;
        RECT 23.615 0.065 23.785 0.235 ;
        RECT 23.975 0.065 24.145 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 24.575 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 1.145 5.515 1.315 7.250 ;
        RECT 2.025 5.515 2.195 7.250 ;
        RECT 1.145 5.345 2.675 5.515 ;
        RECT 1.795 4.940 1.965 5.095 ;
        RECT 1.765 4.765 1.965 4.940 ;
        RECT 1.765 2.055 1.935 4.765 ;
        RECT 0.610 1.805 0.780 1.885 ;
        RECT 1.580 1.805 1.750 1.885 ;
        RECT 2.505 1.880 2.675 5.345 ;
        RECT 4.775 5.470 4.945 7.250 ;
        RECT 5.655 5.470 5.825 7.250 ;
        RECT 6.535 5.470 6.705 7.250 ;
        RECT 9.585 5.470 9.755 7.250 ;
        RECT 10.465 5.470 10.635 7.250 ;
        RECT 11.345 5.470 11.515 7.250 ;
        RECT 14.095 5.515 14.265 7.250 ;
        RECT 14.975 5.515 15.145 7.250 ;
        RECT 17.425 5.515 17.595 7.250 ;
        RECT 18.305 5.515 18.475 7.250 ;
        RECT 4.775 5.300 7.485 5.470 ;
        RECT 9.585 5.300 12.295 5.470 ;
        RECT 14.095 5.345 15.625 5.515 ;
        RECT 17.425 5.345 18.955 5.515 ;
        RECT 4.355 2.055 4.525 5.095 ;
        RECT 6.575 2.055 6.745 5.095 ;
        RECT 7.315 4.605 7.485 5.300 ;
        RECT 7.310 4.275 7.485 4.605 ;
        RECT 0.610 1.635 1.750 1.805 ;
        RECT 0.610 0.505 0.780 1.635 ;
        RECT 1.580 0.755 1.750 1.635 ;
        RECT 2.065 1.710 2.675 1.880 ;
        RECT 3.835 1.815 4.005 1.895 ;
        RECT 4.805 1.815 4.975 1.895 ;
        RECT 5.775 1.815 5.945 1.895 ;
        RECT 2.065 0.975 2.235 1.710 ;
        RECT 3.835 1.645 5.945 1.815 ;
        RECT 2.550 0.755 2.720 1.525 ;
        RECT 1.580 0.585 2.720 0.755 ;
        RECT 1.580 0.505 1.750 0.585 ;
        RECT 2.550 0.505 2.720 0.585 ;
        RECT 3.835 0.515 4.005 1.645 ;
        RECT 4.805 0.765 4.975 1.645 ;
        RECT 5.775 1.565 5.945 1.645 ;
        RECT 5.295 1.220 5.465 1.300 ;
        RECT 6.345 1.220 6.515 1.895 ;
        RECT 7.315 1.890 7.485 4.275 ;
        RECT 9.165 2.055 9.335 5.095 ;
        RECT 11.385 2.055 11.555 5.095 ;
        RECT 5.295 1.050 6.515 1.220 ;
        RECT 5.295 0.970 5.465 1.050 ;
        RECT 5.775 0.765 5.945 0.845 ;
        RECT 4.805 0.595 5.945 0.765 ;
        RECT 4.805 0.515 4.975 0.595 ;
        RECT 5.775 0.515 5.945 0.595 ;
        RECT 6.345 0.765 6.515 1.050 ;
        RECT 6.830 1.720 7.485 1.890 ;
        RECT 8.645 1.815 8.815 1.895 ;
        RECT 9.615 1.815 9.785 1.895 ;
        RECT 10.585 1.815 10.755 1.895 ;
        RECT 6.830 0.985 7.000 1.720 ;
        RECT 8.645 1.645 10.755 1.815 ;
        RECT 7.315 0.765 7.485 1.535 ;
        RECT 6.345 0.595 7.485 0.765 ;
        RECT 6.345 0.515 6.515 0.595 ;
        RECT 7.315 0.515 7.485 0.595 ;
        RECT 8.645 0.515 8.815 1.645 ;
        RECT 9.615 0.765 9.785 1.645 ;
        RECT 10.585 1.565 10.755 1.645 ;
        RECT 10.105 1.220 10.275 1.300 ;
        RECT 11.155 1.220 11.325 1.895 ;
        RECT 12.125 1.890 12.295 5.300 ;
        RECT 13.975 2.055 14.145 5.095 ;
        RECT 10.105 1.050 11.325 1.220 ;
        RECT 10.105 0.970 10.275 1.050 ;
        RECT 10.585 0.765 10.755 0.845 ;
        RECT 9.615 0.595 10.755 0.765 ;
        RECT 9.615 0.515 9.785 0.595 ;
        RECT 10.585 0.515 10.755 0.595 ;
        RECT 11.155 0.765 11.325 1.050 ;
        RECT 11.640 1.720 12.295 1.890 ;
        RECT 13.560 1.805 13.730 1.885 ;
        RECT 14.530 1.805 14.700 1.885 ;
        RECT 15.455 1.880 15.625 5.345 ;
        RECT 17.305 2.055 17.475 5.095 ;
        RECT 11.640 0.985 11.810 1.720 ;
        RECT 13.560 1.635 14.700 1.805 ;
        RECT 12.125 0.765 12.295 1.535 ;
        RECT 11.155 0.595 12.295 0.765 ;
        RECT 11.155 0.515 11.325 0.595 ;
        RECT 12.125 0.515 12.295 0.595 ;
        RECT 13.560 0.505 13.730 1.635 ;
        RECT 14.530 0.755 14.700 1.635 ;
        RECT 15.015 1.710 15.625 1.880 ;
        RECT 16.890 1.805 17.060 1.885 ;
        RECT 17.860 1.805 18.030 1.885 ;
        RECT 18.785 1.880 18.955 5.345 ;
        RECT 20.635 2.055 20.805 5.095 ;
        RECT 22.855 2.055 23.025 5.095 ;
        RECT 15.015 0.975 15.185 1.710 ;
        RECT 16.890 1.635 18.030 1.805 ;
        RECT 15.500 0.755 15.670 1.525 ;
        RECT 14.530 0.585 15.670 0.755 ;
        RECT 14.530 0.505 14.700 0.585 ;
        RECT 15.500 0.505 15.670 0.585 ;
        RECT 16.890 0.505 17.060 1.635 ;
        RECT 17.860 0.755 18.030 1.635 ;
        RECT 18.345 1.710 18.955 1.880 ;
        RECT 20.115 1.815 20.285 1.895 ;
        RECT 21.085 1.815 21.255 1.895 ;
        RECT 22.055 1.815 22.225 1.895 ;
        RECT 18.345 0.975 18.515 1.710 ;
        RECT 20.115 1.645 22.225 1.815 ;
        RECT 18.830 0.755 19.000 1.525 ;
        RECT 17.860 0.585 19.000 0.755 ;
        RECT 17.860 0.505 18.030 0.585 ;
        RECT 18.830 0.505 19.000 0.585 ;
        RECT 20.115 0.515 20.285 1.645 ;
        RECT 21.085 0.765 21.255 1.645 ;
        RECT 22.055 1.565 22.225 1.645 ;
        RECT 21.575 1.220 21.745 1.300 ;
        RECT 22.625 1.220 22.795 1.895 ;
        RECT 21.575 1.050 22.795 1.220 ;
        RECT 21.575 0.970 21.745 1.050 ;
        RECT 22.055 0.765 22.225 0.845 ;
        RECT 21.085 0.595 22.225 0.765 ;
        RECT 21.085 0.515 21.255 0.595 ;
        RECT 22.055 0.515 22.225 0.595 ;
        RECT 22.625 0.765 22.795 1.050 ;
        RECT 23.595 0.765 23.765 1.535 ;
        RECT 22.625 0.595 23.765 0.765 ;
        RECT 22.625 0.515 22.795 0.595 ;
        RECT 23.595 0.515 23.765 0.595 ;
      LAYER mcon ;
        RECT 1.765 4.355 1.935 4.525 ;
        RECT 2.505 2.875 2.675 3.045 ;
        RECT 4.355 2.870 4.525 3.040 ;
        RECT 7.310 4.355 7.480 4.525 ;
        RECT 6.575 3.985 6.745 4.155 ;
        RECT 9.165 2.875 9.335 3.045 ;
        RECT 11.385 3.985 11.555 4.155 ;
        RECT 12.125 2.875 12.295 3.045 ;
        RECT 13.975 2.875 14.145 3.045 ;
        RECT 15.455 3.985 15.625 4.155 ;
        RECT 17.305 4.355 17.475 4.525 ;
        RECT 18.785 3.245 18.955 3.415 ;
        RECT 20.635 3.245 20.805 3.415 ;
        RECT 22.855 3.985 23.025 4.155 ;
      LAYER met1 ;
        RECT 1.735 4.525 1.965 4.555 ;
        RECT 7.280 4.525 7.510 4.555 ;
        RECT 17.275 4.525 17.505 4.555 ;
        RECT 1.705 4.355 17.535 4.525 ;
        RECT 1.735 4.325 1.965 4.355 ;
        RECT 7.280 4.325 7.510 4.355 ;
        RECT 17.275 4.325 17.505 4.355 ;
        RECT 6.545 4.155 6.775 4.185 ;
        RECT 11.355 4.155 11.585 4.185 ;
        RECT 15.425 4.155 15.655 4.185 ;
        RECT 22.825 4.155 23.055 4.185 ;
        RECT 6.515 3.985 23.085 4.155 ;
        RECT 6.545 3.955 6.775 3.985 ;
        RECT 11.355 3.955 11.585 3.985 ;
        RECT 15.425 3.955 15.655 3.985 ;
        RECT 22.825 3.955 23.055 3.985 ;
        RECT 18.755 3.415 18.985 3.445 ;
        RECT 20.605 3.415 20.835 3.445 ;
        RECT 18.725 3.245 20.865 3.415 ;
        RECT 18.755 3.215 18.985 3.245 ;
        RECT 20.605 3.215 20.835 3.245 ;
        RECT 2.475 3.045 2.705 3.075 ;
        RECT 4.325 3.045 4.555 3.070 ;
        RECT 9.135 3.045 9.365 3.075 ;
        RECT 12.095 3.045 12.325 3.075 ;
        RECT 13.945 3.045 14.175 3.075 ;
        RECT 2.445 2.875 9.395 3.045 ;
        RECT 12.065 2.875 14.205 3.045 ;
        RECT 2.475 2.845 2.705 2.875 ;
        RECT 4.295 2.870 4.705 2.875 ;
        RECT 4.325 2.840 4.555 2.870 ;
        RECT 9.135 2.845 9.365 2.875 ;
        RECT 12.095 2.845 12.325 2.875 ;
        RECT 13.945 2.845 14.175 2.875 ;
  END
END DFFSNQX1






MACRO DFFSNRNQNX1
  CLASS BLOCK ;
  FOREIGN DFFSNRNQNX1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 29.700 BY 7.950 ;
  PIN QN
    ANTENNAGATEAREA 1.033250 ;
    ANTENNADIFFAREA 1.931900 ;
    PORT
      LAYER li1 ;
        RECT 20.685 5.470 20.855 7.250 ;
        RECT 21.565 5.470 21.735 7.250 ;
        RECT 22.445 5.470 22.615 7.250 ;
        RECT 20.685 5.300 23.395 5.470 ;
        RECT 23.225 1.890 23.395 5.300 ;
        RECT 25.075 2.055 25.245 5.095 ;
        RECT 22.740 1.720 23.395 1.890 ;
        RECT 22.740 0.985 22.910 1.720 ;
      LAYER mcon ;
        RECT 23.225 3.245 23.395 3.415 ;
        RECT 25.075 3.245 25.245 3.415 ;
      LAYER met1 ;
        RECT 23.195 3.415 23.425 3.445 ;
        RECT 25.045 3.415 25.275 3.445 ;
        RECT 23.165 3.245 25.305 3.415 ;
        RECT 23.195 3.215 23.425 3.245 ;
        RECT 25.045 3.215 25.275 3.245 ;
    END
  END QN
  PIN D
    ANTENNAGATEAREA 1.033250 ;
    PORT
      LAYER li1 ;
        RECT 1.025 2.055 1.195 5.095 ;
      LAYER mcon ;
        RECT 1.025 2.875 1.195 3.045 ;
      LAYER met1 ;
        RECT 0.995 3.045 1.225 3.075 ;
        RECT 0.845 2.875 1.255 3.045 ;
        RECT 0.995 2.845 1.225 2.875 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 2.029700 ;
    PORT
      LAYER li1 ;
        RECT 6.945 2.055 7.115 5.095 ;
        RECT 16.565 2.055 16.735 5.095 ;
      LAYER mcon ;
        RECT 6.945 3.245 7.115 3.415 ;
        RECT 16.565 3.245 16.735 3.415 ;
      LAYER met1 ;
        RECT 6.915 3.415 7.145 3.445 ;
        RECT 16.535 3.415 16.765 3.445 ;
        RECT 6.885 3.245 16.795 3.415 ;
        RECT 6.915 3.215 7.145 3.245 ;
        RECT 16.535 3.215 16.765 3.245 ;
    END
  END CLK
  PIN SN
    ANTENNAGATEAREA 2.029700 ;
    PORT
      LAYER li1 ;
        RECT 11.755 2.055 11.925 5.095 ;
        RECT 26.185 2.055 26.355 5.095 ;
      LAYER mcon ;
        RECT 11.755 2.510 11.925 2.680 ;
        RECT 26.185 2.505 26.355 2.675 ;
      LAYER met1 ;
        RECT 11.725 2.680 11.955 2.710 ;
        RECT 11.695 2.675 12.105 2.680 ;
        RECT 26.155 2.675 26.385 2.705 ;
        RECT 11.695 2.510 26.415 2.675 ;
        RECT 11.725 2.505 26.415 2.510 ;
        RECT 11.725 2.480 11.955 2.505 ;
        RECT 26.155 2.475 26.385 2.505 ;
    END
  END SN
  PIN RN
    ANTENNAGATEAREA 3.056950 ;
    PORT
      LAYER li1 ;
        RECT 2.135 2.055 2.305 5.095 ;
        RECT 17.675 2.055 17.845 5.095 ;
        RECT 21.375 2.055 21.545 5.095 ;
      LAYER mcon ;
        RECT 2.135 4.355 2.305 4.525 ;
        RECT 17.675 4.355 17.845 4.525 ;
        RECT 21.375 4.355 21.545 4.525 ;
      LAYER met1 ;
        RECT 2.105 4.525 2.335 4.555 ;
        RECT 17.645 4.525 17.875 4.555 ;
        RECT 21.345 4.525 21.575 4.555 ;
        RECT 2.075 4.355 21.605 4.525 ;
        RECT 2.105 4.325 2.335 4.355 ;
        RECT 17.645 4.325 17.875 4.355 ;
        RECT 21.345 4.325 21.575 4.355 ;
    END
  END RN
  PIN VDD
    ANTENNADIFFAREA 33.800350 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 29.280 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 29.015 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 1.005 5.445 1.175 7.460 ;
        RECT 1.885 5.785 2.055 7.460 ;
        RECT 2.765 5.785 2.935 7.460 ;
        RECT 3.645 5.785 3.815 7.460 ;
        RECT 4.655 4.340 4.965 7.460 ;
        RECT 5.815 5.445 5.985 7.460 ;
        RECT 6.695 5.785 6.865 7.460 ;
        RECT 7.575 5.785 7.745 7.460 ;
        RECT 8.455 5.785 8.625 7.460 ;
        RECT 9.465 4.340 9.775 7.460 ;
        RECT 10.625 5.445 10.795 7.460 ;
        RECT 11.505 5.785 11.675 7.460 ;
        RECT 12.385 5.785 12.555 7.460 ;
        RECT 13.265 5.785 13.435 7.460 ;
        RECT 14.275 4.340 14.585 7.460 ;
        RECT 15.435 5.445 15.605 7.460 ;
        RECT 16.315 5.785 16.485 7.460 ;
        RECT 17.195 5.785 17.365 7.460 ;
        RECT 18.075 5.785 18.245 7.460 ;
        RECT 19.085 4.340 19.395 7.460 ;
        RECT 20.245 5.445 20.415 7.460 ;
        RECT 21.125 5.785 21.295 7.460 ;
        RECT 22.005 5.785 22.175 7.460 ;
        RECT 22.885 5.785 23.055 7.460 ;
        RECT 23.895 4.340 24.205 7.460 ;
        RECT 25.055 5.445 25.225 7.460 ;
        RECT 25.935 5.785 26.105 7.460 ;
        RECT 26.815 5.785 26.985 7.460 ;
        RECT 27.695 5.785 27.865 7.460 ;
        RECT 28.705 4.340 29.015 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 0.995 7.525 1.165 7.695 ;
        RECT 1.355 7.525 1.525 7.695 ;
        RECT 1.715 7.525 1.885 7.695 ;
        RECT 2.075 7.525 2.245 7.695 ;
        RECT 2.565 7.525 2.735 7.695 ;
        RECT 2.925 7.525 3.095 7.695 ;
        RECT 3.285 7.525 3.455 7.695 ;
        RECT 3.645 7.525 3.815 7.695 ;
        RECT 4.005 7.525 4.175 7.695 ;
        RECT 4.365 7.525 4.535 7.695 ;
        RECT 5.085 7.525 5.255 7.695 ;
        RECT 5.445 7.525 5.615 7.695 ;
        RECT 5.805 7.525 5.975 7.695 ;
        RECT 6.165 7.525 6.335 7.695 ;
        RECT 6.525 7.525 6.695 7.695 ;
        RECT 6.885 7.525 7.055 7.695 ;
        RECT 7.375 7.525 7.545 7.695 ;
        RECT 7.735 7.525 7.905 7.695 ;
        RECT 8.095 7.525 8.265 7.695 ;
        RECT 8.455 7.525 8.625 7.695 ;
        RECT 8.815 7.525 8.985 7.695 ;
        RECT 9.175 7.525 9.345 7.695 ;
        RECT 9.895 7.525 10.065 7.695 ;
        RECT 10.255 7.525 10.425 7.695 ;
        RECT 10.615 7.525 10.785 7.695 ;
        RECT 10.975 7.525 11.145 7.695 ;
        RECT 11.335 7.525 11.505 7.695 ;
        RECT 11.695 7.525 11.865 7.695 ;
        RECT 12.185 7.525 12.355 7.695 ;
        RECT 12.545 7.525 12.715 7.695 ;
        RECT 12.905 7.525 13.075 7.695 ;
        RECT 13.265 7.525 13.435 7.695 ;
        RECT 13.625 7.525 13.795 7.695 ;
        RECT 13.985 7.525 14.155 7.695 ;
        RECT 14.705 7.525 14.875 7.695 ;
        RECT 15.065 7.525 15.235 7.695 ;
        RECT 15.425 7.525 15.595 7.695 ;
        RECT 15.785 7.525 15.955 7.695 ;
        RECT 16.145 7.525 16.315 7.695 ;
        RECT 16.505 7.525 16.675 7.695 ;
        RECT 16.995 7.525 17.165 7.695 ;
        RECT 17.355 7.525 17.525 7.695 ;
        RECT 17.715 7.525 17.885 7.695 ;
        RECT 18.075 7.525 18.245 7.695 ;
        RECT 18.435 7.525 18.605 7.695 ;
        RECT 18.795 7.525 18.965 7.695 ;
        RECT 19.515 7.525 19.685 7.695 ;
        RECT 19.875 7.525 20.045 7.695 ;
        RECT 20.235 7.525 20.405 7.695 ;
        RECT 20.595 7.525 20.765 7.695 ;
        RECT 20.955 7.525 21.125 7.695 ;
        RECT 21.315 7.525 21.485 7.695 ;
        RECT 21.805 7.525 21.975 7.695 ;
        RECT 22.165 7.525 22.335 7.695 ;
        RECT 22.525 7.525 22.695 7.695 ;
        RECT 22.885 7.525 23.055 7.695 ;
        RECT 23.245 7.525 23.415 7.695 ;
        RECT 23.605 7.525 23.775 7.695 ;
        RECT 24.325 7.525 24.495 7.695 ;
        RECT 24.685 7.525 24.855 7.695 ;
        RECT 25.045 7.525 25.215 7.695 ;
        RECT 25.405 7.525 25.575 7.695 ;
        RECT 25.765 7.525 25.935 7.695 ;
        RECT 26.125 7.525 26.295 7.695 ;
        RECT 26.615 7.525 26.785 7.695 ;
        RECT 26.975 7.525 27.145 7.695 ;
        RECT 27.335 7.525 27.505 7.695 ;
        RECT 27.695 7.525 27.865 7.695 ;
        RECT 28.055 7.525 28.225 7.695 ;
        RECT 28.415 7.525 28.585 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 29.015 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 20.198250 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 29.145 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 4.525 -0.075 5.095 -0.065 ;
        RECT 9.335 -0.075 9.905 -0.065 ;
        RECT 14.145 -0.075 14.715 -0.065 ;
        RECT 18.955 -0.075 19.525 -0.065 ;
        RECT 23.765 -0.075 24.335 -0.065 ;
        RECT 28.575 -0.075 29.145 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 0.990 0.310 1.160 1.270 ;
        RECT 4.655 0.310 4.965 2.860 ;
        RECT 5.800 0.310 5.970 1.270 ;
        RECT 9.465 0.310 9.775 2.860 ;
        RECT 10.610 0.310 10.780 1.270 ;
        RECT 14.275 0.310 14.585 2.860 ;
        RECT 15.420 0.310 15.590 1.270 ;
        RECT 19.085 0.310 19.395 2.860 ;
        RECT 20.230 0.310 20.400 1.270 ;
        RECT 23.895 0.310 24.205 2.860 ;
        RECT 25.040 0.310 25.210 1.270 ;
        RECT 28.705 0.310 29.015 2.860 ;
        RECT -0.155 0.000 29.015 0.310 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 0.995 0.065 1.165 0.235 ;
        RECT 1.355 0.065 1.525 0.235 ;
        RECT 1.715 0.065 1.885 0.235 ;
        RECT 2.075 0.065 2.245 0.235 ;
        RECT 2.565 0.065 2.735 0.235 ;
        RECT 2.925 0.065 3.095 0.235 ;
        RECT 3.285 0.065 3.455 0.235 ;
        RECT 3.645 0.065 3.815 0.235 ;
        RECT 4.005 0.065 4.175 0.235 ;
        RECT 4.365 0.065 4.535 0.235 ;
        RECT 5.085 0.065 5.255 0.235 ;
        RECT 5.445 0.065 5.615 0.235 ;
        RECT 5.805 0.065 5.975 0.235 ;
        RECT 6.165 0.065 6.335 0.235 ;
        RECT 6.525 0.065 6.695 0.235 ;
        RECT 6.885 0.065 7.055 0.235 ;
        RECT 7.375 0.065 7.545 0.235 ;
        RECT 7.735 0.065 7.905 0.235 ;
        RECT 8.095 0.065 8.265 0.235 ;
        RECT 8.455 0.065 8.625 0.235 ;
        RECT 8.815 0.065 8.985 0.235 ;
        RECT 9.175 0.065 9.345 0.235 ;
        RECT 9.895 0.065 10.065 0.235 ;
        RECT 10.255 0.065 10.425 0.235 ;
        RECT 10.615 0.065 10.785 0.235 ;
        RECT 10.975 0.065 11.145 0.235 ;
        RECT 11.335 0.065 11.505 0.235 ;
        RECT 11.695 0.065 11.865 0.235 ;
        RECT 12.185 0.065 12.355 0.235 ;
        RECT 12.545 0.065 12.715 0.235 ;
        RECT 12.905 0.065 13.075 0.235 ;
        RECT 13.265 0.065 13.435 0.235 ;
        RECT 13.625 0.065 13.795 0.235 ;
        RECT 13.985 0.065 14.155 0.235 ;
        RECT 14.705 0.065 14.875 0.235 ;
        RECT 15.065 0.065 15.235 0.235 ;
        RECT 15.425 0.065 15.595 0.235 ;
        RECT 15.785 0.065 15.955 0.235 ;
        RECT 16.145 0.065 16.315 0.235 ;
        RECT 16.505 0.065 16.675 0.235 ;
        RECT 16.995 0.065 17.165 0.235 ;
        RECT 17.355 0.065 17.525 0.235 ;
        RECT 17.715 0.065 17.885 0.235 ;
        RECT 18.075 0.065 18.245 0.235 ;
        RECT 18.435 0.065 18.605 0.235 ;
        RECT 18.795 0.065 18.965 0.235 ;
        RECT 19.515 0.065 19.685 0.235 ;
        RECT 19.875 0.065 20.045 0.235 ;
        RECT 20.235 0.065 20.405 0.235 ;
        RECT 20.595 0.065 20.765 0.235 ;
        RECT 20.955 0.065 21.125 0.235 ;
        RECT 21.315 0.065 21.485 0.235 ;
        RECT 21.805 0.065 21.975 0.235 ;
        RECT 22.165 0.065 22.335 0.235 ;
        RECT 22.525 0.065 22.695 0.235 ;
        RECT 22.885 0.065 23.055 0.235 ;
        RECT 23.245 0.065 23.415 0.235 ;
        RECT 23.605 0.065 23.775 0.235 ;
        RECT 24.325 0.065 24.495 0.235 ;
        RECT 24.685 0.065 24.855 0.235 ;
        RECT 25.045 0.065 25.215 0.235 ;
        RECT 25.405 0.065 25.575 0.235 ;
        RECT 25.765 0.065 25.935 0.235 ;
        RECT 26.125 0.065 26.295 0.235 ;
        RECT 26.615 0.065 26.785 0.235 ;
        RECT 26.975 0.065 27.145 0.235 ;
        RECT 27.335 0.065 27.505 0.235 ;
        RECT 27.695 0.065 27.865 0.235 ;
        RECT 28.055 0.065 28.225 0.235 ;
        RECT 28.415 0.065 28.585 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 29.015 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 1.445 5.470 1.615 7.250 ;
        RECT 2.325 5.470 2.495 7.250 ;
        RECT 3.205 5.470 3.375 7.250 ;
        RECT 6.255 5.470 6.425 7.250 ;
        RECT 7.135 5.470 7.305 7.250 ;
        RECT 8.015 5.470 8.185 7.250 ;
        RECT 11.065 5.470 11.235 7.250 ;
        RECT 11.945 5.470 12.115 7.250 ;
        RECT 12.825 5.470 12.995 7.250 ;
        RECT 15.875 5.470 16.045 7.250 ;
        RECT 16.755 5.470 16.925 7.250 ;
        RECT 17.635 5.470 17.805 7.250 ;
        RECT 25.495 5.470 25.665 7.250 ;
        RECT 26.375 5.470 26.545 7.250 ;
        RECT 27.255 5.470 27.425 7.250 ;
        RECT 1.445 5.300 4.155 5.470 ;
        RECT 6.255 5.300 8.965 5.470 ;
        RECT 11.065 5.300 13.775 5.470 ;
        RECT 15.875 5.300 18.585 5.470 ;
        RECT 25.495 5.300 28.205 5.470 ;
        RECT 3.245 2.055 3.415 5.095 ;
        RECT 0.505 1.815 0.675 1.895 ;
        RECT 1.475 1.815 1.645 1.895 ;
        RECT 2.445 1.815 2.615 1.895 ;
        RECT 0.505 1.645 2.615 1.815 ;
        RECT 0.505 0.515 0.675 1.645 ;
        RECT 1.475 0.765 1.645 1.645 ;
        RECT 2.445 1.565 2.615 1.645 ;
        RECT 1.965 1.220 2.135 1.300 ;
        RECT 3.015 1.220 3.185 1.895 ;
        RECT 3.985 1.890 4.155 5.300 ;
        RECT 5.835 2.055 6.005 5.095 ;
        RECT 8.055 4.235 8.225 5.095 ;
        RECT 8.050 3.905 8.225 4.235 ;
        RECT 8.055 2.055 8.225 3.905 ;
        RECT 1.965 1.050 3.185 1.220 ;
        RECT 1.965 0.970 2.135 1.050 ;
        RECT 2.445 0.765 2.615 0.845 ;
        RECT 1.475 0.595 2.615 0.765 ;
        RECT 1.475 0.515 1.645 0.595 ;
        RECT 2.445 0.515 2.615 0.595 ;
        RECT 3.015 0.765 3.185 1.050 ;
        RECT 3.500 1.720 4.155 1.890 ;
        RECT 5.315 1.815 5.485 1.895 ;
        RECT 6.285 1.815 6.455 1.895 ;
        RECT 7.255 1.815 7.425 1.895 ;
        RECT 3.500 0.985 3.670 1.720 ;
        RECT 5.315 1.645 7.425 1.815 ;
        RECT 3.985 0.765 4.155 1.535 ;
        RECT 3.015 0.595 4.155 0.765 ;
        RECT 3.015 0.515 3.185 0.595 ;
        RECT 3.985 0.515 4.155 0.595 ;
        RECT 5.315 0.515 5.485 1.645 ;
        RECT 6.285 0.765 6.455 1.645 ;
        RECT 7.255 1.565 7.425 1.645 ;
        RECT 6.775 1.220 6.945 1.300 ;
        RECT 7.825 1.220 7.995 1.895 ;
        RECT 8.795 1.890 8.965 5.300 ;
        RECT 10.645 2.055 10.815 5.095 ;
        RECT 12.865 2.055 13.035 5.095 ;
        RECT 6.775 1.050 7.995 1.220 ;
        RECT 6.775 0.970 6.945 1.050 ;
        RECT 7.255 0.765 7.425 0.845 ;
        RECT 6.285 0.595 7.425 0.765 ;
        RECT 6.285 0.515 6.455 0.595 ;
        RECT 7.255 0.515 7.425 0.595 ;
        RECT 7.825 0.765 7.995 1.050 ;
        RECT 8.310 1.720 8.965 1.890 ;
        RECT 10.125 1.815 10.295 1.895 ;
        RECT 11.095 1.815 11.265 1.895 ;
        RECT 12.065 1.815 12.235 1.895 ;
        RECT 8.310 0.985 8.480 1.720 ;
        RECT 10.125 1.645 12.235 1.815 ;
        RECT 8.795 0.765 8.965 1.535 ;
        RECT 7.825 0.595 8.965 0.765 ;
        RECT 7.825 0.515 7.995 0.595 ;
        RECT 8.795 0.515 8.965 0.595 ;
        RECT 10.125 0.515 10.295 1.645 ;
        RECT 11.095 0.765 11.265 1.645 ;
        RECT 12.065 1.565 12.235 1.645 ;
        RECT 11.585 1.220 11.755 1.300 ;
        RECT 12.635 1.220 12.805 1.895 ;
        RECT 13.605 1.890 13.775 5.300 ;
        RECT 15.455 2.055 15.625 5.095 ;
        RECT 11.585 1.050 12.805 1.220 ;
        RECT 11.585 0.970 11.755 1.050 ;
        RECT 12.065 0.765 12.235 0.845 ;
        RECT 11.095 0.595 12.235 0.765 ;
        RECT 11.095 0.515 11.265 0.595 ;
        RECT 12.065 0.515 12.235 0.595 ;
        RECT 12.635 0.765 12.805 1.050 ;
        RECT 13.120 1.720 13.775 1.890 ;
        RECT 14.935 1.815 15.105 1.895 ;
        RECT 15.905 1.815 16.075 1.895 ;
        RECT 16.875 1.815 17.045 1.895 ;
        RECT 13.120 0.985 13.290 1.720 ;
        RECT 14.935 1.645 17.045 1.815 ;
        RECT 13.605 0.765 13.775 1.535 ;
        RECT 12.635 0.595 13.775 0.765 ;
        RECT 12.635 0.515 12.805 0.595 ;
        RECT 13.605 0.515 13.775 0.595 ;
        RECT 14.935 0.515 15.105 1.645 ;
        RECT 15.905 0.765 16.075 1.645 ;
        RECT 16.875 1.565 17.045 1.645 ;
        RECT 16.395 1.220 16.565 1.300 ;
        RECT 17.445 1.220 17.615 1.895 ;
        RECT 18.415 1.890 18.585 5.300 ;
        RECT 20.265 2.055 20.435 5.095 ;
        RECT 22.485 2.055 22.655 5.095 ;
        RECT 27.295 2.055 27.465 5.095 ;
        RECT 16.395 1.050 17.615 1.220 ;
        RECT 16.395 0.970 16.565 1.050 ;
        RECT 16.875 0.765 17.045 0.845 ;
        RECT 15.905 0.595 17.045 0.765 ;
        RECT 15.905 0.515 16.075 0.595 ;
        RECT 16.875 0.515 17.045 0.595 ;
        RECT 17.445 0.765 17.615 1.050 ;
        RECT 17.930 1.720 18.585 1.890 ;
        RECT 19.745 1.815 19.915 1.895 ;
        RECT 20.715 1.815 20.885 1.895 ;
        RECT 21.685 1.815 21.855 1.895 ;
        RECT 17.930 0.985 18.100 1.720 ;
        RECT 19.745 1.645 21.855 1.815 ;
        RECT 18.415 0.765 18.585 1.535 ;
        RECT 17.445 0.595 18.585 0.765 ;
        RECT 17.445 0.515 17.615 0.595 ;
        RECT 18.415 0.515 18.585 0.595 ;
        RECT 19.745 0.515 19.915 1.645 ;
        RECT 20.715 0.765 20.885 1.645 ;
        RECT 21.685 1.565 21.855 1.645 ;
        RECT 21.205 1.220 21.375 1.300 ;
        RECT 22.255 1.220 22.425 1.895 ;
        RECT 24.555 1.815 24.725 1.895 ;
        RECT 25.525 1.815 25.695 1.895 ;
        RECT 26.495 1.815 26.665 1.895 ;
        RECT 24.555 1.645 26.665 1.815 ;
        RECT 21.205 1.050 22.425 1.220 ;
        RECT 21.205 0.970 21.375 1.050 ;
        RECT 21.685 0.765 21.855 0.845 ;
        RECT 20.715 0.595 21.855 0.765 ;
        RECT 20.715 0.515 20.885 0.595 ;
        RECT 21.685 0.515 21.855 0.595 ;
        RECT 22.255 0.765 22.425 1.050 ;
        RECT 23.225 0.765 23.395 1.535 ;
        RECT 22.255 0.595 23.395 0.765 ;
        RECT 22.255 0.515 22.425 0.595 ;
        RECT 23.225 0.515 23.395 0.595 ;
        RECT 24.555 0.515 24.725 1.645 ;
        RECT 25.525 0.765 25.695 1.645 ;
        RECT 26.495 1.565 26.665 1.645 ;
        RECT 26.015 1.220 26.185 1.300 ;
        RECT 27.065 1.220 27.235 1.895 ;
        RECT 28.035 1.890 28.205 5.300 ;
        RECT 26.015 1.050 27.235 1.220 ;
        RECT 26.015 0.970 26.185 1.050 ;
        RECT 26.495 0.765 26.665 0.845 ;
        RECT 25.525 0.595 26.665 0.765 ;
        RECT 25.525 0.515 25.695 0.595 ;
        RECT 26.495 0.515 26.665 0.595 ;
        RECT 27.065 0.765 27.235 1.050 ;
        RECT 27.550 1.720 28.205 1.890 ;
        RECT 27.550 0.985 27.720 1.720 ;
        RECT 28.035 0.765 28.205 1.535 ;
        RECT 27.065 0.595 28.205 0.765 ;
        RECT 27.065 0.515 27.235 0.595 ;
        RECT 28.035 0.515 28.205 0.595 ;
      LAYER mcon ;
        RECT 3.245 3.615 3.415 3.785 ;
        RECT 3.985 2.880 4.155 3.050 ;
        RECT 8.050 3.985 8.220 4.155 ;
        RECT 5.835 2.880 6.005 3.050 ;
        RECT 8.795 3.615 8.965 3.785 ;
        RECT 10.645 2.880 10.815 3.050 ;
        RECT 12.865 3.985 13.035 4.155 ;
        RECT 13.605 2.875 13.775 3.045 ;
        RECT 15.455 2.875 15.625 3.045 ;
        RECT 18.415 3.985 18.585 4.155 ;
        RECT 20.265 3.615 20.435 3.785 ;
        RECT 22.485 3.615 22.655 3.785 ;
        RECT 27.295 3.985 27.465 4.155 ;
        RECT 28.035 3.615 28.205 3.785 ;
      LAYER met1 ;
        RECT 8.020 4.155 8.250 4.185 ;
        RECT 12.835 4.155 13.065 4.185 ;
        RECT 18.385 4.155 18.615 4.185 ;
        RECT 27.265 4.155 27.495 4.185 ;
        RECT 7.990 3.985 27.525 4.155 ;
        RECT 8.020 3.955 8.250 3.985 ;
        RECT 12.835 3.955 13.065 3.985 ;
        RECT 18.385 3.955 18.615 3.985 ;
        RECT 27.265 3.955 27.495 3.985 ;
        RECT 3.215 3.785 3.445 3.815 ;
        RECT 8.765 3.785 8.995 3.815 ;
        RECT 20.235 3.785 20.465 3.815 ;
        RECT 22.455 3.785 22.685 3.815 ;
        RECT 28.005 3.785 28.235 3.815 ;
        RECT 3.185 3.615 20.495 3.785 ;
        RECT 22.425 3.615 28.265 3.785 ;
        RECT 3.215 3.585 3.445 3.615 ;
        RECT 8.765 3.585 8.995 3.615 ;
        RECT 20.235 3.585 20.465 3.615 ;
        RECT 22.455 3.585 22.685 3.615 ;
        RECT 28.005 3.585 28.235 3.615 ;
        RECT 3.955 3.050 4.185 3.080 ;
        RECT 5.805 3.050 6.035 3.080 ;
        RECT 10.615 3.050 10.845 3.080 ;
        RECT 3.925 2.880 10.875 3.050 ;
        RECT 13.575 3.045 13.805 3.075 ;
        RECT 15.425 3.045 15.655 3.075 ;
        RECT 3.955 2.850 4.185 2.880 ;
        RECT 5.805 2.850 6.035 2.880 ;
        RECT 10.615 2.850 10.845 2.880 ;
        RECT 13.545 2.875 15.685 3.045 ;
        RECT 13.575 2.845 13.805 2.875 ;
        RECT 15.425 2.845 15.655 2.875 ;
  END
END DFFSNRNQNX1






MACRO DFFSNRNQX1
  CLASS BLOCK ;
  FOREIGN DFFSNRNQX1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 29.700 BY 7.950 ;
  PIN Q
    ANTENNAGATEAREA 1.027250 ;
    ANTENNADIFFAREA 1.931900 ;
    PORT
      LAYER li1 ;
        RECT 25.495 5.470 25.665 7.250 ;
        RECT 26.375 5.470 26.545 7.250 ;
        RECT 27.255 5.470 27.425 7.250 ;
        RECT 25.495 5.300 28.205 5.470 ;
        RECT 22.485 2.055 22.655 5.095 ;
        RECT 28.035 1.890 28.205 5.300 ;
        RECT 27.550 1.720 28.205 1.890 ;
        RECT 27.550 0.985 27.720 1.720 ;
      LAYER mcon ;
        RECT 22.485 3.615 22.655 3.785 ;
        RECT 28.035 3.615 28.205 3.785 ;
      LAYER met1 ;
        RECT 22.455 3.785 22.685 3.815 ;
        RECT 28.005 3.785 28.235 3.815 ;
        RECT 22.425 3.615 28.265 3.785 ;
        RECT 22.455 3.585 22.685 3.615 ;
        RECT 28.005 3.585 28.235 3.615 ;
    END
  END Q
  PIN D
    ANTENNAGATEAREA 1.033250 ;
    PORT
      LAYER li1 ;
        RECT 1.025 2.055 1.195 5.095 ;
      LAYER mcon ;
        RECT 1.025 2.875 1.195 3.045 ;
      LAYER met1 ;
        RECT 0.995 3.045 1.225 3.075 ;
        RECT 0.845 2.875 1.255 3.045 ;
        RECT 0.995 2.845 1.225 2.875 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 2.029700 ;
    PORT
      LAYER li1 ;
        RECT 6.945 2.055 7.115 5.095 ;
        RECT 16.565 2.055 16.735 5.095 ;
      LAYER mcon ;
        RECT 6.945 3.245 7.115 3.415 ;
        RECT 16.565 3.245 16.735 3.415 ;
      LAYER met1 ;
        RECT 6.915 3.415 7.145 3.445 ;
        RECT 16.535 3.415 16.765 3.445 ;
        RECT 6.885 3.245 16.795 3.415 ;
        RECT 6.915 3.215 7.145 3.245 ;
        RECT 16.535 3.215 16.765 3.245 ;
    END
  END CLK
  PIN SN
    ANTENNAGATEAREA 2.029700 ;
    PORT
      LAYER li1 ;
        RECT 11.755 2.055 11.925 5.095 ;
        RECT 26.185 2.055 26.355 5.095 ;
      LAYER mcon ;
        RECT 11.755 2.510 11.925 2.680 ;
        RECT 26.185 2.505 26.355 2.675 ;
      LAYER met1 ;
        RECT 11.725 2.680 11.955 2.710 ;
        RECT 11.695 2.675 12.105 2.680 ;
        RECT 26.155 2.675 26.385 2.705 ;
        RECT 11.695 2.510 26.415 2.675 ;
        RECT 11.725 2.505 26.415 2.510 ;
        RECT 11.725 2.480 11.955 2.505 ;
        RECT 26.155 2.475 26.385 2.505 ;
    END
  END SN
  PIN RN
    ANTENNAGATEAREA 3.056950 ;
    PORT
      LAYER li1 ;
        RECT 2.135 2.055 2.305 5.095 ;
        RECT 17.675 2.055 17.845 5.095 ;
        RECT 21.375 2.055 21.545 5.095 ;
      LAYER mcon ;
        RECT 2.135 4.355 2.305 4.525 ;
        RECT 17.675 4.355 17.845 4.525 ;
        RECT 21.375 4.355 21.545 4.525 ;
      LAYER met1 ;
        RECT 2.105 4.525 2.335 4.555 ;
        RECT 17.645 4.525 17.875 4.555 ;
        RECT 21.345 4.525 21.575 4.555 ;
        RECT 2.075 4.355 21.605 4.525 ;
        RECT 2.105 4.325 2.335 4.355 ;
        RECT 17.645 4.325 17.875 4.355 ;
        RECT 21.345 4.325 21.575 4.355 ;
    END
  END RN
  PIN VDD
    ANTENNADIFFAREA 33.800350 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 29.280 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 29.015 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 1.005 5.445 1.175 7.460 ;
        RECT 1.885 5.785 2.055 7.460 ;
        RECT 2.765 5.785 2.935 7.460 ;
        RECT 3.645 5.785 3.815 7.460 ;
        RECT 4.655 4.340 4.965 7.460 ;
        RECT 5.815 5.445 5.985 7.460 ;
        RECT 6.695 5.785 6.865 7.460 ;
        RECT 7.575 5.785 7.745 7.460 ;
        RECT 8.455 5.785 8.625 7.460 ;
        RECT 9.465 4.340 9.775 7.460 ;
        RECT 10.625 5.445 10.795 7.460 ;
        RECT 11.505 5.785 11.675 7.460 ;
        RECT 12.385 5.785 12.555 7.460 ;
        RECT 13.265 5.785 13.435 7.460 ;
        RECT 14.275 4.340 14.585 7.460 ;
        RECT 15.435 5.445 15.605 7.460 ;
        RECT 16.315 5.785 16.485 7.460 ;
        RECT 17.195 5.785 17.365 7.460 ;
        RECT 18.075 5.785 18.245 7.460 ;
        RECT 19.085 4.340 19.395 7.460 ;
        RECT 20.245 5.445 20.415 7.460 ;
        RECT 21.125 5.785 21.295 7.460 ;
        RECT 22.005 5.785 22.175 7.460 ;
        RECT 22.885 5.785 23.055 7.460 ;
        RECT 23.895 4.340 24.205 7.460 ;
        RECT 25.055 5.445 25.225 7.460 ;
        RECT 25.935 5.785 26.105 7.460 ;
        RECT 26.815 5.785 26.985 7.460 ;
        RECT 27.695 5.785 27.865 7.460 ;
        RECT 28.705 4.340 29.015 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 0.995 7.525 1.165 7.695 ;
        RECT 1.355 7.525 1.525 7.695 ;
        RECT 1.715 7.525 1.885 7.695 ;
        RECT 2.075 7.525 2.245 7.695 ;
        RECT 2.565 7.525 2.735 7.695 ;
        RECT 2.925 7.525 3.095 7.695 ;
        RECT 3.285 7.525 3.455 7.695 ;
        RECT 3.645 7.525 3.815 7.695 ;
        RECT 4.005 7.525 4.175 7.695 ;
        RECT 4.365 7.525 4.535 7.695 ;
        RECT 5.085 7.525 5.255 7.695 ;
        RECT 5.445 7.525 5.615 7.695 ;
        RECT 5.805 7.525 5.975 7.695 ;
        RECT 6.165 7.525 6.335 7.695 ;
        RECT 6.525 7.525 6.695 7.695 ;
        RECT 6.885 7.525 7.055 7.695 ;
        RECT 7.375 7.525 7.545 7.695 ;
        RECT 7.735 7.525 7.905 7.695 ;
        RECT 8.095 7.525 8.265 7.695 ;
        RECT 8.455 7.525 8.625 7.695 ;
        RECT 8.815 7.525 8.985 7.695 ;
        RECT 9.175 7.525 9.345 7.695 ;
        RECT 9.895 7.525 10.065 7.695 ;
        RECT 10.255 7.525 10.425 7.695 ;
        RECT 10.615 7.525 10.785 7.695 ;
        RECT 10.975 7.525 11.145 7.695 ;
        RECT 11.335 7.525 11.505 7.695 ;
        RECT 11.695 7.525 11.865 7.695 ;
        RECT 12.185 7.525 12.355 7.695 ;
        RECT 12.545 7.525 12.715 7.695 ;
        RECT 12.905 7.525 13.075 7.695 ;
        RECT 13.265 7.525 13.435 7.695 ;
        RECT 13.625 7.525 13.795 7.695 ;
        RECT 13.985 7.525 14.155 7.695 ;
        RECT 14.705 7.525 14.875 7.695 ;
        RECT 15.065 7.525 15.235 7.695 ;
        RECT 15.425 7.525 15.595 7.695 ;
        RECT 15.785 7.525 15.955 7.695 ;
        RECT 16.145 7.525 16.315 7.695 ;
        RECT 16.505 7.525 16.675 7.695 ;
        RECT 16.995 7.525 17.165 7.695 ;
        RECT 17.355 7.525 17.525 7.695 ;
        RECT 17.715 7.525 17.885 7.695 ;
        RECT 18.075 7.525 18.245 7.695 ;
        RECT 18.435 7.525 18.605 7.695 ;
        RECT 18.795 7.525 18.965 7.695 ;
        RECT 19.515 7.525 19.685 7.695 ;
        RECT 19.875 7.525 20.045 7.695 ;
        RECT 20.235 7.525 20.405 7.695 ;
        RECT 20.595 7.525 20.765 7.695 ;
        RECT 20.955 7.525 21.125 7.695 ;
        RECT 21.315 7.525 21.485 7.695 ;
        RECT 21.805 7.525 21.975 7.695 ;
        RECT 22.165 7.525 22.335 7.695 ;
        RECT 22.525 7.525 22.695 7.695 ;
        RECT 22.885 7.525 23.055 7.695 ;
        RECT 23.245 7.525 23.415 7.695 ;
        RECT 23.605 7.525 23.775 7.695 ;
        RECT 24.325 7.525 24.495 7.695 ;
        RECT 24.685 7.525 24.855 7.695 ;
        RECT 25.045 7.525 25.215 7.695 ;
        RECT 25.405 7.525 25.575 7.695 ;
        RECT 25.765 7.525 25.935 7.695 ;
        RECT 26.125 7.525 26.295 7.695 ;
        RECT 26.615 7.525 26.785 7.695 ;
        RECT 26.975 7.525 27.145 7.695 ;
        RECT 27.335 7.525 27.505 7.695 ;
        RECT 27.695 7.525 27.865 7.695 ;
        RECT 28.055 7.525 28.225 7.695 ;
        RECT 28.415 7.525 28.585 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 29.015 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 20.198250 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 29.145 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 4.525 -0.075 5.095 -0.065 ;
        RECT 9.335 -0.075 9.905 -0.065 ;
        RECT 14.145 -0.075 14.715 -0.065 ;
        RECT 18.955 -0.075 19.525 -0.065 ;
        RECT 23.765 -0.075 24.335 -0.065 ;
        RECT 28.575 -0.075 29.145 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 0.990 0.310 1.160 1.270 ;
        RECT 4.655 0.310 4.965 2.860 ;
        RECT 5.800 0.310 5.970 1.270 ;
        RECT 9.465 0.310 9.775 2.860 ;
        RECT 10.610 0.310 10.780 1.270 ;
        RECT 14.275 0.310 14.585 2.860 ;
        RECT 15.420 0.310 15.590 1.270 ;
        RECT 19.085 0.310 19.395 2.860 ;
        RECT 20.230 0.310 20.400 1.270 ;
        RECT 23.895 0.310 24.205 2.860 ;
        RECT 25.040 0.310 25.210 1.270 ;
        RECT 28.705 0.310 29.015 2.860 ;
        RECT -0.155 0.000 29.015 0.310 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 0.995 0.065 1.165 0.235 ;
        RECT 1.355 0.065 1.525 0.235 ;
        RECT 1.715 0.065 1.885 0.235 ;
        RECT 2.075 0.065 2.245 0.235 ;
        RECT 2.565 0.065 2.735 0.235 ;
        RECT 2.925 0.065 3.095 0.235 ;
        RECT 3.285 0.065 3.455 0.235 ;
        RECT 3.645 0.065 3.815 0.235 ;
        RECT 4.005 0.065 4.175 0.235 ;
        RECT 4.365 0.065 4.535 0.235 ;
        RECT 5.085 0.065 5.255 0.235 ;
        RECT 5.445 0.065 5.615 0.235 ;
        RECT 5.805 0.065 5.975 0.235 ;
        RECT 6.165 0.065 6.335 0.235 ;
        RECT 6.525 0.065 6.695 0.235 ;
        RECT 6.885 0.065 7.055 0.235 ;
        RECT 7.375 0.065 7.545 0.235 ;
        RECT 7.735 0.065 7.905 0.235 ;
        RECT 8.095 0.065 8.265 0.235 ;
        RECT 8.455 0.065 8.625 0.235 ;
        RECT 8.815 0.065 8.985 0.235 ;
        RECT 9.175 0.065 9.345 0.235 ;
        RECT 9.895 0.065 10.065 0.235 ;
        RECT 10.255 0.065 10.425 0.235 ;
        RECT 10.615 0.065 10.785 0.235 ;
        RECT 10.975 0.065 11.145 0.235 ;
        RECT 11.335 0.065 11.505 0.235 ;
        RECT 11.695 0.065 11.865 0.235 ;
        RECT 12.185 0.065 12.355 0.235 ;
        RECT 12.545 0.065 12.715 0.235 ;
        RECT 12.905 0.065 13.075 0.235 ;
        RECT 13.265 0.065 13.435 0.235 ;
        RECT 13.625 0.065 13.795 0.235 ;
        RECT 13.985 0.065 14.155 0.235 ;
        RECT 14.705 0.065 14.875 0.235 ;
        RECT 15.065 0.065 15.235 0.235 ;
        RECT 15.425 0.065 15.595 0.235 ;
        RECT 15.785 0.065 15.955 0.235 ;
        RECT 16.145 0.065 16.315 0.235 ;
        RECT 16.505 0.065 16.675 0.235 ;
        RECT 16.995 0.065 17.165 0.235 ;
        RECT 17.355 0.065 17.525 0.235 ;
        RECT 17.715 0.065 17.885 0.235 ;
        RECT 18.075 0.065 18.245 0.235 ;
        RECT 18.435 0.065 18.605 0.235 ;
        RECT 18.795 0.065 18.965 0.235 ;
        RECT 19.515 0.065 19.685 0.235 ;
        RECT 19.875 0.065 20.045 0.235 ;
        RECT 20.235 0.065 20.405 0.235 ;
        RECT 20.595 0.065 20.765 0.235 ;
        RECT 20.955 0.065 21.125 0.235 ;
        RECT 21.315 0.065 21.485 0.235 ;
        RECT 21.805 0.065 21.975 0.235 ;
        RECT 22.165 0.065 22.335 0.235 ;
        RECT 22.525 0.065 22.695 0.235 ;
        RECT 22.885 0.065 23.055 0.235 ;
        RECT 23.245 0.065 23.415 0.235 ;
        RECT 23.605 0.065 23.775 0.235 ;
        RECT 24.325 0.065 24.495 0.235 ;
        RECT 24.685 0.065 24.855 0.235 ;
        RECT 25.045 0.065 25.215 0.235 ;
        RECT 25.405 0.065 25.575 0.235 ;
        RECT 25.765 0.065 25.935 0.235 ;
        RECT 26.125 0.065 26.295 0.235 ;
        RECT 26.615 0.065 26.785 0.235 ;
        RECT 26.975 0.065 27.145 0.235 ;
        RECT 27.335 0.065 27.505 0.235 ;
        RECT 27.695 0.065 27.865 0.235 ;
        RECT 28.055 0.065 28.225 0.235 ;
        RECT 28.415 0.065 28.585 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 29.015 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 1.445 5.470 1.615 7.250 ;
        RECT 2.325 5.470 2.495 7.250 ;
        RECT 3.205 5.470 3.375 7.250 ;
        RECT 6.255 5.470 6.425 7.250 ;
        RECT 7.135 5.470 7.305 7.250 ;
        RECT 8.015 5.470 8.185 7.250 ;
        RECT 11.065 5.470 11.235 7.250 ;
        RECT 11.945 5.470 12.115 7.250 ;
        RECT 12.825 5.470 12.995 7.250 ;
        RECT 15.875 5.470 16.045 7.250 ;
        RECT 16.755 5.470 16.925 7.250 ;
        RECT 17.635 5.470 17.805 7.250 ;
        RECT 20.685 5.470 20.855 7.250 ;
        RECT 21.565 5.470 21.735 7.250 ;
        RECT 22.445 5.470 22.615 7.250 ;
        RECT 1.445 5.300 4.155 5.470 ;
        RECT 6.255 5.300 8.965 5.470 ;
        RECT 11.065 5.300 13.775 5.470 ;
        RECT 15.875 5.300 18.585 5.470 ;
        RECT 20.685 5.300 23.395 5.470 ;
        RECT 3.245 2.055 3.415 5.095 ;
        RECT 0.505 1.815 0.675 1.895 ;
        RECT 1.475 1.815 1.645 1.895 ;
        RECT 2.445 1.815 2.615 1.895 ;
        RECT 0.505 1.645 2.615 1.815 ;
        RECT 0.505 0.515 0.675 1.645 ;
        RECT 1.475 0.765 1.645 1.645 ;
        RECT 2.445 1.565 2.615 1.645 ;
        RECT 1.965 1.220 2.135 1.300 ;
        RECT 3.015 1.220 3.185 1.895 ;
        RECT 3.985 1.890 4.155 5.300 ;
        RECT 5.835 2.055 6.005 5.095 ;
        RECT 8.055 4.235 8.225 5.095 ;
        RECT 8.050 3.905 8.225 4.235 ;
        RECT 8.055 2.055 8.225 3.905 ;
        RECT 1.965 1.050 3.185 1.220 ;
        RECT 1.965 0.970 2.135 1.050 ;
        RECT 2.445 0.765 2.615 0.845 ;
        RECT 1.475 0.595 2.615 0.765 ;
        RECT 1.475 0.515 1.645 0.595 ;
        RECT 2.445 0.515 2.615 0.595 ;
        RECT 3.015 0.765 3.185 1.050 ;
        RECT 3.500 1.720 4.155 1.890 ;
        RECT 5.315 1.815 5.485 1.895 ;
        RECT 6.285 1.815 6.455 1.895 ;
        RECT 7.255 1.815 7.425 1.895 ;
        RECT 3.500 0.985 3.670 1.720 ;
        RECT 5.315 1.645 7.425 1.815 ;
        RECT 3.985 0.765 4.155 1.535 ;
        RECT 3.015 0.595 4.155 0.765 ;
        RECT 3.015 0.515 3.185 0.595 ;
        RECT 3.985 0.515 4.155 0.595 ;
        RECT 5.315 0.515 5.485 1.645 ;
        RECT 6.285 0.765 6.455 1.645 ;
        RECT 7.255 1.565 7.425 1.645 ;
        RECT 6.775 1.220 6.945 1.300 ;
        RECT 7.825 1.220 7.995 1.895 ;
        RECT 8.795 1.890 8.965 5.300 ;
        RECT 10.645 2.055 10.815 5.095 ;
        RECT 12.865 2.055 13.035 5.095 ;
        RECT 6.775 1.050 7.995 1.220 ;
        RECT 6.775 0.970 6.945 1.050 ;
        RECT 7.255 0.765 7.425 0.845 ;
        RECT 6.285 0.595 7.425 0.765 ;
        RECT 6.285 0.515 6.455 0.595 ;
        RECT 7.255 0.515 7.425 0.595 ;
        RECT 7.825 0.765 7.995 1.050 ;
        RECT 8.310 1.720 8.965 1.890 ;
        RECT 10.125 1.815 10.295 1.895 ;
        RECT 11.095 1.815 11.265 1.895 ;
        RECT 12.065 1.815 12.235 1.895 ;
        RECT 8.310 0.985 8.480 1.720 ;
        RECT 10.125 1.645 12.235 1.815 ;
        RECT 8.795 0.765 8.965 1.535 ;
        RECT 7.825 0.595 8.965 0.765 ;
        RECT 7.825 0.515 7.995 0.595 ;
        RECT 8.795 0.515 8.965 0.595 ;
        RECT 10.125 0.515 10.295 1.645 ;
        RECT 11.095 0.765 11.265 1.645 ;
        RECT 12.065 1.565 12.235 1.645 ;
        RECT 11.585 1.220 11.755 1.300 ;
        RECT 12.635 1.220 12.805 1.895 ;
        RECT 13.605 1.890 13.775 5.300 ;
        RECT 15.455 2.055 15.625 5.095 ;
        RECT 11.585 1.050 12.805 1.220 ;
        RECT 11.585 0.970 11.755 1.050 ;
        RECT 12.065 0.765 12.235 0.845 ;
        RECT 11.095 0.595 12.235 0.765 ;
        RECT 11.095 0.515 11.265 0.595 ;
        RECT 12.065 0.515 12.235 0.595 ;
        RECT 12.635 0.765 12.805 1.050 ;
        RECT 13.120 1.720 13.775 1.890 ;
        RECT 14.935 1.815 15.105 1.895 ;
        RECT 15.905 1.815 16.075 1.895 ;
        RECT 16.875 1.815 17.045 1.895 ;
        RECT 13.120 0.985 13.290 1.720 ;
        RECT 14.935 1.645 17.045 1.815 ;
        RECT 13.605 0.765 13.775 1.535 ;
        RECT 12.635 0.595 13.775 0.765 ;
        RECT 12.635 0.515 12.805 0.595 ;
        RECT 13.605 0.515 13.775 0.595 ;
        RECT 14.935 0.515 15.105 1.645 ;
        RECT 15.905 0.765 16.075 1.645 ;
        RECT 16.875 1.565 17.045 1.645 ;
        RECT 16.395 1.220 16.565 1.300 ;
        RECT 17.445 1.220 17.615 1.895 ;
        RECT 18.415 1.890 18.585 5.300 ;
        RECT 20.265 2.055 20.435 5.095 ;
        RECT 16.395 1.050 17.615 1.220 ;
        RECT 16.395 0.970 16.565 1.050 ;
        RECT 16.875 0.765 17.045 0.845 ;
        RECT 15.905 0.595 17.045 0.765 ;
        RECT 15.905 0.515 16.075 0.595 ;
        RECT 16.875 0.515 17.045 0.595 ;
        RECT 17.445 0.765 17.615 1.050 ;
        RECT 17.930 1.720 18.585 1.890 ;
        RECT 19.745 1.815 19.915 1.895 ;
        RECT 20.715 1.815 20.885 1.895 ;
        RECT 21.685 1.815 21.855 1.895 ;
        RECT 17.930 0.985 18.100 1.720 ;
        RECT 19.745 1.645 21.855 1.815 ;
        RECT 18.415 0.765 18.585 1.535 ;
        RECT 17.445 0.595 18.585 0.765 ;
        RECT 17.445 0.515 17.615 0.595 ;
        RECT 18.415 0.515 18.585 0.595 ;
        RECT 19.745 0.515 19.915 1.645 ;
        RECT 20.715 0.765 20.885 1.645 ;
        RECT 21.685 1.565 21.855 1.645 ;
        RECT 21.205 1.220 21.375 1.300 ;
        RECT 22.255 1.220 22.425 1.895 ;
        RECT 23.225 1.890 23.395 5.300 ;
        RECT 25.075 2.055 25.245 5.095 ;
        RECT 27.295 2.055 27.465 5.095 ;
        RECT 21.205 1.050 22.425 1.220 ;
        RECT 21.205 0.970 21.375 1.050 ;
        RECT 21.685 0.765 21.855 0.845 ;
        RECT 20.715 0.595 21.855 0.765 ;
        RECT 20.715 0.515 20.885 0.595 ;
        RECT 21.685 0.515 21.855 0.595 ;
        RECT 22.255 0.765 22.425 1.050 ;
        RECT 22.740 1.720 23.395 1.890 ;
        RECT 24.555 1.815 24.725 1.895 ;
        RECT 25.525 1.815 25.695 1.895 ;
        RECT 26.495 1.815 26.665 1.895 ;
        RECT 22.740 0.985 22.910 1.720 ;
        RECT 24.555 1.645 26.665 1.815 ;
        RECT 23.225 0.765 23.395 1.535 ;
        RECT 22.255 0.595 23.395 0.765 ;
        RECT 22.255 0.515 22.425 0.595 ;
        RECT 23.225 0.515 23.395 0.595 ;
        RECT 24.555 0.515 24.725 1.645 ;
        RECT 25.525 0.765 25.695 1.645 ;
        RECT 26.495 1.565 26.665 1.645 ;
        RECT 26.015 1.220 26.185 1.300 ;
        RECT 27.065 1.220 27.235 1.895 ;
        RECT 26.015 1.050 27.235 1.220 ;
        RECT 26.015 0.970 26.185 1.050 ;
        RECT 26.495 0.765 26.665 0.845 ;
        RECT 25.525 0.595 26.665 0.765 ;
        RECT 25.525 0.515 25.695 0.595 ;
        RECT 26.495 0.515 26.665 0.595 ;
        RECT 27.065 0.765 27.235 1.050 ;
        RECT 28.035 0.765 28.205 1.535 ;
        RECT 27.065 0.595 28.205 0.765 ;
        RECT 27.065 0.515 27.235 0.595 ;
        RECT 28.035 0.515 28.205 0.595 ;
      LAYER mcon ;
        RECT 3.245 3.615 3.415 3.785 ;
        RECT 3.985 2.880 4.155 3.050 ;
        RECT 8.050 3.985 8.220 4.155 ;
        RECT 5.835 2.880 6.005 3.050 ;
        RECT 8.795 3.615 8.965 3.785 ;
        RECT 10.645 2.880 10.815 3.050 ;
        RECT 12.865 3.985 13.035 4.155 ;
        RECT 13.605 2.875 13.775 3.045 ;
        RECT 15.455 2.875 15.625 3.045 ;
        RECT 18.415 3.985 18.585 4.155 ;
        RECT 20.265 3.615 20.435 3.785 ;
        RECT 23.225 3.245 23.395 3.415 ;
        RECT 25.075 3.245 25.245 3.415 ;
        RECT 27.295 3.985 27.465 4.155 ;
      LAYER met1 ;
        RECT 8.020 4.155 8.250 4.185 ;
        RECT 12.835 4.155 13.065 4.185 ;
        RECT 18.385 4.155 18.615 4.185 ;
        RECT 27.265 4.155 27.495 4.185 ;
        RECT 7.990 3.985 27.525 4.155 ;
        RECT 8.020 3.955 8.250 3.985 ;
        RECT 12.835 3.955 13.065 3.985 ;
        RECT 18.385 3.955 18.615 3.985 ;
        RECT 27.265 3.955 27.495 3.985 ;
        RECT 3.215 3.785 3.445 3.815 ;
        RECT 8.765 3.785 8.995 3.815 ;
        RECT 20.235 3.785 20.465 3.815 ;
        RECT 3.185 3.615 20.495 3.785 ;
        RECT 3.215 3.585 3.445 3.615 ;
        RECT 8.765 3.585 8.995 3.615 ;
        RECT 20.235 3.585 20.465 3.615 ;
        RECT 23.195 3.415 23.425 3.445 ;
        RECT 25.045 3.415 25.275 3.445 ;
        RECT 23.165 3.245 25.305 3.415 ;
        RECT 23.195 3.215 23.425 3.245 ;
        RECT 25.045 3.215 25.275 3.245 ;
        RECT 3.955 3.050 4.185 3.080 ;
        RECT 5.805 3.050 6.035 3.080 ;
        RECT 10.615 3.050 10.845 3.080 ;
        RECT 3.925 2.880 10.875 3.050 ;
        RECT 13.575 3.045 13.805 3.075 ;
        RECT 15.425 3.045 15.655 3.075 ;
        RECT 3.955 2.850 4.185 2.880 ;
        RECT 5.805 2.850 6.035 2.880 ;
        RECT 10.615 2.850 10.845 2.880 ;
        RECT 13.545 2.875 15.685 3.045 ;
        RECT 13.575 2.845 13.805 2.875 ;
        RECT 15.425 2.845 15.655 2.875 ;
  END
END DFFSNRNQX1






MACRO DFFSNRNX1
  CLASS BLOCK ;
  FOREIGN DFFSNRNX1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 29.700 BY 7.950 ;
  PIN Q
    ANTENNAGATEAREA 1.027250 ;
    ANTENNADIFFAREA 1.931900 ;
    PORT
      LAYER li1 ;
        RECT 25.495 5.470 25.665 7.250 ;
        RECT 26.375 5.470 26.545 7.250 ;
        RECT 27.255 5.470 27.425 7.250 ;
        RECT 25.495 5.300 28.205 5.470 ;
        RECT 22.485 2.055 22.655 5.095 ;
        RECT 28.035 1.890 28.205 5.300 ;
        RECT 27.550 1.720 28.205 1.890 ;
        RECT 27.550 0.985 27.720 1.720 ;
      LAYER mcon ;
        RECT 22.485 3.615 22.655 3.785 ;
        RECT 28.035 3.615 28.205 3.785 ;
      LAYER met1 ;
        RECT 22.455 3.785 22.685 3.815 ;
        RECT 28.005 3.785 28.235 3.815 ;
        RECT 22.425 3.615 28.265 3.785 ;
        RECT 22.455 3.585 22.685 3.615 ;
        RECT 28.005 3.585 28.235 3.615 ;
    END
  END Q
  PIN QN
    ANTENNAGATEAREA 1.033250 ;
    ANTENNADIFFAREA 1.931900 ;
    PORT
      LAYER li1 ;
        RECT 20.685 5.470 20.855 7.250 ;
        RECT 21.565 5.470 21.735 7.250 ;
        RECT 22.445 5.470 22.615 7.250 ;
        RECT 20.685 5.300 23.395 5.470 ;
        RECT 23.225 1.890 23.395 5.300 ;
        RECT 25.075 2.055 25.245 5.095 ;
        RECT 22.740 1.720 23.395 1.890 ;
        RECT 22.740 0.985 22.910 1.720 ;
      LAYER mcon ;
        RECT 23.225 3.245 23.395 3.415 ;
        RECT 25.075 3.245 25.245 3.415 ;
      LAYER met1 ;
        RECT 23.195 3.415 23.425 3.445 ;
        RECT 25.045 3.415 25.275 3.445 ;
        RECT 23.165 3.245 25.305 3.415 ;
        RECT 23.195 3.215 23.425 3.245 ;
        RECT 25.045 3.215 25.275 3.245 ;
    END
  END QN
  PIN D
    ANTENNAGATEAREA 1.033250 ;
    PORT
      LAYER li1 ;
        RECT 1.025 2.055 1.195 5.095 ;
      LAYER mcon ;
        RECT 1.025 2.875 1.195 3.045 ;
      LAYER met1 ;
        RECT 0.995 3.045 1.225 3.075 ;
        RECT 0.845 2.875 1.255 3.045 ;
        RECT 0.995 2.845 1.225 2.875 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 2.029700 ;
    PORT
      LAYER li1 ;
        RECT 6.945 2.055 7.115 5.095 ;
        RECT 16.565 2.055 16.735 5.095 ;
      LAYER mcon ;
        RECT 6.945 3.245 7.115 3.415 ;
        RECT 16.565 3.245 16.735 3.415 ;
      LAYER met1 ;
        RECT 6.915 3.415 7.145 3.445 ;
        RECT 16.535 3.415 16.765 3.445 ;
        RECT 6.885 3.245 16.795 3.415 ;
        RECT 6.915 3.215 7.145 3.245 ;
        RECT 16.535 3.215 16.765 3.245 ;
    END
  END CLK
  PIN SN
    ANTENNAGATEAREA 2.029700 ;
    PORT
      LAYER li1 ;
        RECT 11.755 2.055 11.925 5.095 ;
        RECT 26.185 2.055 26.355 5.095 ;
      LAYER mcon ;
        RECT 11.755 2.510 11.925 2.680 ;
        RECT 26.185 2.505 26.355 2.675 ;
      LAYER met1 ;
        RECT 11.725 2.680 11.955 2.710 ;
        RECT 11.695 2.675 12.105 2.680 ;
        RECT 26.155 2.675 26.385 2.705 ;
        RECT 11.695 2.510 26.415 2.675 ;
        RECT 11.725 2.505 26.415 2.510 ;
        RECT 11.725 2.480 11.955 2.505 ;
        RECT 26.155 2.475 26.385 2.505 ;
    END
  END SN
  PIN RN
    ANTENNAGATEAREA 3.056950 ;
    PORT
      LAYER li1 ;
        RECT 2.135 2.055 2.305 5.095 ;
        RECT 17.675 2.055 17.845 5.095 ;
        RECT 21.375 2.055 21.545 5.095 ;
      LAYER mcon ;
        RECT 2.135 4.355 2.305 4.525 ;
        RECT 17.675 4.355 17.845 4.525 ;
        RECT 21.375 4.355 21.545 4.525 ;
      LAYER met1 ;
        RECT 2.105 4.525 2.335 4.555 ;
        RECT 17.645 4.525 17.875 4.555 ;
        RECT 21.345 4.525 21.575 4.555 ;
        RECT 2.075 4.355 21.605 4.525 ;
        RECT 2.105 4.325 2.335 4.355 ;
        RECT 17.645 4.325 17.875 4.355 ;
        RECT 21.345 4.325 21.575 4.355 ;
    END
  END RN
  PIN VDD
    ANTENNADIFFAREA 33.800350 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 29.280 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 29.015 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 1.005 5.445 1.175 7.460 ;
        RECT 1.885 5.785 2.055 7.460 ;
        RECT 2.765 5.785 2.935 7.460 ;
        RECT 3.645 5.785 3.815 7.460 ;
        RECT 4.655 4.340 4.965 7.460 ;
        RECT 5.815 5.445 5.985 7.460 ;
        RECT 6.695 5.785 6.865 7.460 ;
        RECT 7.575 5.785 7.745 7.460 ;
        RECT 8.455 5.785 8.625 7.460 ;
        RECT 9.465 4.340 9.775 7.460 ;
        RECT 10.625 5.445 10.795 7.460 ;
        RECT 11.505 5.785 11.675 7.460 ;
        RECT 12.385 5.785 12.555 7.460 ;
        RECT 13.265 5.785 13.435 7.460 ;
        RECT 14.275 4.340 14.585 7.460 ;
        RECT 15.435 5.445 15.605 7.460 ;
        RECT 16.315 5.785 16.485 7.460 ;
        RECT 17.195 5.785 17.365 7.460 ;
        RECT 18.075 5.785 18.245 7.460 ;
        RECT 19.085 4.340 19.395 7.460 ;
        RECT 20.245 5.445 20.415 7.460 ;
        RECT 21.125 5.785 21.295 7.460 ;
        RECT 22.005 5.785 22.175 7.460 ;
        RECT 22.885 5.785 23.055 7.460 ;
        RECT 23.895 4.340 24.205 7.460 ;
        RECT 25.055 5.445 25.225 7.460 ;
        RECT 25.935 5.785 26.105 7.460 ;
        RECT 26.815 5.785 26.985 7.460 ;
        RECT 27.695 5.785 27.865 7.460 ;
        RECT 28.705 4.340 29.015 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 0.995 7.525 1.165 7.695 ;
        RECT 1.355 7.525 1.525 7.695 ;
        RECT 1.715 7.525 1.885 7.695 ;
        RECT 2.075 7.525 2.245 7.695 ;
        RECT 2.565 7.525 2.735 7.695 ;
        RECT 2.925 7.525 3.095 7.695 ;
        RECT 3.285 7.525 3.455 7.695 ;
        RECT 3.645 7.525 3.815 7.695 ;
        RECT 4.005 7.525 4.175 7.695 ;
        RECT 4.365 7.525 4.535 7.695 ;
        RECT 5.085 7.525 5.255 7.695 ;
        RECT 5.445 7.525 5.615 7.695 ;
        RECT 5.805 7.525 5.975 7.695 ;
        RECT 6.165 7.525 6.335 7.695 ;
        RECT 6.525 7.525 6.695 7.695 ;
        RECT 6.885 7.525 7.055 7.695 ;
        RECT 7.375 7.525 7.545 7.695 ;
        RECT 7.735 7.525 7.905 7.695 ;
        RECT 8.095 7.525 8.265 7.695 ;
        RECT 8.455 7.525 8.625 7.695 ;
        RECT 8.815 7.525 8.985 7.695 ;
        RECT 9.175 7.525 9.345 7.695 ;
        RECT 9.895 7.525 10.065 7.695 ;
        RECT 10.255 7.525 10.425 7.695 ;
        RECT 10.615 7.525 10.785 7.695 ;
        RECT 10.975 7.525 11.145 7.695 ;
        RECT 11.335 7.525 11.505 7.695 ;
        RECT 11.695 7.525 11.865 7.695 ;
        RECT 12.185 7.525 12.355 7.695 ;
        RECT 12.545 7.525 12.715 7.695 ;
        RECT 12.905 7.525 13.075 7.695 ;
        RECT 13.265 7.525 13.435 7.695 ;
        RECT 13.625 7.525 13.795 7.695 ;
        RECT 13.985 7.525 14.155 7.695 ;
        RECT 14.705 7.525 14.875 7.695 ;
        RECT 15.065 7.525 15.235 7.695 ;
        RECT 15.425 7.525 15.595 7.695 ;
        RECT 15.785 7.525 15.955 7.695 ;
        RECT 16.145 7.525 16.315 7.695 ;
        RECT 16.505 7.525 16.675 7.695 ;
        RECT 16.995 7.525 17.165 7.695 ;
        RECT 17.355 7.525 17.525 7.695 ;
        RECT 17.715 7.525 17.885 7.695 ;
        RECT 18.075 7.525 18.245 7.695 ;
        RECT 18.435 7.525 18.605 7.695 ;
        RECT 18.795 7.525 18.965 7.695 ;
        RECT 19.515 7.525 19.685 7.695 ;
        RECT 19.875 7.525 20.045 7.695 ;
        RECT 20.235 7.525 20.405 7.695 ;
        RECT 20.595 7.525 20.765 7.695 ;
        RECT 20.955 7.525 21.125 7.695 ;
        RECT 21.315 7.525 21.485 7.695 ;
        RECT 21.805 7.525 21.975 7.695 ;
        RECT 22.165 7.525 22.335 7.695 ;
        RECT 22.525 7.525 22.695 7.695 ;
        RECT 22.885 7.525 23.055 7.695 ;
        RECT 23.245 7.525 23.415 7.695 ;
        RECT 23.605 7.525 23.775 7.695 ;
        RECT 24.325 7.525 24.495 7.695 ;
        RECT 24.685 7.525 24.855 7.695 ;
        RECT 25.045 7.525 25.215 7.695 ;
        RECT 25.405 7.525 25.575 7.695 ;
        RECT 25.765 7.525 25.935 7.695 ;
        RECT 26.125 7.525 26.295 7.695 ;
        RECT 26.615 7.525 26.785 7.695 ;
        RECT 26.975 7.525 27.145 7.695 ;
        RECT 27.335 7.525 27.505 7.695 ;
        RECT 27.695 7.525 27.865 7.695 ;
        RECT 28.055 7.525 28.225 7.695 ;
        RECT 28.415 7.525 28.585 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 29.015 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 20.198250 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 29.145 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 4.525 -0.075 5.095 -0.065 ;
        RECT 9.335 -0.075 9.905 -0.065 ;
        RECT 14.145 -0.075 14.715 -0.065 ;
        RECT 18.955 -0.075 19.525 -0.065 ;
        RECT 23.765 -0.075 24.335 -0.065 ;
        RECT 28.575 -0.075 29.145 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 0.990 0.310 1.160 1.270 ;
        RECT 4.655 0.310 4.965 2.860 ;
        RECT 5.800 0.310 5.970 1.270 ;
        RECT 9.465 0.310 9.775 2.860 ;
        RECT 10.610 0.310 10.780 1.270 ;
        RECT 14.275 0.310 14.585 2.860 ;
        RECT 15.420 0.310 15.590 1.270 ;
        RECT 19.085 0.310 19.395 2.860 ;
        RECT 20.230 0.310 20.400 1.270 ;
        RECT 23.895 0.310 24.205 2.860 ;
        RECT 25.040 0.310 25.210 1.270 ;
        RECT 28.705 0.310 29.015 2.860 ;
        RECT -0.155 0.000 29.015 0.310 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 0.995 0.065 1.165 0.235 ;
        RECT 1.355 0.065 1.525 0.235 ;
        RECT 1.715 0.065 1.885 0.235 ;
        RECT 2.075 0.065 2.245 0.235 ;
        RECT 2.565 0.065 2.735 0.235 ;
        RECT 2.925 0.065 3.095 0.235 ;
        RECT 3.285 0.065 3.455 0.235 ;
        RECT 3.645 0.065 3.815 0.235 ;
        RECT 4.005 0.065 4.175 0.235 ;
        RECT 4.365 0.065 4.535 0.235 ;
        RECT 5.085 0.065 5.255 0.235 ;
        RECT 5.445 0.065 5.615 0.235 ;
        RECT 5.805 0.065 5.975 0.235 ;
        RECT 6.165 0.065 6.335 0.235 ;
        RECT 6.525 0.065 6.695 0.235 ;
        RECT 6.885 0.065 7.055 0.235 ;
        RECT 7.375 0.065 7.545 0.235 ;
        RECT 7.735 0.065 7.905 0.235 ;
        RECT 8.095 0.065 8.265 0.235 ;
        RECT 8.455 0.065 8.625 0.235 ;
        RECT 8.815 0.065 8.985 0.235 ;
        RECT 9.175 0.065 9.345 0.235 ;
        RECT 9.895 0.065 10.065 0.235 ;
        RECT 10.255 0.065 10.425 0.235 ;
        RECT 10.615 0.065 10.785 0.235 ;
        RECT 10.975 0.065 11.145 0.235 ;
        RECT 11.335 0.065 11.505 0.235 ;
        RECT 11.695 0.065 11.865 0.235 ;
        RECT 12.185 0.065 12.355 0.235 ;
        RECT 12.545 0.065 12.715 0.235 ;
        RECT 12.905 0.065 13.075 0.235 ;
        RECT 13.265 0.065 13.435 0.235 ;
        RECT 13.625 0.065 13.795 0.235 ;
        RECT 13.985 0.065 14.155 0.235 ;
        RECT 14.705 0.065 14.875 0.235 ;
        RECT 15.065 0.065 15.235 0.235 ;
        RECT 15.425 0.065 15.595 0.235 ;
        RECT 15.785 0.065 15.955 0.235 ;
        RECT 16.145 0.065 16.315 0.235 ;
        RECT 16.505 0.065 16.675 0.235 ;
        RECT 16.995 0.065 17.165 0.235 ;
        RECT 17.355 0.065 17.525 0.235 ;
        RECT 17.715 0.065 17.885 0.235 ;
        RECT 18.075 0.065 18.245 0.235 ;
        RECT 18.435 0.065 18.605 0.235 ;
        RECT 18.795 0.065 18.965 0.235 ;
        RECT 19.515 0.065 19.685 0.235 ;
        RECT 19.875 0.065 20.045 0.235 ;
        RECT 20.235 0.065 20.405 0.235 ;
        RECT 20.595 0.065 20.765 0.235 ;
        RECT 20.955 0.065 21.125 0.235 ;
        RECT 21.315 0.065 21.485 0.235 ;
        RECT 21.805 0.065 21.975 0.235 ;
        RECT 22.165 0.065 22.335 0.235 ;
        RECT 22.525 0.065 22.695 0.235 ;
        RECT 22.885 0.065 23.055 0.235 ;
        RECT 23.245 0.065 23.415 0.235 ;
        RECT 23.605 0.065 23.775 0.235 ;
        RECT 24.325 0.065 24.495 0.235 ;
        RECT 24.685 0.065 24.855 0.235 ;
        RECT 25.045 0.065 25.215 0.235 ;
        RECT 25.405 0.065 25.575 0.235 ;
        RECT 25.765 0.065 25.935 0.235 ;
        RECT 26.125 0.065 26.295 0.235 ;
        RECT 26.615 0.065 26.785 0.235 ;
        RECT 26.975 0.065 27.145 0.235 ;
        RECT 27.335 0.065 27.505 0.235 ;
        RECT 27.695 0.065 27.865 0.235 ;
        RECT 28.055 0.065 28.225 0.235 ;
        RECT 28.415 0.065 28.585 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 29.015 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 1.445 5.470 1.615 7.250 ;
        RECT 2.325 5.470 2.495 7.250 ;
        RECT 3.205 5.470 3.375 7.250 ;
        RECT 6.255 5.470 6.425 7.250 ;
        RECT 7.135 5.470 7.305 7.250 ;
        RECT 8.015 5.470 8.185 7.250 ;
        RECT 11.065 5.470 11.235 7.250 ;
        RECT 11.945 5.470 12.115 7.250 ;
        RECT 12.825 5.470 12.995 7.250 ;
        RECT 15.875 5.470 16.045 7.250 ;
        RECT 16.755 5.470 16.925 7.250 ;
        RECT 17.635 5.470 17.805 7.250 ;
        RECT 1.445 5.300 4.155 5.470 ;
        RECT 6.255 5.300 8.965 5.470 ;
        RECT 11.065 5.300 13.775 5.470 ;
        RECT 15.875 5.300 18.585 5.470 ;
        RECT 3.245 2.055 3.415 5.095 ;
        RECT 0.505 1.815 0.675 1.895 ;
        RECT 1.475 1.815 1.645 1.895 ;
        RECT 2.445 1.815 2.615 1.895 ;
        RECT 0.505 1.645 2.615 1.815 ;
        RECT 0.505 0.515 0.675 1.645 ;
        RECT 1.475 0.765 1.645 1.645 ;
        RECT 2.445 1.565 2.615 1.645 ;
        RECT 1.965 1.220 2.135 1.300 ;
        RECT 3.015 1.220 3.185 1.895 ;
        RECT 3.985 1.890 4.155 5.300 ;
        RECT 5.835 2.055 6.005 5.095 ;
        RECT 8.055 4.235 8.225 5.095 ;
        RECT 8.050 3.905 8.225 4.235 ;
        RECT 8.055 2.055 8.225 3.905 ;
        RECT 1.965 1.050 3.185 1.220 ;
        RECT 1.965 0.970 2.135 1.050 ;
        RECT 2.445 0.765 2.615 0.845 ;
        RECT 1.475 0.595 2.615 0.765 ;
        RECT 1.475 0.515 1.645 0.595 ;
        RECT 2.445 0.515 2.615 0.595 ;
        RECT 3.015 0.765 3.185 1.050 ;
        RECT 3.500 1.720 4.155 1.890 ;
        RECT 5.315 1.815 5.485 1.895 ;
        RECT 6.285 1.815 6.455 1.895 ;
        RECT 7.255 1.815 7.425 1.895 ;
        RECT 3.500 0.985 3.670 1.720 ;
        RECT 5.315 1.645 7.425 1.815 ;
        RECT 3.985 0.765 4.155 1.535 ;
        RECT 3.015 0.595 4.155 0.765 ;
        RECT 3.015 0.515 3.185 0.595 ;
        RECT 3.985 0.515 4.155 0.595 ;
        RECT 5.315 0.515 5.485 1.645 ;
        RECT 6.285 0.765 6.455 1.645 ;
        RECT 7.255 1.565 7.425 1.645 ;
        RECT 6.775 1.220 6.945 1.300 ;
        RECT 7.825 1.220 7.995 1.895 ;
        RECT 8.795 1.890 8.965 5.300 ;
        RECT 10.645 2.055 10.815 5.095 ;
        RECT 12.865 2.055 13.035 5.095 ;
        RECT 6.775 1.050 7.995 1.220 ;
        RECT 6.775 0.970 6.945 1.050 ;
        RECT 7.255 0.765 7.425 0.845 ;
        RECT 6.285 0.595 7.425 0.765 ;
        RECT 6.285 0.515 6.455 0.595 ;
        RECT 7.255 0.515 7.425 0.595 ;
        RECT 7.825 0.765 7.995 1.050 ;
        RECT 8.310 1.720 8.965 1.890 ;
        RECT 10.125 1.815 10.295 1.895 ;
        RECT 11.095 1.815 11.265 1.895 ;
        RECT 12.065 1.815 12.235 1.895 ;
        RECT 8.310 0.985 8.480 1.720 ;
        RECT 10.125 1.645 12.235 1.815 ;
        RECT 8.795 0.765 8.965 1.535 ;
        RECT 7.825 0.595 8.965 0.765 ;
        RECT 7.825 0.515 7.995 0.595 ;
        RECT 8.795 0.515 8.965 0.595 ;
        RECT 10.125 0.515 10.295 1.645 ;
        RECT 11.095 0.765 11.265 1.645 ;
        RECT 12.065 1.565 12.235 1.645 ;
        RECT 11.585 1.220 11.755 1.300 ;
        RECT 12.635 1.220 12.805 1.895 ;
        RECT 13.605 1.890 13.775 5.300 ;
        RECT 15.455 2.055 15.625 5.095 ;
        RECT 11.585 1.050 12.805 1.220 ;
        RECT 11.585 0.970 11.755 1.050 ;
        RECT 12.065 0.765 12.235 0.845 ;
        RECT 11.095 0.595 12.235 0.765 ;
        RECT 11.095 0.515 11.265 0.595 ;
        RECT 12.065 0.515 12.235 0.595 ;
        RECT 12.635 0.765 12.805 1.050 ;
        RECT 13.120 1.720 13.775 1.890 ;
        RECT 14.935 1.815 15.105 1.895 ;
        RECT 15.905 1.815 16.075 1.895 ;
        RECT 16.875 1.815 17.045 1.895 ;
        RECT 13.120 0.985 13.290 1.720 ;
        RECT 14.935 1.645 17.045 1.815 ;
        RECT 13.605 0.765 13.775 1.535 ;
        RECT 12.635 0.595 13.775 0.765 ;
        RECT 12.635 0.515 12.805 0.595 ;
        RECT 13.605 0.515 13.775 0.595 ;
        RECT 14.935 0.515 15.105 1.645 ;
        RECT 15.905 0.765 16.075 1.645 ;
        RECT 16.875 1.565 17.045 1.645 ;
        RECT 16.395 1.220 16.565 1.300 ;
        RECT 17.445 1.220 17.615 1.895 ;
        RECT 18.415 1.890 18.585 5.300 ;
        RECT 20.265 2.055 20.435 5.095 ;
        RECT 27.295 2.055 27.465 5.095 ;
        RECT 16.395 1.050 17.615 1.220 ;
        RECT 16.395 0.970 16.565 1.050 ;
        RECT 16.875 0.765 17.045 0.845 ;
        RECT 15.905 0.595 17.045 0.765 ;
        RECT 15.905 0.515 16.075 0.595 ;
        RECT 16.875 0.515 17.045 0.595 ;
        RECT 17.445 0.765 17.615 1.050 ;
        RECT 17.930 1.720 18.585 1.890 ;
        RECT 19.745 1.815 19.915 1.895 ;
        RECT 20.715 1.815 20.885 1.895 ;
        RECT 21.685 1.815 21.855 1.895 ;
        RECT 17.930 0.985 18.100 1.720 ;
        RECT 19.745 1.645 21.855 1.815 ;
        RECT 18.415 0.765 18.585 1.535 ;
        RECT 17.445 0.595 18.585 0.765 ;
        RECT 17.445 0.515 17.615 0.595 ;
        RECT 18.415 0.515 18.585 0.595 ;
        RECT 19.745 0.515 19.915 1.645 ;
        RECT 20.715 0.765 20.885 1.645 ;
        RECT 21.685 1.565 21.855 1.645 ;
        RECT 21.205 1.220 21.375 1.300 ;
        RECT 22.255 1.220 22.425 1.895 ;
        RECT 24.555 1.815 24.725 1.895 ;
        RECT 25.525 1.815 25.695 1.895 ;
        RECT 26.495 1.815 26.665 1.895 ;
        RECT 24.555 1.645 26.665 1.815 ;
        RECT 21.205 1.050 22.425 1.220 ;
        RECT 21.205 0.970 21.375 1.050 ;
        RECT 21.685 0.765 21.855 0.845 ;
        RECT 20.715 0.595 21.855 0.765 ;
        RECT 20.715 0.515 20.885 0.595 ;
        RECT 21.685 0.515 21.855 0.595 ;
        RECT 22.255 0.765 22.425 1.050 ;
        RECT 23.225 0.765 23.395 1.535 ;
        RECT 22.255 0.595 23.395 0.765 ;
        RECT 22.255 0.515 22.425 0.595 ;
        RECT 23.225 0.515 23.395 0.595 ;
        RECT 24.555 0.515 24.725 1.645 ;
        RECT 25.525 0.765 25.695 1.645 ;
        RECT 26.495 1.565 26.665 1.645 ;
        RECT 26.015 1.220 26.185 1.300 ;
        RECT 27.065 1.220 27.235 1.895 ;
        RECT 26.015 1.050 27.235 1.220 ;
        RECT 26.015 0.970 26.185 1.050 ;
        RECT 26.495 0.765 26.665 0.845 ;
        RECT 25.525 0.595 26.665 0.765 ;
        RECT 25.525 0.515 25.695 0.595 ;
        RECT 26.495 0.515 26.665 0.595 ;
        RECT 27.065 0.765 27.235 1.050 ;
        RECT 28.035 0.765 28.205 1.535 ;
        RECT 27.065 0.595 28.205 0.765 ;
        RECT 27.065 0.515 27.235 0.595 ;
        RECT 28.035 0.515 28.205 0.595 ;
      LAYER mcon ;
        RECT 3.245 3.615 3.415 3.785 ;
        RECT 3.985 2.880 4.155 3.050 ;
        RECT 8.050 3.985 8.220 4.155 ;
        RECT 5.835 2.880 6.005 3.050 ;
        RECT 8.795 3.615 8.965 3.785 ;
        RECT 10.645 2.880 10.815 3.050 ;
        RECT 12.865 3.985 13.035 4.155 ;
        RECT 13.605 2.875 13.775 3.045 ;
        RECT 15.455 2.875 15.625 3.045 ;
        RECT 18.415 3.985 18.585 4.155 ;
        RECT 20.265 3.615 20.435 3.785 ;
        RECT 27.295 3.985 27.465 4.155 ;
      LAYER met1 ;
        RECT 8.020 4.155 8.250 4.185 ;
        RECT 12.835 4.155 13.065 4.185 ;
        RECT 18.385 4.155 18.615 4.185 ;
        RECT 27.265 4.155 27.495 4.185 ;
        RECT 7.990 3.985 27.525 4.155 ;
        RECT 8.020 3.955 8.250 3.985 ;
        RECT 12.835 3.955 13.065 3.985 ;
        RECT 18.385 3.955 18.615 3.985 ;
        RECT 27.265 3.955 27.495 3.985 ;
        RECT 3.215 3.785 3.445 3.815 ;
        RECT 8.765 3.785 8.995 3.815 ;
        RECT 20.235 3.785 20.465 3.815 ;
        RECT 3.185 3.615 20.495 3.785 ;
        RECT 3.215 3.585 3.445 3.615 ;
        RECT 8.765 3.585 8.995 3.615 ;
        RECT 20.235 3.585 20.465 3.615 ;
        RECT 3.955 3.050 4.185 3.080 ;
        RECT 5.805 3.050 6.035 3.080 ;
        RECT 10.615 3.050 10.845 3.080 ;
        RECT 3.925 2.880 10.875 3.050 ;
        RECT 13.575 3.045 13.805 3.075 ;
        RECT 15.425 3.045 15.655 3.075 ;
        RECT 3.955 2.850 4.185 2.880 ;
        RECT 5.805 2.850 6.035 2.880 ;
        RECT 10.615 2.850 10.845 2.880 ;
        RECT 13.545 2.875 15.685 3.045 ;
        RECT 13.575 2.845 13.805 2.875 ;
        RECT 15.425 2.845 15.655 2.875 ;
  END
END DFFSNRNX1






MACRO DFFSNX1
  CLASS BLOCK ;
  FOREIGN DFFSNX1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 25.260 BY 7.950 ;
  PIN Q
    ANTENNAGATEAREA 1.027250 ;
    ANTENNADIFFAREA 1.931900 ;
    PORT
      LAYER li1 ;
        RECT 21.055 5.470 21.225 7.250 ;
        RECT 21.935 5.470 22.105 7.250 ;
        RECT 22.815 5.470 22.985 7.250 ;
        RECT 21.055 5.300 23.765 5.470 ;
        RECT 18.075 4.940 18.245 5.095 ;
        RECT 18.045 4.765 18.245 4.940 ;
        RECT 18.045 2.055 18.215 4.765 ;
        RECT 23.595 1.890 23.765 5.300 ;
        RECT 23.110 1.720 23.765 1.890 ;
        RECT 23.110 0.985 23.280 1.720 ;
      LAYER mcon ;
        RECT 18.045 3.615 18.215 3.785 ;
        RECT 23.595 3.615 23.765 3.785 ;
      LAYER met1 ;
        RECT 18.015 3.785 18.245 3.815 ;
        RECT 23.565 3.785 23.795 3.815 ;
        RECT 17.985 3.615 23.825 3.785 ;
        RECT 18.015 3.585 18.245 3.615 ;
        RECT 23.565 3.585 23.795 3.615 ;
    END
  END Q
  PIN QN
    ANTENNAGATEAREA 1.033250 ;
    ANTENNADIFFAREA 1.351900 ;
    PORT
      LAYER li1 ;
        RECT 17.425 5.515 17.595 7.250 ;
        RECT 18.305 5.515 18.475 7.250 ;
        RECT 17.425 5.345 18.955 5.515 ;
        RECT 18.785 1.880 18.955 5.345 ;
        RECT 20.635 2.055 20.805 5.095 ;
        RECT 18.345 1.710 18.955 1.880 ;
        RECT 18.345 0.975 18.515 1.710 ;
      LAYER mcon ;
        RECT 18.785 3.245 18.955 3.415 ;
        RECT 20.635 3.245 20.805 3.415 ;
      LAYER met1 ;
        RECT 18.755 3.415 18.985 3.445 ;
        RECT 20.605 3.415 20.835 3.445 ;
        RECT 18.725 3.245 20.865 3.415 ;
        RECT 18.755 3.215 18.985 3.245 ;
        RECT 20.605 3.215 20.835 3.245 ;
    END
  END QN
  PIN D
    ANTENNAGATEAREA 1.033250 ;
    PORT
      LAYER li1 ;
        RECT 1.025 2.055 1.195 5.095 ;
      LAYER mcon ;
        RECT 1.025 3.985 1.195 4.155 ;
      LAYER met1 ;
        RECT 0.995 4.155 1.225 4.185 ;
        RECT 0.845 3.985 1.255 4.155 ;
        RECT 0.995 3.955 1.225 3.985 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 2.042100 ;
    PORT
      LAYER li1 ;
        RECT 5.465 2.055 5.635 5.095 ;
        RECT 14.745 4.975 14.915 5.095 ;
        RECT 14.715 4.765 14.915 4.975 ;
        RECT 14.715 2.055 14.885 4.765 ;
      LAYER mcon ;
        RECT 5.465 4.725 5.635 4.895 ;
        RECT 14.715 4.725 14.885 4.895 ;
      LAYER met1 ;
        RECT 5.435 4.895 5.665 4.925 ;
        RECT 14.685 4.895 14.915 4.925 ;
        RECT 5.405 4.725 14.945 4.895 ;
        RECT 5.435 4.695 5.665 4.725 ;
        RECT 14.685 4.695 14.915 4.725 ;
    END
  END CLK
  PIN SN
    ANTENNAGATEAREA 2.029700 ;
    PORT
      LAYER li1 ;
        RECT 10.275 2.055 10.445 5.095 ;
        RECT 21.745 2.055 21.915 5.095 ;
      LAYER mcon ;
        RECT 10.275 2.505 10.445 2.675 ;
        RECT 21.745 2.505 21.915 2.675 ;
      LAYER met1 ;
        RECT 10.245 2.675 10.475 2.705 ;
        RECT 21.715 2.675 21.945 2.705 ;
        RECT 10.215 2.505 21.975 2.675 ;
        RECT 10.245 2.475 10.475 2.505 ;
        RECT 21.715 2.475 21.945 2.505 ;
    END
  END SN
  PIN VDD
    ANTENNADIFFAREA 29.929150 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 24.840 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 24.575 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 0.705 5.365 0.875 7.460 ;
        RECT 1.585 5.785 1.755 7.460 ;
        RECT 2.465 5.785 2.635 7.460 ;
        RECT 3.175 4.340 3.485 7.460 ;
        RECT 4.335 5.445 4.505 7.460 ;
        RECT 5.215 5.785 5.385 7.460 ;
        RECT 6.095 5.785 6.265 7.460 ;
        RECT 6.975 5.785 7.145 7.460 ;
        RECT 7.985 4.340 8.295 7.460 ;
        RECT 9.145 5.445 9.315 7.460 ;
        RECT 10.025 5.785 10.195 7.460 ;
        RECT 10.905 5.785 11.075 7.460 ;
        RECT 11.785 5.785 11.955 7.460 ;
        RECT 12.795 4.340 13.105 7.460 ;
        RECT 13.655 5.365 13.825 7.460 ;
        RECT 14.535 5.785 14.705 7.460 ;
        RECT 15.415 5.785 15.585 7.460 ;
        RECT 16.125 4.340 16.435 7.460 ;
        RECT 16.985 5.365 17.155 7.460 ;
        RECT 17.865 5.785 18.035 7.460 ;
        RECT 18.745 5.785 18.915 7.460 ;
        RECT 19.455 4.340 19.765 7.460 ;
        RECT 20.615 5.445 20.785 7.460 ;
        RECT 21.495 5.785 21.665 7.460 ;
        RECT 22.375 5.785 22.545 7.460 ;
        RECT 23.255 5.785 23.425 7.460 ;
        RECT 24.265 4.340 24.575 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 0.995 7.525 1.165 7.695 ;
        RECT 1.355 7.525 1.525 7.695 ;
        RECT 1.805 7.525 1.975 7.695 ;
        RECT 2.165 7.525 2.335 7.695 ;
        RECT 2.525 7.525 2.695 7.695 ;
        RECT 2.885 7.525 3.055 7.695 ;
        RECT 3.605 7.525 3.775 7.695 ;
        RECT 3.965 7.525 4.135 7.695 ;
        RECT 4.325 7.525 4.495 7.695 ;
        RECT 4.685 7.525 4.855 7.695 ;
        RECT 5.045 7.525 5.215 7.695 ;
        RECT 5.405 7.525 5.575 7.695 ;
        RECT 5.895 7.525 6.065 7.695 ;
        RECT 6.255 7.525 6.425 7.695 ;
        RECT 6.615 7.525 6.785 7.695 ;
        RECT 6.975 7.525 7.145 7.695 ;
        RECT 7.335 7.525 7.505 7.695 ;
        RECT 7.695 7.525 7.865 7.695 ;
        RECT 8.415 7.525 8.585 7.695 ;
        RECT 8.775 7.525 8.945 7.695 ;
        RECT 9.135 7.525 9.305 7.695 ;
        RECT 9.495 7.525 9.665 7.695 ;
        RECT 9.855 7.525 10.025 7.695 ;
        RECT 10.215 7.525 10.385 7.695 ;
        RECT 10.705 7.525 10.875 7.695 ;
        RECT 11.065 7.525 11.235 7.695 ;
        RECT 11.425 7.525 11.595 7.695 ;
        RECT 11.785 7.525 11.955 7.695 ;
        RECT 12.145 7.525 12.315 7.695 ;
        RECT 12.505 7.525 12.675 7.695 ;
        RECT 13.225 7.525 13.395 7.695 ;
        RECT 13.585 7.525 13.755 7.695 ;
        RECT 13.945 7.525 14.115 7.695 ;
        RECT 14.305 7.525 14.475 7.695 ;
        RECT 14.755 7.525 14.925 7.695 ;
        RECT 15.115 7.525 15.285 7.695 ;
        RECT 15.475 7.525 15.645 7.695 ;
        RECT 15.835 7.525 16.005 7.695 ;
        RECT 16.555 7.525 16.725 7.695 ;
        RECT 16.915 7.525 17.085 7.695 ;
        RECT 17.275 7.525 17.445 7.695 ;
        RECT 17.635 7.525 17.805 7.695 ;
        RECT 18.085 7.525 18.255 7.695 ;
        RECT 18.445 7.525 18.615 7.695 ;
        RECT 18.805 7.525 18.975 7.695 ;
        RECT 19.165 7.525 19.335 7.695 ;
        RECT 19.885 7.525 20.055 7.695 ;
        RECT 20.245 7.525 20.415 7.695 ;
        RECT 20.605 7.525 20.775 7.695 ;
        RECT 20.965 7.525 21.135 7.695 ;
        RECT 21.325 7.525 21.495 7.695 ;
        RECT 21.685 7.525 21.855 7.695 ;
        RECT 22.175 7.525 22.345 7.695 ;
        RECT 22.535 7.525 22.705 7.695 ;
        RECT 22.895 7.525 23.065 7.695 ;
        RECT 23.255 7.525 23.425 7.695 ;
        RECT 23.615 7.525 23.785 7.695 ;
        RECT 23.975 7.525 24.145 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 24.575 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 18.067049 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 24.705 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 3.045 -0.075 3.615 -0.065 ;
        RECT 7.855 -0.075 8.425 -0.065 ;
        RECT 12.665 -0.075 13.235 -0.065 ;
        RECT 15.995 -0.075 16.565 -0.065 ;
        RECT 19.325 -0.075 19.895 -0.065 ;
        RECT 24.135 -0.075 24.705 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 1.095 0.310 1.265 1.260 ;
        RECT 3.175 0.310 3.485 2.860 ;
        RECT 4.320 0.310 4.490 1.270 ;
        RECT 7.985 0.310 8.295 2.860 ;
        RECT 9.130 0.310 9.300 1.270 ;
        RECT 12.795 0.310 13.105 2.860 ;
        RECT 14.045 0.310 14.215 1.260 ;
        RECT 16.125 0.310 16.435 2.860 ;
        RECT 17.375 0.310 17.545 1.260 ;
        RECT 19.455 0.310 19.765 2.860 ;
        RECT 20.600 0.310 20.770 1.270 ;
        RECT 24.265 0.310 24.575 2.860 ;
        RECT -0.155 0.000 24.575 0.310 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 0.995 0.065 1.165 0.235 ;
        RECT 1.355 0.065 1.525 0.235 ;
        RECT 1.805 0.065 1.975 0.235 ;
        RECT 2.165 0.065 2.335 0.235 ;
        RECT 2.525 0.065 2.695 0.235 ;
        RECT 2.885 0.065 3.055 0.235 ;
        RECT 3.605 0.065 3.775 0.235 ;
        RECT 3.965 0.065 4.135 0.235 ;
        RECT 4.325 0.065 4.495 0.235 ;
        RECT 4.685 0.065 4.855 0.235 ;
        RECT 5.045 0.065 5.215 0.235 ;
        RECT 5.405 0.065 5.575 0.235 ;
        RECT 5.895 0.065 6.065 0.235 ;
        RECT 6.255 0.065 6.425 0.235 ;
        RECT 6.615 0.065 6.785 0.235 ;
        RECT 6.975 0.065 7.145 0.235 ;
        RECT 7.335 0.065 7.505 0.235 ;
        RECT 7.695 0.065 7.865 0.235 ;
        RECT 8.415 0.065 8.585 0.235 ;
        RECT 8.775 0.065 8.945 0.235 ;
        RECT 9.135 0.065 9.305 0.235 ;
        RECT 9.495 0.065 9.665 0.235 ;
        RECT 9.855 0.065 10.025 0.235 ;
        RECT 10.215 0.065 10.385 0.235 ;
        RECT 10.705 0.065 10.875 0.235 ;
        RECT 11.065 0.065 11.235 0.235 ;
        RECT 11.425 0.065 11.595 0.235 ;
        RECT 11.785 0.065 11.955 0.235 ;
        RECT 12.145 0.065 12.315 0.235 ;
        RECT 12.505 0.065 12.675 0.235 ;
        RECT 13.225 0.065 13.395 0.235 ;
        RECT 13.585 0.065 13.755 0.235 ;
        RECT 13.945 0.065 14.115 0.235 ;
        RECT 14.305 0.065 14.475 0.235 ;
        RECT 14.755 0.065 14.925 0.235 ;
        RECT 15.115 0.065 15.285 0.235 ;
        RECT 15.475 0.065 15.645 0.235 ;
        RECT 15.835 0.065 16.005 0.235 ;
        RECT 16.555 0.065 16.725 0.235 ;
        RECT 16.915 0.065 17.085 0.235 ;
        RECT 17.275 0.065 17.445 0.235 ;
        RECT 17.635 0.065 17.805 0.235 ;
        RECT 18.085 0.065 18.255 0.235 ;
        RECT 18.445 0.065 18.615 0.235 ;
        RECT 18.805 0.065 18.975 0.235 ;
        RECT 19.165 0.065 19.335 0.235 ;
        RECT 19.885 0.065 20.055 0.235 ;
        RECT 20.245 0.065 20.415 0.235 ;
        RECT 20.605 0.065 20.775 0.235 ;
        RECT 20.965 0.065 21.135 0.235 ;
        RECT 21.325 0.065 21.495 0.235 ;
        RECT 21.685 0.065 21.855 0.235 ;
        RECT 22.175 0.065 22.345 0.235 ;
        RECT 22.535 0.065 22.705 0.235 ;
        RECT 22.895 0.065 23.065 0.235 ;
        RECT 23.255 0.065 23.425 0.235 ;
        RECT 23.615 0.065 23.785 0.235 ;
        RECT 23.975 0.065 24.145 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 24.575 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 1.145 5.515 1.315 7.250 ;
        RECT 2.025 5.515 2.195 7.250 ;
        RECT 1.145 5.345 2.675 5.515 ;
        RECT 1.795 4.940 1.965 5.095 ;
        RECT 1.765 4.765 1.965 4.940 ;
        RECT 1.765 2.055 1.935 4.765 ;
        RECT 0.610 1.805 0.780 1.885 ;
        RECT 1.580 1.805 1.750 1.885 ;
        RECT 2.505 1.880 2.675 5.345 ;
        RECT 4.775 5.470 4.945 7.250 ;
        RECT 5.655 5.470 5.825 7.250 ;
        RECT 6.535 5.470 6.705 7.250 ;
        RECT 9.585 5.470 9.755 7.250 ;
        RECT 10.465 5.470 10.635 7.250 ;
        RECT 11.345 5.470 11.515 7.250 ;
        RECT 14.095 5.515 14.265 7.250 ;
        RECT 14.975 5.515 15.145 7.250 ;
        RECT 4.775 5.300 7.485 5.470 ;
        RECT 9.585 5.300 12.295 5.470 ;
        RECT 14.095 5.345 15.625 5.515 ;
        RECT 4.355 2.055 4.525 5.095 ;
        RECT 6.575 2.055 6.745 5.095 ;
        RECT 7.315 4.605 7.485 5.300 ;
        RECT 7.310 4.275 7.485 4.605 ;
        RECT 0.610 1.635 1.750 1.805 ;
        RECT 0.610 0.505 0.780 1.635 ;
        RECT 1.580 0.755 1.750 1.635 ;
        RECT 2.065 1.710 2.675 1.880 ;
        RECT 3.835 1.815 4.005 1.895 ;
        RECT 4.805 1.815 4.975 1.895 ;
        RECT 5.775 1.815 5.945 1.895 ;
        RECT 2.065 0.975 2.235 1.710 ;
        RECT 3.835 1.645 5.945 1.815 ;
        RECT 2.550 0.755 2.720 1.525 ;
        RECT 1.580 0.585 2.720 0.755 ;
        RECT 1.580 0.505 1.750 0.585 ;
        RECT 2.550 0.505 2.720 0.585 ;
        RECT 3.835 0.515 4.005 1.645 ;
        RECT 4.805 0.765 4.975 1.645 ;
        RECT 5.775 1.565 5.945 1.645 ;
        RECT 5.295 1.220 5.465 1.300 ;
        RECT 6.345 1.220 6.515 1.895 ;
        RECT 7.315 1.890 7.485 4.275 ;
        RECT 9.165 2.055 9.335 5.095 ;
        RECT 11.385 2.055 11.555 5.095 ;
        RECT 5.295 1.050 6.515 1.220 ;
        RECT 5.295 0.970 5.465 1.050 ;
        RECT 5.775 0.765 5.945 0.845 ;
        RECT 4.805 0.595 5.945 0.765 ;
        RECT 4.805 0.515 4.975 0.595 ;
        RECT 5.775 0.515 5.945 0.595 ;
        RECT 6.345 0.765 6.515 1.050 ;
        RECT 6.830 1.720 7.485 1.890 ;
        RECT 8.645 1.815 8.815 1.895 ;
        RECT 9.615 1.815 9.785 1.895 ;
        RECT 10.585 1.815 10.755 1.895 ;
        RECT 6.830 0.985 7.000 1.720 ;
        RECT 8.645 1.645 10.755 1.815 ;
        RECT 7.315 0.765 7.485 1.535 ;
        RECT 6.345 0.595 7.485 0.765 ;
        RECT 6.345 0.515 6.515 0.595 ;
        RECT 7.315 0.515 7.485 0.595 ;
        RECT 8.645 0.515 8.815 1.645 ;
        RECT 9.615 0.765 9.785 1.645 ;
        RECT 10.585 1.565 10.755 1.645 ;
        RECT 10.105 1.220 10.275 1.300 ;
        RECT 11.155 1.220 11.325 1.895 ;
        RECT 12.125 1.890 12.295 5.300 ;
        RECT 13.975 2.055 14.145 5.095 ;
        RECT 10.105 1.050 11.325 1.220 ;
        RECT 10.105 0.970 10.275 1.050 ;
        RECT 10.585 0.765 10.755 0.845 ;
        RECT 9.615 0.595 10.755 0.765 ;
        RECT 9.615 0.515 9.785 0.595 ;
        RECT 10.585 0.515 10.755 0.595 ;
        RECT 11.155 0.765 11.325 1.050 ;
        RECT 11.640 1.720 12.295 1.890 ;
        RECT 13.560 1.805 13.730 1.885 ;
        RECT 14.530 1.805 14.700 1.885 ;
        RECT 15.455 1.880 15.625 5.345 ;
        RECT 17.305 2.055 17.475 5.095 ;
        RECT 22.855 2.055 23.025 5.095 ;
        RECT 11.640 0.985 11.810 1.720 ;
        RECT 13.560 1.635 14.700 1.805 ;
        RECT 12.125 0.765 12.295 1.535 ;
        RECT 11.155 0.595 12.295 0.765 ;
        RECT 11.155 0.515 11.325 0.595 ;
        RECT 12.125 0.515 12.295 0.595 ;
        RECT 13.560 0.505 13.730 1.635 ;
        RECT 14.530 0.755 14.700 1.635 ;
        RECT 15.015 1.710 15.625 1.880 ;
        RECT 16.890 1.805 17.060 1.885 ;
        RECT 17.860 1.805 18.030 1.885 ;
        RECT 15.015 0.975 15.185 1.710 ;
        RECT 16.890 1.635 18.030 1.805 ;
        RECT 15.500 0.755 15.670 1.525 ;
        RECT 14.530 0.585 15.670 0.755 ;
        RECT 14.530 0.505 14.700 0.585 ;
        RECT 15.500 0.505 15.670 0.585 ;
        RECT 16.890 0.505 17.060 1.635 ;
        RECT 17.860 0.755 18.030 1.635 ;
        RECT 20.115 1.815 20.285 1.895 ;
        RECT 21.085 1.815 21.255 1.895 ;
        RECT 22.055 1.815 22.225 1.895 ;
        RECT 20.115 1.645 22.225 1.815 ;
        RECT 18.830 0.755 19.000 1.525 ;
        RECT 17.860 0.585 19.000 0.755 ;
        RECT 17.860 0.505 18.030 0.585 ;
        RECT 18.830 0.505 19.000 0.585 ;
        RECT 20.115 0.515 20.285 1.645 ;
        RECT 21.085 0.765 21.255 1.645 ;
        RECT 22.055 1.565 22.225 1.645 ;
        RECT 21.575 1.220 21.745 1.300 ;
        RECT 22.625 1.220 22.795 1.895 ;
        RECT 21.575 1.050 22.795 1.220 ;
        RECT 21.575 0.970 21.745 1.050 ;
        RECT 22.055 0.765 22.225 0.845 ;
        RECT 21.085 0.595 22.225 0.765 ;
        RECT 21.085 0.515 21.255 0.595 ;
        RECT 22.055 0.515 22.225 0.595 ;
        RECT 22.625 0.765 22.795 1.050 ;
        RECT 23.595 0.765 23.765 1.535 ;
        RECT 22.625 0.595 23.765 0.765 ;
        RECT 22.625 0.515 22.795 0.595 ;
        RECT 23.595 0.515 23.765 0.595 ;
      LAYER mcon ;
        RECT 1.765 4.355 1.935 4.525 ;
        RECT 2.505 2.875 2.675 3.045 ;
        RECT 4.355 2.870 4.525 3.040 ;
        RECT 7.310 4.355 7.480 4.525 ;
        RECT 6.575 3.985 6.745 4.155 ;
        RECT 9.165 2.875 9.335 3.045 ;
        RECT 11.385 3.985 11.555 4.155 ;
        RECT 12.125 2.875 12.295 3.045 ;
        RECT 13.975 2.875 14.145 3.045 ;
        RECT 15.455 3.985 15.625 4.155 ;
        RECT 17.305 4.355 17.475 4.525 ;
        RECT 22.855 3.985 23.025 4.155 ;
      LAYER met1 ;
        RECT 1.735 4.525 1.965 4.555 ;
        RECT 7.280 4.525 7.510 4.555 ;
        RECT 17.275 4.525 17.505 4.555 ;
        RECT 1.705 4.355 17.535 4.525 ;
        RECT 1.735 4.325 1.965 4.355 ;
        RECT 7.280 4.325 7.510 4.355 ;
        RECT 17.275 4.325 17.505 4.355 ;
        RECT 6.545 4.155 6.775 4.185 ;
        RECT 11.355 4.155 11.585 4.185 ;
        RECT 15.425 4.155 15.655 4.185 ;
        RECT 22.825 4.155 23.055 4.185 ;
        RECT 6.515 3.985 23.085 4.155 ;
        RECT 6.545 3.955 6.775 3.985 ;
        RECT 11.355 3.955 11.585 3.985 ;
        RECT 15.425 3.955 15.655 3.985 ;
        RECT 22.825 3.955 23.055 3.985 ;
        RECT 2.475 3.045 2.705 3.075 ;
        RECT 4.325 3.045 4.555 3.070 ;
        RECT 9.135 3.045 9.365 3.075 ;
        RECT 12.095 3.045 12.325 3.075 ;
        RECT 13.945 3.045 14.175 3.075 ;
        RECT 2.445 2.875 9.395 3.045 ;
        RECT 12.065 2.875 14.205 3.045 ;
        RECT 2.475 2.845 2.705 2.875 ;
        RECT 4.295 2.870 4.705 2.875 ;
        RECT 4.325 2.840 4.555 2.870 ;
        RECT 9.135 2.845 9.365 2.875 ;
        RECT 12.095 2.845 12.325 2.875 ;
        RECT 13.945 2.845 14.175 2.875 ;
  END
END DFFSNX1






MACRO DFFX1
  CLASS BLOCK ;
  FOREIGN DFFX1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 22.300 BY 7.950 ;
  PIN Q
    ANTENNAGATEAREA 1.027250 ;
    ANTENNADIFFAREA 1.351900 ;
    PORT
      LAYER li1 ;
        RECT 19.275 5.515 19.445 7.250 ;
        RECT 20.155 5.515 20.325 7.250 ;
        RECT 19.275 5.345 20.805 5.515 ;
        RECT 16.595 4.940 16.765 5.095 ;
        RECT 16.565 4.765 16.765 4.940 ;
        RECT 16.565 2.055 16.735 4.765 ;
        RECT 20.635 1.880 20.805 5.345 ;
        RECT 20.195 1.710 20.805 1.880 ;
        RECT 20.195 0.975 20.365 1.710 ;
      LAYER mcon ;
        RECT 16.565 3.985 16.735 4.155 ;
        RECT 20.635 3.985 20.805 4.155 ;
      LAYER met1 ;
        RECT 16.535 4.155 16.765 4.185 ;
        RECT 20.605 4.155 20.835 4.185 ;
        RECT 16.505 3.985 20.865 4.155 ;
        RECT 16.535 3.955 16.765 3.985 ;
        RECT 20.605 3.955 20.835 3.985 ;
    END
  END Q
  PIN QN
    ANTENNAGATEAREA 1.033250 ;
    ANTENNADIFFAREA 1.351900 ;
    PORT
      LAYER li1 ;
        RECT 15.945 5.515 16.115 7.250 ;
        RECT 16.825 5.515 16.995 7.250 ;
        RECT 15.945 5.345 17.475 5.515 ;
        RECT 17.305 1.880 17.475 5.345 ;
        RECT 19.155 2.055 19.325 5.095 ;
        RECT 16.865 1.710 17.475 1.880 ;
        RECT 16.865 0.975 17.035 1.710 ;
      LAYER mcon ;
        RECT 17.305 3.615 17.475 3.785 ;
        RECT 19.155 3.615 19.325 3.785 ;
      LAYER met1 ;
        RECT 17.275 3.785 17.505 3.815 ;
        RECT 19.125 3.785 19.355 3.815 ;
        RECT 17.245 3.615 19.385 3.785 ;
        RECT 17.275 3.585 17.505 3.615 ;
        RECT 19.125 3.585 19.355 3.615 ;
    END
  END QN
  PIN D
    ANTENNAGATEAREA 1.027250 ;
    PORT
      LAYER li1 ;
        RECT 6.605 4.940 6.775 5.095 ;
        RECT 6.575 4.765 6.775 4.940 ;
        RECT 6.575 2.055 6.745 4.765 ;
      LAYER mcon ;
        RECT 6.575 3.245 6.745 3.415 ;
        RECT 6.575 2.135 6.745 2.305 ;
      LAYER met1 ;
        RECT 6.545 3.415 6.775 3.445 ;
        RECT 6.395 3.245 6.805 3.415 ;
        RECT 6.545 3.215 6.775 3.245 ;
        RECT 6.545 2.305 6.775 2.335 ;
        RECT 6.395 2.135 6.805 2.305 ;
        RECT 6.545 2.105 6.775 2.135 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 2.042100 ;
    PORT
      LAYER li1 ;
        RECT 2.135 2.055 2.305 5.095 ;
        RECT 13.265 4.975 13.435 5.095 ;
        RECT 13.235 4.765 13.435 4.975 ;
        RECT 13.235 2.055 13.405 4.765 ;
      LAYER mcon ;
        RECT 2.135 4.725 2.305 4.895 ;
        RECT 13.235 4.725 13.405 4.895 ;
      LAYER met1 ;
        RECT 2.105 4.895 2.335 4.925 ;
        RECT 13.205 4.895 13.435 4.925 ;
        RECT 2.075 4.725 13.465 4.895 ;
        RECT 2.105 4.695 2.335 4.725 ;
        RECT 13.205 4.695 13.435 4.725 ;
    END
  END CLK
  PIN VDD
    ANTENNADIFFAREA 27.348349 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 21.880 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 21.615 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 1.005 5.445 1.175 7.460 ;
        RECT 1.885 5.785 2.055 7.460 ;
        RECT 2.765 5.785 2.935 7.460 ;
        RECT 3.645 5.785 3.815 7.460 ;
        RECT 4.655 4.340 4.965 7.460 ;
        RECT 5.515 5.365 5.685 7.460 ;
        RECT 6.395 5.785 6.565 7.460 ;
        RECT 7.275 5.785 7.445 7.460 ;
        RECT 7.985 4.340 8.295 7.460 ;
        RECT 8.845 5.365 9.015 7.460 ;
        RECT 9.725 5.785 9.895 7.460 ;
        RECT 10.605 5.785 10.775 7.460 ;
        RECT 11.315 4.340 11.625 7.460 ;
        RECT 12.175 5.365 12.345 7.460 ;
        RECT 13.055 5.785 13.225 7.460 ;
        RECT 13.935 5.785 14.105 7.460 ;
        RECT 14.645 4.340 14.955 7.460 ;
        RECT 15.505 5.365 15.675 7.460 ;
        RECT 16.385 5.785 16.555 7.460 ;
        RECT 17.265 5.785 17.435 7.460 ;
        RECT 17.975 4.340 18.285 7.460 ;
        RECT 18.835 5.365 19.005 7.460 ;
        RECT 19.715 5.785 19.885 7.460 ;
        RECT 20.595 5.785 20.765 7.460 ;
        RECT 21.305 4.340 21.615 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 0.995 7.525 1.165 7.695 ;
        RECT 1.355 7.525 1.525 7.695 ;
        RECT 1.715 7.525 1.885 7.695 ;
        RECT 2.075 7.525 2.245 7.695 ;
        RECT 2.565 7.525 2.735 7.695 ;
        RECT 2.925 7.525 3.095 7.695 ;
        RECT 3.285 7.525 3.455 7.695 ;
        RECT 3.645 7.525 3.815 7.695 ;
        RECT 4.005 7.525 4.175 7.695 ;
        RECT 4.365 7.525 4.535 7.695 ;
        RECT 5.085 7.525 5.255 7.695 ;
        RECT 5.445 7.525 5.615 7.695 ;
        RECT 5.805 7.525 5.975 7.695 ;
        RECT 6.165 7.525 6.335 7.695 ;
        RECT 6.615 7.525 6.785 7.695 ;
        RECT 6.975 7.525 7.145 7.695 ;
        RECT 7.335 7.525 7.505 7.695 ;
        RECT 7.695 7.525 7.865 7.695 ;
        RECT 8.415 7.525 8.585 7.695 ;
        RECT 8.775 7.525 8.945 7.695 ;
        RECT 9.135 7.525 9.305 7.695 ;
        RECT 9.495 7.525 9.665 7.695 ;
        RECT 9.945 7.525 10.115 7.695 ;
        RECT 10.305 7.525 10.475 7.695 ;
        RECT 10.665 7.525 10.835 7.695 ;
        RECT 11.025 7.525 11.195 7.695 ;
        RECT 11.745 7.525 11.915 7.695 ;
        RECT 12.105 7.525 12.275 7.695 ;
        RECT 12.465 7.525 12.635 7.695 ;
        RECT 12.825 7.525 12.995 7.695 ;
        RECT 13.275 7.525 13.445 7.695 ;
        RECT 13.635 7.525 13.805 7.695 ;
        RECT 13.995 7.525 14.165 7.695 ;
        RECT 14.355 7.525 14.525 7.695 ;
        RECT 15.075 7.525 15.245 7.695 ;
        RECT 15.435 7.525 15.605 7.695 ;
        RECT 15.795 7.525 15.965 7.695 ;
        RECT 16.155 7.525 16.325 7.695 ;
        RECT 16.605 7.525 16.775 7.695 ;
        RECT 16.965 7.525 17.135 7.695 ;
        RECT 17.325 7.525 17.495 7.695 ;
        RECT 17.685 7.525 17.855 7.695 ;
        RECT 18.405 7.525 18.575 7.695 ;
        RECT 18.765 7.525 18.935 7.695 ;
        RECT 19.125 7.525 19.295 7.695 ;
        RECT 19.485 7.525 19.655 7.695 ;
        RECT 19.935 7.525 20.105 7.695 ;
        RECT 20.295 7.525 20.465 7.695 ;
        RECT 20.655 7.525 20.825 7.695 ;
        RECT 21.015 7.525 21.185 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 21.615 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 16.646250 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 21.745 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 4.525 -0.075 5.095 -0.065 ;
        RECT 7.855 -0.075 8.425 -0.065 ;
        RECT 11.185 -0.075 11.755 -0.065 ;
        RECT 14.515 -0.075 15.085 -0.065 ;
        RECT 17.845 -0.075 18.415 -0.065 ;
        RECT 21.175 -0.075 21.745 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 0.990 0.310 1.160 1.270 ;
        RECT 4.655 0.310 4.965 2.860 ;
        RECT 5.905 0.310 6.075 1.260 ;
        RECT 7.985 0.310 8.295 2.860 ;
        RECT 9.235 0.310 9.405 1.260 ;
        RECT 11.315 0.310 11.625 2.860 ;
        RECT 12.565 0.310 12.735 1.260 ;
        RECT 14.645 0.310 14.955 2.860 ;
        RECT 15.895 0.310 16.065 1.260 ;
        RECT 17.975 0.310 18.285 2.860 ;
        RECT 19.225 0.310 19.395 1.260 ;
        RECT 21.305 0.310 21.615 2.860 ;
        RECT -0.155 0.000 21.615 0.310 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 0.995 0.065 1.165 0.235 ;
        RECT 1.355 0.065 1.525 0.235 ;
        RECT 1.715 0.065 1.885 0.235 ;
        RECT 2.075 0.065 2.245 0.235 ;
        RECT 2.565 0.065 2.735 0.235 ;
        RECT 2.925 0.065 3.095 0.235 ;
        RECT 3.285 0.065 3.455 0.235 ;
        RECT 3.645 0.065 3.815 0.235 ;
        RECT 4.005 0.065 4.175 0.235 ;
        RECT 4.365 0.065 4.535 0.235 ;
        RECT 5.085 0.065 5.255 0.235 ;
        RECT 5.445 0.065 5.615 0.235 ;
        RECT 5.805 0.065 5.975 0.235 ;
        RECT 6.165 0.065 6.335 0.235 ;
        RECT 6.615 0.065 6.785 0.235 ;
        RECT 6.975 0.065 7.145 0.235 ;
        RECT 7.335 0.065 7.505 0.235 ;
        RECT 7.695 0.065 7.865 0.235 ;
        RECT 8.415 0.065 8.585 0.235 ;
        RECT 8.775 0.065 8.945 0.235 ;
        RECT 9.135 0.065 9.305 0.235 ;
        RECT 9.495 0.065 9.665 0.235 ;
        RECT 9.945 0.065 10.115 0.235 ;
        RECT 10.305 0.065 10.475 0.235 ;
        RECT 10.665 0.065 10.835 0.235 ;
        RECT 11.025 0.065 11.195 0.235 ;
        RECT 11.745 0.065 11.915 0.235 ;
        RECT 12.105 0.065 12.275 0.235 ;
        RECT 12.465 0.065 12.635 0.235 ;
        RECT 12.825 0.065 12.995 0.235 ;
        RECT 13.275 0.065 13.445 0.235 ;
        RECT 13.635 0.065 13.805 0.235 ;
        RECT 13.995 0.065 14.165 0.235 ;
        RECT 14.355 0.065 14.525 0.235 ;
        RECT 15.075 0.065 15.245 0.235 ;
        RECT 15.435 0.065 15.605 0.235 ;
        RECT 15.795 0.065 15.965 0.235 ;
        RECT 16.155 0.065 16.325 0.235 ;
        RECT 16.605 0.065 16.775 0.235 ;
        RECT 16.965 0.065 17.135 0.235 ;
        RECT 17.325 0.065 17.495 0.235 ;
        RECT 17.685 0.065 17.855 0.235 ;
        RECT 18.405 0.065 18.575 0.235 ;
        RECT 18.765 0.065 18.935 0.235 ;
        RECT 19.125 0.065 19.295 0.235 ;
        RECT 19.485 0.065 19.655 0.235 ;
        RECT 19.935 0.065 20.105 0.235 ;
        RECT 20.295 0.065 20.465 0.235 ;
        RECT 20.655 0.065 20.825 0.235 ;
        RECT 21.015 0.065 21.185 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 21.615 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 1.445 5.470 1.615 7.250 ;
        RECT 2.325 5.470 2.495 7.250 ;
        RECT 3.205 5.470 3.375 7.250 ;
        RECT 5.955 5.515 6.125 7.250 ;
        RECT 6.835 5.515 7.005 7.250 ;
        RECT 9.285 5.515 9.455 7.250 ;
        RECT 10.165 5.515 10.335 7.250 ;
        RECT 12.615 5.515 12.785 7.250 ;
        RECT 13.495 5.515 13.665 7.250 ;
        RECT 1.445 5.300 4.155 5.470 ;
        RECT 5.955 5.345 7.485 5.515 ;
        RECT 9.285 5.345 10.815 5.515 ;
        RECT 12.615 5.345 14.145 5.515 ;
        RECT 1.025 2.055 1.195 5.095 ;
        RECT 3.245 2.055 3.415 5.095 ;
        RECT 0.505 1.815 0.675 1.895 ;
        RECT 1.475 1.815 1.645 1.895 ;
        RECT 2.445 1.815 2.615 1.895 ;
        RECT 0.505 1.645 2.615 1.815 ;
        RECT 0.505 0.515 0.675 1.645 ;
        RECT 1.475 0.765 1.645 1.645 ;
        RECT 2.445 1.565 2.615 1.645 ;
        RECT 1.965 1.220 2.135 1.300 ;
        RECT 3.015 1.220 3.185 1.895 ;
        RECT 3.985 1.890 4.155 5.300 ;
        RECT 5.835 2.055 6.005 5.095 ;
        RECT 1.965 1.050 3.185 1.220 ;
        RECT 1.965 0.970 2.135 1.050 ;
        RECT 2.445 0.765 2.615 0.845 ;
        RECT 1.475 0.595 2.615 0.765 ;
        RECT 1.475 0.515 1.645 0.595 ;
        RECT 2.445 0.515 2.615 0.595 ;
        RECT 3.015 0.765 3.185 1.050 ;
        RECT 3.500 1.720 4.155 1.890 ;
        RECT 5.420 1.805 5.590 1.885 ;
        RECT 6.390 1.805 6.560 1.885 ;
        RECT 7.315 1.880 7.485 5.345 ;
        RECT 9.165 2.055 9.335 5.095 ;
        RECT 9.935 4.940 10.105 5.095 ;
        RECT 9.905 4.765 10.105 4.940 ;
        RECT 9.905 2.055 10.075 4.765 ;
        RECT 3.500 0.985 3.670 1.720 ;
        RECT 5.420 1.635 6.560 1.805 ;
        RECT 3.985 0.765 4.155 1.535 ;
        RECT 3.015 0.595 4.155 0.765 ;
        RECT 3.015 0.515 3.185 0.595 ;
        RECT 3.985 0.515 4.155 0.595 ;
        RECT 5.420 0.505 5.590 1.635 ;
        RECT 6.390 0.755 6.560 1.635 ;
        RECT 6.875 1.710 7.485 1.880 ;
        RECT 8.750 1.805 8.920 1.885 ;
        RECT 9.720 1.805 9.890 1.885 ;
        RECT 10.645 1.880 10.815 5.345 ;
        RECT 12.495 2.055 12.665 5.095 ;
        RECT 6.875 0.975 7.045 1.710 ;
        RECT 8.750 1.635 9.890 1.805 ;
        RECT 7.360 0.755 7.530 1.525 ;
        RECT 6.390 0.585 7.530 0.755 ;
        RECT 6.390 0.505 6.560 0.585 ;
        RECT 7.360 0.505 7.530 0.585 ;
        RECT 8.750 0.505 8.920 1.635 ;
        RECT 9.720 0.755 9.890 1.635 ;
        RECT 10.205 1.710 10.815 1.880 ;
        RECT 12.080 1.805 12.250 1.885 ;
        RECT 13.050 1.805 13.220 1.885 ;
        RECT 13.975 1.880 14.145 5.345 ;
        RECT 15.825 2.055 15.995 5.095 ;
        RECT 19.925 4.940 20.095 5.095 ;
        RECT 19.895 4.765 20.095 4.940 ;
        RECT 19.895 2.055 20.065 4.765 ;
        RECT 10.205 0.975 10.375 1.710 ;
        RECT 12.080 1.635 13.220 1.805 ;
        RECT 10.690 0.755 10.860 1.525 ;
        RECT 9.720 0.585 10.860 0.755 ;
        RECT 9.720 0.505 9.890 0.585 ;
        RECT 10.690 0.505 10.860 0.585 ;
        RECT 12.080 0.505 12.250 1.635 ;
        RECT 13.050 0.755 13.220 1.635 ;
        RECT 13.535 1.710 14.145 1.880 ;
        RECT 15.410 1.805 15.580 1.885 ;
        RECT 16.380 1.805 16.550 1.885 ;
        RECT 13.535 0.975 13.705 1.710 ;
        RECT 15.410 1.635 16.550 1.805 ;
        RECT 14.020 0.755 14.190 1.525 ;
        RECT 13.050 0.585 14.190 0.755 ;
        RECT 13.050 0.505 13.220 0.585 ;
        RECT 14.020 0.505 14.190 0.585 ;
        RECT 15.410 0.505 15.580 1.635 ;
        RECT 16.380 0.755 16.550 1.635 ;
        RECT 18.740 1.805 18.910 1.885 ;
        RECT 19.710 1.805 19.880 1.885 ;
        RECT 18.740 1.635 19.880 1.805 ;
        RECT 17.350 0.755 17.520 1.525 ;
        RECT 16.380 0.585 17.520 0.755 ;
        RECT 16.380 0.505 16.550 0.585 ;
        RECT 17.350 0.505 17.520 0.585 ;
        RECT 18.740 0.505 18.910 1.635 ;
        RECT 19.710 0.755 19.880 1.635 ;
        RECT 20.680 0.755 20.850 1.525 ;
        RECT 19.710 0.585 20.850 0.755 ;
        RECT 19.710 0.505 19.880 0.585 ;
        RECT 20.680 0.505 20.850 0.585 ;
      LAYER mcon ;
        RECT 1.025 4.355 1.195 4.525 ;
        RECT 3.245 3.615 3.415 3.785 ;
        RECT 3.985 3.985 4.155 4.155 ;
        RECT 5.835 3.985 6.005 4.155 ;
        RECT 7.315 3.615 7.485 3.785 ;
        RECT 9.165 3.615 9.335 3.785 ;
        RECT 9.905 4.355 10.075 4.525 ;
        RECT 10.645 3.615 10.815 3.785 ;
        RECT 12.495 3.615 12.665 3.785 ;
        RECT 13.975 4.355 14.145 4.525 ;
        RECT 15.825 3.985 15.995 4.155 ;
        RECT 19.895 4.355 20.065 4.525 ;
      LAYER met1 ;
        RECT 0.995 4.525 1.225 4.555 ;
        RECT 9.875 4.525 10.105 4.555 ;
        RECT 13.945 4.525 14.175 4.555 ;
        RECT 19.865 4.525 20.095 4.555 ;
        RECT 0.965 4.355 20.125 4.525 ;
        RECT 0.995 4.325 1.225 4.355 ;
        RECT 9.875 4.325 10.105 4.355 ;
        RECT 13.945 4.325 14.175 4.355 ;
        RECT 19.865 4.325 20.095 4.355 ;
        RECT 3.955 4.155 4.185 4.185 ;
        RECT 5.805 4.155 6.035 4.185 ;
        RECT 15.795 4.155 16.025 4.185 ;
        RECT 3.925 3.985 16.055 4.155 ;
        RECT 3.955 3.955 4.185 3.985 ;
        RECT 5.805 3.955 6.035 3.985 ;
        RECT 15.795 3.955 16.025 3.985 ;
        RECT 3.215 3.785 3.445 3.815 ;
        RECT 7.285 3.785 7.515 3.815 ;
        RECT 9.135 3.785 9.365 3.815 ;
        RECT 10.615 3.785 10.845 3.815 ;
        RECT 12.465 3.785 12.695 3.815 ;
        RECT 3.185 3.615 9.395 3.785 ;
        RECT 10.585 3.615 12.725 3.785 ;
        RECT 3.215 3.585 3.445 3.615 ;
        RECT 7.285 3.585 7.515 3.615 ;
        RECT 9.135 3.585 9.365 3.615 ;
        RECT 10.615 3.585 10.845 3.615 ;
        RECT 12.465 3.585 12.695 3.615 ;
  END
END DFFX1






MACRO DLATCH
  CLASS BLOCK ;
  FOREIGN DLATCH ;
  ORIGIN 0.420 0.075 ;
  SIZE 20.820 BY 7.950 ;
  PIN Q
    ANTENNAGATEAREA 1.027250 ;
    ANTENNADIFFAREA 0.963050 ;
    PORT
      LAYER li1 ;
        RECT 15.345 5.525 15.515 6.795 ;
        RECT 15.345 5.355 15.995 5.525 ;
        RECT 15.825 1.880 15.995 5.355 ;
        RECT 17.520 4.940 17.690 5.100 ;
        RECT 17.520 4.770 17.845 4.940 ;
        RECT 17.675 2.055 17.845 4.770 ;
        RECT 14.415 1.710 15.995 1.880 ;
        RECT 14.415 0.975 14.585 1.710 ;
        RECT 15.385 0.975 15.555 1.710 ;
      LAYER mcon ;
        RECT 15.825 3.245 15.995 3.415 ;
        RECT 17.675 3.245 17.845 3.415 ;
      LAYER met1 ;
        RECT 15.795 3.415 16.025 3.445 ;
        RECT 17.645 3.415 17.875 3.445 ;
        RECT 15.765 3.245 17.905 3.415 ;
        RECT 15.795 3.215 16.025 3.245 ;
        RECT 17.645 3.215 17.875 3.245 ;
    END
  END Q
  PIN D
    ANTENNAGATEAREA 2.054500 ;
    PORT
      LAYER li1 ;
        RECT 0.655 2.055 0.825 5.095 ;
        RECT 9.565 4.940 9.735 5.095 ;
        RECT 9.535 4.765 9.735 4.940 ;
        RECT 9.535 2.055 9.705 4.765 ;
      LAYER mcon ;
        RECT 0.655 3.985 0.825 4.155 ;
        RECT 9.535 3.985 9.705 4.155 ;
      LAYER met1 ;
        RECT 0.625 4.155 0.855 4.185 ;
        RECT 9.505 4.155 9.735 4.185 ;
        RECT 0.595 3.985 9.765 4.155 ;
        RECT 0.625 3.955 0.855 3.985 ;
        RECT 9.505 3.955 9.735 3.985 ;
    END
  END D
  PIN GATE
    ANTENNAGATEAREA 2.060500 ;
    PORT
      LAYER li1 ;
        RECT 4.015 4.940 4.185 5.095 ;
        RECT 3.985 4.765 4.185 4.940 ;
        RECT 3.985 2.055 4.155 4.765 ;
        RECT 8.795 2.055 8.965 5.095 ;
      LAYER mcon ;
        RECT 3.985 2.875 4.155 3.045 ;
        RECT 8.795 2.875 8.965 3.045 ;
      LAYER met1 ;
        RECT 3.955 3.045 4.185 3.075 ;
        RECT 8.765 3.045 8.995 3.075 ;
        RECT 3.925 2.875 9.025 3.045 ;
        RECT 3.955 2.845 4.185 2.875 ;
        RECT 8.765 2.845 8.995 2.875 ;
    END
  END GATE
  PIN VDD
    ANTENNADIFFAREA 24.689199 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 20.400 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 20.135 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 0.585 5.415 0.755 7.460 ;
        RECT 1.465 5.415 1.635 7.460 ;
        RECT 2.065 4.340 2.375 7.460 ;
        RECT 2.925 5.365 3.095 7.460 ;
        RECT 3.805 5.785 3.975 7.460 ;
        RECT 4.685 5.785 4.855 7.460 ;
        RECT 5.395 4.340 5.705 7.460 ;
        RECT 6.135 5.415 6.305 7.460 ;
        RECT 7.015 5.415 7.185 7.460 ;
        RECT 7.615 4.340 7.925 7.460 ;
        RECT 8.475 5.365 8.645 7.460 ;
        RECT 9.355 5.785 9.525 7.460 ;
        RECT 10.235 5.785 10.405 7.460 ;
        RECT 10.945 4.340 11.255 7.460 ;
        RECT 11.685 5.415 11.855 7.460 ;
        RECT 12.565 5.415 12.735 7.460 ;
        RECT 13.165 4.340 13.475 7.460 ;
        RECT 14.465 5.785 14.635 7.460 ;
        RECT 16.495 4.340 16.805 7.460 ;
        RECT 17.795 5.785 17.965 7.460 ;
        RECT 19.825 4.340 20.135 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 1.025 7.525 1.195 7.695 ;
        RECT 1.415 7.525 1.585 7.695 ;
        RECT 1.775 7.525 1.945 7.695 ;
        RECT 2.495 7.525 2.665 7.695 ;
        RECT 2.855 7.525 3.025 7.695 ;
        RECT 3.215 7.525 3.385 7.695 ;
        RECT 3.575 7.525 3.745 7.695 ;
        RECT 4.025 7.525 4.195 7.695 ;
        RECT 4.385 7.525 4.555 7.695 ;
        RECT 4.745 7.525 4.915 7.695 ;
        RECT 5.105 7.525 5.275 7.695 ;
        RECT 5.825 7.525 5.995 7.695 ;
        RECT 6.185 7.525 6.355 7.695 ;
        RECT 6.575 7.525 6.745 7.695 ;
        RECT 6.965 7.525 7.135 7.695 ;
        RECT 7.325 7.525 7.495 7.695 ;
        RECT 8.045 7.525 8.215 7.695 ;
        RECT 8.405 7.525 8.575 7.695 ;
        RECT 8.765 7.525 8.935 7.695 ;
        RECT 9.125 7.525 9.295 7.695 ;
        RECT 9.575 7.525 9.745 7.695 ;
        RECT 9.935 7.525 10.105 7.695 ;
        RECT 10.295 7.525 10.465 7.695 ;
        RECT 10.655 7.525 10.825 7.695 ;
        RECT 11.375 7.525 11.545 7.695 ;
        RECT 11.735 7.525 11.905 7.695 ;
        RECT 12.125 7.525 12.295 7.695 ;
        RECT 12.515 7.525 12.685 7.695 ;
        RECT 12.875 7.525 13.045 7.695 ;
        RECT 13.595 7.525 13.765 7.695 ;
        RECT 13.955 7.525 14.125 7.695 ;
        RECT 14.315 7.525 14.485 7.695 ;
        RECT 14.675 7.525 14.845 7.695 ;
        RECT 15.125 7.525 15.295 7.695 ;
        RECT 15.485 7.525 15.655 7.695 ;
        RECT 15.845 7.525 16.015 7.695 ;
        RECT 16.205 7.525 16.375 7.695 ;
        RECT 16.925 7.525 17.095 7.695 ;
        RECT 17.285 7.525 17.455 7.695 ;
        RECT 17.645 7.525 17.815 7.695 ;
        RECT 18.005 7.525 18.175 7.695 ;
        RECT 18.455 7.525 18.625 7.695 ;
        RECT 18.815 7.525 18.985 7.695 ;
        RECT 19.175 7.525 19.345 7.695 ;
        RECT 19.535 7.525 19.705 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 20.135 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 23.443249 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 20.265 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 1.935 -0.075 2.505 -0.065 ;
        RECT 5.265 -0.075 5.835 -0.065 ;
        RECT 7.485 -0.075 8.055 -0.065 ;
        RECT 10.815 -0.075 11.385 -0.065 ;
        RECT 13.035 -0.075 13.605 -0.065 ;
        RECT 16.365 -0.075 16.935 -0.065 ;
        RECT 19.695 -0.075 20.265 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 0.545 0.755 0.715 1.885 ;
        RECT 1.515 0.755 1.685 1.885 ;
        RECT 0.545 0.585 1.685 0.755 ;
        RECT 0.545 0.310 0.715 0.585 ;
        RECT 1.030 0.310 1.200 0.585 ;
        RECT 1.515 0.310 1.685 0.585 ;
        RECT 2.065 0.310 2.375 2.860 ;
        RECT 3.315 0.310 3.485 1.260 ;
        RECT 5.395 0.310 5.705 2.860 ;
        RECT 6.095 0.755 6.265 1.885 ;
        RECT 7.065 0.755 7.235 1.885 ;
        RECT 6.095 0.585 7.235 0.755 ;
        RECT 6.095 0.310 6.265 0.585 ;
        RECT 6.580 0.310 6.750 0.585 ;
        RECT 7.065 0.310 7.235 0.585 ;
        RECT 7.615 0.310 7.925 2.860 ;
        RECT 8.865 0.310 9.035 1.260 ;
        RECT 10.945 0.310 11.255 2.860 ;
        RECT 11.645 0.755 11.815 1.885 ;
        RECT 12.615 0.755 12.785 1.885 ;
        RECT 11.645 0.585 12.785 0.755 ;
        RECT 11.645 0.310 11.815 0.585 ;
        RECT 12.130 0.310 12.300 0.585 ;
        RECT 12.615 0.310 12.785 0.585 ;
        RECT 13.165 0.310 13.475 2.860 ;
        RECT 13.930 0.755 14.100 1.885 ;
        RECT 14.900 0.755 15.070 1.530 ;
        RECT 15.870 0.755 16.040 1.530 ;
        RECT 13.930 0.585 16.040 0.755 ;
        RECT 13.930 0.310 14.100 0.585 ;
        RECT 14.415 0.310 14.585 0.585 ;
        RECT 14.900 0.310 15.070 0.585 ;
        RECT 15.385 0.310 15.555 0.585 ;
        RECT 15.870 0.310 16.040 0.585 ;
        RECT 16.495 0.310 16.805 2.860 ;
        RECT 17.260 0.755 17.430 1.885 ;
        RECT 18.230 0.755 18.400 1.530 ;
        RECT 19.200 0.755 19.370 1.530 ;
        RECT 17.260 0.585 19.370 0.755 ;
        RECT 17.260 0.310 17.430 0.585 ;
        RECT 17.745 0.310 17.915 0.585 ;
        RECT 18.230 0.310 18.400 0.585 ;
        RECT 18.715 0.310 18.885 0.585 ;
        RECT 19.200 0.310 19.370 0.585 ;
        RECT 19.825 0.310 20.135 2.860 ;
        RECT -0.155 0.000 20.135 0.310 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 1.025 0.065 1.195 0.235 ;
        RECT 1.415 0.065 1.585 0.235 ;
        RECT 1.775 0.065 1.945 0.235 ;
        RECT 2.495 0.065 2.665 0.235 ;
        RECT 2.855 0.065 3.025 0.235 ;
        RECT 3.215 0.065 3.385 0.235 ;
        RECT 3.575 0.065 3.745 0.235 ;
        RECT 4.025 0.065 4.195 0.235 ;
        RECT 4.385 0.065 4.555 0.235 ;
        RECT 4.745 0.065 4.915 0.235 ;
        RECT 5.105 0.065 5.275 0.235 ;
        RECT 5.825 0.065 5.995 0.235 ;
        RECT 6.185 0.065 6.355 0.235 ;
        RECT 6.575 0.065 6.745 0.235 ;
        RECT 6.965 0.065 7.135 0.235 ;
        RECT 7.325 0.065 7.495 0.235 ;
        RECT 8.045 0.065 8.215 0.235 ;
        RECT 8.405 0.065 8.575 0.235 ;
        RECT 8.765 0.065 8.935 0.235 ;
        RECT 9.125 0.065 9.295 0.235 ;
        RECT 9.575 0.065 9.745 0.235 ;
        RECT 9.935 0.065 10.105 0.235 ;
        RECT 10.295 0.065 10.465 0.235 ;
        RECT 10.655 0.065 10.825 0.235 ;
        RECT 11.375 0.065 11.545 0.235 ;
        RECT 11.735 0.065 11.905 0.235 ;
        RECT 12.125 0.065 12.295 0.235 ;
        RECT 12.515 0.065 12.685 0.235 ;
        RECT 12.875 0.065 13.045 0.235 ;
        RECT 13.595 0.065 13.765 0.235 ;
        RECT 13.955 0.065 14.125 0.235 ;
        RECT 14.315 0.065 14.485 0.235 ;
        RECT 14.675 0.065 14.845 0.235 ;
        RECT 15.125 0.065 15.295 0.235 ;
        RECT 15.485 0.065 15.655 0.235 ;
        RECT 15.845 0.065 16.015 0.235 ;
        RECT 16.205 0.065 16.375 0.235 ;
        RECT 16.925 0.065 17.095 0.235 ;
        RECT 17.285 0.065 17.455 0.235 ;
        RECT 17.645 0.065 17.815 0.235 ;
        RECT 18.005 0.065 18.175 0.235 ;
        RECT 18.455 0.065 18.625 0.235 ;
        RECT 18.815 0.065 18.985 0.235 ;
        RECT 19.175 0.065 19.345 0.235 ;
        RECT 19.535 0.065 19.705 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 20.135 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 1.025 4.895 1.195 7.250 ;
        RECT 3.365 5.515 3.535 7.250 ;
        RECT 4.245 5.515 4.415 7.250 ;
        RECT 3.365 5.345 4.895 5.515 ;
        RECT 1.025 4.725 1.565 4.895 ;
        RECT 1.395 2.305 1.565 4.725 ;
        RECT 1.025 2.135 1.565 2.305 ;
        RECT 1.025 0.975 1.195 2.135 ;
        RECT 3.245 2.055 3.415 5.095 ;
        RECT 2.830 1.805 3.000 1.885 ;
        RECT 3.800 1.805 3.970 1.885 ;
        RECT 4.725 1.880 4.895 5.345 ;
        RECT 6.205 2.055 6.375 5.095 ;
        RECT 6.575 4.895 6.745 7.250 ;
        RECT 8.915 5.515 9.085 7.250 ;
        RECT 9.795 5.515 9.965 7.250 ;
        RECT 8.915 5.345 10.445 5.515 ;
        RECT 6.575 4.725 7.115 4.895 ;
        RECT 6.945 2.305 7.115 4.725 ;
        RECT 6.575 2.135 7.115 2.305 ;
        RECT 2.830 1.635 3.970 1.805 ;
        RECT 2.830 0.505 3.000 1.635 ;
        RECT 3.800 0.755 3.970 1.635 ;
        RECT 4.285 1.710 4.895 1.880 ;
        RECT 4.285 0.975 4.455 1.710 ;
        RECT 4.770 0.755 4.940 1.525 ;
        RECT 6.575 0.975 6.745 2.135 ;
        RECT 8.380 1.805 8.550 1.885 ;
        RECT 9.350 1.805 9.520 1.885 ;
        RECT 10.275 1.880 10.445 5.345 ;
        RECT 11.755 2.055 11.925 5.095 ;
        RECT 12.125 4.895 12.295 7.250 ;
        RECT 14.025 5.525 14.195 7.255 ;
        RECT 14.905 7.055 15.955 7.225 ;
        RECT 14.905 5.525 15.075 7.055 ;
        RECT 15.785 5.785 15.955 7.055 ;
        RECT 14.025 5.355 15.075 5.525 ;
        RECT 17.355 5.525 17.525 7.255 ;
        RECT 18.235 7.055 19.285 7.225 ;
        RECT 18.235 5.525 18.405 7.055 ;
        RECT 17.355 5.355 18.405 5.525 ;
        RECT 18.675 5.525 18.845 6.795 ;
        RECT 19.115 5.785 19.285 7.055 ;
        RECT 18.675 5.355 19.325 5.525 ;
        RECT 14.190 4.940 14.360 5.100 ;
        RECT 15.120 4.940 15.290 5.100 ;
        RECT 18.450 4.940 18.620 5.100 ;
        RECT 12.125 4.725 12.665 4.895 ;
        RECT 14.190 4.770 14.515 4.940 ;
        RECT 12.495 2.305 12.665 4.725 ;
        RECT 12.125 2.135 12.665 2.305 ;
        RECT 8.380 1.635 9.520 1.805 ;
        RECT 3.800 0.585 4.940 0.755 ;
        RECT 3.800 0.505 3.970 0.585 ;
        RECT 4.770 0.505 4.940 0.585 ;
        RECT 8.380 0.505 8.550 1.635 ;
        RECT 9.350 0.755 9.520 1.635 ;
        RECT 9.835 1.710 10.445 1.880 ;
        RECT 9.835 0.975 10.005 1.710 ;
        RECT 10.320 0.755 10.490 1.525 ;
        RECT 12.125 0.975 12.295 2.135 ;
        RECT 14.345 2.055 14.515 4.770 ;
        RECT 15.085 4.770 15.290 4.940 ;
        RECT 18.415 4.770 18.620 4.940 ;
        RECT 15.085 2.055 15.255 4.770 ;
        RECT 18.415 2.055 18.585 4.770 ;
        RECT 19.155 1.880 19.325 5.355 ;
        RECT 17.745 1.710 19.325 1.880 ;
        RECT 17.745 0.975 17.915 1.710 ;
        RECT 18.715 0.975 18.885 1.710 ;
        RECT 9.350 0.585 10.490 0.755 ;
        RECT 9.350 0.505 9.520 0.585 ;
        RECT 10.320 0.505 10.490 0.585 ;
      LAYER mcon ;
        RECT 1.395 3.615 1.565 3.785 ;
        RECT 3.245 3.615 3.415 3.785 ;
        RECT 4.725 3.245 4.895 3.415 ;
        RECT 6.205 3.245 6.375 3.415 ;
        RECT 6.945 3.615 7.115 3.785 ;
        RECT 10.275 3.245 10.445 3.415 ;
        RECT 11.755 3.245 11.925 3.415 ;
        RECT 12.495 3.985 12.665 4.155 ;
        RECT 14.345 3.615 14.515 3.785 ;
        RECT 15.085 3.615 15.255 3.785 ;
        RECT 18.415 3.985 18.585 4.155 ;
        RECT 19.155 3.615 19.325 3.785 ;
      LAYER met1 ;
        RECT 12.465 4.155 12.695 4.185 ;
        RECT 18.385 4.155 18.615 4.185 ;
        RECT 12.435 3.985 18.645 4.155 ;
        RECT 12.465 3.955 12.695 3.985 ;
        RECT 18.385 3.955 18.615 3.985 ;
        RECT 1.365 3.785 1.595 3.815 ;
        RECT 3.215 3.785 3.445 3.815 ;
        RECT 6.915 3.785 7.145 3.815 ;
        RECT 14.315 3.785 14.545 3.815 ;
        RECT 15.055 3.785 15.285 3.815 ;
        RECT 19.125 3.785 19.355 3.815 ;
        RECT 1.335 3.615 3.475 3.785 ;
        RECT 6.885 3.615 14.575 3.785 ;
        RECT 15.025 3.615 19.385 3.785 ;
        RECT 1.365 3.585 1.595 3.615 ;
        RECT 3.215 3.585 3.445 3.615 ;
        RECT 6.915 3.585 7.145 3.615 ;
        RECT 14.315 3.585 14.545 3.615 ;
        RECT 15.055 3.585 15.285 3.615 ;
        RECT 19.125 3.585 19.355 3.615 ;
        RECT 4.695 3.415 4.925 3.445 ;
        RECT 6.175 3.415 6.405 3.445 ;
        RECT 10.245 3.415 10.475 3.445 ;
        RECT 11.725 3.415 11.955 3.445 ;
        RECT 4.665 3.245 6.435 3.415 ;
        RECT 10.215 3.245 11.985 3.415 ;
        RECT 4.695 3.215 4.925 3.245 ;
        RECT 6.175 3.215 6.405 3.245 ;
        RECT 10.245 3.215 10.475 3.245 ;
        RECT 11.725 3.215 11.955 3.245 ;
  END
END DLATCH






MACRO DLATCHN
  CLASS BLOCK ;
  FOREIGN DLATCHN ;
  ORIGIN 2.640 0.075 ;
  SIZE 23.040 BY 7.950 ;
  PIN Q
    ANTENNAGATEAREA 1.027250 ;
    ANTENNADIFFAREA 0.963050 ;
    PORT
      LAYER li1 ;
        RECT 15.345 5.525 15.515 6.795 ;
        RECT 15.345 5.355 15.995 5.525 ;
        RECT 15.825 1.880 15.995 5.355 ;
        RECT 17.520 4.940 17.690 5.100 ;
        RECT 17.520 4.770 17.845 4.940 ;
        RECT 17.675 2.055 17.845 4.770 ;
        RECT 14.415 1.710 15.995 1.880 ;
        RECT 14.415 0.975 14.585 1.710 ;
        RECT 15.385 0.975 15.555 1.710 ;
      LAYER mcon ;
        RECT 15.825 3.245 15.995 3.415 ;
        RECT 17.675 3.245 17.845 3.415 ;
      LAYER met1 ;
        RECT 15.795 3.415 16.025 3.445 ;
        RECT 17.645 3.415 17.875 3.445 ;
        RECT 15.765 3.245 17.905 3.415 ;
        RECT 15.795 3.215 16.025 3.245 ;
        RECT 17.645 3.215 17.875 3.245 ;
    END
  END Q
  PIN D
    ANTENNAGATEAREA 2.054500 ;
    PORT
      LAYER li1 ;
        RECT 0.655 2.055 0.825 5.095 ;
        RECT 9.565 4.940 9.735 5.095 ;
        RECT 9.535 4.765 9.735 4.940 ;
        RECT 9.535 2.055 9.705 4.765 ;
      LAYER mcon ;
        RECT 0.655 3.985 0.825 4.155 ;
        RECT 9.535 3.985 9.705 4.155 ;
      LAYER met1 ;
        RECT 0.625 4.155 0.855 4.185 ;
        RECT 9.505 4.155 9.735 4.185 ;
        RECT 0.595 3.985 9.765 4.155 ;
        RECT 0.625 3.955 0.855 3.985 ;
        RECT 9.505 3.955 9.735 3.985 ;
    END
  END D
  PIN GATE_N
    ANTENNAGATEAREA 1.027250 ;
    PORT
      LAYER li1 ;
        RECT -1.565 2.055 -1.395 5.095 ;
      LAYER mcon ;
        RECT -1.565 2.875 -1.395 3.045 ;
      LAYER met1 ;
        RECT -1.595 3.045 -1.365 3.075 ;
        RECT -1.745 2.875 -1.335 3.045 ;
        RECT -1.595 2.845 -1.365 2.875 ;
    END
  END GATE_N
  PIN VDD
    ANTENNADIFFAREA 27.746050 ;
    PORT
      LAYER nwell ;
        RECT -2.640 4.160 20.400 7.875 ;
      LAYER li1 ;
        RECT -2.375 7.460 20.135 7.770 ;
        RECT -2.375 4.340 -2.065 7.460 ;
        RECT -1.635 5.415 -1.465 7.460 ;
        RECT -0.755 5.415 -0.585 7.460 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 0.585 5.415 0.755 7.460 ;
        RECT 1.465 5.415 1.635 7.460 ;
        RECT 2.065 4.340 2.375 7.460 ;
        RECT 2.925 5.365 3.095 7.460 ;
        RECT 3.805 5.785 3.975 7.460 ;
        RECT 4.685 5.785 4.855 7.460 ;
        RECT 5.395 4.340 5.705 7.460 ;
        RECT 6.135 5.415 6.305 7.460 ;
        RECT 7.015 5.415 7.185 7.460 ;
        RECT 7.615 4.340 7.925 7.460 ;
        RECT 8.475 5.365 8.645 7.460 ;
        RECT 9.355 5.785 9.525 7.460 ;
        RECT 10.235 5.785 10.405 7.460 ;
        RECT 10.945 4.340 11.255 7.460 ;
        RECT 11.685 5.415 11.855 7.460 ;
        RECT 12.565 5.415 12.735 7.460 ;
        RECT 13.165 4.340 13.475 7.460 ;
        RECT 14.465 5.785 14.635 7.460 ;
        RECT 16.495 4.340 16.805 7.460 ;
        RECT 17.795 5.785 17.965 7.460 ;
        RECT 19.825 4.340 20.135 7.460 ;
      LAYER mcon ;
        RECT -1.945 7.525 -1.775 7.695 ;
        RECT -1.585 7.525 -1.415 7.695 ;
        RECT -1.195 7.525 -1.025 7.695 ;
        RECT -0.805 7.525 -0.635 7.695 ;
        RECT -0.445 7.525 -0.275 7.695 ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 1.025 7.525 1.195 7.695 ;
        RECT 1.415 7.525 1.585 7.695 ;
        RECT 1.775 7.525 1.945 7.695 ;
        RECT 2.495 7.525 2.665 7.695 ;
        RECT 2.855 7.525 3.025 7.695 ;
        RECT 3.215 7.525 3.385 7.695 ;
        RECT 3.575 7.525 3.745 7.695 ;
        RECT 4.025 7.525 4.195 7.695 ;
        RECT 4.385 7.525 4.555 7.695 ;
        RECT 4.745 7.525 4.915 7.695 ;
        RECT 5.105 7.525 5.275 7.695 ;
        RECT 5.825 7.525 5.995 7.695 ;
        RECT 6.185 7.525 6.355 7.695 ;
        RECT 6.575 7.525 6.745 7.695 ;
        RECT 6.965 7.525 7.135 7.695 ;
        RECT 7.325 7.525 7.495 7.695 ;
        RECT 8.045 7.525 8.215 7.695 ;
        RECT 8.405 7.525 8.575 7.695 ;
        RECT 8.765 7.525 8.935 7.695 ;
        RECT 9.125 7.525 9.295 7.695 ;
        RECT 9.575 7.525 9.745 7.695 ;
        RECT 9.935 7.525 10.105 7.695 ;
        RECT 10.295 7.525 10.465 7.695 ;
        RECT 10.655 7.525 10.825 7.695 ;
        RECT 11.375 7.525 11.545 7.695 ;
        RECT 11.735 7.525 11.905 7.695 ;
        RECT 12.125 7.525 12.295 7.695 ;
        RECT 12.515 7.525 12.685 7.695 ;
        RECT 12.875 7.525 13.045 7.695 ;
        RECT 13.595 7.525 13.765 7.695 ;
        RECT 13.955 7.525 14.125 7.695 ;
        RECT 14.315 7.525 14.485 7.695 ;
        RECT 14.675 7.525 14.845 7.695 ;
        RECT 15.125 7.525 15.295 7.695 ;
        RECT 15.485 7.525 15.655 7.695 ;
        RECT 15.845 7.525 16.015 7.695 ;
        RECT 16.205 7.525 16.375 7.695 ;
        RECT 16.925 7.525 17.095 7.695 ;
        RECT 17.285 7.525 17.455 7.695 ;
        RECT 17.645 7.525 17.815 7.695 ;
        RECT 18.005 7.525 18.175 7.695 ;
        RECT 18.455 7.525 18.625 7.695 ;
        RECT 18.815 7.525 18.985 7.695 ;
        RECT 19.175 7.525 19.345 7.695 ;
        RECT 19.535 7.525 19.705 7.695 ;
      LAYER met1 ;
        RECT -2.375 7.460 20.135 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 26.407349 ;
    PORT
      LAYER pwell ;
        RECT -2.505 -0.065 20.265 2.990 ;
        RECT -2.505 -0.075 -1.935 -0.065 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 1.935 -0.075 2.505 -0.065 ;
        RECT 5.265 -0.075 5.835 -0.065 ;
        RECT 7.485 -0.075 8.055 -0.065 ;
        RECT 10.815 -0.075 11.385 -0.065 ;
        RECT 13.035 -0.075 13.605 -0.065 ;
        RECT 16.365 -0.075 16.935 -0.065 ;
        RECT 19.695 -0.075 20.265 -0.065 ;
      LAYER li1 ;
        RECT -2.375 0.310 -2.065 2.860 ;
        RECT -1.675 0.755 -1.505 1.885 ;
        RECT -0.705 0.755 -0.535 1.885 ;
        RECT -1.675 0.585 -0.535 0.755 ;
        RECT -1.675 0.310 -1.505 0.585 ;
        RECT -1.190 0.310 -1.020 0.585 ;
        RECT -0.705 0.310 -0.535 0.585 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 0.545 0.755 0.715 1.885 ;
        RECT 1.515 0.755 1.685 1.885 ;
        RECT 0.545 0.585 1.685 0.755 ;
        RECT 0.545 0.310 0.715 0.585 ;
        RECT 1.030 0.310 1.200 0.585 ;
        RECT 1.515 0.310 1.685 0.585 ;
        RECT 2.065 0.310 2.375 2.860 ;
        RECT 3.315 0.310 3.485 1.260 ;
        RECT 5.395 0.310 5.705 2.860 ;
        RECT 6.095 0.755 6.265 1.885 ;
        RECT 7.065 0.755 7.235 1.885 ;
        RECT 6.095 0.585 7.235 0.755 ;
        RECT 6.095 0.310 6.265 0.585 ;
        RECT 6.580 0.310 6.750 0.585 ;
        RECT 7.065 0.310 7.235 0.585 ;
        RECT 7.615 0.310 7.925 2.860 ;
        RECT 8.865 0.310 9.035 1.260 ;
        RECT 10.945 0.310 11.255 2.860 ;
        RECT 11.645 0.755 11.815 1.885 ;
        RECT 12.615 0.755 12.785 1.885 ;
        RECT 11.645 0.585 12.785 0.755 ;
        RECT 11.645 0.310 11.815 0.585 ;
        RECT 12.130 0.310 12.300 0.585 ;
        RECT 12.615 0.310 12.785 0.585 ;
        RECT 13.165 0.310 13.475 2.860 ;
        RECT 13.930 0.755 14.100 1.885 ;
        RECT 14.900 0.755 15.070 1.530 ;
        RECT 15.870 0.755 16.040 1.530 ;
        RECT 13.930 0.585 16.040 0.755 ;
        RECT 13.930 0.310 14.100 0.585 ;
        RECT 14.415 0.310 14.585 0.585 ;
        RECT 14.900 0.310 15.070 0.585 ;
        RECT 15.385 0.310 15.555 0.585 ;
        RECT 15.870 0.310 16.040 0.585 ;
        RECT 16.495 0.310 16.805 2.860 ;
        RECT 17.260 0.755 17.430 1.885 ;
        RECT 18.230 0.755 18.400 1.530 ;
        RECT 19.200 0.755 19.370 1.530 ;
        RECT 17.260 0.585 19.370 0.755 ;
        RECT 17.260 0.310 17.430 0.585 ;
        RECT 17.745 0.310 17.915 0.585 ;
        RECT 18.230 0.310 18.400 0.585 ;
        RECT 18.715 0.310 18.885 0.585 ;
        RECT 19.200 0.310 19.370 0.585 ;
        RECT 19.825 0.310 20.135 2.860 ;
        RECT -2.375 0.000 20.135 0.310 ;
      LAYER mcon ;
        RECT -1.945 0.065 -1.775 0.235 ;
        RECT -1.585 0.065 -1.415 0.235 ;
        RECT -1.195 0.065 -1.025 0.235 ;
        RECT -0.805 0.065 -0.635 0.235 ;
        RECT -0.445 0.065 -0.275 0.235 ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 1.025 0.065 1.195 0.235 ;
        RECT 1.415 0.065 1.585 0.235 ;
        RECT 1.775 0.065 1.945 0.235 ;
        RECT 2.495 0.065 2.665 0.235 ;
        RECT 2.855 0.065 3.025 0.235 ;
        RECT 3.215 0.065 3.385 0.235 ;
        RECT 3.575 0.065 3.745 0.235 ;
        RECT 4.025 0.065 4.195 0.235 ;
        RECT 4.385 0.065 4.555 0.235 ;
        RECT 4.745 0.065 4.915 0.235 ;
        RECT 5.105 0.065 5.275 0.235 ;
        RECT 5.825 0.065 5.995 0.235 ;
        RECT 6.185 0.065 6.355 0.235 ;
        RECT 6.575 0.065 6.745 0.235 ;
        RECT 6.965 0.065 7.135 0.235 ;
        RECT 7.325 0.065 7.495 0.235 ;
        RECT 8.045 0.065 8.215 0.235 ;
        RECT 8.405 0.065 8.575 0.235 ;
        RECT 8.765 0.065 8.935 0.235 ;
        RECT 9.125 0.065 9.295 0.235 ;
        RECT 9.575 0.065 9.745 0.235 ;
        RECT 9.935 0.065 10.105 0.235 ;
        RECT 10.295 0.065 10.465 0.235 ;
        RECT 10.655 0.065 10.825 0.235 ;
        RECT 11.375 0.065 11.545 0.235 ;
        RECT 11.735 0.065 11.905 0.235 ;
        RECT 12.125 0.065 12.295 0.235 ;
        RECT 12.515 0.065 12.685 0.235 ;
        RECT 12.875 0.065 13.045 0.235 ;
        RECT 13.595 0.065 13.765 0.235 ;
        RECT 13.955 0.065 14.125 0.235 ;
        RECT 14.315 0.065 14.485 0.235 ;
        RECT 14.675 0.065 14.845 0.235 ;
        RECT 15.125 0.065 15.295 0.235 ;
        RECT 15.485 0.065 15.655 0.235 ;
        RECT 15.845 0.065 16.015 0.235 ;
        RECT 16.205 0.065 16.375 0.235 ;
        RECT 16.925 0.065 17.095 0.235 ;
        RECT 17.285 0.065 17.455 0.235 ;
        RECT 17.645 0.065 17.815 0.235 ;
        RECT 18.005 0.065 18.175 0.235 ;
        RECT 18.455 0.065 18.625 0.235 ;
        RECT 18.815 0.065 18.985 0.235 ;
        RECT 19.175 0.065 19.345 0.235 ;
        RECT 19.535 0.065 19.705 0.235 ;
      LAYER met1 ;
        RECT -2.375 0.000 20.135 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT -1.195 4.895 -1.025 7.250 ;
        RECT 1.025 4.895 1.195 7.250 ;
        RECT 3.365 5.515 3.535 7.250 ;
        RECT 4.245 5.515 4.415 7.250 ;
        RECT 3.365 5.345 4.895 5.515 ;
        RECT -1.195 4.725 -0.655 4.895 ;
        RECT 1.025 4.725 1.565 4.895 ;
        RECT -0.825 2.305 -0.655 4.725 ;
        RECT 1.395 2.305 1.565 4.725 ;
        RECT -1.195 2.135 -0.655 2.305 ;
        RECT 1.025 2.135 1.565 2.305 ;
        RECT -1.195 0.975 -1.025 2.135 ;
        RECT 1.025 0.975 1.195 2.135 ;
        RECT 3.245 2.055 3.415 5.095 ;
        RECT 4.015 4.940 4.185 5.095 ;
        RECT 3.985 4.765 4.185 4.940 ;
        RECT 3.985 2.055 4.155 4.765 ;
        RECT 2.830 1.805 3.000 1.885 ;
        RECT 3.800 1.805 3.970 1.885 ;
        RECT 4.725 1.880 4.895 5.345 ;
        RECT 6.205 2.055 6.375 5.095 ;
        RECT 6.575 4.895 6.745 7.250 ;
        RECT 8.915 5.515 9.085 7.250 ;
        RECT 9.795 5.515 9.965 7.250 ;
        RECT 8.915 5.345 10.445 5.515 ;
        RECT 6.575 4.725 7.115 4.895 ;
        RECT 6.945 2.305 7.115 4.725 ;
        RECT 6.575 2.135 7.115 2.305 ;
        RECT 2.830 1.635 3.970 1.805 ;
        RECT 2.830 0.505 3.000 1.635 ;
        RECT 3.800 0.755 3.970 1.635 ;
        RECT 4.285 1.710 4.895 1.880 ;
        RECT 4.285 0.975 4.455 1.710 ;
        RECT 4.770 0.755 4.940 1.525 ;
        RECT 6.575 0.975 6.745 2.135 ;
        RECT 8.795 2.055 8.965 5.095 ;
        RECT 8.380 1.805 8.550 1.885 ;
        RECT 9.350 1.805 9.520 1.885 ;
        RECT 10.275 1.880 10.445 5.345 ;
        RECT 11.755 2.055 11.925 5.095 ;
        RECT 12.125 4.895 12.295 7.250 ;
        RECT 14.025 5.525 14.195 7.255 ;
        RECT 14.905 7.055 15.955 7.225 ;
        RECT 14.905 5.525 15.075 7.055 ;
        RECT 15.785 5.785 15.955 7.055 ;
        RECT 14.025 5.355 15.075 5.525 ;
        RECT 17.355 5.525 17.525 7.255 ;
        RECT 18.235 7.055 19.285 7.225 ;
        RECT 18.235 5.525 18.405 7.055 ;
        RECT 17.355 5.355 18.405 5.525 ;
        RECT 18.675 5.525 18.845 6.795 ;
        RECT 19.115 5.785 19.285 7.055 ;
        RECT 18.675 5.355 19.325 5.525 ;
        RECT 14.190 4.940 14.360 5.100 ;
        RECT 15.120 4.940 15.290 5.100 ;
        RECT 18.450 4.940 18.620 5.100 ;
        RECT 12.125 4.725 12.665 4.895 ;
        RECT 14.190 4.770 14.515 4.940 ;
        RECT 12.495 2.305 12.665 4.725 ;
        RECT 12.125 2.135 12.665 2.305 ;
        RECT 8.380 1.635 9.520 1.805 ;
        RECT 3.800 0.585 4.940 0.755 ;
        RECT 3.800 0.505 3.970 0.585 ;
        RECT 4.770 0.505 4.940 0.585 ;
        RECT 8.380 0.505 8.550 1.635 ;
        RECT 9.350 0.755 9.520 1.635 ;
        RECT 9.835 1.710 10.445 1.880 ;
        RECT 9.835 0.975 10.005 1.710 ;
        RECT 10.320 0.755 10.490 1.525 ;
        RECT 12.125 0.975 12.295 2.135 ;
        RECT 14.345 2.055 14.515 4.770 ;
        RECT 15.085 4.770 15.290 4.940 ;
        RECT 18.415 4.770 18.620 4.940 ;
        RECT 15.085 2.055 15.255 4.770 ;
        RECT 18.415 2.055 18.585 4.770 ;
        RECT 19.155 1.880 19.325 5.355 ;
        RECT 17.745 1.710 19.325 1.880 ;
        RECT 17.745 0.975 17.915 1.710 ;
        RECT 18.715 0.975 18.885 1.710 ;
        RECT 9.350 0.585 10.490 0.755 ;
        RECT 9.350 0.505 9.520 0.585 ;
        RECT 10.320 0.505 10.490 0.585 ;
      LAYER mcon ;
        RECT -0.825 2.875 -0.655 3.045 ;
        RECT 1.395 3.615 1.565 3.785 ;
        RECT 3.245 3.615 3.415 3.785 ;
        RECT 3.985 2.875 4.155 3.045 ;
        RECT 4.725 3.245 4.895 3.415 ;
        RECT 6.205 3.245 6.375 3.415 ;
        RECT 6.945 3.615 7.115 3.785 ;
        RECT 8.795 2.875 8.965 3.045 ;
        RECT 10.275 3.245 10.445 3.415 ;
        RECT 11.755 3.245 11.925 3.415 ;
        RECT 12.495 3.985 12.665 4.155 ;
        RECT 14.345 3.615 14.515 3.785 ;
        RECT 15.085 3.615 15.255 3.785 ;
        RECT 18.415 3.985 18.585 4.155 ;
        RECT 19.155 3.615 19.325 3.785 ;
      LAYER met1 ;
        RECT 12.465 4.155 12.695 4.185 ;
        RECT 18.385 4.155 18.615 4.185 ;
        RECT 12.435 3.985 18.645 4.155 ;
        RECT 12.465 3.955 12.695 3.985 ;
        RECT 18.385 3.955 18.615 3.985 ;
        RECT 1.365 3.785 1.595 3.815 ;
        RECT 3.215 3.785 3.445 3.815 ;
        RECT 6.915 3.785 7.145 3.815 ;
        RECT 14.315 3.785 14.545 3.815 ;
        RECT 15.055 3.785 15.285 3.815 ;
        RECT 19.125 3.785 19.355 3.815 ;
        RECT 1.335 3.615 3.475 3.785 ;
        RECT 6.885 3.615 14.575 3.785 ;
        RECT 15.025 3.615 19.385 3.785 ;
        RECT 1.365 3.585 1.595 3.615 ;
        RECT 3.215 3.585 3.445 3.615 ;
        RECT 6.915 3.585 7.145 3.615 ;
        RECT 14.315 3.585 14.545 3.615 ;
        RECT 15.055 3.585 15.285 3.615 ;
        RECT 19.125 3.585 19.355 3.615 ;
        RECT 4.695 3.415 4.925 3.445 ;
        RECT 6.175 3.415 6.405 3.445 ;
        RECT 10.245 3.415 10.475 3.445 ;
        RECT 11.725 3.415 11.955 3.445 ;
        RECT 4.665 3.245 6.435 3.415 ;
        RECT 10.215 3.245 11.985 3.415 ;
        RECT 4.695 3.215 4.925 3.245 ;
        RECT 6.175 3.215 6.405 3.245 ;
        RECT 10.245 3.215 10.475 3.245 ;
        RECT 11.725 3.215 11.955 3.245 ;
        RECT -0.855 3.045 -0.625 3.075 ;
        RECT 3.955 3.045 4.185 3.075 ;
        RECT 8.765 3.045 8.995 3.075 ;
        RECT -0.885 2.875 9.025 3.045 ;
        RECT -0.855 2.845 -0.625 2.875 ;
        RECT 3.955 2.845 4.185 2.875 ;
        RECT 8.765 2.845 8.995 2.875 ;
  END
END DLATCHN






MACRO FA
  CLASS BLOCK ;
  FOREIGN FA ;
  ORIGIN 0.420 0.075 ;
  SIZE 39.690 BY 7.950 ;
  PIN SUM
    ANTENNADIFFAREA 1.543800 ;
    PORT
      LAYER li1 ;
        RECT 15.345 5.525 15.515 6.795 ;
        RECT 18.675 5.525 18.845 6.795 ;
        RECT 15.345 5.355 15.995 5.525 ;
        RECT 18.675 5.355 19.325 5.525 ;
        RECT 15.825 1.875 15.995 5.355 ;
        RECT 19.155 1.875 19.325 5.355 ;
        RECT 15.385 1.705 15.995 1.875 ;
        RECT 18.715 1.705 19.325 1.875 ;
        RECT 15.385 0.975 15.555 1.705 ;
        RECT 18.715 0.975 18.885 1.705 ;
      LAYER mcon ;
        RECT 15.825 3.615 15.995 3.785 ;
        RECT 19.155 3.615 19.325 3.785 ;
      LAYER met1 ;
        RECT 15.795 3.785 16.025 3.815 ;
        RECT 19.125 3.785 19.355 3.815 ;
        RECT 15.765 3.615 19.385 3.785 ;
        RECT 15.795 3.585 16.025 3.615 ;
        RECT 19.125 3.585 19.355 3.615 ;
    END
  END SUM
  PIN COUT
    ANTENNADIFFAREA 0.771900 ;
    PORT
      LAYER li1 ;
        RECT 37.655 4.895 37.825 7.250 ;
        RECT 37.655 4.725 38.195 4.895 ;
        RECT 38.025 2.305 38.195 4.725 ;
        RECT 37.655 2.135 38.195 2.305 ;
        RECT 37.655 0.975 37.825 2.135 ;
      LAYER mcon ;
        RECT 38.025 3.245 38.195 3.415 ;
      LAYER met1 ;
        RECT 37.995 3.415 38.225 3.445 ;
        RECT 37.965 3.245 38.375 3.415 ;
        RECT 37.995 3.215 38.225 3.245 ;
    END
  END COUT
  PIN A
    ANTENNAGATEAREA 3.087750 ;
    PORT
      LAYER li1 ;
        RECT 0.655 2.055 0.825 5.095 ;
        RECT 3.245 2.305 3.415 5.100 ;
        RECT 29.545 4.940 29.715 5.095 ;
        RECT 29.515 4.765 29.715 4.940 ;
        RECT 29.515 2.305 29.685 4.765 ;
        RECT 3.165 2.135 3.495 2.305 ;
        RECT 29.435 2.135 29.765 2.305 ;
        RECT 3.245 2.055 3.415 2.135 ;
        RECT 29.515 2.055 29.685 2.135 ;
      LAYER mcon ;
        RECT 0.655 4.355 0.825 4.525 ;
        RECT 3.245 4.355 3.415 4.525 ;
        RECT 3.245 2.135 3.415 2.305 ;
        RECT 29.515 2.135 29.685 2.305 ;
      LAYER met1 ;
        RECT 0.625 4.525 0.855 4.555 ;
        RECT 3.215 4.525 3.445 4.555 ;
        RECT 0.595 4.355 3.475 4.525 ;
        RECT 0.625 4.325 0.855 4.355 ;
        RECT 3.215 4.325 3.445 4.355 ;
        RECT 3.245 2.335 3.415 2.365 ;
        RECT 29.515 2.335 29.685 2.365 ;
        RECT 3.215 2.105 3.445 2.335 ;
        RECT 29.485 2.105 29.715 2.335 ;
        RECT 3.245 1.935 3.415 2.105 ;
        RECT 29.515 1.935 29.685 2.105 ;
        RECT 3.245 1.765 29.685 1.935 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 3.087750 ;
    PORT
      LAYER li1 ;
        RECT 6.575 4.275 6.745 5.100 ;
        RECT 4.355 2.055 4.525 2.755 ;
        RECT 10.275 2.055 10.445 5.095 ;
        RECT 28.775 2.055 28.945 5.095 ;
      LAYER mcon ;
        RECT 6.575 4.355 6.745 4.525 ;
        RECT 10.275 4.725 10.445 4.895 ;
        RECT 10.275 4.355 10.445 4.525 ;
        RECT 4.355 2.505 4.525 2.675 ;
        RECT 10.275 2.505 10.445 2.675 ;
        RECT 28.775 4.725 28.945 4.895 ;
      LAYER met1 ;
        RECT 10.245 4.895 10.475 4.925 ;
        RECT 28.745 4.895 28.975 4.925 ;
        RECT 10.215 4.725 29.005 4.895 ;
        RECT 10.245 4.695 10.475 4.725 ;
        RECT 28.745 4.695 28.975 4.725 ;
        RECT 6.545 4.525 6.775 4.555 ;
        RECT 10.245 4.525 10.475 4.555 ;
        RECT 6.515 4.355 10.505 4.525 ;
        RECT 6.545 4.325 6.775 4.355 ;
        RECT 10.245 4.325 10.475 4.355 ;
        RECT 4.325 2.675 4.555 2.705 ;
        RECT 10.245 2.675 10.475 2.705 ;
        RECT 4.295 2.505 10.505 2.675 ;
        RECT 4.325 2.475 4.555 2.505 ;
        RECT 10.245 2.475 10.475 2.505 ;
    END
  END B
  PIN CIN
    ANTENNAGATEAREA 3.087750 ;
    PORT
      LAYER li1 ;
        RECT 17.675 4.275 17.845 5.100 ;
        RECT 15.455 2.055 15.625 2.755 ;
        RECT 21.375 2.055 21.545 5.095 ;
        RECT 23.225 2.055 23.395 5.095 ;
      LAYER mcon ;
        RECT 17.675 4.355 17.845 4.525 ;
        RECT 21.375 4.355 21.545 4.525 ;
        RECT 15.455 2.505 15.625 2.675 ;
        RECT 21.375 2.505 21.545 2.675 ;
        RECT 23.225 4.355 23.395 4.525 ;
      LAYER met1 ;
        RECT 17.645 4.525 17.875 4.555 ;
        RECT 21.345 4.525 21.575 4.555 ;
        RECT 23.195 4.525 23.425 4.555 ;
        RECT 17.615 4.355 23.455 4.525 ;
        RECT 17.645 4.325 17.875 4.355 ;
        RECT 21.345 4.325 21.575 4.355 ;
        RECT 23.195 4.325 23.425 4.355 ;
        RECT 15.425 2.675 15.655 2.705 ;
        RECT 21.345 2.675 21.575 2.705 ;
        RECT 15.395 2.505 21.605 2.675 ;
        RECT 15.425 2.475 15.655 2.505 ;
        RECT 21.345 2.475 21.575 2.505 ;
    END
  END CIN
  PIN VDD
    ANTENNADIFFAREA 46.125549 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 39.270 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 39.005 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 0.585 5.415 0.755 7.460 ;
        RECT 1.465 5.415 1.635 7.460 ;
        RECT 2.065 4.340 2.375 7.460 ;
        RECT 3.365 5.785 3.535 7.460 ;
        RECT 5.395 4.340 5.705 7.460 ;
        RECT 6.695 5.785 6.865 7.460 ;
        RECT 8.725 4.340 9.035 7.460 ;
        RECT 9.465 5.415 9.635 7.460 ;
        RECT 10.345 5.415 10.515 7.460 ;
        RECT 10.945 4.340 11.255 7.460 ;
        RECT 11.685 5.415 11.855 7.460 ;
        RECT 12.565 5.415 12.735 7.460 ;
        RECT 13.165 4.340 13.475 7.460 ;
        RECT 14.465 5.785 14.635 7.460 ;
        RECT 16.495 4.340 16.805 7.460 ;
        RECT 17.795 5.785 17.965 7.460 ;
        RECT 19.825 4.340 20.135 7.460 ;
        RECT 20.565 5.415 20.735 7.460 ;
        RECT 21.445 5.415 21.615 7.460 ;
        RECT 22.045 4.340 22.355 7.460 ;
        RECT 22.905 5.365 23.075 7.460 ;
        RECT 23.785 5.785 23.955 7.460 ;
        RECT 24.665 5.785 24.835 7.460 ;
        RECT 25.375 4.340 25.685 7.460 ;
        RECT 26.115 5.415 26.285 7.460 ;
        RECT 26.995 5.415 27.165 7.460 ;
        RECT 27.595 4.340 27.905 7.460 ;
        RECT 28.455 5.365 28.625 7.460 ;
        RECT 29.335 5.785 29.505 7.460 ;
        RECT 30.215 5.785 30.385 7.460 ;
        RECT 30.925 4.340 31.235 7.460 ;
        RECT 31.665 5.415 31.835 7.460 ;
        RECT 32.545 5.415 32.715 7.460 ;
        RECT 33.145 4.340 33.455 7.460 ;
        RECT 34.445 5.785 34.615 7.460 ;
        RECT 36.475 4.340 36.785 7.460 ;
        RECT 37.215 5.415 37.385 7.460 ;
        RECT 38.095 5.415 38.265 7.460 ;
        RECT 38.695 4.340 39.005 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 1.025 7.525 1.195 7.695 ;
        RECT 1.415 7.525 1.585 7.695 ;
        RECT 1.775 7.525 1.945 7.695 ;
        RECT 2.495 7.525 2.665 7.695 ;
        RECT 2.855 7.525 3.025 7.695 ;
        RECT 3.215 7.525 3.385 7.695 ;
        RECT 3.575 7.525 3.745 7.695 ;
        RECT 4.025 7.525 4.195 7.695 ;
        RECT 4.385 7.525 4.555 7.695 ;
        RECT 4.745 7.525 4.915 7.695 ;
        RECT 5.105 7.525 5.275 7.695 ;
        RECT 5.825 7.525 5.995 7.695 ;
        RECT 6.185 7.525 6.355 7.695 ;
        RECT 6.545 7.525 6.715 7.695 ;
        RECT 6.905 7.525 7.075 7.695 ;
        RECT 7.355 7.525 7.525 7.695 ;
        RECT 7.715 7.525 7.885 7.695 ;
        RECT 8.075 7.525 8.245 7.695 ;
        RECT 8.435 7.525 8.605 7.695 ;
        RECT 9.155 7.525 9.325 7.695 ;
        RECT 9.515 7.525 9.685 7.695 ;
        RECT 9.905 7.525 10.075 7.695 ;
        RECT 10.295 7.525 10.465 7.695 ;
        RECT 10.655 7.525 10.825 7.695 ;
        RECT 11.375 7.525 11.545 7.695 ;
        RECT 11.735 7.525 11.905 7.695 ;
        RECT 12.125 7.525 12.295 7.695 ;
        RECT 12.515 7.525 12.685 7.695 ;
        RECT 12.875 7.525 13.045 7.695 ;
        RECT 13.595 7.525 13.765 7.695 ;
        RECT 13.955 7.525 14.125 7.695 ;
        RECT 14.315 7.525 14.485 7.695 ;
        RECT 14.675 7.525 14.845 7.695 ;
        RECT 15.125 7.525 15.295 7.695 ;
        RECT 15.485 7.525 15.655 7.695 ;
        RECT 15.845 7.525 16.015 7.695 ;
        RECT 16.205 7.525 16.375 7.695 ;
        RECT 16.925 7.525 17.095 7.695 ;
        RECT 17.285 7.525 17.455 7.695 ;
        RECT 17.645 7.525 17.815 7.695 ;
        RECT 18.005 7.525 18.175 7.695 ;
        RECT 18.455 7.525 18.625 7.695 ;
        RECT 18.815 7.525 18.985 7.695 ;
        RECT 19.175 7.525 19.345 7.695 ;
        RECT 19.535 7.525 19.705 7.695 ;
        RECT 20.255 7.525 20.425 7.695 ;
        RECT 20.615 7.525 20.785 7.695 ;
        RECT 21.005 7.525 21.175 7.695 ;
        RECT 21.395 7.525 21.565 7.695 ;
        RECT 21.755 7.525 21.925 7.695 ;
        RECT 22.475 7.525 22.645 7.695 ;
        RECT 22.835 7.525 23.005 7.695 ;
        RECT 23.195 7.525 23.365 7.695 ;
        RECT 23.555 7.525 23.725 7.695 ;
        RECT 24.005 7.525 24.175 7.695 ;
        RECT 24.365 7.525 24.535 7.695 ;
        RECT 24.725 7.525 24.895 7.695 ;
        RECT 25.085 7.525 25.255 7.695 ;
        RECT 25.805 7.525 25.975 7.695 ;
        RECT 26.165 7.525 26.335 7.695 ;
        RECT 26.555 7.525 26.725 7.695 ;
        RECT 26.945 7.525 27.115 7.695 ;
        RECT 27.305 7.525 27.475 7.695 ;
        RECT 28.025 7.525 28.195 7.695 ;
        RECT 28.385 7.525 28.555 7.695 ;
        RECT 28.745 7.525 28.915 7.695 ;
        RECT 29.105 7.525 29.275 7.695 ;
        RECT 29.555 7.525 29.725 7.695 ;
        RECT 29.915 7.525 30.085 7.695 ;
        RECT 30.275 7.525 30.445 7.695 ;
        RECT 30.635 7.525 30.805 7.695 ;
        RECT 31.355 7.525 31.525 7.695 ;
        RECT 31.715 7.525 31.885 7.695 ;
        RECT 32.105 7.525 32.275 7.695 ;
        RECT 32.495 7.525 32.665 7.695 ;
        RECT 32.855 7.525 33.025 7.695 ;
        RECT 33.575 7.525 33.745 7.695 ;
        RECT 33.935 7.525 34.105 7.695 ;
        RECT 34.295 7.525 34.465 7.695 ;
        RECT 34.655 7.525 34.825 7.695 ;
        RECT 35.105 7.525 35.275 7.695 ;
        RECT 35.465 7.525 35.635 7.695 ;
        RECT 35.825 7.525 35.995 7.695 ;
        RECT 36.185 7.525 36.355 7.695 ;
        RECT 36.905 7.525 37.075 7.695 ;
        RECT 37.265 7.525 37.435 7.695 ;
        RECT 37.655 7.525 37.825 7.695 ;
        RECT 38.045 7.525 38.215 7.695 ;
        RECT 38.405 7.525 38.575 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 39.005 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 41.014198 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 39.135 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 1.935 -0.075 2.505 -0.065 ;
        RECT 5.265 -0.075 5.835 -0.065 ;
        RECT 8.595 -0.075 9.165 -0.065 ;
        RECT 10.815 -0.075 11.385 -0.065 ;
        RECT 13.035 -0.075 13.605 -0.065 ;
        RECT 16.365 -0.075 16.935 -0.065 ;
        RECT 19.695 -0.075 20.265 -0.065 ;
        RECT 21.915 -0.075 22.485 -0.065 ;
        RECT 25.245 -0.075 25.815 -0.065 ;
        RECT 27.465 -0.075 28.035 -0.065 ;
        RECT 30.795 -0.075 31.365 -0.065 ;
        RECT 33.015 -0.075 33.585 -0.065 ;
        RECT 36.345 -0.075 36.915 -0.065 ;
        RECT 38.565 -0.075 39.135 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 0.545 0.755 0.715 1.885 ;
        RECT 1.515 0.755 1.685 1.885 ;
        RECT 0.545 0.585 1.685 0.755 ;
        RECT 0.545 0.310 0.715 0.585 ;
        RECT 1.030 0.310 1.200 0.585 ;
        RECT 1.515 0.310 1.685 0.585 ;
        RECT 2.065 0.310 2.375 2.860 ;
        RECT 3.315 0.310 3.485 1.260 ;
        RECT 5.395 0.310 5.705 2.860 ;
        RECT 6.645 0.310 6.815 1.260 ;
        RECT 8.725 0.310 9.035 2.860 ;
        RECT 9.415 0.755 9.585 1.885 ;
        RECT 10.385 0.755 10.555 1.885 ;
        RECT 9.415 0.585 10.555 0.755 ;
        RECT 9.415 0.310 9.585 0.585 ;
        RECT 9.900 0.310 10.070 0.585 ;
        RECT 10.385 0.310 10.555 0.585 ;
        RECT 10.945 0.310 11.255 2.860 ;
        RECT 11.645 0.755 11.815 1.885 ;
        RECT 12.615 0.755 12.785 1.885 ;
        RECT 11.645 0.585 12.785 0.755 ;
        RECT 11.645 0.310 11.815 0.585 ;
        RECT 12.130 0.310 12.300 0.585 ;
        RECT 12.615 0.310 12.785 0.585 ;
        RECT 13.165 0.310 13.475 2.860 ;
        RECT 14.415 0.310 14.585 1.260 ;
        RECT 16.495 0.310 16.805 2.860 ;
        RECT 17.745 0.310 17.915 1.260 ;
        RECT 19.825 0.310 20.135 2.860 ;
        RECT 20.515 0.755 20.685 1.885 ;
        RECT 21.485 0.755 21.655 1.885 ;
        RECT 20.515 0.585 21.655 0.755 ;
        RECT 20.515 0.310 20.685 0.585 ;
        RECT 21.000 0.310 21.170 0.585 ;
        RECT 21.485 0.310 21.655 0.585 ;
        RECT 22.045 0.310 22.355 2.860 ;
        RECT 23.295 0.310 23.465 1.260 ;
        RECT 25.375 0.310 25.685 2.860 ;
        RECT 26.075 0.755 26.245 1.885 ;
        RECT 27.045 0.755 27.215 1.885 ;
        RECT 26.075 0.585 27.215 0.755 ;
        RECT 26.075 0.310 26.245 0.585 ;
        RECT 26.560 0.310 26.730 0.585 ;
        RECT 27.045 0.310 27.215 0.585 ;
        RECT 27.595 0.310 27.905 2.860 ;
        RECT 28.845 0.310 29.015 1.260 ;
        RECT 30.925 0.310 31.235 2.860 ;
        RECT 31.625 0.755 31.795 1.885 ;
        RECT 32.595 0.755 32.765 1.885 ;
        RECT 31.625 0.585 32.765 0.755 ;
        RECT 31.625 0.310 31.795 0.585 ;
        RECT 32.110 0.310 32.280 0.585 ;
        RECT 32.595 0.310 32.765 0.585 ;
        RECT 33.145 0.310 33.455 2.860 ;
        RECT 33.910 0.755 34.080 1.885 ;
        RECT 34.880 0.755 35.050 1.530 ;
        RECT 35.850 0.755 36.020 1.530 ;
        RECT 33.910 0.585 36.020 0.755 ;
        RECT 33.910 0.310 34.080 0.585 ;
        RECT 34.395 0.310 34.565 0.585 ;
        RECT 34.880 0.310 35.050 0.585 ;
        RECT 35.365 0.310 35.535 0.585 ;
        RECT 35.850 0.310 36.020 0.585 ;
        RECT 36.475 0.310 36.785 2.860 ;
        RECT 37.175 0.755 37.345 1.885 ;
        RECT 38.145 0.755 38.315 1.885 ;
        RECT 37.175 0.585 38.315 0.755 ;
        RECT 37.175 0.310 37.345 0.585 ;
        RECT 37.660 0.310 37.830 0.585 ;
        RECT 38.145 0.310 38.315 0.585 ;
        RECT 38.695 0.310 39.005 2.860 ;
        RECT -0.155 0.000 39.005 0.310 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 1.025 0.065 1.195 0.235 ;
        RECT 1.415 0.065 1.585 0.235 ;
        RECT 1.775 0.065 1.945 0.235 ;
        RECT 2.495 0.065 2.665 0.235 ;
        RECT 2.855 0.065 3.025 0.235 ;
        RECT 3.215 0.065 3.385 0.235 ;
        RECT 3.575 0.065 3.745 0.235 ;
        RECT 4.025 0.065 4.195 0.235 ;
        RECT 4.385 0.065 4.555 0.235 ;
        RECT 4.745 0.065 4.915 0.235 ;
        RECT 5.105 0.065 5.275 0.235 ;
        RECT 5.825 0.065 5.995 0.235 ;
        RECT 6.185 0.065 6.355 0.235 ;
        RECT 6.545 0.065 6.715 0.235 ;
        RECT 6.905 0.065 7.075 0.235 ;
        RECT 7.355 0.065 7.525 0.235 ;
        RECT 7.715 0.065 7.885 0.235 ;
        RECT 8.075 0.065 8.245 0.235 ;
        RECT 8.435 0.065 8.605 0.235 ;
        RECT 9.155 0.065 9.325 0.235 ;
        RECT 9.515 0.065 9.685 0.235 ;
        RECT 9.905 0.065 10.075 0.235 ;
        RECT 10.295 0.065 10.465 0.235 ;
        RECT 10.655 0.065 10.825 0.235 ;
        RECT 11.375 0.065 11.545 0.235 ;
        RECT 11.735 0.065 11.905 0.235 ;
        RECT 12.125 0.065 12.295 0.235 ;
        RECT 12.515 0.065 12.685 0.235 ;
        RECT 12.875 0.065 13.045 0.235 ;
        RECT 13.595 0.065 13.765 0.235 ;
        RECT 13.955 0.065 14.125 0.235 ;
        RECT 14.315 0.065 14.485 0.235 ;
        RECT 14.675 0.065 14.845 0.235 ;
        RECT 15.125 0.065 15.295 0.235 ;
        RECT 15.485 0.065 15.655 0.235 ;
        RECT 15.845 0.065 16.015 0.235 ;
        RECT 16.205 0.065 16.375 0.235 ;
        RECT 16.925 0.065 17.095 0.235 ;
        RECT 17.285 0.065 17.455 0.235 ;
        RECT 17.645 0.065 17.815 0.235 ;
        RECT 18.005 0.065 18.175 0.235 ;
        RECT 18.455 0.065 18.625 0.235 ;
        RECT 18.815 0.065 18.985 0.235 ;
        RECT 19.175 0.065 19.345 0.235 ;
        RECT 19.535 0.065 19.705 0.235 ;
        RECT 20.255 0.065 20.425 0.235 ;
        RECT 20.615 0.065 20.785 0.235 ;
        RECT 21.005 0.065 21.175 0.235 ;
        RECT 21.395 0.065 21.565 0.235 ;
        RECT 21.755 0.065 21.925 0.235 ;
        RECT 22.475 0.065 22.645 0.235 ;
        RECT 22.835 0.065 23.005 0.235 ;
        RECT 23.195 0.065 23.365 0.235 ;
        RECT 23.555 0.065 23.725 0.235 ;
        RECT 24.005 0.065 24.175 0.235 ;
        RECT 24.365 0.065 24.535 0.235 ;
        RECT 24.725 0.065 24.895 0.235 ;
        RECT 25.085 0.065 25.255 0.235 ;
        RECT 25.805 0.065 25.975 0.235 ;
        RECT 26.165 0.065 26.335 0.235 ;
        RECT 26.555 0.065 26.725 0.235 ;
        RECT 26.945 0.065 27.115 0.235 ;
        RECT 27.305 0.065 27.475 0.235 ;
        RECT 28.025 0.065 28.195 0.235 ;
        RECT 28.385 0.065 28.555 0.235 ;
        RECT 28.745 0.065 28.915 0.235 ;
        RECT 29.105 0.065 29.275 0.235 ;
        RECT 29.555 0.065 29.725 0.235 ;
        RECT 29.915 0.065 30.085 0.235 ;
        RECT 30.275 0.065 30.445 0.235 ;
        RECT 30.635 0.065 30.805 0.235 ;
        RECT 31.355 0.065 31.525 0.235 ;
        RECT 31.715 0.065 31.885 0.235 ;
        RECT 32.105 0.065 32.275 0.235 ;
        RECT 32.495 0.065 32.665 0.235 ;
        RECT 32.855 0.065 33.025 0.235 ;
        RECT 33.575 0.065 33.745 0.235 ;
        RECT 33.935 0.065 34.105 0.235 ;
        RECT 34.295 0.065 34.465 0.235 ;
        RECT 34.655 0.065 34.825 0.235 ;
        RECT 35.105 0.065 35.275 0.235 ;
        RECT 35.465 0.065 35.635 0.235 ;
        RECT 35.825 0.065 35.995 0.235 ;
        RECT 36.185 0.065 36.355 0.235 ;
        RECT 36.905 0.065 37.075 0.235 ;
        RECT 37.265 0.065 37.435 0.235 ;
        RECT 37.655 0.065 37.825 0.235 ;
        RECT 38.045 0.065 38.215 0.235 ;
        RECT 38.405 0.065 38.575 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 39.005 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 1.025 4.895 1.195 7.250 ;
        RECT 2.925 5.525 3.095 7.135 ;
        RECT 3.805 7.055 4.855 7.225 ;
        RECT 3.805 5.525 3.975 7.055 ;
        RECT 2.925 5.355 3.975 5.525 ;
        RECT 4.245 5.525 4.415 6.795 ;
        RECT 4.685 5.785 4.855 7.055 ;
        RECT 6.255 5.525 6.425 7.135 ;
        RECT 7.135 7.055 8.185 7.225 ;
        RECT 7.135 5.525 7.305 7.055 ;
        RECT 4.245 5.355 4.895 5.525 ;
        RECT 6.255 5.355 7.305 5.525 ;
        RECT 7.575 5.525 7.745 6.795 ;
        RECT 8.015 5.785 8.185 7.055 ;
        RECT 7.575 5.355 8.225 5.525 ;
        RECT 1.025 4.725 1.565 4.895 ;
        RECT 1.395 2.305 1.565 4.725 ;
        RECT 4.355 3.905 4.525 5.100 ;
        RECT 1.025 2.135 1.565 2.305 ;
        RECT 1.025 0.975 1.195 2.135 ;
        RECT 2.830 1.805 3.000 1.885 ;
        RECT 3.800 1.805 3.970 1.885 ;
        RECT 4.725 1.875 4.895 5.355 ;
        RECT 6.575 2.055 6.745 3.125 ;
        RECT 7.685 2.055 7.855 5.100 ;
        RECT 2.830 1.635 3.970 1.805 ;
        RECT 2.830 0.505 3.000 1.635 ;
        RECT 3.800 0.755 3.970 1.635 ;
        RECT 4.285 1.705 4.895 1.875 ;
        RECT 6.160 1.805 6.330 1.885 ;
        RECT 7.130 1.805 7.300 1.885 ;
        RECT 8.055 1.875 8.225 5.355 ;
        RECT 9.905 4.895 10.075 7.250 ;
        RECT 9.535 4.725 10.075 4.895 ;
        RECT 9.535 2.305 9.705 4.725 ;
        RECT 9.535 2.135 10.075 2.305 ;
        RECT 4.285 0.975 4.455 1.705 ;
        RECT 6.160 1.635 7.300 1.805 ;
        RECT 4.770 0.755 4.940 1.525 ;
        RECT 3.800 0.585 4.940 0.755 ;
        RECT 3.800 0.505 3.970 0.585 ;
        RECT 4.770 0.505 4.940 0.585 ;
        RECT 6.160 0.505 6.330 1.635 ;
        RECT 7.130 0.755 7.300 1.635 ;
        RECT 7.615 1.705 8.225 1.875 ;
        RECT 7.615 0.975 7.785 1.705 ;
        RECT 8.100 0.755 8.270 1.525 ;
        RECT 9.905 0.975 10.075 2.135 ;
        RECT 11.755 2.055 11.925 5.095 ;
        RECT 12.125 4.895 12.295 7.250 ;
        RECT 14.025 5.525 14.195 7.135 ;
        RECT 14.905 7.055 15.955 7.225 ;
        RECT 14.905 5.525 15.075 7.055 ;
        RECT 15.785 5.785 15.955 7.055 ;
        RECT 14.025 5.355 15.075 5.525 ;
        RECT 17.355 5.525 17.525 7.135 ;
        RECT 18.235 7.055 19.285 7.225 ;
        RECT 18.235 5.525 18.405 7.055 ;
        RECT 19.115 5.785 19.285 7.055 ;
        RECT 17.355 5.355 18.405 5.525 ;
        RECT 12.125 4.725 12.665 4.895 ;
        RECT 12.495 2.305 12.665 4.725 ;
        RECT 12.125 2.135 12.665 2.305 ;
        RECT 12.125 0.975 12.295 2.135 ;
        RECT 14.345 2.055 14.515 5.100 ;
        RECT 15.455 3.905 15.625 5.100 ;
        RECT 17.675 2.055 17.845 3.125 ;
        RECT 18.785 2.055 18.955 5.100 ;
        RECT 21.005 4.895 21.175 7.250 ;
        RECT 23.345 5.515 23.515 7.250 ;
        RECT 24.225 5.515 24.395 7.250 ;
        RECT 23.345 5.345 24.875 5.515 ;
        RECT 23.995 4.940 24.165 5.095 ;
        RECT 20.635 4.725 21.175 4.895 ;
        RECT 23.965 4.765 24.165 4.940 ;
        RECT 20.635 2.305 20.805 4.725 ;
        RECT 20.635 2.135 21.175 2.305 ;
        RECT 13.930 1.805 14.100 1.885 ;
        RECT 14.900 1.805 15.070 1.885 ;
        RECT 13.930 1.635 15.070 1.805 ;
        RECT 7.130 0.585 8.270 0.755 ;
        RECT 7.130 0.505 7.300 0.585 ;
        RECT 8.100 0.505 8.270 0.585 ;
        RECT 13.930 0.505 14.100 1.635 ;
        RECT 14.900 0.755 15.070 1.635 ;
        RECT 17.260 1.805 17.430 1.885 ;
        RECT 18.230 1.805 18.400 1.885 ;
        RECT 17.260 1.635 18.400 1.805 ;
        RECT 15.870 0.755 16.040 1.525 ;
        RECT 14.900 0.585 16.040 0.755 ;
        RECT 14.900 0.505 15.070 0.585 ;
        RECT 15.870 0.505 16.040 0.585 ;
        RECT 17.260 0.505 17.430 1.635 ;
        RECT 18.230 0.755 18.400 1.635 ;
        RECT 19.200 0.755 19.370 1.525 ;
        RECT 21.005 0.975 21.175 2.135 ;
        RECT 23.965 2.055 24.135 4.765 ;
        RECT 22.810 1.805 22.980 1.885 ;
        RECT 23.780 1.805 23.950 1.885 ;
        RECT 24.705 1.880 24.875 5.345 ;
        RECT 26.185 2.055 26.355 5.095 ;
        RECT 26.555 4.895 26.725 7.250 ;
        RECT 28.895 5.515 29.065 7.250 ;
        RECT 29.775 5.515 29.945 7.250 ;
        RECT 28.895 5.345 30.425 5.515 ;
        RECT 26.555 4.725 27.095 4.895 ;
        RECT 26.925 2.305 27.095 4.725 ;
        RECT 26.555 2.135 27.095 2.305 ;
        RECT 22.810 1.635 23.950 1.805 ;
        RECT 18.230 0.585 19.370 0.755 ;
        RECT 18.230 0.505 18.400 0.585 ;
        RECT 19.200 0.505 19.370 0.585 ;
        RECT 22.810 0.505 22.980 1.635 ;
        RECT 23.780 0.755 23.950 1.635 ;
        RECT 24.265 1.710 24.875 1.880 ;
        RECT 24.265 0.975 24.435 1.710 ;
        RECT 24.750 0.755 24.920 1.525 ;
        RECT 26.555 0.975 26.725 2.135 ;
        RECT 28.360 1.805 28.530 1.885 ;
        RECT 29.330 1.805 29.500 1.885 ;
        RECT 30.255 1.880 30.425 5.345 ;
        RECT 31.735 2.055 31.905 5.095 ;
        RECT 32.105 4.895 32.275 7.250 ;
        RECT 34.005 5.525 34.175 7.255 ;
        RECT 34.885 7.055 35.935 7.225 ;
        RECT 34.885 5.525 35.055 7.055 ;
        RECT 34.005 5.355 35.055 5.525 ;
        RECT 35.325 5.525 35.495 6.795 ;
        RECT 35.765 5.785 35.935 7.055 ;
        RECT 35.325 5.355 35.975 5.525 ;
        RECT 34.170 4.940 34.340 5.100 ;
        RECT 35.100 4.940 35.270 5.100 ;
        RECT 32.105 4.725 32.645 4.895 ;
        RECT 34.170 4.770 34.495 4.940 ;
        RECT 32.475 2.305 32.645 4.725 ;
        RECT 32.105 2.135 32.645 2.305 ;
        RECT 28.360 1.635 29.500 1.805 ;
        RECT 23.780 0.585 24.920 0.755 ;
        RECT 23.780 0.505 23.950 0.585 ;
        RECT 24.750 0.505 24.920 0.585 ;
        RECT 28.360 0.505 28.530 1.635 ;
        RECT 29.330 0.755 29.500 1.635 ;
        RECT 29.815 1.710 30.425 1.880 ;
        RECT 29.815 0.975 29.985 1.710 ;
        RECT 30.300 0.755 30.470 1.525 ;
        RECT 32.105 0.975 32.275 2.135 ;
        RECT 34.325 2.055 34.495 4.770 ;
        RECT 35.065 4.770 35.270 4.940 ;
        RECT 35.065 2.055 35.235 4.770 ;
        RECT 35.805 1.880 35.975 5.355 ;
        RECT 37.285 2.055 37.455 5.095 ;
        RECT 34.395 1.710 35.975 1.880 ;
        RECT 34.395 0.975 34.565 1.710 ;
        RECT 35.365 0.975 35.535 1.710 ;
        RECT 29.330 0.585 30.470 0.755 ;
        RECT 29.330 0.505 29.500 0.585 ;
        RECT 30.300 0.505 30.470 0.585 ;
      LAYER mcon ;
        RECT 4.355 3.985 4.525 4.155 ;
        RECT 1.395 3.245 1.565 3.415 ;
        RECT 4.725 3.615 4.895 3.785 ;
        RECT 7.685 3.245 7.855 3.415 ;
        RECT 6.575 2.875 6.745 3.045 ;
        RECT 8.055 3.615 8.225 3.785 ;
        RECT 9.535 3.985 9.705 4.155 ;
        RECT 9.535 2.875 9.705 3.045 ;
        RECT 11.755 4.355 11.925 4.525 ;
        RECT 11.755 3.615 11.925 3.785 ;
        RECT 12.495 3.245 12.665 3.415 ;
        RECT 11.755 2.135 11.925 2.305 ;
        RECT 14.345 4.355 14.515 4.525 ;
        RECT 15.455 3.985 15.625 4.155 ;
        RECT 18.785 3.245 18.955 3.415 ;
        RECT 17.675 2.875 17.845 3.045 ;
        RECT 20.635 3.985 20.805 4.155 ;
        RECT 20.635 2.875 20.805 3.045 ;
        RECT 23.965 2.135 24.135 2.305 ;
        RECT 24.705 3.245 24.875 3.415 ;
        RECT 26.185 3.245 26.355 3.415 ;
        RECT 26.925 2.875 27.095 3.045 ;
        RECT 30.255 3.245 30.425 3.415 ;
        RECT 31.735 3.245 31.905 3.415 ;
        RECT 32.475 3.245 32.645 3.415 ;
        RECT 34.325 2.875 34.495 3.045 ;
        RECT 35.065 3.245 35.235 3.415 ;
        RECT 35.805 3.245 35.975 3.415 ;
        RECT 37.285 3.245 37.455 3.415 ;
      LAYER met1 ;
        RECT 11.725 4.525 11.955 4.555 ;
        RECT 14.315 4.525 14.545 4.555 ;
        RECT 11.695 4.355 14.575 4.525 ;
        RECT 11.725 4.325 11.955 4.355 ;
        RECT 14.315 4.325 14.545 4.355 ;
        RECT 4.325 4.155 4.555 4.185 ;
        RECT 9.505 4.155 9.735 4.185 ;
        RECT 15.425 4.155 15.655 4.185 ;
        RECT 20.605 4.155 20.835 4.185 ;
        RECT 4.295 3.985 9.765 4.155 ;
        RECT 15.395 3.985 20.865 4.155 ;
        RECT 4.325 3.955 4.555 3.985 ;
        RECT 9.505 3.955 9.735 3.985 ;
        RECT 15.425 3.955 15.655 3.985 ;
        RECT 20.605 3.955 20.835 3.985 ;
        RECT 4.695 3.785 4.925 3.815 ;
        RECT 8.025 3.785 8.255 3.815 ;
        RECT 11.725 3.785 11.955 3.815 ;
        RECT 4.665 3.615 11.985 3.785 ;
        RECT 4.695 3.585 4.925 3.615 ;
        RECT 8.025 3.585 8.255 3.615 ;
        RECT 11.725 3.585 11.955 3.615 ;
        RECT 1.365 3.415 1.595 3.445 ;
        RECT 7.655 3.415 7.885 3.445 ;
        RECT 12.465 3.415 12.695 3.445 ;
        RECT 18.755 3.415 18.985 3.445 ;
        RECT 24.675 3.415 24.905 3.445 ;
        RECT 26.155 3.415 26.385 3.445 ;
        RECT 30.225 3.415 30.455 3.445 ;
        RECT 31.705 3.415 31.935 3.445 ;
        RECT 32.445 3.415 32.675 3.445 ;
        RECT 35.035 3.415 35.265 3.445 ;
        RECT 35.775 3.415 36.005 3.445 ;
        RECT 37.255 3.415 37.485 3.445 ;
        RECT 1.335 3.245 7.915 3.415 ;
        RECT 12.435 3.245 19.015 3.415 ;
        RECT 24.645 3.245 26.415 3.415 ;
        RECT 30.195 3.245 31.965 3.415 ;
        RECT 32.415 3.245 35.295 3.415 ;
        RECT 35.745 3.245 37.515 3.415 ;
        RECT 1.365 3.215 1.595 3.245 ;
        RECT 7.655 3.215 7.885 3.245 ;
        RECT 12.465 3.215 12.695 3.245 ;
        RECT 18.755 3.215 18.985 3.245 ;
        RECT 24.675 3.215 24.905 3.245 ;
        RECT 26.155 3.215 26.385 3.245 ;
        RECT 30.225 3.215 30.455 3.245 ;
        RECT 31.705 3.215 31.935 3.245 ;
        RECT 32.445 3.215 32.675 3.245 ;
        RECT 35.035 3.215 35.265 3.245 ;
        RECT 35.775 3.215 36.005 3.245 ;
        RECT 37.255 3.215 37.485 3.245 ;
        RECT 6.545 3.045 6.775 3.075 ;
        RECT 9.505 3.045 9.735 3.075 ;
        RECT 17.645 3.045 17.875 3.075 ;
        RECT 20.605 3.045 20.835 3.075 ;
        RECT 26.895 3.045 27.125 3.075 ;
        RECT 34.295 3.045 34.525 3.075 ;
        RECT 6.515 2.875 9.765 3.045 ;
        RECT 17.615 2.875 20.865 3.045 ;
        RECT 26.865 2.875 34.555 3.045 ;
        RECT 6.545 2.845 6.775 2.875 ;
        RECT 9.505 2.845 9.735 2.875 ;
        RECT 17.645 2.845 17.875 2.875 ;
        RECT 20.605 2.845 20.835 2.875 ;
        RECT 26.895 2.845 27.125 2.875 ;
        RECT 34.295 2.845 34.525 2.875 ;
        RECT 11.725 2.305 11.955 2.335 ;
        RECT 23.935 2.305 24.165 2.335 ;
        RECT 11.695 2.135 24.195 2.305 ;
        RECT 11.725 2.105 11.955 2.135 ;
        RECT 23.935 2.105 24.165 2.135 ;
  END
END FA






MACRO FILL1
  CLASS BLOCK ;
  FOREIGN FILL1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 1.580 BY 7.950 ;
  OBS
      LAYER nwell ;
        RECT -0.420 4.160 1.160 7.875 ;
      LAYER pwell ;
        RECT -0.285 -0.075 1.025 2.990 ;
      LAYER li1 ;
        RECT -0.155 7.460 0.895 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 0.585 4.340 0.895 7.460 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 0.585 0.310 0.895 2.860 ;
        RECT -0.155 0.000 0.895 0.310 ;
      LAYER met1 ;
        RECT -0.155 7.460 0.895 7.770 ;
        RECT -0.155 0.000 0.895 0.310 ;
  END
END FILL1






MACRO HA
  CLASS BLOCK ;
  FOREIGN HA ;
  ORIGIN 0.420 0.075 ;
  SIZE 17.490 BY 7.950 ;
  PIN SUM
    ANTENNADIFFAREA 1.543800 ;
    PORT
      LAYER li1 ;
        RECT 9.795 5.525 9.965 6.795 ;
        RECT 13.125 5.525 13.295 6.795 ;
        RECT 9.795 5.355 10.445 5.525 ;
        RECT 13.125 5.355 13.775 5.525 ;
        RECT 10.275 1.875 10.445 5.355 ;
        RECT 13.605 1.875 13.775 5.355 ;
        RECT 9.835 1.705 10.445 1.875 ;
        RECT 13.165 1.705 13.775 1.875 ;
        RECT 9.835 0.975 10.005 1.705 ;
        RECT 13.165 0.975 13.335 1.705 ;
      LAYER mcon ;
        RECT 10.275 3.615 10.445 3.785 ;
        RECT 13.605 3.615 13.775 3.785 ;
      LAYER met1 ;
        RECT 10.245 3.785 10.475 3.815 ;
        RECT 13.575 3.785 13.805 3.815 ;
        RECT 10.215 3.615 13.835 3.785 ;
        RECT 10.245 3.585 10.475 3.615 ;
        RECT 13.575 3.585 13.805 3.615 ;
    END
  END SUM
  PIN COUT
    ANTENNADIFFAREA 0.771900 ;
    PORT
      LAYER li1 ;
        RECT 4.355 4.895 4.525 7.250 ;
        RECT 4.355 4.725 4.895 4.895 ;
        RECT 4.725 2.305 4.895 4.725 ;
        RECT 4.355 2.135 4.895 2.305 ;
        RECT 4.355 0.975 4.525 2.135 ;
      LAYER mcon ;
        RECT 4.725 2.875 4.895 3.045 ;
      LAYER met1 ;
        RECT 4.695 3.045 4.925 3.075 ;
        RECT 4.545 2.875 4.955 3.045 ;
        RECT 4.695 2.845 4.925 2.875 ;
    END
  END COUT
  PIN A
    ANTENNAGATEAREA 3.093750 ;
    PORT
      LAYER li1 ;
        RECT 1.025 2.055 1.195 5.095 ;
        RECT 6.205 2.055 6.375 5.095 ;
        RECT 8.795 2.055 8.965 5.100 ;
      LAYER mcon ;
        RECT 1.025 4.355 1.195 4.525 ;
        RECT 6.205 4.355 6.375 4.525 ;
        RECT 8.795 4.355 8.965 4.525 ;
      LAYER met1 ;
        RECT 0.995 4.525 1.225 4.555 ;
        RECT 6.175 4.525 6.405 4.555 ;
        RECT 8.765 4.525 8.995 4.555 ;
        RECT 0.965 4.355 9.025 4.525 ;
        RECT 0.995 4.325 1.225 4.355 ;
        RECT 6.175 4.325 6.405 4.355 ;
        RECT 8.765 4.325 8.995 4.355 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 3.081750 ;
    PORT
      LAYER li1 ;
        RECT 1.795 4.940 1.965 5.095 ;
        RECT 1.765 4.765 1.965 4.940 ;
        RECT 1.765 2.055 1.935 4.765 ;
        RECT 9.535 3.535 9.705 4.605 ;
        RECT 12.125 4.275 12.295 5.100 ;
        RECT 9.905 2.055 10.075 2.755 ;
        RECT 15.825 2.055 15.995 5.095 ;
      LAYER mcon ;
        RECT 1.765 3.615 1.935 3.785 ;
        RECT 9.535 4.355 9.705 4.525 ;
        RECT 12.125 4.355 12.295 4.525 ;
        RECT 15.825 4.355 15.995 4.525 ;
        RECT 9.535 3.615 9.705 3.785 ;
        RECT 9.905 2.505 10.075 2.675 ;
        RECT 15.825 2.505 15.995 2.675 ;
      LAYER met1 ;
        RECT 9.505 4.525 9.735 4.555 ;
        RECT 12.095 4.525 12.325 4.555 ;
        RECT 15.795 4.525 16.025 4.555 ;
        RECT 9.475 4.355 16.055 4.525 ;
        RECT 9.505 4.325 9.735 4.355 ;
        RECT 12.095 4.325 12.325 4.355 ;
        RECT 15.795 4.325 16.025 4.355 ;
        RECT 1.735 3.785 1.965 3.815 ;
        RECT 9.505 3.785 9.735 3.815 ;
        RECT 1.705 3.615 9.765 3.785 ;
        RECT 1.735 3.585 1.965 3.615 ;
        RECT 9.505 3.585 9.735 3.615 ;
        RECT 9.875 2.675 10.105 2.705 ;
        RECT 15.795 2.675 16.025 2.705 ;
        RECT 9.845 2.505 16.055 2.675 ;
        RECT 9.875 2.475 10.105 2.505 ;
        RECT 15.795 2.475 16.025 2.505 ;
    END
  END B
  PIN VDD
    ANTENNADIFFAREA 20.519550 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 17.070 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 16.805 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 0.705 5.365 0.875 7.460 ;
        RECT 1.585 5.785 1.755 7.460 ;
        RECT 2.465 5.785 2.635 7.460 ;
        RECT 3.175 4.340 3.485 7.460 ;
        RECT 3.915 5.415 4.085 7.460 ;
        RECT 4.795 5.415 4.965 7.460 ;
        RECT 5.395 4.340 5.705 7.460 ;
        RECT 6.135 5.415 6.305 7.460 ;
        RECT 7.015 5.415 7.185 7.460 ;
        RECT 7.615 4.340 7.925 7.460 ;
        RECT 8.915 5.785 9.085 7.460 ;
        RECT 10.945 4.340 11.255 7.460 ;
        RECT 12.245 5.785 12.415 7.460 ;
        RECT 14.275 4.340 14.585 7.460 ;
        RECT 15.015 5.415 15.185 7.460 ;
        RECT 15.895 5.415 16.065 7.460 ;
        RECT 16.495 4.340 16.805 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 0.995 7.525 1.165 7.695 ;
        RECT 1.355 7.525 1.525 7.695 ;
        RECT 1.805 7.525 1.975 7.695 ;
        RECT 2.165 7.525 2.335 7.695 ;
        RECT 2.525 7.525 2.695 7.695 ;
        RECT 2.885 7.525 3.055 7.695 ;
        RECT 3.605 7.525 3.775 7.695 ;
        RECT 3.965 7.525 4.135 7.695 ;
        RECT 4.355 7.525 4.525 7.695 ;
        RECT 4.745 7.525 4.915 7.695 ;
        RECT 5.105 7.525 5.275 7.695 ;
        RECT 5.825 7.525 5.995 7.695 ;
        RECT 6.185 7.525 6.355 7.695 ;
        RECT 6.575 7.525 6.745 7.695 ;
        RECT 6.965 7.525 7.135 7.695 ;
        RECT 7.325 7.525 7.495 7.695 ;
        RECT 8.045 7.525 8.215 7.695 ;
        RECT 8.405 7.525 8.575 7.695 ;
        RECT 8.765 7.525 8.935 7.695 ;
        RECT 9.125 7.525 9.295 7.695 ;
        RECT 9.575 7.525 9.745 7.695 ;
        RECT 9.935 7.525 10.105 7.695 ;
        RECT 10.295 7.525 10.465 7.695 ;
        RECT 10.655 7.525 10.825 7.695 ;
        RECT 11.375 7.525 11.545 7.695 ;
        RECT 11.735 7.525 11.905 7.695 ;
        RECT 12.095 7.525 12.265 7.695 ;
        RECT 12.455 7.525 12.625 7.695 ;
        RECT 12.905 7.525 13.075 7.695 ;
        RECT 13.265 7.525 13.435 7.695 ;
        RECT 13.625 7.525 13.795 7.695 ;
        RECT 13.985 7.525 14.155 7.695 ;
        RECT 14.705 7.525 14.875 7.695 ;
        RECT 15.065 7.525 15.235 7.695 ;
        RECT 15.455 7.525 15.625 7.695 ;
        RECT 15.845 7.525 16.015 7.695 ;
        RECT 16.205 7.525 16.375 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 16.805 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 17.295000 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 16.935 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 3.045 -0.075 3.615 -0.065 ;
        RECT 5.265 -0.075 5.835 -0.065 ;
        RECT 7.485 -0.075 8.055 -0.065 ;
        RECT 10.815 -0.075 11.385 -0.065 ;
        RECT 14.145 -0.075 14.715 -0.065 ;
        RECT 16.365 -0.075 16.935 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 1.095 0.310 1.265 1.260 ;
        RECT 3.175 0.310 3.485 2.860 ;
        RECT 3.875 0.755 4.045 1.885 ;
        RECT 4.845 0.755 5.015 1.885 ;
        RECT 3.875 0.585 5.015 0.755 ;
        RECT 3.875 0.310 4.045 0.585 ;
        RECT 4.360 0.310 4.530 0.585 ;
        RECT 4.845 0.310 5.015 0.585 ;
        RECT 5.395 0.310 5.705 2.860 ;
        RECT 6.095 0.755 6.265 1.885 ;
        RECT 7.065 0.755 7.235 1.885 ;
        RECT 6.095 0.585 7.235 0.755 ;
        RECT 6.095 0.310 6.265 0.585 ;
        RECT 6.580 0.310 6.750 0.585 ;
        RECT 7.065 0.310 7.235 0.585 ;
        RECT 7.615 0.310 7.925 2.860 ;
        RECT 8.865 0.310 9.035 1.260 ;
        RECT 10.945 0.310 11.255 2.860 ;
        RECT 12.195 0.310 12.365 1.260 ;
        RECT 14.275 0.310 14.585 2.860 ;
        RECT 14.965 0.755 15.135 1.885 ;
        RECT 15.935 0.755 16.105 1.885 ;
        RECT 14.965 0.585 16.105 0.755 ;
        RECT 14.965 0.310 15.135 0.585 ;
        RECT 15.450 0.310 15.620 0.585 ;
        RECT 15.935 0.310 16.105 0.585 ;
        RECT 16.495 0.310 16.805 2.860 ;
        RECT -0.155 0.000 16.805 0.310 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 0.995 0.065 1.165 0.235 ;
        RECT 1.355 0.065 1.525 0.235 ;
        RECT 1.805 0.065 1.975 0.235 ;
        RECT 2.165 0.065 2.335 0.235 ;
        RECT 2.525 0.065 2.695 0.235 ;
        RECT 2.885 0.065 3.055 0.235 ;
        RECT 3.605 0.065 3.775 0.235 ;
        RECT 3.965 0.065 4.135 0.235 ;
        RECT 4.355 0.065 4.525 0.235 ;
        RECT 4.745 0.065 4.915 0.235 ;
        RECT 5.105 0.065 5.275 0.235 ;
        RECT 5.825 0.065 5.995 0.235 ;
        RECT 6.185 0.065 6.355 0.235 ;
        RECT 6.575 0.065 6.745 0.235 ;
        RECT 6.965 0.065 7.135 0.235 ;
        RECT 7.325 0.065 7.495 0.235 ;
        RECT 8.045 0.065 8.215 0.235 ;
        RECT 8.405 0.065 8.575 0.235 ;
        RECT 8.765 0.065 8.935 0.235 ;
        RECT 9.125 0.065 9.295 0.235 ;
        RECT 9.575 0.065 9.745 0.235 ;
        RECT 9.935 0.065 10.105 0.235 ;
        RECT 10.295 0.065 10.465 0.235 ;
        RECT 10.655 0.065 10.825 0.235 ;
        RECT 11.375 0.065 11.545 0.235 ;
        RECT 11.735 0.065 11.905 0.235 ;
        RECT 12.095 0.065 12.265 0.235 ;
        RECT 12.455 0.065 12.625 0.235 ;
        RECT 12.905 0.065 13.075 0.235 ;
        RECT 13.265 0.065 13.435 0.235 ;
        RECT 13.625 0.065 13.795 0.235 ;
        RECT 13.985 0.065 14.155 0.235 ;
        RECT 14.705 0.065 14.875 0.235 ;
        RECT 15.065 0.065 15.235 0.235 ;
        RECT 15.455 0.065 15.625 0.235 ;
        RECT 15.845 0.065 16.015 0.235 ;
        RECT 16.205 0.065 16.375 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 16.805 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 1.145 5.515 1.315 7.250 ;
        RECT 2.025 5.515 2.195 7.250 ;
        RECT 1.145 5.345 2.675 5.515 ;
        RECT 0.610 1.805 0.780 1.885 ;
        RECT 1.580 1.805 1.750 1.885 ;
        RECT 2.505 1.880 2.675 5.345 ;
        RECT 3.985 2.055 4.155 5.095 ;
        RECT 6.575 4.895 6.745 7.250 ;
        RECT 8.475 5.525 8.645 7.135 ;
        RECT 9.355 7.055 10.405 7.225 ;
        RECT 9.355 5.525 9.525 7.055 ;
        RECT 10.235 5.785 10.405 7.055 ;
        RECT 8.475 5.355 9.525 5.525 ;
        RECT 11.805 5.525 11.975 7.135 ;
        RECT 12.685 7.055 13.735 7.225 ;
        RECT 12.685 5.525 12.855 7.055 ;
        RECT 13.565 5.785 13.735 7.055 ;
        RECT 11.805 5.355 12.855 5.525 ;
        RECT 6.575 4.725 7.115 4.895 ;
        RECT 6.945 2.305 7.115 4.725 ;
        RECT 9.905 3.905 10.075 5.100 ;
        RECT 6.575 2.135 7.115 2.305 ;
        RECT 0.610 1.635 1.750 1.805 ;
        RECT 0.610 0.505 0.780 1.635 ;
        RECT 1.580 0.755 1.750 1.635 ;
        RECT 2.065 1.710 2.675 1.880 ;
        RECT 2.065 0.975 2.235 1.710 ;
        RECT 2.550 0.755 2.720 1.525 ;
        RECT 6.575 0.975 6.745 2.135 ;
        RECT 12.125 2.055 12.295 3.125 ;
        RECT 13.235 2.055 13.405 5.100 ;
        RECT 15.455 4.895 15.625 7.250 ;
        RECT 15.085 4.725 15.625 4.895 ;
        RECT 15.085 2.305 15.255 4.725 ;
        RECT 15.085 2.135 15.625 2.305 ;
        RECT 8.380 1.805 8.550 1.885 ;
        RECT 9.350 1.805 9.520 1.885 ;
        RECT 8.380 1.635 9.520 1.805 ;
        RECT 1.580 0.585 2.720 0.755 ;
        RECT 1.580 0.505 1.750 0.585 ;
        RECT 2.550 0.505 2.720 0.585 ;
        RECT 8.380 0.505 8.550 1.635 ;
        RECT 9.350 0.755 9.520 1.635 ;
        RECT 11.710 1.805 11.880 1.885 ;
        RECT 12.680 1.805 12.850 1.885 ;
        RECT 11.710 1.635 12.850 1.805 ;
        RECT 10.320 0.755 10.490 1.525 ;
        RECT 9.350 0.585 10.490 0.755 ;
        RECT 9.350 0.505 9.520 0.585 ;
        RECT 10.320 0.505 10.490 0.585 ;
        RECT 11.710 0.505 11.880 1.635 ;
        RECT 12.680 0.755 12.850 1.635 ;
        RECT 13.650 0.755 13.820 1.525 ;
        RECT 15.455 0.975 15.625 2.135 ;
        RECT 12.680 0.585 13.820 0.755 ;
        RECT 12.680 0.505 12.850 0.585 ;
        RECT 13.650 0.505 13.820 0.585 ;
      LAYER mcon ;
        RECT 2.505 3.245 2.675 3.415 ;
        RECT 3.985 3.245 4.155 3.415 ;
        RECT 9.905 3.985 10.075 4.155 ;
        RECT 6.945 3.245 7.115 3.415 ;
        RECT 13.235 3.245 13.405 3.415 ;
        RECT 12.125 2.875 12.295 3.045 ;
        RECT 15.085 3.985 15.255 4.155 ;
        RECT 15.085 2.875 15.255 3.045 ;
      LAYER met1 ;
        RECT 9.875 4.155 10.105 4.185 ;
        RECT 15.055 4.155 15.285 4.185 ;
        RECT 9.845 3.985 15.315 4.155 ;
        RECT 9.875 3.955 10.105 3.985 ;
        RECT 15.055 3.955 15.285 3.985 ;
        RECT 2.475 3.415 2.705 3.445 ;
        RECT 3.955 3.415 4.185 3.445 ;
        RECT 6.915 3.415 7.145 3.445 ;
        RECT 13.205 3.415 13.435 3.445 ;
        RECT 2.445 3.245 4.215 3.415 ;
        RECT 6.885 3.245 13.465 3.415 ;
        RECT 2.475 3.215 2.705 3.245 ;
        RECT 3.955 3.215 4.185 3.245 ;
        RECT 6.915 3.215 7.145 3.245 ;
        RECT 13.205 3.215 13.435 3.245 ;
        RECT 12.095 3.045 12.325 3.075 ;
        RECT 15.055 3.045 15.285 3.075 ;
        RECT 12.065 2.875 15.315 3.045 ;
        RECT 12.095 2.845 12.325 2.875 ;
        RECT 15.055 2.845 15.285 2.875 ;
  END
END HA






MACRO INVX1
  CLASS BLOCK ;
  FOREIGN INVX1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 3.060 BY 7.950 ;
  PIN Y
    ANTENNADIFFAREA 0.771900 ;
    PORT
      LAYER li1 ;
        RECT 1.025 4.895 1.195 7.250 ;
        RECT 1.025 4.725 1.565 4.895 ;
        RECT 1.395 2.305 1.565 4.725 ;
        RECT 1.025 2.135 1.565 2.305 ;
        RECT 1.025 0.975 1.195 2.135 ;
      LAYER mcon ;
        RECT 1.395 3.245 1.565 3.415 ;
      LAYER met1 ;
        RECT 1.365 3.415 1.595 3.445 ;
        RECT 1.335 3.245 1.745 3.415 ;
        RECT 1.365 3.215 1.595 3.245 ;
    END
  END Y
  PIN A
    ANTENNAGATEAREA 1.027250 ;
    PORT
      LAYER li1 ;
        RECT 0.655 2.055 0.825 5.095 ;
      LAYER mcon ;
        RECT 0.655 3.245 0.825 3.415 ;
      LAYER met1 ;
        RECT 0.625 3.415 0.855 3.445 ;
        RECT 0.475 3.245 0.885 3.415 ;
        RECT 0.625 3.215 0.855 3.245 ;
    END
  END A
  PIN VDD
    ANTENNADIFFAREA 4.096900 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 2.640 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 2.375 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 0.585 5.415 0.755 7.460 ;
        RECT 1.465 5.415 1.635 7.460 ;
        RECT 2.065 4.340 2.375 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 1.025 7.525 1.195 7.695 ;
        RECT 1.415 7.525 1.585 7.695 ;
        RECT 1.775 7.525 1.945 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 2.375 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 3.833650 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 2.505 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 1.935 -0.075 2.505 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 0.545 0.755 0.715 1.885 ;
        RECT 1.515 0.755 1.685 1.885 ;
        RECT 0.545 0.585 1.685 0.755 ;
        RECT 0.545 0.310 0.715 0.585 ;
        RECT 1.030 0.310 1.200 0.585 ;
        RECT 1.515 0.310 1.685 0.585 ;
        RECT 2.065 0.310 2.375 2.860 ;
        RECT -0.155 0.000 2.375 0.310 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 1.025 0.065 1.195 0.235 ;
        RECT 1.415 0.065 1.585 0.235 ;
        RECT 1.775 0.065 1.945 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 2.375 0.310 ;
    END
  END VSS
END INVX1






MACRO Mod4Counter
  CLASS BLOCK ;
  FOREIGN Mod4Counter ;
  ORIGIN 0.420 0.075 ;
  SIZE 43.760 BY 7.950 ;
  PIN y0
    ANTENNAGATEAREA 2.060500 ;
    ANTENNADIFFAREA 1.351900 ;
    PORT
      LAYER li1 ;
        RECT 15.945 5.515 16.115 7.250 ;
        RECT 16.825 5.515 16.995 7.250 ;
        RECT 15.945 5.345 17.475 5.515 ;
        RECT 6.605 4.940 6.775 5.095 ;
        RECT 6.575 4.765 6.775 4.940 ;
        RECT 6.575 2.055 6.745 4.765 ;
        RECT 17.305 1.880 17.475 5.345 ;
        RECT 19.155 2.055 19.325 5.095 ;
        RECT 16.865 1.710 17.475 1.880 ;
        RECT 16.865 0.975 17.035 1.710 ;
      LAYER mcon ;
        RECT 6.575 3.245 6.745 3.415 ;
        RECT 6.575 2.135 6.745 2.305 ;
        RECT 17.305 3.245 17.475 3.415 ;
        RECT 19.155 3.245 19.325 3.415 ;
      LAYER met1 ;
        RECT 6.545 3.415 6.775 3.445 ;
        RECT 17.275 3.415 17.505 3.445 ;
        RECT 19.125 3.415 19.355 3.445 ;
        RECT 6.395 3.245 19.385 3.415 ;
        RECT 6.545 3.215 6.775 3.245 ;
        RECT 17.275 3.215 17.505 3.245 ;
        RECT 19.125 3.215 19.355 3.245 ;
        RECT 6.545 2.305 6.775 2.335 ;
        RECT 6.395 2.135 6.805 2.305 ;
        RECT 6.545 2.105 6.775 2.135 ;
    END
  END y0
  PIN y1
    ANTENNAGATEAREA 2.060500 ;
    ANTENNADIFFAREA 1.351900 ;
    PORT
      LAYER li1 ;
        RECT 37.405 5.515 37.575 7.250 ;
        RECT 38.285 5.515 38.455 7.250 ;
        RECT 37.405 5.345 38.935 5.515 ;
        RECT 28.065 4.940 28.235 5.095 ;
        RECT 28.035 4.765 28.235 4.940 ;
        RECT 28.035 2.055 28.205 4.765 ;
        RECT 38.765 1.880 38.935 5.345 ;
        RECT 40.615 2.055 40.785 5.095 ;
        RECT 38.325 1.710 38.935 1.880 ;
        RECT 38.325 0.975 38.495 1.710 ;
      LAYER mcon ;
        RECT 28.035 3.245 28.205 3.415 ;
        RECT 28.035 2.135 28.205 2.305 ;
        RECT 38.765 3.245 38.935 3.415 ;
        RECT 40.615 3.245 40.785 3.415 ;
      LAYER met1 ;
        RECT 28.005 3.415 28.235 3.445 ;
        RECT 38.735 3.415 38.965 3.445 ;
        RECT 40.585 3.415 40.815 3.445 ;
        RECT 27.855 3.245 40.845 3.415 ;
        RECT 28.005 3.215 28.235 3.245 ;
        RECT 38.735 3.215 38.965 3.245 ;
        RECT 40.585 3.215 40.815 3.245 ;
        RECT 28.005 2.305 28.235 2.335 ;
        RECT 27.855 2.135 28.265 2.305 ;
        RECT 28.005 2.105 28.235 2.135 ;
    END
  END y1
  PIN CLK
    ANTENNAGATEAREA 2.042100 ;
    PORT
      LAYER li1 ;
        RECT 2.135 2.055 2.305 5.095 ;
        RECT 13.265 4.975 13.435 5.095 ;
        RECT 13.235 4.765 13.435 4.975 ;
        RECT 13.235 2.055 13.405 4.765 ;
      LAYER mcon ;
        RECT 2.135 4.725 2.305 4.895 ;
        RECT 13.235 4.725 13.405 4.895 ;
      LAYER met1 ;
        RECT 2.105 4.895 2.335 4.925 ;
        RECT 13.205 4.895 13.435 4.925 ;
        RECT 2.075 4.725 13.465 4.895 ;
        RECT 2.105 4.695 2.335 4.725 ;
        RECT 13.205 4.695 13.435 4.725 ;
    END
  END CLK
  PIN VDD
    ANTENNADIFFAREA 53.656651 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 43.340 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 43.075 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 1.005 5.445 1.175 7.460 ;
        RECT 1.885 5.785 2.055 7.460 ;
        RECT 2.765 5.785 2.935 7.460 ;
        RECT 3.645 5.785 3.815 7.460 ;
        RECT 4.655 4.340 4.965 7.460 ;
        RECT 5.515 5.365 5.685 7.460 ;
        RECT 6.395 5.785 6.565 7.460 ;
        RECT 7.275 5.785 7.445 7.460 ;
        RECT 7.985 4.340 8.295 7.460 ;
        RECT 8.845 5.365 9.015 7.460 ;
        RECT 9.725 5.785 9.895 7.460 ;
        RECT 10.605 5.785 10.775 7.460 ;
        RECT 11.315 4.340 11.625 7.460 ;
        RECT 12.175 5.365 12.345 7.460 ;
        RECT 13.055 5.785 13.225 7.460 ;
        RECT 13.935 5.785 14.105 7.460 ;
        RECT 14.645 4.340 14.955 7.460 ;
        RECT 15.505 5.365 15.675 7.460 ;
        RECT 16.385 5.785 16.555 7.460 ;
        RECT 17.265 5.785 17.435 7.460 ;
        RECT 17.975 4.340 18.285 7.460 ;
        RECT 18.835 5.365 19.005 7.460 ;
        RECT 19.715 5.785 19.885 7.460 ;
        RECT 20.595 5.785 20.765 7.460 ;
        RECT 21.305 4.340 21.615 7.460 ;
        RECT 22.465 5.445 22.635 7.460 ;
        RECT 23.345 5.785 23.515 7.460 ;
        RECT 24.225 5.785 24.395 7.460 ;
        RECT 25.105 5.785 25.275 7.460 ;
        RECT 26.115 4.340 26.425 7.460 ;
        RECT 26.975 5.365 27.145 7.460 ;
        RECT 27.855 5.785 28.025 7.460 ;
        RECT 28.735 5.785 28.905 7.460 ;
        RECT 29.445 4.340 29.755 7.460 ;
        RECT 30.305 5.365 30.475 7.460 ;
        RECT 31.185 5.785 31.355 7.460 ;
        RECT 32.065 5.785 32.235 7.460 ;
        RECT 32.775 4.340 33.085 7.460 ;
        RECT 33.635 5.365 33.805 7.460 ;
        RECT 34.515 5.785 34.685 7.460 ;
        RECT 35.395 5.785 35.565 7.460 ;
        RECT 36.105 4.340 36.415 7.460 ;
        RECT 36.965 5.365 37.135 7.460 ;
        RECT 37.845 5.785 38.015 7.460 ;
        RECT 38.725 5.785 38.895 7.460 ;
        RECT 39.435 4.340 39.745 7.460 ;
        RECT 40.295 5.365 40.465 7.460 ;
        RECT 41.175 5.785 41.345 7.460 ;
        RECT 42.055 5.785 42.225 7.460 ;
        RECT 42.765 4.340 43.075 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 0.995 7.525 1.165 7.695 ;
        RECT 1.355 7.525 1.525 7.695 ;
        RECT 1.715 7.525 1.885 7.695 ;
        RECT 2.075 7.525 2.245 7.695 ;
        RECT 2.565 7.525 2.735 7.695 ;
        RECT 2.925 7.525 3.095 7.695 ;
        RECT 3.285 7.525 3.455 7.695 ;
        RECT 3.645 7.525 3.815 7.695 ;
        RECT 4.005 7.525 4.175 7.695 ;
        RECT 4.365 7.525 4.535 7.695 ;
        RECT 5.085 7.525 5.255 7.695 ;
        RECT 5.445 7.525 5.615 7.695 ;
        RECT 5.805 7.525 5.975 7.695 ;
        RECT 6.165 7.525 6.335 7.695 ;
        RECT 6.615 7.525 6.785 7.695 ;
        RECT 6.975 7.525 7.145 7.695 ;
        RECT 7.335 7.525 7.505 7.695 ;
        RECT 7.695 7.525 7.865 7.695 ;
        RECT 8.415 7.525 8.585 7.695 ;
        RECT 8.775 7.525 8.945 7.695 ;
        RECT 9.135 7.525 9.305 7.695 ;
        RECT 9.495 7.525 9.665 7.695 ;
        RECT 9.945 7.525 10.115 7.695 ;
        RECT 10.305 7.525 10.475 7.695 ;
        RECT 10.665 7.525 10.835 7.695 ;
        RECT 11.025 7.525 11.195 7.695 ;
        RECT 11.745 7.525 11.915 7.695 ;
        RECT 12.105 7.525 12.275 7.695 ;
        RECT 12.465 7.525 12.635 7.695 ;
        RECT 12.825 7.525 12.995 7.695 ;
        RECT 13.275 7.525 13.445 7.695 ;
        RECT 13.635 7.525 13.805 7.695 ;
        RECT 13.995 7.525 14.165 7.695 ;
        RECT 14.355 7.525 14.525 7.695 ;
        RECT 15.075 7.525 15.245 7.695 ;
        RECT 15.435 7.525 15.605 7.695 ;
        RECT 15.795 7.525 15.965 7.695 ;
        RECT 16.155 7.525 16.325 7.695 ;
        RECT 16.605 7.525 16.775 7.695 ;
        RECT 16.965 7.525 17.135 7.695 ;
        RECT 17.325 7.525 17.495 7.695 ;
        RECT 17.685 7.525 17.855 7.695 ;
        RECT 18.405 7.525 18.575 7.695 ;
        RECT 18.765 7.525 18.935 7.695 ;
        RECT 19.125 7.525 19.295 7.695 ;
        RECT 19.485 7.525 19.655 7.695 ;
        RECT 19.935 7.525 20.105 7.695 ;
        RECT 20.295 7.525 20.465 7.695 ;
        RECT 20.655 7.525 20.825 7.695 ;
        RECT 21.015 7.525 21.185 7.695 ;
        RECT 21.735 7.525 21.905 7.695 ;
        RECT 22.095 7.525 22.265 7.695 ;
        RECT 22.455 7.525 22.625 7.695 ;
        RECT 22.815 7.525 22.985 7.695 ;
        RECT 23.175 7.525 23.345 7.695 ;
        RECT 23.535 7.525 23.705 7.695 ;
        RECT 24.025 7.525 24.195 7.695 ;
        RECT 24.385 7.525 24.555 7.695 ;
        RECT 24.745 7.525 24.915 7.695 ;
        RECT 25.105 7.525 25.275 7.695 ;
        RECT 25.465 7.525 25.635 7.695 ;
        RECT 25.825 7.525 25.995 7.695 ;
        RECT 26.545 7.525 26.715 7.695 ;
        RECT 26.905 7.525 27.075 7.695 ;
        RECT 27.265 7.525 27.435 7.695 ;
        RECT 27.625 7.525 27.795 7.695 ;
        RECT 28.075 7.525 28.245 7.695 ;
        RECT 28.435 7.525 28.605 7.695 ;
        RECT 28.795 7.525 28.965 7.695 ;
        RECT 29.155 7.525 29.325 7.695 ;
        RECT 29.875 7.525 30.045 7.695 ;
        RECT 30.235 7.525 30.405 7.695 ;
        RECT 30.595 7.525 30.765 7.695 ;
        RECT 30.955 7.525 31.125 7.695 ;
        RECT 31.405 7.525 31.575 7.695 ;
        RECT 31.765 7.525 31.935 7.695 ;
        RECT 32.125 7.525 32.295 7.695 ;
        RECT 32.485 7.525 32.655 7.695 ;
        RECT 33.205 7.525 33.375 7.695 ;
        RECT 33.565 7.525 33.735 7.695 ;
        RECT 33.925 7.525 34.095 7.695 ;
        RECT 34.285 7.525 34.455 7.695 ;
        RECT 34.735 7.525 34.905 7.695 ;
        RECT 35.095 7.525 35.265 7.695 ;
        RECT 35.455 7.525 35.625 7.695 ;
        RECT 35.815 7.525 35.985 7.695 ;
        RECT 36.535 7.525 36.705 7.695 ;
        RECT 36.895 7.525 37.065 7.695 ;
        RECT 37.255 7.525 37.425 7.695 ;
        RECT 37.615 7.525 37.785 7.695 ;
        RECT 38.065 7.525 38.235 7.695 ;
        RECT 38.425 7.525 38.595 7.695 ;
        RECT 38.785 7.525 38.955 7.695 ;
        RECT 39.145 7.525 39.315 7.695 ;
        RECT 39.865 7.525 40.035 7.695 ;
        RECT 40.225 7.525 40.395 7.695 ;
        RECT 40.585 7.525 40.755 7.695 ;
        RECT 40.945 7.525 41.115 7.695 ;
        RECT 41.395 7.525 41.565 7.695 ;
        RECT 41.755 7.525 41.925 7.695 ;
        RECT 42.115 7.525 42.285 7.695 ;
        RECT 42.475 7.525 42.645 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 43.075 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 32.422951 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 43.205 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 4.525 -0.075 5.095 -0.065 ;
        RECT 7.855 -0.075 8.425 -0.065 ;
        RECT 11.185 -0.075 11.755 -0.065 ;
        RECT 14.515 -0.075 15.085 -0.065 ;
        RECT 17.845 -0.075 18.415 -0.065 ;
        RECT 21.175 -0.075 21.745 -0.065 ;
        RECT 25.985 -0.075 26.555 -0.065 ;
        RECT 29.315 -0.075 29.885 -0.065 ;
        RECT 32.645 -0.075 33.215 -0.065 ;
        RECT 35.975 -0.075 36.545 -0.065 ;
        RECT 39.305 -0.075 39.875 -0.065 ;
        RECT 42.635 -0.075 43.205 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 0.990 0.310 1.160 1.270 ;
        RECT 4.655 0.310 4.965 2.860 ;
        RECT 5.905 0.310 6.075 1.260 ;
        RECT 7.985 0.310 8.295 2.860 ;
        RECT 9.235 0.310 9.405 1.260 ;
        RECT 11.315 0.310 11.625 2.860 ;
        RECT 12.565 0.310 12.735 1.260 ;
        RECT 14.645 0.310 14.955 2.860 ;
        RECT 15.895 0.310 16.065 1.260 ;
        RECT 17.975 0.310 18.285 2.860 ;
        RECT 19.225 0.310 19.395 1.260 ;
        RECT 21.305 0.310 21.615 2.860 ;
        RECT 22.450 0.310 22.620 1.270 ;
        RECT 26.115 0.310 26.425 2.860 ;
        RECT 27.365 0.310 27.535 1.260 ;
        RECT 29.445 0.310 29.755 2.860 ;
        RECT 30.695 0.310 30.865 1.260 ;
        RECT 32.775 0.310 33.085 2.860 ;
        RECT 34.025 0.310 34.195 1.260 ;
        RECT 36.105 0.310 36.415 2.860 ;
        RECT 37.355 0.310 37.525 1.260 ;
        RECT 39.435 0.310 39.745 2.860 ;
        RECT 40.685 0.310 40.855 1.260 ;
        RECT 42.765 0.310 43.075 2.860 ;
        RECT -0.155 0.000 43.075 0.310 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 0.995 0.065 1.165 0.235 ;
        RECT 1.355 0.065 1.525 0.235 ;
        RECT 1.715 0.065 1.885 0.235 ;
        RECT 2.075 0.065 2.245 0.235 ;
        RECT 2.565 0.065 2.735 0.235 ;
        RECT 2.925 0.065 3.095 0.235 ;
        RECT 3.285 0.065 3.455 0.235 ;
        RECT 3.645 0.065 3.815 0.235 ;
        RECT 4.005 0.065 4.175 0.235 ;
        RECT 4.365 0.065 4.535 0.235 ;
        RECT 5.085 0.065 5.255 0.235 ;
        RECT 5.445 0.065 5.615 0.235 ;
        RECT 5.805 0.065 5.975 0.235 ;
        RECT 6.165 0.065 6.335 0.235 ;
        RECT 6.615 0.065 6.785 0.235 ;
        RECT 6.975 0.065 7.145 0.235 ;
        RECT 7.335 0.065 7.505 0.235 ;
        RECT 7.695 0.065 7.865 0.235 ;
        RECT 8.415 0.065 8.585 0.235 ;
        RECT 8.775 0.065 8.945 0.235 ;
        RECT 9.135 0.065 9.305 0.235 ;
        RECT 9.495 0.065 9.665 0.235 ;
        RECT 9.945 0.065 10.115 0.235 ;
        RECT 10.305 0.065 10.475 0.235 ;
        RECT 10.665 0.065 10.835 0.235 ;
        RECT 11.025 0.065 11.195 0.235 ;
        RECT 11.745 0.065 11.915 0.235 ;
        RECT 12.105 0.065 12.275 0.235 ;
        RECT 12.465 0.065 12.635 0.235 ;
        RECT 12.825 0.065 12.995 0.235 ;
        RECT 13.275 0.065 13.445 0.235 ;
        RECT 13.635 0.065 13.805 0.235 ;
        RECT 13.995 0.065 14.165 0.235 ;
        RECT 14.355 0.065 14.525 0.235 ;
        RECT 15.075 0.065 15.245 0.235 ;
        RECT 15.435 0.065 15.605 0.235 ;
        RECT 15.795 0.065 15.965 0.235 ;
        RECT 16.155 0.065 16.325 0.235 ;
        RECT 16.605 0.065 16.775 0.235 ;
        RECT 16.965 0.065 17.135 0.235 ;
        RECT 17.325 0.065 17.495 0.235 ;
        RECT 17.685 0.065 17.855 0.235 ;
        RECT 18.405 0.065 18.575 0.235 ;
        RECT 18.765 0.065 18.935 0.235 ;
        RECT 19.125 0.065 19.295 0.235 ;
        RECT 19.485 0.065 19.655 0.235 ;
        RECT 19.935 0.065 20.105 0.235 ;
        RECT 20.295 0.065 20.465 0.235 ;
        RECT 20.655 0.065 20.825 0.235 ;
        RECT 21.015 0.065 21.185 0.235 ;
        RECT 21.735 0.065 21.905 0.235 ;
        RECT 22.095 0.065 22.265 0.235 ;
        RECT 22.455 0.065 22.625 0.235 ;
        RECT 22.815 0.065 22.985 0.235 ;
        RECT 23.175 0.065 23.345 0.235 ;
        RECT 23.535 0.065 23.705 0.235 ;
        RECT 24.025 0.065 24.195 0.235 ;
        RECT 24.385 0.065 24.555 0.235 ;
        RECT 24.745 0.065 24.915 0.235 ;
        RECT 25.105 0.065 25.275 0.235 ;
        RECT 25.465 0.065 25.635 0.235 ;
        RECT 25.825 0.065 25.995 0.235 ;
        RECT 26.545 0.065 26.715 0.235 ;
        RECT 26.905 0.065 27.075 0.235 ;
        RECT 27.265 0.065 27.435 0.235 ;
        RECT 27.625 0.065 27.795 0.235 ;
        RECT 28.075 0.065 28.245 0.235 ;
        RECT 28.435 0.065 28.605 0.235 ;
        RECT 28.795 0.065 28.965 0.235 ;
        RECT 29.155 0.065 29.325 0.235 ;
        RECT 29.875 0.065 30.045 0.235 ;
        RECT 30.235 0.065 30.405 0.235 ;
        RECT 30.595 0.065 30.765 0.235 ;
        RECT 30.955 0.065 31.125 0.235 ;
        RECT 31.405 0.065 31.575 0.235 ;
        RECT 31.765 0.065 31.935 0.235 ;
        RECT 32.125 0.065 32.295 0.235 ;
        RECT 32.485 0.065 32.655 0.235 ;
        RECT 33.205 0.065 33.375 0.235 ;
        RECT 33.565 0.065 33.735 0.235 ;
        RECT 33.925 0.065 34.095 0.235 ;
        RECT 34.285 0.065 34.455 0.235 ;
        RECT 34.735 0.065 34.905 0.235 ;
        RECT 35.095 0.065 35.265 0.235 ;
        RECT 35.455 0.065 35.625 0.235 ;
        RECT 35.815 0.065 35.985 0.235 ;
        RECT 36.535 0.065 36.705 0.235 ;
        RECT 36.895 0.065 37.065 0.235 ;
        RECT 37.255 0.065 37.425 0.235 ;
        RECT 37.615 0.065 37.785 0.235 ;
        RECT 38.065 0.065 38.235 0.235 ;
        RECT 38.425 0.065 38.595 0.235 ;
        RECT 38.785 0.065 38.955 0.235 ;
        RECT 39.145 0.065 39.315 0.235 ;
        RECT 39.865 0.065 40.035 0.235 ;
        RECT 40.225 0.065 40.395 0.235 ;
        RECT 40.585 0.065 40.755 0.235 ;
        RECT 40.945 0.065 41.115 0.235 ;
        RECT 41.395 0.065 41.565 0.235 ;
        RECT 41.755 0.065 41.925 0.235 ;
        RECT 42.115 0.065 42.285 0.235 ;
        RECT 42.475 0.065 42.645 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 43.075 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 1.445 5.470 1.615 7.250 ;
        RECT 2.325 5.470 2.495 7.250 ;
        RECT 3.205 5.470 3.375 7.250 ;
        RECT 5.955 5.515 6.125 7.250 ;
        RECT 6.835 5.515 7.005 7.250 ;
        RECT 9.285 5.515 9.455 7.250 ;
        RECT 10.165 5.515 10.335 7.250 ;
        RECT 12.615 5.515 12.785 7.250 ;
        RECT 13.495 5.515 13.665 7.250 ;
        RECT 19.275 5.515 19.445 7.250 ;
        RECT 20.155 5.515 20.325 7.250 ;
        RECT 1.445 5.300 4.155 5.470 ;
        RECT 5.955 5.345 7.485 5.515 ;
        RECT 9.285 5.345 10.815 5.515 ;
        RECT 12.615 5.345 14.145 5.515 ;
        RECT 19.275 5.345 20.805 5.515 ;
        RECT 1.025 2.055 1.195 5.095 ;
        RECT 3.245 2.055 3.415 5.095 ;
        RECT 0.505 1.815 0.675 1.895 ;
        RECT 1.475 1.815 1.645 1.895 ;
        RECT 2.445 1.815 2.615 1.895 ;
        RECT 0.505 1.645 2.615 1.815 ;
        RECT 0.505 0.515 0.675 1.645 ;
        RECT 1.475 0.765 1.645 1.645 ;
        RECT 2.445 1.565 2.615 1.645 ;
        RECT 1.965 1.220 2.135 1.300 ;
        RECT 3.015 1.220 3.185 1.895 ;
        RECT 3.985 1.890 4.155 5.300 ;
        RECT 5.835 2.055 6.005 5.095 ;
        RECT 1.965 1.050 3.185 1.220 ;
        RECT 1.965 0.970 2.135 1.050 ;
        RECT 2.445 0.765 2.615 0.845 ;
        RECT 1.475 0.595 2.615 0.765 ;
        RECT 1.475 0.515 1.645 0.595 ;
        RECT 2.445 0.515 2.615 0.595 ;
        RECT 3.015 0.765 3.185 1.050 ;
        RECT 3.500 1.720 4.155 1.890 ;
        RECT 5.420 1.805 5.590 1.885 ;
        RECT 6.390 1.805 6.560 1.885 ;
        RECT 7.315 1.880 7.485 5.345 ;
        RECT 9.165 2.055 9.335 5.095 ;
        RECT 9.935 4.940 10.105 5.095 ;
        RECT 9.905 4.765 10.105 4.940 ;
        RECT 9.905 2.055 10.075 4.765 ;
        RECT 3.500 0.985 3.670 1.720 ;
        RECT 5.420 1.635 6.560 1.805 ;
        RECT 3.985 0.765 4.155 1.535 ;
        RECT 3.015 0.595 4.155 0.765 ;
        RECT 3.015 0.515 3.185 0.595 ;
        RECT 3.985 0.515 4.155 0.595 ;
        RECT 5.420 0.505 5.590 1.635 ;
        RECT 6.390 0.755 6.560 1.635 ;
        RECT 6.875 1.710 7.485 1.880 ;
        RECT 8.750 1.805 8.920 1.885 ;
        RECT 9.720 1.805 9.890 1.885 ;
        RECT 10.645 1.880 10.815 5.345 ;
        RECT 12.495 2.055 12.665 5.095 ;
        RECT 6.875 0.975 7.045 1.710 ;
        RECT 8.750 1.635 9.890 1.805 ;
        RECT 7.360 0.755 7.530 1.525 ;
        RECT 6.390 0.585 7.530 0.755 ;
        RECT 6.390 0.505 6.560 0.585 ;
        RECT 7.360 0.505 7.530 0.585 ;
        RECT 8.750 0.505 8.920 1.635 ;
        RECT 9.720 0.755 9.890 1.635 ;
        RECT 10.205 1.710 10.815 1.880 ;
        RECT 12.080 1.805 12.250 1.885 ;
        RECT 13.050 1.805 13.220 1.885 ;
        RECT 13.975 1.880 14.145 5.345 ;
        RECT 15.825 2.055 15.995 5.095 ;
        RECT 16.595 4.940 16.765 5.095 ;
        RECT 19.925 4.940 20.095 5.095 ;
        RECT 16.565 4.765 16.765 4.940 ;
        RECT 19.895 4.765 20.095 4.940 ;
        RECT 16.565 2.055 16.735 4.765 ;
        RECT 19.895 2.055 20.065 4.765 ;
        RECT 10.205 0.975 10.375 1.710 ;
        RECT 12.080 1.635 13.220 1.805 ;
        RECT 10.690 0.755 10.860 1.525 ;
        RECT 9.720 0.585 10.860 0.755 ;
        RECT 9.720 0.505 9.890 0.585 ;
        RECT 10.690 0.505 10.860 0.585 ;
        RECT 12.080 0.505 12.250 1.635 ;
        RECT 13.050 0.755 13.220 1.635 ;
        RECT 13.535 1.710 14.145 1.880 ;
        RECT 15.410 1.805 15.580 1.885 ;
        RECT 16.380 1.805 16.550 1.885 ;
        RECT 13.535 0.975 13.705 1.710 ;
        RECT 15.410 1.635 16.550 1.805 ;
        RECT 14.020 0.755 14.190 1.525 ;
        RECT 13.050 0.585 14.190 0.755 ;
        RECT 13.050 0.505 13.220 0.585 ;
        RECT 14.020 0.505 14.190 0.585 ;
        RECT 15.410 0.505 15.580 1.635 ;
        RECT 16.380 0.755 16.550 1.635 ;
        RECT 18.740 1.805 18.910 1.885 ;
        RECT 19.710 1.805 19.880 1.885 ;
        RECT 20.635 1.880 20.805 5.345 ;
        RECT 22.905 5.470 23.075 7.250 ;
        RECT 23.785 5.470 23.955 7.250 ;
        RECT 24.665 5.470 24.835 7.250 ;
        RECT 27.415 5.515 27.585 7.250 ;
        RECT 28.295 5.515 28.465 7.250 ;
        RECT 30.745 5.515 30.915 7.250 ;
        RECT 31.625 5.515 31.795 7.250 ;
        RECT 34.075 5.515 34.245 7.250 ;
        RECT 34.955 5.515 35.125 7.250 ;
        RECT 40.735 5.515 40.905 7.250 ;
        RECT 41.615 5.515 41.785 7.250 ;
        RECT 22.905 5.300 25.615 5.470 ;
        RECT 27.415 5.345 28.945 5.515 ;
        RECT 30.745 5.345 32.275 5.515 ;
        RECT 34.075 5.345 35.605 5.515 ;
        RECT 40.735 5.345 42.265 5.515 ;
        RECT 22.485 2.055 22.655 5.095 ;
        RECT 23.595 2.055 23.765 5.095 ;
        RECT 24.705 2.055 24.875 5.095 ;
        RECT 18.740 1.635 19.880 1.805 ;
        RECT 17.350 0.755 17.520 1.525 ;
        RECT 16.380 0.585 17.520 0.755 ;
        RECT 16.380 0.505 16.550 0.585 ;
        RECT 17.350 0.505 17.520 0.585 ;
        RECT 18.740 0.505 18.910 1.635 ;
        RECT 19.710 0.755 19.880 1.635 ;
        RECT 20.195 1.710 20.805 1.880 ;
        RECT 21.965 1.815 22.135 1.895 ;
        RECT 22.935 1.815 23.105 1.895 ;
        RECT 23.905 1.815 24.075 1.895 ;
        RECT 20.195 0.975 20.365 1.710 ;
        RECT 21.965 1.645 24.075 1.815 ;
        RECT 20.680 0.755 20.850 1.525 ;
        RECT 19.710 0.585 20.850 0.755 ;
        RECT 19.710 0.505 19.880 0.585 ;
        RECT 20.680 0.505 20.850 0.585 ;
        RECT 21.965 0.515 22.135 1.645 ;
        RECT 22.935 0.765 23.105 1.645 ;
        RECT 23.905 1.565 24.075 1.645 ;
        RECT 23.425 1.220 23.595 1.300 ;
        RECT 24.475 1.220 24.645 1.895 ;
        RECT 25.445 1.890 25.615 5.300 ;
        RECT 27.295 2.055 27.465 5.095 ;
        RECT 23.425 1.050 24.645 1.220 ;
        RECT 23.425 0.970 23.595 1.050 ;
        RECT 23.905 0.765 24.075 0.845 ;
        RECT 22.935 0.595 24.075 0.765 ;
        RECT 22.935 0.515 23.105 0.595 ;
        RECT 23.905 0.515 24.075 0.595 ;
        RECT 24.475 0.765 24.645 1.050 ;
        RECT 24.960 1.720 25.615 1.890 ;
        RECT 26.880 1.805 27.050 1.885 ;
        RECT 27.850 1.805 28.020 1.885 ;
        RECT 28.775 1.880 28.945 5.345 ;
        RECT 30.625 2.055 30.795 5.095 ;
        RECT 31.395 4.940 31.565 5.095 ;
        RECT 31.365 4.765 31.565 4.940 ;
        RECT 31.365 2.055 31.535 4.765 ;
        RECT 24.960 0.985 25.130 1.720 ;
        RECT 26.880 1.635 28.020 1.805 ;
        RECT 25.445 0.765 25.615 1.535 ;
        RECT 24.475 0.595 25.615 0.765 ;
        RECT 24.475 0.515 24.645 0.595 ;
        RECT 25.445 0.515 25.615 0.595 ;
        RECT 26.880 0.505 27.050 1.635 ;
        RECT 27.850 0.755 28.020 1.635 ;
        RECT 28.335 1.710 28.945 1.880 ;
        RECT 30.210 1.805 30.380 1.885 ;
        RECT 31.180 1.805 31.350 1.885 ;
        RECT 32.105 1.880 32.275 5.345 ;
        RECT 33.955 2.055 34.125 5.095 ;
        RECT 34.725 4.975 34.895 5.095 ;
        RECT 34.695 4.765 34.895 4.975 ;
        RECT 34.695 2.055 34.865 4.765 ;
        RECT 28.335 0.975 28.505 1.710 ;
        RECT 30.210 1.635 31.350 1.805 ;
        RECT 28.820 0.755 28.990 1.525 ;
        RECT 27.850 0.585 28.990 0.755 ;
        RECT 27.850 0.505 28.020 0.585 ;
        RECT 28.820 0.505 28.990 0.585 ;
        RECT 30.210 0.505 30.380 1.635 ;
        RECT 31.180 0.755 31.350 1.635 ;
        RECT 31.665 1.710 32.275 1.880 ;
        RECT 33.540 1.805 33.710 1.885 ;
        RECT 34.510 1.805 34.680 1.885 ;
        RECT 35.435 1.880 35.605 5.345 ;
        RECT 37.285 2.055 37.455 5.095 ;
        RECT 38.055 4.940 38.225 5.095 ;
        RECT 41.385 4.940 41.555 5.095 ;
        RECT 38.025 4.765 38.225 4.940 ;
        RECT 41.355 4.765 41.555 4.940 ;
        RECT 38.025 2.055 38.195 4.765 ;
        RECT 41.355 2.055 41.525 4.765 ;
        RECT 31.665 0.975 31.835 1.710 ;
        RECT 33.540 1.635 34.680 1.805 ;
        RECT 32.150 0.755 32.320 1.525 ;
        RECT 31.180 0.585 32.320 0.755 ;
        RECT 31.180 0.505 31.350 0.585 ;
        RECT 32.150 0.505 32.320 0.585 ;
        RECT 33.540 0.505 33.710 1.635 ;
        RECT 34.510 0.755 34.680 1.635 ;
        RECT 34.995 1.710 35.605 1.880 ;
        RECT 36.870 1.805 37.040 1.885 ;
        RECT 37.840 1.805 38.010 1.885 ;
        RECT 34.995 0.975 35.165 1.710 ;
        RECT 36.870 1.635 38.010 1.805 ;
        RECT 35.480 0.755 35.650 1.525 ;
        RECT 34.510 0.585 35.650 0.755 ;
        RECT 34.510 0.505 34.680 0.585 ;
        RECT 35.480 0.505 35.650 0.585 ;
        RECT 36.870 0.505 37.040 1.635 ;
        RECT 37.840 0.755 38.010 1.635 ;
        RECT 40.200 1.805 40.370 1.885 ;
        RECT 41.170 1.805 41.340 1.885 ;
        RECT 42.095 1.880 42.265 5.345 ;
        RECT 40.200 1.635 41.340 1.805 ;
        RECT 38.810 0.755 38.980 1.525 ;
        RECT 37.840 0.585 38.980 0.755 ;
        RECT 37.840 0.505 38.010 0.585 ;
        RECT 38.810 0.505 38.980 0.585 ;
        RECT 40.200 0.505 40.370 1.635 ;
        RECT 41.170 0.755 41.340 1.635 ;
        RECT 41.655 1.710 42.265 1.880 ;
        RECT 41.655 0.975 41.825 1.710 ;
        RECT 42.140 0.755 42.310 1.525 ;
        RECT 41.170 0.585 42.310 0.755 ;
        RECT 41.170 0.505 41.340 0.585 ;
        RECT 42.140 0.505 42.310 0.585 ;
      LAYER mcon ;
        RECT 1.025 4.355 1.195 4.525 ;
        RECT 3.245 3.615 3.415 3.785 ;
        RECT 3.985 3.985 4.155 4.155 ;
        RECT 5.835 3.985 6.005 4.155 ;
        RECT 7.315 3.615 7.485 3.785 ;
        RECT 9.165 3.615 9.335 3.785 ;
        RECT 9.905 4.355 10.075 4.525 ;
        RECT 10.645 3.615 10.815 3.785 ;
        RECT 12.495 3.615 12.665 3.785 ;
        RECT 13.975 4.355 14.145 4.525 ;
        RECT 15.825 3.985 15.995 4.155 ;
        RECT 16.565 3.985 16.735 4.155 ;
        RECT 19.895 4.355 20.065 4.525 ;
        RECT 20.635 3.985 20.805 4.155 ;
        RECT 22.485 4.355 22.655 4.525 ;
        RECT 23.595 4.725 23.765 4.895 ;
        RECT 23.595 3.985 23.765 4.155 ;
        RECT 24.705 3.615 24.875 3.785 ;
        RECT 25.445 3.985 25.615 4.155 ;
        RECT 27.295 3.985 27.465 4.155 ;
        RECT 28.775 3.615 28.945 3.785 ;
        RECT 30.625 3.615 30.795 3.785 ;
        RECT 31.365 4.355 31.535 4.525 ;
        RECT 32.105 3.615 32.275 3.785 ;
        RECT 33.955 3.615 34.125 3.785 ;
        RECT 34.695 4.725 34.865 4.895 ;
        RECT 35.435 4.355 35.605 4.525 ;
        RECT 37.285 3.985 37.455 4.155 ;
        RECT 38.025 3.985 38.195 4.155 ;
        RECT 41.355 4.355 41.525 4.525 ;
        RECT 42.095 3.985 42.265 4.155 ;
      LAYER met1 ;
        RECT 23.565 4.895 23.795 4.925 ;
        RECT 34.665 4.895 34.895 4.925 ;
        RECT 23.535 4.725 34.925 4.895 ;
        RECT 23.565 4.695 23.795 4.725 ;
        RECT 34.665 4.695 34.895 4.725 ;
        RECT 0.995 4.525 1.225 4.555 ;
        RECT 9.875 4.525 10.105 4.555 ;
        RECT 13.945 4.525 14.175 4.555 ;
        RECT 19.865 4.525 20.095 4.555 ;
        RECT 22.455 4.525 22.685 4.555 ;
        RECT 31.335 4.525 31.565 4.555 ;
        RECT 35.405 4.525 35.635 4.555 ;
        RECT 41.325 4.525 41.555 4.555 ;
        RECT 0.965 4.355 20.125 4.525 ;
        RECT 22.425 4.355 41.585 4.525 ;
        RECT 0.995 4.325 1.225 4.355 ;
        RECT 9.875 4.325 10.105 4.355 ;
        RECT 13.945 4.325 14.175 4.355 ;
        RECT 19.865 4.325 20.095 4.355 ;
        RECT 22.455 4.325 22.685 4.355 ;
        RECT 31.335 4.325 31.565 4.355 ;
        RECT 35.405 4.325 35.635 4.355 ;
        RECT 41.325 4.325 41.555 4.355 ;
        RECT 3.955 4.155 4.185 4.185 ;
        RECT 5.805 4.155 6.035 4.185 ;
        RECT 15.795 4.155 16.025 4.185 ;
        RECT 16.535 4.155 16.765 4.185 ;
        RECT 20.605 4.155 20.835 4.185 ;
        RECT 23.565 4.155 23.795 4.185 ;
        RECT 25.415 4.155 25.645 4.185 ;
        RECT 27.265 4.155 27.495 4.185 ;
        RECT 37.255 4.155 37.485 4.185 ;
        RECT 37.995 4.155 38.225 4.185 ;
        RECT 42.065 4.155 42.295 4.185 ;
        RECT 3.925 3.985 16.055 4.155 ;
        RECT 16.505 3.985 23.825 4.155 ;
        RECT 25.385 3.985 37.515 4.155 ;
        RECT 37.965 3.985 42.325 4.155 ;
        RECT 3.955 3.955 4.185 3.985 ;
        RECT 5.805 3.955 6.035 3.985 ;
        RECT 15.795 3.955 16.025 3.985 ;
        RECT 16.535 3.955 16.765 3.985 ;
        RECT 20.605 3.955 20.835 3.985 ;
        RECT 23.565 3.955 23.795 3.985 ;
        RECT 25.415 3.955 25.645 3.985 ;
        RECT 27.265 3.955 27.495 3.985 ;
        RECT 37.255 3.955 37.485 3.985 ;
        RECT 37.995 3.955 38.225 3.985 ;
        RECT 42.065 3.955 42.295 3.985 ;
        RECT 3.215 3.785 3.445 3.815 ;
        RECT 7.285 3.785 7.515 3.815 ;
        RECT 9.135 3.785 9.365 3.815 ;
        RECT 10.615 3.785 10.845 3.815 ;
        RECT 12.465 3.785 12.695 3.815 ;
        RECT 24.675 3.785 24.905 3.815 ;
        RECT 28.745 3.785 28.975 3.815 ;
        RECT 30.595 3.785 30.825 3.815 ;
        RECT 32.075 3.785 32.305 3.815 ;
        RECT 33.925 3.785 34.155 3.815 ;
        RECT 3.185 3.615 9.395 3.785 ;
        RECT 10.585 3.615 12.725 3.785 ;
        RECT 24.645 3.615 30.855 3.785 ;
        RECT 32.045 3.615 34.185 3.785 ;
        RECT 3.215 3.585 3.445 3.615 ;
        RECT 7.285 3.585 7.515 3.615 ;
        RECT 9.135 3.585 9.365 3.615 ;
        RECT 10.615 3.585 10.845 3.615 ;
        RECT 12.465 3.585 12.695 3.615 ;
        RECT 24.675 3.585 24.905 3.615 ;
        RECT 28.745 3.585 28.975 3.615 ;
        RECT 30.595 3.585 30.825 3.615 ;
        RECT 32.075 3.585 32.305 3.615 ;
        RECT 33.925 3.585 34.155 3.615 ;
  END
END Mod4Counter






MACRO MUX2X1
  CLASS BLOCK ;
  FOREIGN MUX2X1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 13.050 BY 7.950 ;
  PIN Y
    ANTENNADIFFAREA 1.351900 ;
    PORT
      LAYER li1 ;
        RECT 10.025 5.515 10.195 7.250 ;
        RECT 10.905 5.515 11.075 7.250 ;
        RECT 10.025 5.345 11.555 5.515 ;
        RECT 11.385 1.880 11.555 5.345 ;
        RECT 10.945 1.710 11.555 1.880 ;
        RECT 10.945 0.975 11.115 1.710 ;
      LAYER mcon ;
        RECT 11.385 3.245 11.555 3.415 ;
      LAYER met1 ;
        RECT 11.355 3.415 11.585 3.445 ;
        RECT 11.325 3.245 11.735 3.415 ;
        RECT 11.355 3.215 11.585 3.245 ;
    END
  END Y
  PIN A0
    ANTENNAGATEAREA 1.027250 ;
    PORT
      LAYER li1 ;
        RECT 4.015 4.940 4.185 5.095 ;
        RECT 3.985 4.765 4.185 4.940 ;
        RECT 3.985 2.055 4.155 4.765 ;
      LAYER mcon ;
        RECT 3.985 3.615 4.155 3.785 ;
      LAYER met1 ;
        RECT 3.955 3.785 4.185 3.815 ;
        RECT 3.805 3.615 4.215 3.785 ;
        RECT 3.955 3.585 4.185 3.615 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA 1.027250 ;
    PORT
      LAYER li1 ;
        RECT 7.345 4.940 7.515 5.095 ;
        RECT 7.315 4.765 7.515 4.940 ;
        RECT 7.315 2.055 7.485 4.765 ;
      LAYER mcon ;
        RECT 7.315 3.985 7.485 4.155 ;
      LAYER met1 ;
        RECT 7.285 4.155 7.515 4.185 ;
        RECT 7.135 3.985 7.545 4.155 ;
        RECT 7.285 3.955 7.515 3.985 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA 2.060500 ;
    PORT
      LAYER li1 ;
        RECT 0.655 2.055 0.825 5.095 ;
        RECT 3.245 2.055 3.415 5.095 ;
      LAYER mcon ;
        RECT 0.655 2.875 0.825 3.045 ;
        RECT 3.245 2.875 3.415 3.045 ;
      LAYER met1 ;
        RECT 0.625 3.045 0.855 3.075 ;
        RECT 3.215 3.045 3.445 3.075 ;
        RECT 0.475 2.875 3.475 3.045 ;
        RECT 0.625 2.845 0.855 2.875 ;
        RECT 3.215 2.845 3.445 2.875 ;
    END
  END S
  PIN VDD
    ANTENNADIFFAREA 16.605850 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 12.630 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 12.365 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 0.585 5.415 0.755 7.460 ;
        RECT 1.465 5.415 1.635 7.460 ;
        RECT 2.065 4.340 2.375 7.460 ;
        RECT 2.925 5.365 3.095 7.460 ;
        RECT 3.805 5.785 3.975 7.460 ;
        RECT 4.685 5.785 4.855 7.460 ;
        RECT 5.395 4.340 5.705 7.460 ;
        RECT 6.255 5.365 6.425 7.460 ;
        RECT 7.135 5.785 7.305 7.460 ;
        RECT 8.015 5.785 8.185 7.460 ;
        RECT 8.725 4.340 9.035 7.460 ;
        RECT 9.585 5.365 9.755 7.460 ;
        RECT 10.465 5.785 10.635 7.460 ;
        RECT 11.345 5.785 11.515 7.460 ;
        RECT 12.055 4.340 12.365 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 1.025 7.525 1.195 7.695 ;
        RECT 1.415 7.525 1.585 7.695 ;
        RECT 1.775 7.525 1.945 7.695 ;
        RECT 2.495 7.525 2.665 7.695 ;
        RECT 2.855 7.525 3.025 7.695 ;
        RECT 3.215 7.525 3.385 7.695 ;
        RECT 3.575 7.525 3.745 7.695 ;
        RECT 4.025 7.525 4.195 7.695 ;
        RECT 4.385 7.525 4.555 7.695 ;
        RECT 4.745 7.525 4.915 7.695 ;
        RECT 5.105 7.525 5.275 7.695 ;
        RECT 5.825 7.525 5.995 7.695 ;
        RECT 6.185 7.525 6.355 7.695 ;
        RECT 6.545 7.525 6.715 7.695 ;
        RECT 6.905 7.525 7.075 7.695 ;
        RECT 7.355 7.525 7.525 7.695 ;
        RECT 7.715 7.525 7.885 7.695 ;
        RECT 8.075 7.525 8.245 7.695 ;
        RECT 8.435 7.525 8.605 7.695 ;
        RECT 9.155 7.525 9.325 7.695 ;
        RECT 9.515 7.525 9.685 7.695 ;
        RECT 9.875 7.525 10.045 7.695 ;
        RECT 10.235 7.525 10.405 7.695 ;
        RECT 10.685 7.525 10.855 7.695 ;
        RECT 11.045 7.525 11.215 7.695 ;
        RECT 11.405 7.525 11.575 7.695 ;
        RECT 11.765 7.525 11.935 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 12.365 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 11.366799 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 12.495 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 1.935 -0.075 2.505 -0.065 ;
        RECT 5.265 -0.075 5.835 -0.065 ;
        RECT 8.595 -0.075 9.165 -0.065 ;
        RECT 11.925 -0.075 12.495 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 0.545 0.755 0.715 1.885 ;
        RECT 1.515 0.755 1.685 1.885 ;
        RECT 0.545 0.585 1.685 0.755 ;
        RECT 0.545 0.310 0.715 0.585 ;
        RECT 1.030 0.310 1.200 0.585 ;
        RECT 1.515 0.310 1.685 0.585 ;
        RECT 2.065 0.310 2.375 2.860 ;
        RECT 3.315 0.310 3.485 1.260 ;
        RECT 5.395 0.310 5.705 2.860 ;
        RECT 6.645 0.310 6.815 1.260 ;
        RECT 8.725 0.310 9.035 2.860 ;
        RECT 9.975 0.310 10.145 1.260 ;
        RECT 12.055 0.310 12.365 2.860 ;
        RECT -0.155 0.000 12.365 0.310 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 1.025 0.065 1.195 0.235 ;
        RECT 1.415 0.065 1.585 0.235 ;
        RECT 1.775 0.065 1.945 0.235 ;
        RECT 2.495 0.065 2.665 0.235 ;
        RECT 2.855 0.065 3.025 0.235 ;
        RECT 3.215 0.065 3.385 0.235 ;
        RECT 3.575 0.065 3.745 0.235 ;
        RECT 4.025 0.065 4.195 0.235 ;
        RECT 4.385 0.065 4.555 0.235 ;
        RECT 4.745 0.065 4.915 0.235 ;
        RECT 5.105 0.065 5.275 0.235 ;
        RECT 5.825 0.065 5.995 0.235 ;
        RECT 6.185 0.065 6.355 0.235 ;
        RECT 6.545 0.065 6.715 0.235 ;
        RECT 6.905 0.065 7.075 0.235 ;
        RECT 7.355 0.065 7.525 0.235 ;
        RECT 7.715 0.065 7.885 0.235 ;
        RECT 8.075 0.065 8.245 0.235 ;
        RECT 8.435 0.065 8.605 0.235 ;
        RECT 9.155 0.065 9.325 0.235 ;
        RECT 9.515 0.065 9.685 0.235 ;
        RECT 9.875 0.065 10.045 0.235 ;
        RECT 10.235 0.065 10.405 0.235 ;
        RECT 10.685 0.065 10.855 0.235 ;
        RECT 11.045 0.065 11.215 0.235 ;
        RECT 11.405 0.065 11.575 0.235 ;
        RECT 11.765 0.065 11.935 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 12.365 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 1.025 4.895 1.195 7.250 ;
        RECT 3.365 5.515 3.535 7.250 ;
        RECT 4.245 5.515 4.415 7.250 ;
        RECT 6.695 5.515 6.865 7.250 ;
        RECT 7.575 5.515 7.745 7.250 ;
        RECT 3.365 5.345 4.895 5.515 ;
        RECT 6.695 5.345 8.225 5.515 ;
        RECT 1.025 4.725 1.565 4.895 ;
        RECT 1.395 2.305 1.565 4.725 ;
        RECT 1.025 2.135 1.565 2.305 ;
        RECT 1.025 0.975 1.195 2.135 ;
        RECT 2.830 1.805 3.000 1.885 ;
        RECT 3.800 1.805 3.970 1.885 ;
        RECT 4.725 1.880 4.895 5.345 ;
        RECT 6.575 2.055 6.745 5.095 ;
        RECT 2.830 1.635 3.970 1.805 ;
        RECT 2.830 0.505 3.000 1.635 ;
        RECT 3.800 0.755 3.970 1.635 ;
        RECT 4.285 1.710 4.895 1.880 ;
        RECT 6.160 1.805 6.330 1.885 ;
        RECT 7.130 1.805 7.300 1.885 ;
        RECT 8.055 1.880 8.225 5.345 ;
        RECT 9.905 2.055 10.075 5.095 ;
        RECT 10.675 4.940 10.845 5.095 ;
        RECT 10.645 4.765 10.845 4.940 ;
        RECT 10.645 2.055 10.815 4.765 ;
        RECT 4.285 0.975 4.455 1.710 ;
        RECT 6.160 1.635 7.300 1.805 ;
        RECT 4.770 0.755 4.940 1.525 ;
        RECT 3.800 0.585 4.940 0.755 ;
        RECT 3.800 0.505 3.970 0.585 ;
        RECT 4.770 0.505 4.940 0.585 ;
        RECT 6.160 0.505 6.330 1.635 ;
        RECT 7.130 0.755 7.300 1.635 ;
        RECT 7.615 1.710 8.225 1.880 ;
        RECT 9.490 1.805 9.660 1.885 ;
        RECT 10.460 1.805 10.630 1.885 ;
        RECT 7.615 0.975 7.785 1.710 ;
        RECT 9.490 1.635 10.630 1.805 ;
        RECT 8.100 0.755 8.270 1.525 ;
        RECT 7.130 0.585 8.270 0.755 ;
        RECT 7.130 0.505 7.300 0.585 ;
        RECT 8.100 0.505 8.270 0.585 ;
        RECT 9.490 0.505 9.660 1.635 ;
        RECT 10.460 0.755 10.630 1.635 ;
        RECT 11.430 0.755 11.600 1.525 ;
        RECT 10.460 0.585 11.600 0.755 ;
        RECT 10.460 0.505 10.630 0.585 ;
        RECT 11.430 0.505 11.600 0.585 ;
      LAYER mcon ;
        RECT 1.395 3.245 1.565 3.415 ;
        RECT 4.725 2.875 4.895 3.045 ;
        RECT 6.575 3.245 6.745 3.415 ;
        RECT 8.055 3.245 8.225 3.415 ;
        RECT 9.905 2.875 10.075 3.045 ;
        RECT 10.645 3.245 10.815 3.415 ;
      LAYER met1 ;
        RECT 1.365 3.415 1.595 3.445 ;
        RECT 6.545 3.415 6.775 3.445 ;
        RECT 8.025 3.415 8.255 3.445 ;
        RECT 10.615 3.415 10.845 3.445 ;
        RECT 1.335 3.245 6.805 3.415 ;
        RECT 7.995 3.245 10.875 3.415 ;
        RECT 1.365 3.215 1.595 3.245 ;
        RECT 6.545 3.215 6.775 3.245 ;
        RECT 8.025 3.215 8.255 3.245 ;
        RECT 10.615 3.215 10.845 3.245 ;
        RECT 4.695 3.045 4.925 3.075 ;
        RECT 9.875 3.045 10.105 3.075 ;
        RECT 4.665 2.875 10.135 3.045 ;
        RECT 4.695 2.845 4.925 2.875 ;
        RECT 9.875 2.845 10.105 2.875 ;
  END
END MUX2X1






MACRO NAND2X1
  CLASS BLOCK ;
  FOREIGN NAND2X1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 4.170 BY 7.950 ;
  PIN Y
    ANTENNADIFFAREA 1.351900 ;
    PORT
      LAYER li1 ;
        RECT 1.145 5.515 1.315 7.250 ;
        RECT 2.025 5.515 2.195 7.250 ;
        RECT 1.145 5.345 2.675 5.515 ;
        RECT 2.505 1.880 2.675 5.345 ;
        RECT 2.065 1.710 2.675 1.880 ;
        RECT 2.065 0.975 2.235 1.710 ;
      LAYER mcon ;
        RECT 2.505 3.245 2.675 3.415 ;
      LAYER met1 ;
        RECT 2.475 3.415 2.705 3.445 ;
        RECT 2.445 3.245 2.855 3.415 ;
        RECT 2.475 3.215 2.705 3.245 ;
    END
  END Y
  PIN A
    ANTENNAGATEAREA 1.033250 ;
    PORT
      LAYER li1 ;
        RECT 1.025 2.055 1.195 5.095 ;
      LAYER mcon ;
        RECT 1.025 3.985 1.195 4.155 ;
      LAYER met1 ;
        RECT 0.995 4.155 1.225 4.185 ;
        RECT 0.845 3.985 1.255 4.155 ;
        RECT 0.995 3.955 1.225 3.985 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 1.027250 ;
    PORT
      LAYER li1 ;
        RECT 1.795 4.940 1.965 5.095 ;
        RECT 1.765 4.765 1.965 4.940 ;
        RECT 1.765 2.055 1.935 4.765 ;
      LAYER mcon ;
        RECT 1.765 3.615 1.935 3.785 ;
      LAYER met1 ;
        RECT 1.735 3.785 1.965 3.815 ;
        RECT 1.585 3.615 1.995 3.785 ;
        RECT 1.735 3.585 1.965 3.615 ;
    END
  END B
  PIN VDD
    ANTENNADIFFAREA 5.209700 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 3.750 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 3.485 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 0.705 5.365 0.875 7.460 ;
        RECT 1.585 5.785 1.755 7.460 ;
        RECT 2.465 5.785 2.635 7.460 ;
        RECT 3.175 4.340 3.485 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 0.995 7.525 1.165 7.695 ;
        RECT 1.355 7.525 1.525 7.695 ;
        RECT 1.805 7.525 1.975 7.695 ;
        RECT 2.165 7.525 2.335 7.695 ;
        RECT 2.525 7.525 2.695 7.695 ;
        RECT 2.885 7.525 3.055 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 3.485 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 3.380600 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 3.615 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 3.045 -0.075 3.615 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 1.095 0.310 1.265 1.260 ;
        RECT 3.175 0.310 3.485 2.860 ;
        RECT -0.155 0.000 3.485 0.310 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 0.995 0.065 1.165 0.235 ;
        RECT 1.355 0.065 1.525 0.235 ;
        RECT 1.805 0.065 1.975 0.235 ;
        RECT 2.165 0.065 2.335 0.235 ;
        RECT 2.525 0.065 2.695 0.235 ;
        RECT 2.885 0.065 3.055 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 3.485 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 0.610 1.805 0.780 1.885 ;
        RECT 1.580 1.805 1.750 1.885 ;
        RECT 0.610 1.635 1.750 1.805 ;
        RECT 0.610 0.505 0.780 1.635 ;
        RECT 1.580 0.755 1.750 1.635 ;
        RECT 2.550 0.755 2.720 1.525 ;
        RECT 1.580 0.585 2.720 0.755 ;
        RECT 1.580 0.505 1.750 0.585 ;
        RECT 2.550 0.505 2.720 0.585 ;
  END
END NAND2X1






MACRO NAND3X1
  CLASS BLOCK ;
  FOREIGN NAND3X1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 5.650 BY 7.950 ;
  PIN Y
    ANTENNADIFFAREA 1.931900 ;
    PORT
      LAYER li1 ;
        RECT 1.445 5.470 1.615 7.250 ;
        RECT 2.325 5.470 2.495 7.250 ;
        RECT 3.205 5.470 3.375 7.250 ;
        RECT 1.445 5.300 4.155 5.470 ;
        RECT 3.985 1.890 4.155 5.300 ;
        RECT 3.500 1.720 4.155 1.890 ;
        RECT 3.500 0.985 3.670 1.720 ;
      LAYER mcon ;
        RECT 3.985 3.245 4.155 3.415 ;
      LAYER met1 ;
        RECT 3.955 3.415 4.185 3.445 ;
        RECT 3.925 3.245 4.335 3.415 ;
        RECT 3.955 3.215 4.185 3.245 ;
    END
  END Y
  PIN A
    ANTENNAGATEAREA 1.033250 ;
    PORT
      LAYER li1 ;
        RECT 1.025 2.055 1.195 5.095 ;
      LAYER mcon ;
        RECT 1.025 3.615 1.195 3.785 ;
      LAYER met1 ;
        RECT 0.995 3.785 1.225 3.815 ;
        RECT 0.845 3.615 1.255 3.785 ;
        RECT 0.995 3.585 1.225 3.615 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 1.014850 ;
    PORT
      LAYER li1 ;
        RECT 2.135 2.055 2.305 5.095 ;
      LAYER mcon ;
        RECT 2.135 3.985 2.305 4.155 ;
      LAYER met1 ;
        RECT 2.105 4.155 2.335 4.185 ;
        RECT 1.955 3.985 2.365 4.155 ;
        RECT 2.105 3.955 2.335 3.985 ;
    END
  END B
  PIN VDD
    ANTENNADIFFAREA 6.500100 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 5.230 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 4.965 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 1.005 5.445 1.175 7.460 ;
        RECT 1.885 5.785 2.055 7.460 ;
        RECT 2.765 5.785 2.935 7.460 ;
        RECT 3.645 5.785 3.815 7.460 ;
        RECT 4.655 4.340 4.965 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 0.995 7.525 1.165 7.695 ;
        RECT 1.355 7.525 1.525 7.695 ;
        RECT 1.715 7.525 1.885 7.695 ;
        RECT 2.075 7.525 2.245 7.695 ;
        RECT 2.565 7.525 2.735 7.695 ;
        RECT 2.925 7.525 3.095 7.695 ;
        RECT 3.285 7.525 3.455 7.695 ;
        RECT 3.645 7.525 3.815 7.695 ;
        RECT 4.005 7.525 4.175 7.695 ;
        RECT 4.365 7.525 4.535 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 4.965 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 4.091000 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 5.095 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 4.525 -0.075 5.095 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 0.990 0.310 1.160 1.270 ;
        RECT 4.655 0.310 4.965 2.860 ;
        RECT -0.155 0.000 4.965 0.310 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 0.995 0.065 1.165 0.235 ;
        RECT 1.355 0.065 1.525 0.235 ;
        RECT 1.715 0.065 1.885 0.235 ;
        RECT 2.075 0.065 2.245 0.235 ;
        RECT 2.565 0.065 2.735 0.235 ;
        RECT 2.925 0.065 3.095 0.235 ;
        RECT 3.285 0.065 3.455 0.235 ;
        RECT 3.645 0.065 3.815 0.235 ;
        RECT 4.005 0.065 4.175 0.235 ;
        RECT 4.365 0.065 4.535 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 4.965 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 3.245 2.055 3.415 5.095 ;
        RECT 0.505 1.815 0.675 1.895 ;
        RECT 1.475 1.815 1.645 1.895 ;
        RECT 2.445 1.815 2.615 1.895 ;
        RECT 0.505 1.645 2.615 1.815 ;
        RECT 0.505 0.515 0.675 1.645 ;
        RECT 1.475 0.765 1.645 1.645 ;
        RECT 2.445 1.565 2.615 1.645 ;
        RECT 1.965 1.220 2.135 1.300 ;
        RECT 3.015 1.220 3.185 1.895 ;
        RECT 1.965 1.050 3.185 1.220 ;
        RECT 1.965 0.970 2.135 1.050 ;
        RECT 2.445 0.765 2.615 0.845 ;
        RECT 1.475 0.595 2.615 0.765 ;
        RECT 1.475 0.515 1.645 0.595 ;
        RECT 2.445 0.515 2.615 0.595 ;
        RECT 3.015 0.765 3.185 1.050 ;
        RECT 3.985 0.765 4.155 1.535 ;
        RECT 3.015 0.595 4.155 0.765 ;
        RECT 3.015 0.515 3.185 0.595 ;
        RECT 3.985 0.515 4.155 0.595 ;
  END
END NAND3X1






MACRO NOR2X1
  CLASS BLOCK ;
  FOREIGN NOR2X1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 4.170 BY 7.950 ;
  PIN Y
    ANTENNADIFFAREA 0.963050 ;
    PORT
      LAYER li1 ;
        RECT 2.025 5.525 2.195 6.795 ;
        RECT 2.025 5.355 2.675 5.525 ;
        RECT 2.505 3.865 2.675 5.355 ;
        RECT 2.500 3.535 2.675 3.865 ;
        RECT 2.505 1.880 2.675 3.535 ;
        RECT 1.095 1.710 2.675 1.880 ;
        RECT 1.095 0.975 1.265 1.710 ;
        RECT 2.065 0.975 2.235 1.710 ;
      LAYER mcon ;
        RECT 2.500 3.615 2.670 3.785 ;
      LAYER met1 ;
        RECT 2.470 3.785 2.700 3.815 ;
        RECT 2.440 3.615 2.850 3.785 ;
        RECT 2.470 3.585 2.700 3.615 ;
    END
  END Y
  PIN A
    ANTENNAGATEAREA 1.027250 ;
    PORT
      LAYER li1 ;
        RECT 0.870 4.940 1.040 5.100 ;
        RECT 0.870 4.770 1.195 4.940 ;
        RECT 1.025 2.055 1.195 4.770 ;
      LAYER mcon ;
        RECT 1.025 3.985 1.195 4.155 ;
      LAYER met1 ;
        RECT 0.995 4.155 1.225 4.185 ;
        RECT 0.845 3.985 1.255 4.155 ;
        RECT 0.995 3.955 1.225 3.985 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 1.026450 ;
    PORT
      LAYER li1 ;
        RECT 1.800 4.940 1.970 5.100 ;
        RECT 1.765 4.770 1.970 4.940 ;
        RECT 1.765 2.055 1.935 4.770 ;
      LAYER mcon ;
        RECT 1.765 3.615 1.935 3.785 ;
      LAYER met1 ;
        RECT 1.735 3.785 1.965 3.815 ;
        RECT 1.585 3.615 1.995 3.785 ;
        RECT 1.735 3.585 1.965 3.615 ;
    END
  END B
  PIN VDD
    ANTENNADIFFAREA 4.109700 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 3.750 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 3.485 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 1.145 5.785 1.315 7.460 ;
        RECT 3.175 4.340 3.485 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 0.995 7.525 1.165 7.695 ;
        RECT 1.355 7.525 1.525 7.695 ;
        RECT 1.805 7.525 1.975 7.695 ;
        RECT 2.165 7.525 2.335 7.695 ;
        RECT 2.525 7.525 2.695 7.695 ;
        RECT 2.885 7.525 3.055 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 3.485 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 5.199200 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 3.615 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 3.045 -0.075 3.615 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 0.610 0.755 0.780 1.885 ;
        RECT 1.580 0.755 1.750 1.530 ;
        RECT 2.550 0.755 2.720 1.530 ;
        RECT 0.610 0.585 2.720 0.755 ;
        RECT 0.610 0.310 0.780 0.585 ;
        RECT 1.095 0.310 1.265 0.585 ;
        RECT 1.580 0.310 1.750 0.585 ;
        RECT 2.065 0.310 2.235 0.585 ;
        RECT 2.550 0.310 2.720 0.585 ;
        RECT 3.175 0.310 3.485 2.860 ;
        RECT -0.155 0.000 3.485 0.310 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 0.995 0.065 1.165 0.235 ;
        RECT 1.355 0.065 1.525 0.235 ;
        RECT 1.805 0.065 1.975 0.235 ;
        RECT 2.165 0.065 2.335 0.235 ;
        RECT 2.525 0.065 2.695 0.235 ;
        RECT 2.885 0.065 3.055 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 3.485 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 0.705 5.525 0.875 7.255 ;
        RECT 1.585 7.055 2.635 7.225 ;
        RECT 1.585 5.525 1.755 7.055 ;
        RECT 2.465 5.785 2.635 7.055 ;
        RECT 0.705 5.355 1.755 5.525 ;
  END
END NOR2X1






MACRO OR2X1
  CLASS BLOCK ;
  FOREIGN OR2X1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 6.390 BY 7.950 ;
  PIN Y
    ANTENNADIFFAREA 0.771900 ;
    PORT
      LAYER li1 ;
        RECT 4.355 4.895 4.525 7.250 ;
        RECT 4.355 4.725 4.895 4.895 ;
        RECT 4.725 2.305 4.895 4.725 ;
        RECT 4.355 2.135 4.895 2.305 ;
        RECT 4.355 0.975 4.525 2.135 ;
      LAYER mcon ;
        RECT 4.725 3.245 4.895 3.415 ;
      LAYER met1 ;
        RECT 4.695 3.415 4.925 3.445 ;
        RECT 4.665 3.245 5.075 3.415 ;
        RECT 4.695 3.215 4.925 3.245 ;
    END
  END Y
  PIN A
    ANTENNAGATEAREA 1.027250 ;
    PORT
      LAYER li1 ;
        RECT 0.870 4.940 1.040 5.100 ;
        RECT 0.870 4.770 1.195 4.940 ;
        RECT 1.025 2.055 1.195 4.770 ;
      LAYER mcon ;
        RECT 1.025 3.985 1.195 4.155 ;
      LAYER met1 ;
        RECT 0.995 4.155 1.225 4.185 ;
        RECT 0.845 3.985 1.255 4.155 ;
        RECT 0.995 3.955 1.225 3.985 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 1.026450 ;
    PORT
      LAYER li1 ;
        RECT 1.800 4.940 1.970 5.100 ;
        RECT 1.765 4.770 1.970 4.940 ;
        RECT 1.765 2.055 1.935 4.770 ;
      LAYER mcon ;
        RECT 1.765 3.615 1.935 3.785 ;
      LAYER met1 ;
        RECT 1.735 3.785 1.965 3.815 ;
        RECT 1.585 3.615 1.995 3.785 ;
        RECT 1.735 3.585 1.965 3.615 ;
    END
  END B
  PIN VDD
    ANTENNADIFFAREA 7.166550 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 5.970 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 5.705 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 1.145 5.785 1.315 7.460 ;
        RECT 3.175 4.340 3.485 7.460 ;
        RECT 3.915 5.415 4.085 7.460 ;
        RECT 4.795 5.415 4.965 7.460 ;
        RECT 5.395 4.340 5.705 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 0.995 7.525 1.165 7.695 ;
        RECT 1.355 7.525 1.525 7.695 ;
        RECT 1.805 7.525 1.975 7.695 ;
        RECT 2.165 7.525 2.335 7.695 ;
        RECT 2.525 7.525 2.695 7.695 ;
        RECT 2.885 7.525 3.055 7.695 ;
        RECT 3.605 7.525 3.775 7.695 ;
        RECT 3.965 7.525 4.135 7.695 ;
        RECT 4.355 7.525 4.525 7.695 ;
        RECT 4.745 7.525 4.915 7.695 ;
        RECT 5.105 7.525 5.275 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 5.705 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 8.163300 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 5.835 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 3.045 -0.075 3.615 -0.065 ;
        RECT 5.265 -0.075 5.835 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 0.610 0.755 0.780 1.885 ;
        RECT 1.580 0.755 1.750 1.530 ;
        RECT 2.550 0.755 2.720 1.530 ;
        RECT 0.610 0.585 2.720 0.755 ;
        RECT 0.610 0.310 0.780 0.585 ;
        RECT 1.095 0.310 1.265 0.585 ;
        RECT 1.580 0.310 1.750 0.585 ;
        RECT 2.065 0.310 2.235 0.585 ;
        RECT 2.550 0.310 2.720 0.585 ;
        RECT 3.175 0.310 3.485 2.860 ;
        RECT 3.875 0.755 4.045 1.885 ;
        RECT 4.845 0.755 5.015 1.885 ;
        RECT 3.875 0.585 5.015 0.755 ;
        RECT 3.875 0.310 4.045 0.585 ;
        RECT 4.360 0.310 4.530 0.585 ;
        RECT 4.845 0.310 5.015 0.585 ;
        RECT 5.395 0.310 5.705 2.860 ;
        RECT -0.155 0.000 5.705 0.310 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 0.995 0.065 1.165 0.235 ;
        RECT 1.355 0.065 1.525 0.235 ;
        RECT 1.805 0.065 1.975 0.235 ;
        RECT 2.165 0.065 2.335 0.235 ;
        RECT 2.525 0.065 2.695 0.235 ;
        RECT 2.885 0.065 3.055 0.235 ;
        RECT 3.605 0.065 3.775 0.235 ;
        RECT 3.965 0.065 4.135 0.235 ;
        RECT 4.355 0.065 4.525 0.235 ;
        RECT 4.745 0.065 4.915 0.235 ;
        RECT 5.105 0.065 5.275 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 5.705 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 0.705 5.525 0.875 7.255 ;
        RECT 1.585 7.055 2.635 7.225 ;
        RECT 1.585 5.525 1.755 7.055 ;
        RECT 0.705 5.355 1.755 5.525 ;
        RECT 2.025 5.525 2.195 6.795 ;
        RECT 2.465 5.785 2.635 7.055 ;
        RECT 2.025 5.355 2.675 5.525 ;
        RECT 2.505 1.880 2.675 5.355 ;
        RECT 3.985 2.055 4.155 5.095 ;
        RECT 1.095 1.710 2.675 1.880 ;
        RECT 1.095 0.975 1.265 1.710 ;
        RECT 2.065 0.975 2.235 1.710 ;
      LAYER mcon ;
        RECT 2.505 3.245 2.675 3.415 ;
        RECT 3.985 3.245 4.155 3.415 ;
      LAYER met1 ;
        RECT 2.475 3.415 2.705 3.445 ;
        RECT 3.955 3.415 4.185 3.445 ;
        RECT 2.445 3.245 4.215 3.415 ;
        RECT 2.475 3.215 2.705 3.245 ;
        RECT 3.955 3.215 4.185 3.245 ;
  END
END OR2X1






MACRO TMRDFFQNX1
  CLASS BLOCK ;
  FOREIGN TMRDFFQNX1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 75.210 BY 7.950 ;
  PIN QN
    ANTENNADIFFAREA 1.734950 ;
    PORT
      LAYER li1 ;
        RECT 72.185 5.525 72.355 6.795 ;
        RECT 73.065 5.525 73.235 6.795 ;
        RECT 72.185 5.355 73.715 5.525 ;
        RECT 73.545 1.870 73.715 5.355 ;
        RECT 73.105 1.700 73.715 1.870 ;
        RECT 66.445 1.310 66.615 1.485 ;
        RECT 66.440 1.155 66.615 1.310 ;
        RECT 66.440 0.975 66.610 1.155 ;
        RECT 69.775 0.975 69.945 1.485 ;
        RECT 73.105 0.975 73.275 1.700 ;
      LAYER mcon ;
        RECT 73.545 3.985 73.715 4.155 ;
        RECT 66.445 1.235 66.615 1.405 ;
        RECT 69.775 1.235 69.945 1.405 ;
        RECT 73.105 1.235 73.275 1.405 ;
      LAYER met1 ;
        RECT 73.515 4.155 73.745 4.185 ;
        RECT 73.485 3.985 73.895 4.155 ;
        RECT 73.515 3.955 73.745 3.985 ;
        RECT 66.415 1.405 66.645 1.435 ;
        RECT 69.745 1.405 69.975 1.435 ;
        RECT 73.075 1.405 73.305 1.435 ;
        RECT 66.385 1.235 73.335 1.405 ;
        RECT 66.415 1.205 66.645 1.235 ;
        RECT 69.745 1.205 69.975 1.235 ;
        RECT 73.075 1.205 73.305 1.235 ;
    END
  END QN
  PIN D
    ANTENNAGATEAREA 3.081750 ;
    PORT
      LAYER li1 ;
        RECT 6.605 4.940 6.775 5.095 ;
        RECT 28.065 4.940 28.235 5.095 ;
        RECT 49.525 4.940 49.695 5.095 ;
        RECT 6.575 4.765 6.775 4.940 ;
        RECT 28.035 4.765 28.235 4.940 ;
        RECT 49.495 4.765 49.695 4.940 ;
        RECT 6.575 2.055 6.745 4.765 ;
        RECT 28.035 2.055 28.205 4.765 ;
        RECT 49.495 2.055 49.665 4.765 ;
      LAYER mcon ;
        RECT 6.575 2.135 6.745 2.305 ;
        RECT 28.035 2.135 28.205 2.305 ;
        RECT 49.495 2.135 49.665 2.305 ;
      LAYER met1 ;
        RECT 6.545 2.305 6.775 2.335 ;
        RECT 28.005 2.305 28.235 2.335 ;
        RECT 49.465 2.305 49.695 2.335 ;
        RECT 6.395 2.135 49.725 2.305 ;
        RECT 6.545 2.105 6.775 2.135 ;
        RECT 28.005 2.105 28.235 2.135 ;
        RECT 49.465 2.105 49.695 2.135 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 6.126300 ;
    PORT
      LAYER li1 ;
        RECT 2.135 2.055 2.305 5.095 ;
        RECT 13.265 4.975 13.435 5.095 ;
        RECT 13.235 4.765 13.435 4.975 ;
        RECT 13.235 2.055 13.405 4.765 ;
        RECT 23.595 2.055 23.765 5.095 ;
        RECT 34.725 4.975 34.895 5.095 ;
        RECT 34.695 4.765 34.895 4.975 ;
        RECT 34.695 2.055 34.865 4.765 ;
        RECT 45.055 2.055 45.225 5.095 ;
        RECT 56.185 4.975 56.355 5.095 ;
        RECT 56.155 4.765 56.355 4.975 ;
        RECT 56.155 2.055 56.325 4.765 ;
      LAYER mcon ;
        RECT 2.135 4.725 2.305 4.895 ;
        RECT 13.235 4.725 13.405 4.895 ;
        RECT 23.595 4.725 23.765 4.895 ;
        RECT 34.695 4.725 34.865 4.895 ;
        RECT 45.055 4.725 45.225 4.895 ;
        RECT 56.155 4.725 56.325 4.895 ;
      LAYER met1 ;
        RECT 2.105 4.895 2.335 4.925 ;
        RECT 13.205 4.895 13.435 4.925 ;
        RECT 23.565 4.895 23.795 4.925 ;
        RECT 34.665 4.895 34.895 4.925 ;
        RECT 45.025 4.895 45.255 4.925 ;
        RECT 56.125 4.895 56.355 4.925 ;
        RECT 2.075 4.890 13.465 4.895 ;
        RECT 16.745 4.890 56.385 4.895 ;
        RECT 2.075 4.735 56.385 4.890 ;
        RECT 2.075 4.725 13.465 4.735 ;
        RECT 16.745 4.725 56.385 4.735 ;
        RECT 2.105 4.695 2.335 4.725 ;
        RECT 13.205 4.695 13.435 4.725 ;
        RECT 23.565 4.695 23.795 4.725 ;
        RECT 34.665 4.695 34.895 4.725 ;
        RECT 45.025 4.695 45.255 4.725 ;
        RECT 56.125 4.695 56.355 4.725 ;
    END
  END CLK
  PIN VDD
    ANTENNADIFFAREA 89.113899 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 74.790 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 74.525 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 1.005 5.445 1.175 7.460 ;
        RECT 1.885 5.785 2.055 7.460 ;
        RECT 2.765 5.785 2.935 7.460 ;
        RECT 3.645 5.785 3.815 7.460 ;
        RECT 4.655 4.340 4.965 7.460 ;
        RECT 5.515 5.365 5.685 7.460 ;
        RECT 6.395 5.785 6.565 7.460 ;
        RECT 7.275 5.785 7.445 7.460 ;
        RECT 7.985 4.340 8.295 7.460 ;
        RECT 8.845 5.365 9.015 7.460 ;
        RECT 9.725 5.785 9.895 7.460 ;
        RECT 10.605 5.785 10.775 7.460 ;
        RECT 11.315 4.340 11.625 7.460 ;
        RECT 12.175 5.365 12.345 7.460 ;
        RECT 13.055 5.785 13.225 7.460 ;
        RECT 13.935 5.785 14.105 7.460 ;
        RECT 14.645 4.340 14.955 7.460 ;
        RECT 15.505 5.365 15.675 7.460 ;
        RECT 16.385 5.785 16.555 7.460 ;
        RECT 17.265 5.785 17.435 7.460 ;
        RECT 17.975 4.340 18.285 7.460 ;
        RECT 18.835 5.365 19.005 7.460 ;
        RECT 19.715 5.785 19.885 7.460 ;
        RECT 20.595 5.785 20.765 7.460 ;
        RECT 21.305 4.340 21.615 7.460 ;
        RECT 22.465 5.445 22.635 7.460 ;
        RECT 23.345 5.785 23.515 7.460 ;
        RECT 24.225 5.785 24.395 7.460 ;
        RECT 25.105 5.785 25.275 7.460 ;
        RECT 26.115 4.340 26.425 7.460 ;
        RECT 26.975 5.365 27.145 7.460 ;
        RECT 27.855 5.785 28.025 7.460 ;
        RECT 28.735 5.785 28.905 7.460 ;
        RECT 29.445 4.340 29.755 7.460 ;
        RECT 30.305 5.365 30.475 7.460 ;
        RECT 31.185 5.785 31.355 7.460 ;
        RECT 32.065 5.785 32.235 7.460 ;
        RECT 32.775 4.340 33.085 7.460 ;
        RECT 33.635 5.365 33.805 7.460 ;
        RECT 34.515 5.785 34.685 7.460 ;
        RECT 35.395 5.785 35.565 7.460 ;
        RECT 36.105 4.340 36.415 7.460 ;
        RECT 36.965 5.365 37.135 7.460 ;
        RECT 37.845 5.785 38.015 7.460 ;
        RECT 38.725 5.785 38.895 7.460 ;
        RECT 39.435 4.340 39.745 7.460 ;
        RECT 40.295 5.365 40.465 7.460 ;
        RECT 41.175 5.785 41.345 7.460 ;
        RECT 42.055 5.785 42.225 7.460 ;
        RECT 42.765 4.340 43.075 7.460 ;
        RECT 43.925 5.445 44.095 7.460 ;
        RECT 44.805 5.785 44.975 7.460 ;
        RECT 45.685 5.785 45.855 7.460 ;
        RECT 46.565 5.785 46.735 7.460 ;
        RECT 47.575 4.340 47.885 7.460 ;
        RECT 48.435 5.365 48.605 7.460 ;
        RECT 49.315 5.785 49.485 7.460 ;
        RECT 50.195 5.785 50.365 7.460 ;
        RECT 50.905 4.340 51.215 7.460 ;
        RECT 51.765 5.365 51.935 7.460 ;
        RECT 52.645 5.785 52.815 7.460 ;
        RECT 53.525 5.785 53.695 7.460 ;
        RECT 54.235 4.340 54.545 7.460 ;
        RECT 55.095 5.365 55.265 7.460 ;
        RECT 55.975 5.785 56.145 7.460 ;
        RECT 56.855 5.785 57.025 7.460 ;
        RECT 57.565 4.340 57.875 7.460 ;
        RECT 58.425 5.365 58.595 7.460 ;
        RECT 59.305 5.785 59.475 7.460 ;
        RECT 60.185 5.785 60.355 7.460 ;
        RECT 60.895 4.340 61.205 7.460 ;
        RECT 61.755 5.365 61.925 7.460 ;
        RECT 62.635 5.785 62.805 7.460 ;
        RECT 63.515 5.785 63.685 7.460 ;
        RECT 64.225 4.340 64.535 7.460 ;
        RECT 65.085 5.355 65.255 7.460 ;
        RECT 65.965 5.785 66.135 7.460 ;
        RECT 66.845 5.355 67.015 7.460 ;
        RECT 67.555 4.340 67.865 7.460 ;
        RECT 70.885 4.340 71.195 7.460 ;
        RECT 74.215 4.340 74.525 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 0.995 7.525 1.165 7.695 ;
        RECT 1.355 7.525 1.525 7.695 ;
        RECT 1.715 7.525 1.885 7.695 ;
        RECT 2.075 7.525 2.245 7.695 ;
        RECT 2.565 7.525 2.735 7.695 ;
        RECT 2.925 7.525 3.095 7.695 ;
        RECT 3.285 7.525 3.455 7.695 ;
        RECT 3.645 7.525 3.815 7.695 ;
        RECT 4.005 7.525 4.175 7.695 ;
        RECT 4.365 7.525 4.535 7.695 ;
        RECT 5.085 7.525 5.255 7.695 ;
        RECT 5.445 7.525 5.615 7.695 ;
        RECT 5.805 7.525 5.975 7.695 ;
        RECT 6.165 7.525 6.335 7.695 ;
        RECT 6.615 7.525 6.785 7.695 ;
        RECT 6.975 7.525 7.145 7.695 ;
        RECT 7.335 7.525 7.505 7.695 ;
        RECT 7.695 7.525 7.865 7.695 ;
        RECT 8.415 7.525 8.585 7.695 ;
        RECT 8.775 7.525 8.945 7.695 ;
        RECT 9.135 7.525 9.305 7.695 ;
        RECT 9.495 7.525 9.665 7.695 ;
        RECT 9.945 7.525 10.115 7.695 ;
        RECT 10.305 7.525 10.475 7.695 ;
        RECT 10.665 7.525 10.835 7.695 ;
        RECT 11.025 7.525 11.195 7.695 ;
        RECT 11.745 7.525 11.915 7.695 ;
        RECT 12.105 7.525 12.275 7.695 ;
        RECT 12.465 7.525 12.635 7.695 ;
        RECT 12.825 7.525 12.995 7.695 ;
        RECT 13.275 7.525 13.445 7.695 ;
        RECT 13.635 7.525 13.805 7.695 ;
        RECT 13.995 7.525 14.165 7.695 ;
        RECT 14.355 7.525 14.525 7.695 ;
        RECT 15.075 7.525 15.245 7.695 ;
        RECT 15.435 7.525 15.605 7.695 ;
        RECT 15.795 7.525 15.965 7.695 ;
        RECT 16.155 7.525 16.325 7.695 ;
        RECT 16.605 7.525 16.775 7.695 ;
        RECT 16.965 7.525 17.135 7.695 ;
        RECT 17.325 7.525 17.495 7.695 ;
        RECT 17.685 7.525 17.855 7.695 ;
        RECT 18.405 7.525 18.575 7.695 ;
        RECT 18.765 7.525 18.935 7.695 ;
        RECT 19.125 7.525 19.295 7.695 ;
        RECT 19.485 7.525 19.655 7.695 ;
        RECT 19.935 7.525 20.105 7.695 ;
        RECT 20.295 7.525 20.465 7.695 ;
        RECT 20.655 7.525 20.825 7.695 ;
        RECT 21.015 7.525 21.185 7.695 ;
        RECT 21.735 7.525 21.905 7.695 ;
        RECT 22.095 7.525 22.265 7.695 ;
        RECT 22.455 7.525 22.625 7.695 ;
        RECT 22.815 7.525 22.985 7.695 ;
        RECT 23.175 7.525 23.345 7.695 ;
        RECT 23.535 7.525 23.705 7.695 ;
        RECT 24.025 7.525 24.195 7.695 ;
        RECT 24.385 7.525 24.555 7.695 ;
        RECT 24.745 7.525 24.915 7.695 ;
        RECT 25.105 7.525 25.275 7.695 ;
        RECT 25.465 7.525 25.635 7.695 ;
        RECT 25.825 7.525 25.995 7.695 ;
        RECT 26.545 7.525 26.715 7.695 ;
        RECT 26.905 7.525 27.075 7.695 ;
        RECT 27.265 7.525 27.435 7.695 ;
        RECT 27.625 7.525 27.795 7.695 ;
        RECT 28.075 7.525 28.245 7.695 ;
        RECT 28.435 7.525 28.605 7.695 ;
        RECT 28.795 7.525 28.965 7.695 ;
        RECT 29.155 7.525 29.325 7.695 ;
        RECT 29.875 7.525 30.045 7.695 ;
        RECT 30.235 7.525 30.405 7.695 ;
        RECT 30.595 7.525 30.765 7.695 ;
        RECT 30.955 7.525 31.125 7.695 ;
        RECT 31.405 7.525 31.575 7.695 ;
        RECT 31.765 7.525 31.935 7.695 ;
        RECT 32.125 7.525 32.295 7.695 ;
        RECT 32.485 7.525 32.655 7.695 ;
        RECT 33.205 7.525 33.375 7.695 ;
        RECT 33.565 7.525 33.735 7.695 ;
        RECT 33.925 7.525 34.095 7.695 ;
        RECT 34.285 7.525 34.455 7.695 ;
        RECT 34.735 7.525 34.905 7.695 ;
        RECT 35.095 7.525 35.265 7.695 ;
        RECT 35.455 7.525 35.625 7.695 ;
        RECT 35.815 7.525 35.985 7.695 ;
        RECT 36.535 7.525 36.705 7.695 ;
        RECT 36.895 7.525 37.065 7.695 ;
        RECT 37.255 7.525 37.425 7.695 ;
        RECT 37.615 7.525 37.785 7.695 ;
        RECT 38.065 7.525 38.235 7.695 ;
        RECT 38.425 7.525 38.595 7.695 ;
        RECT 38.785 7.525 38.955 7.695 ;
        RECT 39.145 7.525 39.315 7.695 ;
        RECT 39.865 7.525 40.035 7.695 ;
        RECT 40.225 7.525 40.395 7.695 ;
        RECT 40.585 7.525 40.755 7.695 ;
        RECT 40.945 7.525 41.115 7.695 ;
        RECT 41.395 7.525 41.565 7.695 ;
        RECT 41.755 7.525 41.925 7.695 ;
        RECT 42.115 7.525 42.285 7.695 ;
        RECT 42.475 7.525 42.645 7.695 ;
        RECT 43.195 7.525 43.365 7.695 ;
        RECT 43.555 7.525 43.725 7.695 ;
        RECT 43.915 7.525 44.085 7.695 ;
        RECT 44.275 7.525 44.445 7.695 ;
        RECT 44.635 7.525 44.805 7.695 ;
        RECT 44.995 7.525 45.165 7.695 ;
        RECT 45.485 7.525 45.655 7.695 ;
        RECT 45.845 7.525 46.015 7.695 ;
        RECT 46.205 7.525 46.375 7.695 ;
        RECT 46.565 7.525 46.735 7.695 ;
        RECT 46.925 7.525 47.095 7.695 ;
        RECT 47.285 7.525 47.455 7.695 ;
        RECT 48.005 7.525 48.175 7.695 ;
        RECT 48.365 7.525 48.535 7.695 ;
        RECT 48.725 7.525 48.895 7.695 ;
        RECT 49.085 7.525 49.255 7.695 ;
        RECT 49.535 7.525 49.705 7.695 ;
        RECT 49.895 7.525 50.065 7.695 ;
        RECT 50.255 7.525 50.425 7.695 ;
        RECT 50.615 7.525 50.785 7.695 ;
        RECT 51.335 7.525 51.505 7.695 ;
        RECT 51.695 7.525 51.865 7.695 ;
        RECT 52.055 7.525 52.225 7.695 ;
        RECT 52.415 7.525 52.585 7.695 ;
        RECT 52.865 7.525 53.035 7.695 ;
        RECT 53.225 7.525 53.395 7.695 ;
        RECT 53.585 7.525 53.755 7.695 ;
        RECT 53.945 7.525 54.115 7.695 ;
        RECT 54.665 7.525 54.835 7.695 ;
        RECT 55.025 7.525 55.195 7.695 ;
        RECT 55.385 7.525 55.555 7.695 ;
        RECT 55.745 7.525 55.915 7.695 ;
        RECT 56.195 7.525 56.365 7.695 ;
        RECT 56.555 7.525 56.725 7.695 ;
        RECT 56.915 7.525 57.085 7.695 ;
        RECT 57.275 7.525 57.445 7.695 ;
        RECT 57.995 7.525 58.165 7.695 ;
        RECT 58.355 7.525 58.525 7.695 ;
        RECT 58.715 7.525 58.885 7.695 ;
        RECT 59.075 7.525 59.245 7.695 ;
        RECT 59.525 7.525 59.695 7.695 ;
        RECT 59.885 7.525 60.055 7.695 ;
        RECT 60.245 7.525 60.415 7.695 ;
        RECT 60.605 7.525 60.775 7.695 ;
        RECT 61.325 7.525 61.495 7.695 ;
        RECT 61.685 7.525 61.855 7.695 ;
        RECT 62.045 7.525 62.215 7.695 ;
        RECT 62.405 7.525 62.575 7.695 ;
        RECT 62.855 7.525 63.025 7.695 ;
        RECT 63.215 7.525 63.385 7.695 ;
        RECT 63.575 7.525 63.745 7.695 ;
        RECT 63.935 7.525 64.105 7.695 ;
        RECT 64.655 7.525 64.825 7.695 ;
        RECT 65.015 7.525 65.185 7.695 ;
        RECT 65.375 7.525 65.545 7.695 ;
        RECT 65.735 7.525 65.905 7.695 ;
        RECT 66.185 7.525 66.355 7.695 ;
        RECT 66.545 7.525 66.715 7.695 ;
        RECT 66.905 7.525 67.075 7.695 ;
        RECT 67.265 7.525 67.435 7.695 ;
        RECT 67.985 7.525 68.155 7.695 ;
        RECT 68.345 7.525 68.515 7.695 ;
        RECT 68.705 7.525 68.875 7.695 ;
        RECT 69.065 7.525 69.235 7.695 ;
        RECT 69.515 7.525 69.685 7.695 ;
        RECT 69.875 7.525 70.045 7.695 ;
        RECT 70.235 7.525 70.405 7.695 ;
        RECT 70.595 7.525 70.765 7.695 ;
        RECT 71.315 7.525 71.485 7.695 ;
        RECT 71.675 7.525 71.845 7.695 ;
        RECT 72.035 7.525 72.205 7.695 ;
        RECT 72.395 7.525 72.565 7.695 ;
        RECT 72.845 7.525 73.015 7.695 ;
        RECT 73.205 7.525 73.375 7.695 ;
        RECT 73.565 7.525 73.735 7.695 ;
        RECT 73.925 7.525 74.095 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 74.525 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 55.732800 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 74.655 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 4.525 -0.075 5.095 -0.065 ;
        RECT 7.855 -0.075 8.425 -0.065 ;
        RECT 11.185 -0.075 11.755 -0.065 ;
        RECT 14.515 -0.075 15.085 -0.065 ;
        RECT 17.845 -0.075 18.415 -0.065 ;
        RECT 21.175 -0.075 21.745 -0.065 ;
        RECT 25.985 -0.075 26.555 -0.065 ;
        RECT 29.315 -0.075 29.885 -0.065 ;
        RECT 32.645 -0.075 33.215 -0.065 ;
        RECT 35.975 -0.075 36.545 -0.065 ;
        RECT 39.305 -0.075 39.875 -0.065 ;
        RECT 42.635 -0.075 43.205 -0.065 ;
        RECT 47.445 -0.075 48.015 -0.065 ;
        RECT 50.775 -0.075 51.345 -0.065 ;
        RECT 54.105 -0.075 54.675 -0.065 ;
        RECT 57.435 -0.075 58.005 -0.065 ;
        RECT 60.765 -0.075 61.335 -0.065 ;
        RECT 64.095 -0.075 64.665 -0.065 ;
        RECT 67.425 -0.075 67.995 -0.065 ;
        RECT 70.755 -0.075 71.325 -0.065 ;
        RECT 74.085 -0.075 74.655 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 0.990 0.310 1.160 1.270 ;
        RECT 4.655 0.310 4.965 2.860 ;
        RECT 5.905 0.310 6.075 1.260 ;
        RECT 7.985 0.310 8.295 2.860 ;
        RECT 9.235 0.310 9.405 1.260 ;
        RECT 11.315 0.310 11.625 2.860 ;
        RECT 12.565 0.310 12.735 1.260 ;
        RECT 14.645 0.310 14.955 2.860 ;
        RECT 15.895 0.310 16.065 1.260 ;
        RECT 17.975 0.310 18.285 2.860 ;
        RECT 19.225 0.310 19.395 1.260 ;
        RECT 21.305 0.310 21.615 2.860 ;
        RECT 22.450 0.310 22.620 1.270 ;
        RECT 26.115 0.310 26.425 2.860 ;
        RECT 27.365 0.310 27.535 1.260 ;
        RECT 29.445 0.310 29.755 2.860 ;
        RECT 30.695 0.310 30.865 1.260 ;
        RECT 32.775 0.310 33.085 2.860 ;
        RECT 34.025 0.310 34.195 1.260 ;
        RECT 36.105 0.310 36.415 2.860 ;
        RECT 37.355 0.310 37.525 1.260 ;
        RECT 39.435 0.310 39.745 2.860 ;
        RECT 40.685 0.310 40.855 1.260 ;
        RECT 42.765 0.310 43.075 2.860 ;
        RECT 43.910 0.310 44.080 1.270 ;
        RECT 47.575 0.310 47.885 2.860 ;
        RECT 48.825 0.310 48.995 1.260 ;
        RECT 50.905 0.310 51.215 2.860 ;
        RECT 52.155 0.310 52.325 1.260 ;
        RECT 54.235 0.310 54.545 2.860 ;
        RECT 55.485 0.310 55.655 1.260 ;
        RECT 57.565 0.310 57.875 2.860 ;
        RECT 58.815 0.310 58.985 1.260 ;
        RECT 60.895 0.310 61.205 2.860 ;
        RECT 62.145 0.310 62.315 1.260 ;
        RECT 64.225 0.310 64.535 2.860 ;
        RECT 65.475 0.310 65.645 1.260 ;
        RECT 67.555 0.310 67.865 2.860 ;
        RECT 68.805 0.310 68.975 1.260 ;
        RECT 70.885 0.310 71.195 2.860 ;
        RECT 72.135 0.310 72.305 1.260 ;
        RECT 74.215 0.310 74.525 2.860 ;
        RECT -0.155 0.235 69.775 0.310 ;
        RECT 69.945 0.235 74.525 0.310 ;
        RECT -0.155 0.000 74.525 0.235 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 0.995 0.065 1.165 0.235 ;
        RECT 1.355 0.065 1.525 0.235 ;
        RECT 1.715 0.065 1.885 0.235 ;
        RECT 2.075 0.065 2.245 0.235 ;
        RECT 2.565 0.065 2.735 0.235 ;
        RECT 2.925 0.065 3.095 0.235 ;
        RECT 3.285 0.065 3.455 0.235 ;
        RECT 3.645 0.065 3.815 0.235 ;
        RECT 4.005 0.065 4.175 0.235 ;
        RECT 4.365 0.065 4.535 0.235 ;
        RECT 5.085 0.065 5.255 0.235 ;
        RECT 5.445 0.065 5.615 0.235 ;
        RECT 5.805 0.065 5.975 0.235 ;
        RECT 6.165 0.065 6.335 0.235 ;
        RECT 6.615 0.065 6.785 0.235 ;
        RECT 6.975 0.065 7.145 0.235 ;
        RECT 7.335 0.065 7.505 0.235 ;
        RECT 7.695 0.065 7.865 0.235 ;
        RECT 8.415 0.065 8.585 0.235 ;
        RECT 8.775 0.065 8.945 0.235 ;
        RECT 9.135 0.065 9.305 0.235 ;
        RECT 9.495 0.065 9.665 0.235 ;
        RECT 9.945 0.065 10.115 0.235 ;
        RECT 10.305 0.065 10.475 0.235 ;
        RECT 10.665 0.065 10.835 0.235 ;
        RECT 11.025 0.065 11.195 0.235 ;
        RECT 11.745 0.065 11.915 0.235 ;
        RECT 12.105 0.065 12.275 0.235 ;
        RECT 12.465 0.065 12.635 0.235 ;
        RECT 12.825 0.065 12.995 0.235 ;
        RECT 13.275 0.065 13.445 0.235 ;
        RECT 13.635 0.065 13.805 0.235 ;
        RECT 13.995 0.065 14.165 0.235 ;
        RECT 14.355 0.065 14.525 0.235 ;
        RECT 15.075 0.065 15.245 0.235 ;
        RECT 15.435 0.065 15.605 0.235 ;
        RECT 15.795 0.065 15.965 0.235 ;
        RECT 16.155 0.065 16.325 0.235 ;
        RECT 16.605 0.065 16.775 0.235 ;
        RECT 16.965 0.065 17.135 0.235 ;
        RECT 17.325 0.065 17.495 0.235 ;
        RECT 17.685 0.065 17.855 0.235 ;
        RECT 18.405 0.065 18.575 0.235 ;
        RECT 18.765 0.065 18.935 0.235 ;
        RECT 19.125 0.065 19.295 0.235 ;
        RECT 19.485 0.065 19.655 0.235 ;
        RECT 19.935 0.065 20.105 0.235 ;
        RECT 20.295 0.065 20.465 0.235 ;
        RECT 20.655 0.065 20.825 0.235 ;
        RECT 21.015 0.065 21.185 0.235 ;
        RECT 21.735 0.065 21.905 0.235 ;
        RECT 22.095 0.065 22.265 0.235 ;
        RECT 22.455 0.065 22.625 0.235 ;
        RECT 22.815 0.065 22.985 0.235 ;
        RECT 23.175 0.065 23.345 0.235 ;
        RECT 23.535 0.065 23.705 0.235 ;
        RECT 24.025 0.065 24.195 0.235 ;
        RECT 24.385 0.065 24.555 0.235 ;
        RECT 24.745 0.065 24.915 0.235 ;
        RECT 25.105 0.065 25.275 0.235 ;
        RECT 25.465 0.065 25.635 0.235 ;
        RECT 25.825 0.065 25.995 0.235 ;
        RECT 26.545 0.065 26.715 0.235 ;
        RECT 26.905 0.065 27.075 0.235 ;
        RECT 27.265 0.065 27.435 0.235 ;
        RECT 27.625 0.065 27.795 0.235 ;
        RECT 28.075 0.065 28.245 0.235 ;
        RECT 28.435 0.065 28.605 0.235 ;
        RECT 28.795 0.065 28.965 0.235 ;
        RECT 29.155 0.065 29.325 0.235 ;
        RECT 29.875 0.065 30.045 0.235 ;
        RECT 30.235 0.065 30.405 0.235 ;
        RECT 30.595 0.065 30.765 0.235 ;
        RECT 30.955 0.065 31.125 0.235 ;
        RECT 31.405 0.065 31.575 0.235 ;
        RECT 31.765 0.065 31.935 0.235 ;
        RECT 32.125 0.065 32.295 0.235 ;
        RECT 32.485 0.065 32.655 0.235 ;
        RECT 33.205 0.065 33.375 0.235 ;
        RECT 33.565 0.065 33.735 0.235 ;
        RECT 33.925 0.065 34.095 0.235 ;
        RECT 34.285 0.065 34.455 0.235 ;
        RECT 34.735 0.065 34.905 0.235 ;
        RECT 35.095 0.065 35.265 0.235 ;
        RECT 35.455 0.065 35.625 0.235 ;
        RECT 35.815 0.065 35.985 0.235 ;
        RECT 36.535 0.065 36.705 0.235 ;
        RECT 36.895 0.065 37.065 0.235 ;
        RECT 37.255 0.065 37.425 0.235 ;
        RECT 37.615 0.065 37.785 0.235 ;
        RECT 38.065 0.065 38.235 0.235 ;
        RECT 38.425 0.065 38.595 0.235 ;
        RECT 38.785 0.065 38.955 0.235 ;
        RECT 39.145 0.065 39.315 0.235 ;
        RECT 39.865 0.065 40.035 0.235 ;
        RECT 40.225 0.065 40.395 0.235 ;
        RECT 40.585 0.065 40.755 0.235 ;
        RECT 40.945 0.065 41.115 0.235 ;
        RECT 41.395 0.065 41.565 0.235 ;
        RECT 41.755 0.065 41.925 0.235 ;
        RECT 42.115 0.065 42.285 0.235 ;
        RECT 42.475 0.065 42.645 0.235 ;
        RECT 43.195 0.065 43.365 0.235 ;
        RECT 43.555 0.065 43.725 0.235 ;
        RECT 43.915 0.065 44.085 0.235 ;
        RECT 44.275 0.065 44.445 0.235 ;
        RECT 44.635 0.065 44.805 0.235 ;
        RECT 44.995 0.065 45.165 0.235 ;
        RECT 45.485 0.065 45.655 0.235 ;
        RECT 45.845 0.065 46.015 0.235 ;
        RECT 46.205 0.065 46.375 0.235 ;
        RECT 46.565 0.065 46.735 0.235 ;
        RECT 46.925 0.065 47.095 0.235 ;
        RECT 47.285 0.065 47.455 0.235 ;
        RECT 48.005 0.065 48.175 0.235 ;
        RECT 48.365 0.065 48.535 0.235 ;
        RECT 48.725 0.065 48.895 0.235 ;
        RECT 49.085 0.065 49.255 0.235 ;
        RECT 49.535 0.065 49.705 0.235 ;
        RECT 49.895 0.065 50.065 0.235 ;
        RECT 50.255 0.065 50.425 0.235 ;
        RECT 50.615 0.065 50.785 0.235 ;
        RECT 51.335 0.065 51.505 0.235 ;
        RECT 51.695 0.065 51.865 0.235 ;
        RECT 52.055 0.065 52.225 0.235 ;
        RECT 52.415 0.065 52.585 0.235 ;
        RECT 52.865 0.065 53.035 0.235 ;
        RECT 53.225 0.065 53.395 0.235 ;
        RECT 53.585 0.065 53.755 0.235 ;
        RECT 53.945 0.065 54.115 0.235 ;
        RECT 54.665 0.065 54.835 0.235 ;
        RECT 55.025 0.065 55.195 0.235 ;
        RECT 55.385 0.065 55.555 0.235 ;
        RECT 55.745 0.065 55.915 0.235 ;
        RECT 56.195 0.065 56.365 0.235 ;
        RECT 56.555 0.065 56.725 0.235 ;
        RECT 56.915 0.065 57.085 0.235 ;
        RECT 57.275 0.065 57.445 0.235 ;
        RECT 57.995 0.065 58.165 0.235 ;
        RECT 58.355 0.065 58.525 0.235 ;
        RECT 58.715 0.065 58.885 0.235 ;
        RECT 59.075 0.065 59.245 0.235 ;
        RECT 59.525 0.065 59.695 0.235 ;
        RECT 59.885 0.065 60.055 0.235 ;
        RECT 60.245 0.065 60.415 0.235 ;
        RECT 60.605 0.065 60.775 0.235 ;
        RECT 61.325 0.065 61.495 0.235 ;
        RECT 61.685 0.065 61.855 0.235 ;
        RECT 62.045 0.065 62.215 0.235 ;
        RECT 62.405 0.065 62.575 0.235 ;
        RECT 62.855 0.065 63.025 0.235 ;
        RECT 63.215 0.065 63.385 0.235 ;
        RECT 63.575 0.065 63.745 0.235 ;
        RECT 63.935 0.065 64.105 0.235 ;
        RECT 64.655 0.065 64.825 0.235 ;
        RECT 65.015 0.065 65.185 0.235 ;
        RECT 65.375 0.065 65.545 0.235 ;
        RECT 65.735 0.065 65.905 0.235 ;
        RECT 66.185 0.065 66.355 0.235 ;
        RECT 66.545 0.065 66.715 0.235 ;
        RECT 66.905 0.065 67.075 0.235 ;
        RECT 67.265 0.065 67.435 0.235 ;
        RECT 67.985 0.065 68.155 0.235 ;
        RECT 68.345 0.065 68.515 0.235 ;
        RECT 68.705 0.065 68.875 0.235 ;
        RECT 69.065 0.065 69.235 0.235 ;
        RECT 69.515 0.065 69.685 0.235 ;
        RECT 69.875 0.065 70.045 0.235 ;
        RECT 70.235 0.065 70.405 0.235 ;
        RECT 70.595 0.065 70.765 0.235 ;
        RECT 71.315 0.065 71.485 0.235 ;
        RECT 71.675 0.065 71.845 0.235 ;
        RECT 72.035 0.065 72.205 0.235 ;
        RECT 72.395 0.065 72.565 0.235 ;
        RECT 72.845 0.065 73.015 0.235 ;
        RECT 73.205 0.065 73.375 0.235 ;
        RECT 73.565 0.065 73.735 0.235 ;
        RECT 73.925 0.065 74.095 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 74.525 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 1.445 5.470 1.615 7.250 ;
        RECT 2.325 5.470 2.495 7.250 ;
        RECT 3.205 5.470 3.375 7.250 ;
        RECT 5.955 5.515 6.125 7.250 ;
        RECT 6.835 5.515 7.005 7.250 ;
        RECT 9.285 5.515 9.455 7.250 ;
        RECT 10.165 5.515 10.335 7.250 ;
        RECT 12.615 5.515 12.785 7.250 ;
        RECT 13.495 5.515 13.665 7.250 ;
        RECT 15.945 5.515 16.115 7.250 ;
        RECT 16.825 5.515 16.995 7.250 ;
        RECT 19.275 5.515 19.445 7.250 ;
        RECT 20.155 5.515 20.325 7.250 ;
        RECT 1.445 5.300 4.155 5.470 ;
        RECT 5.955 5.345 7.485 5.515 ;
        RECT 9.285 5.345 10.815 5.515 ;
        RECT 12.615 5.345 14.145 5.515 ;
        RECT 15.945 5.345 17.475 5.515 ;
        RECT 19.275 5.345 20.805 5.515 ;
        RECT 1.025 2.055 1.195 5.095 ;
        RECT 3.245 2.055 3.415 5.095 ;
        RECT 0.505 1.815 0.675 1.895 ;
        RECT 1.475 1.815 1.645 1.895 ;
        RECT 2.445 1.815 2.615 1.895 ;
        RECT 0.505 1.645 2.615 1.815 ;
        RECT 0.505 0.515 0.675 1.645 ;
        RECT 1.475 0.765 1.645 1.645 ;
        RECT 2.445 1.565 2.615 1.645 ;
        RECT 1.965 1.220 2.135 1.300 ;
        RECT 3.015 1.220 3.185 1.895 ;
        RECT 3.985 1.890 4.155 5.300 ;
        RECT 5.835 2.055 6.005 5.095 ;
        RECT 1.965 1.050 3.185 1.220 ;
        RECT 1.965 0.970 2.135 1.050 ;
        RECT 2.445 0.765 2.615 0.845 ;
        RECT 1.475 0.595 2.615 0.765 ;
        RECT 1.475 0.515 1.645 0.595 ;
        RECT 2.445 0.515 2.615 0.595 ;
        RECT 3.015 0.765 3.185 1.050 ;
        RECT 3.500 1.720 4.155 1.890 ;
        RECT 5.420 1.805 5.590 1.885 ;
        RECT 6.390 1.805 6.560 1.885 ;
        RECT 7.315 1.880 7.485 5.345 ;
        RECT 9.165 2.055 9.335 5.095 ;
        RECT 9.935 4.940 10.105 5.095 ;
        RECT 9.905 4.765 10.105 4.940 ;
        RECT 9.905 2.055 10.075 4.765 ;
        RECT 3.500 0.985 3.670 1.720 ;
        RECT 5.420 1.635 6.560 1.805 ;
        RECT 3.985 0.765 4.155 1.535 ;
        RECT 3.015 0.595 4.155 0.765 ;
        RECT 3.015 0.515 3.185 0.595 ;
        RECT 3.985 0.515 4.155 0.595 ;
        RECT 5.420 0.505 5.590 1.635 ;
        RECT 6.390 0.755 6.560 1.635 ;
        RECT 6.875 1.710 7.485 1.880 ;
        RECT 8.750 1.805 8.920 1.885 ;
        RECT 9.720 1.805 9.890 1.885 ;
        RECT 10.645 1.880 10.815 5.345 ;
        RECT 12.495 2.055 12.665 5.095 ;
        RECT 6.875 0.975 7.045 1.710 ;
        RECT 8.750 1.635 9.890 1.805 ;
        RECT 7.360 0.755 7.530 1.525 ;
        RECT 6.390 0.585 7.530 0.755 ;
        RECT 6.390 0.505 6.560 0.585 ;
        RECT 7.360 0.505 7.530 0.585 ;
        RECT 8.750 0.505 8.920 1.635 ;
        RECT 9.720 0.755 9.890 1.635 ;
        RECT 10.205 1.710 10.815 1.880 ;
        RECT 12.080 1.805 12.250 1.885 ;
        RECT 13.050 1.805 13.220 1.885 ;
        RECT 13.975 1.880 14.145 5.345 ;
        RECT 15.825 2.055 15.995 5.095 ;
        RECT 16.595 4.940 16.765 5.095 ;
        RECT 16.565 4.765 16.765 4.940 ;
        RECT 16.565 2.055 16.735 4.765 ;
        RECT 10.205 0.975 10.375 1.710 ;
        RECT 12.080 1.635 13.220 1.805 ;
        RECT 10.690 0.755 10.860 1.525 ;
        RECT 9.720 0.585 10.860 0.755 ;
        RECT 9.720 0.505 9.890 0.585 ;
        RECT 10.690 0.505 10.860 0.585 ;
        RECT 12.080 0.505 12.250 1.635 ;
        RECT 13.050 0.755 13.220 1.635 ;
        RECT 13.535 1.710 14.145 1.880 ;
        RECT 15.410 1.805 15.580 1.885 ;
        RECT 16.380 1.805 16.550 1.885 ;
        RECT 17.305 1.880 17.475 5.345 ;
        RECT 19.155 2.055 19.325 5.095 ;
        RECT 19.925 4.940 20.095 5.095 ;
        RECT 19.895 4.765 20.095 4.940 ;
        RECT 19.895 2.055 20.065 4.765 ;
        RECT 13.535 0.975 13.705 1.710 ;
        RECT 15.410 1.635 16.550 1.805 ;
        RECT 14.020 0.755 14.190 1.525 ;
        RECT 13.050 0.585 14.190 0.755 ;
        RECT 13.050 0.505 13.220 0.585 ;
        RECT 14.020 0.505 14.190 0.585 ;
        RECT 15.410 0.505 15.580 1.635 ;
        RECT 16.380 0.755 16.550 1.635 ;
        RECT 16.865 1.710 17.475 1.880 ;
        RECT 18.740 1.805 18.910 1.885 ;
        RECT 19.710 1.805 19.880 1.885 ;
        RECT 20.635 1.880 20.805 5.345 ;
        RECT 22.905 5.470 23.075 7.250 ;
        RECT 23.785 5.470 23.955 7.250 ;
        RECT 24.665 5.470 24.835 7.250 ;
        RECT 27.415 5.515 27.585 7.250 ;
        RECT 28.295 5.515 28.465 7.250 ;
        RECT 30.745 5.515 30.915 7.250 ;
        RECT 31.625 5.515 31.795 7.250 ;
        RECT 34.075 5.515 34.245 7.250 ;
        RECT 34.955 5.515 35.125 7.250 ;
        RECT 37.405 5.515 37.575 7.250 ;
        RECT 38.285 5.515 38.455 7.250 ;
        RECT 40.735 5.515 40.905 7.250 ;
        RECT 41.615 5.515 41.785 7.250 ;
        RECT 22.905 5.300 25.615 5.470 ;
        RECT 27.415 5.345 28.945 5.515 ;
        RECT 30.745 5.345 32.275 5.515 ;
        RECT 34.075 5.345 35.605 5.515 ;
        RECT 37.405 5.345 38.935 5.515 ;
        RECT 40.735 5.345 42.265 5.515 ;
        RECT 22.485 2.055 22.655 5.095 ;
        RECT 24.705 2.055 24.875 5.095 ;
        RECT 16.865 0.975 17.035 1.710 ;
        RECT 18.740 1.635 19.880 1.805 ;
        RECT 17.350 0.755 17.520 1.525 ;
        RECT 16.380 0.585 17.520 0.755 ;
        RECT 16.380 0.505 16.550 0.585 ;
        RECT 17.350 0.505 17.520 0.585 ;
        RECT 18.740 0.505 18.910 1.635 ;
        RECT 19.710 0.755 19.880 1.635 ;
        RECT 20.195 1.710 20.805 1.880 ;
        RECT 21.965 1.815 22.135 1.895 ;
        RECT 22.935 1.815 23.105 1.895 ;
        RECT 23.905 1.815 24.075 1.895 ;
        RECT 20.195 0.975 20.365 1.710 ;
        RECT 21.965 1.645 24.075 1.815 ;
        RECT 20.680 0.755 20.850 1.525 ;
        RECT 19.710 0.585 20.850 0.755 ;
        RECT 19.710 0.505 19.880 0.585 ;
        RECT 20.680 0.505 20.850 0.585 ;
        RECT 21.965 0.515 22.135 1.645 ;
        RECT 22.935 0.765 23.105 1.645 ;
        RECT 23.905 1.565 24.075 1.645 ;
        RECT 23.425 1.220 23.595 1.300 ;
        RECT 24.475 1.220 24.645 1.895 ;
        RECT 25.445 1.890 25.615 5.300 ;
        RECT 27.295 2.055 27.465 5.095 ;
        RECT 23.425 1.050 24.645 1.220 ;
        RECT 23.425 0.970 23.595 1.050 ;
        RECT 23.905 0.765 24.075 0.845 ;
        RECT 22.935 0.595 24.075 0.765 ;
        RECT 22.935 0.515 23.105 0.595 ;
        RECT 23.905 0.515 24.075 0.595 ;
        RECT 24.475 0.765 24.645 1.050 ;
        RECT 24.960 1.720 25.615 1.890 ;
        RECT 26.880 1.805 27.050 1.885 ;
        RECT 27.850 1.805 28.020 1.885 ;
        RECT 28.775 1.880 28.945 5.345 ;
        RECT 30.625 2.055 30.795 5.095 ;
        RECT 31.395 4.940 31.565 5.095 ;
        RECT 31.365 4.765 31.565 4.940 ;
        RECT 31.365 2.055 31.535 4.765 ;
        RECT 24.960 0.985 25.130 1.720 ;
        RECT 26.880 1.635 28.020 1.805 ;
        RECT 25.445 0.765 25.615 1.535 ;
        RECT 24.475 0.595 25.615 0.765 ;
        RECT 24.475 0.515 24.645 0.595 ;
        RECT 25.445 0.515 25.615 0.595 ;
        RECT 26.880 0.505 27.050 1.635 ;
        RECT 27.850 0.755 28.020 1.635 ;
        RECT 28.335 1.710 28.945 1.880 ;
        RECT 30.210 1.805 30.380 1.885 ;
        RECT 31.180 1.805 31.350 1.885 ;
        RECT 32.105 1.880 32.275 5.345 ;
        RECT 33.955 2.055 34.125 5.095 ;
        RECT 28.335 0.975 28.505 1.710 ;
        RECT 30.210 1.635 31.350 1.805 ;
        RECT 28.820 0.755 28.990 1.525 ;
        RECT 27.850 0.585 28.990 0.755 ;
        RECT 27.850 0.505 28.020 0.585 ;
        RECT 28.820 0.505 28.990 0.585 ;
        RECT 30.210 0.505 30.380 1.635 ;
        RECT 31.180 0.755 31.350 1.635 ;
        RECT 31.665 1.710 32.275 1.880 ;
        RECT 33.540 1.805 33.710 1.885 ;
        RECT 34.510 1.805 34.680 1.885 ;
        RECT 35.435 1.880 35.605 5.345 ;
        RECT 37.285 2.055 37.455 5.095 ;
        RECT 38.055 4.940 38.225 5.095 ;
        RECT 38.025 4.765 38.225 4.940 ;
        RECT 38.025 2.055 38.195 4.765 ;
        RECT 31.665 0.975 31.835 1.710 ;
        RECT 33.540 1.635 34.680 1.805 ;
        RECT 32.150 0.755 32.320 1.525 ;
        RECT 31.180 0.585 32.320 0.755 ;
        RECT 31.180 0.505 31.350 0.585 ;
        RECT 32.150 0.505 32.320 0.585 ;
        RECT 33.540 0.505 33.710 1.635 ;
        RECT 34.510 0.755 34.680 1.635 ;
        RECT 34.995 1.710 35.605 1.880 ;
        RECT 36.870 1.805 37.040 1.885 ;
        RECT 37.840 1.805 38.010 1.885 ;
        RECT 38.765 1.880 38.935 5.345 ;
        RECT 40.615 2.055 40.785 5.095 ;
        RECT 41.385 4.940 41.555 5.095 ;
        RECT 41.355 4.765 41.555 4.940 ;
        RECT 41.355 2.055 41.525 4.765 ;
        RECT 34.995 0.975 35.165 1.710 ;
        RECT 36.870 1.635 38.010 1.805 ;
        RECT 35.480 0.755 35.650 1.525 ;
        RECT 34.510 0.585 35.650 0.755 ;
        RECT 34.510 0.505 34.680 0.585 ;
        RECT 35.480 0.505 35.650 0.585 ;
        RECT 36.870 0.505 37.040 1.635 ;
        RECT 37.840 0.755 38.010 1.635 ;
        RECT 38.325 1.710 38.935 1.880 ;
        RECT 40.200 1.805 40.370 1.885 ;
        RECT 41.170 1.805 41.340 1.885 ;
        RECT 42.095 1.880 42.265 5.345 ;
        RECT 44.365 5.470 44.535 7.250 ;
        RECT 45.245 5.470 45.415 7.250 ;
        RECT 46.125 5.470 46.295 7.250 ;
        RECT 48.875 5.515 49.045 7.250 ;
        RECT 49.755 5.515 49.925 7.250 ;
        RECT 52.205 5.515 52.375 7.250 ;
        RECT 53.085 5.515 53.255 7.250 ;
        RECT 55.535 5.515 55.705 7.250 ;
        RECT 56.415 5.515 56.585 7.250 ;
        RECT 58.865 5.515 59.035 7.250 ;
        RECT 59.745 5.515 59.915 7.250 ;
        RECT 62.195 5.515 62.365 7.250 ;
        RECT 63.075 5.515 63.245 7.250 ;
        RECT 65.525 7.055 65.705 7.225 ;
        RECT 65.525 5.525 65.695 7.055 ;
        RECT 66.405 5.525 66.575 7.225 ;
        RECT 44.365 5.300 47.075 5.470 ;
        RECT 48.875 5.345 50.405 5.515 ;
        RECT 52.205 5.345 53.735 5.515 ;
        RECT 55.535 5.345 57.065 5.515 ;
        RECT 58.865 5.345 60.395 5.515 ;
        RECT 62.195 5.345 63.725 5.515 ;
        RECT 65.525 5.355 66.575 5.525 ;
        RECT 43.945 2.055 44.115 5.095 ;
        RECT 46.165 2.055 46.335 5.095 ;
        RECT 38.325 0.975 38.495 1.710 ;
        RECT 40.200 1.635 41.340 1.805 ;
        RECT 38.810 0.755 38.980 1.525 ;
        RECT 37.840 0.585 38.980 0.755 ;
        RECT 37.840 0.505 38.010 0.585 ;
        RECT 38.810 0.505 38.980 0.585 ;
        RECT 40.200 0.505 40.370 1.635 ;
        RECT 41.170 0.755 41.340 1.635 ;
        RECT 41.655 1.710 42.265 1.880 ;
        RECT 43.425 1.815 43.595 1.895 ;
        RECT 44.395 1.815 44.565 1.895 ;
        RECT 45.365 1.815 45.535 1.895 ;
        RECT 41.655 0.975 41.825 1.710 ;
        RECT 43.425 1.645 45.535 1.815 ;
        RECT 42.140 0.755 42.310 1.525 ;
        RECT 41.170 0.585 42.310 0.755 ;
        RECT 41.170 0.505 41.340 0.585 ;
        RECT 42.140 0.505 42.310 0.585 ;
        RECT 43.425 0.515 43.595 1.645 ;
        RECT 44.395 0.765 44.565 1.645 ;
        RECT 45.365 1.565 45.535 1.645 ;
        RECT 44.885 1.220 45.055 1.300 ;
        RECT 45.935 1.220 46.105 1.895 ;
        RECT 46.905 1.890 47.075 5.300 ;
        RECT 48.755 2.055 48.925 5.095 ;
        RECT 44.885 1.050 46.105 1.220 ;
        RECT 44.885 0.970 45.055 1.050 ;
        RECT 45.365 0.765 45.535 0.845 ;
        RECT 44.395 0.595 45.535 0.765 ;
        RECT 44.395 0.515 44.565 0.595 ;
        RECT 45.365 0.515 45.535 0.595 ;
        RECT 45.935 0.765 46.105 1.050 ;
        RECT 46.420 1.720 47.075 1.890 ;
        RECT 48.340 1.805 48.510 1.885 ;
        RECT 49.310 1.805 49.480 1.885 ;
        RECT 50.235 1.880 50.405 5.345 ;
        RECT 52.085 2.055 52.255 5.095 ;
        RECT 52.855 4.940 53.025 5.095 ;
        RECT 52.825 4.765 53.025 4.940 ;
        RECT 52.825 2.055 52.995 4.765 ;
        RECT 46.420 0.985 46.590 1.720 ;
        RECT 48.340 1.635 49.480 1.805 ;
        RECT 46.905 0.765 47.075 1.535 ;
        RECT 45.935 0.595 47.075 0.765 ;
        RECT 45.935 0.515 46.105 0.595 ;
        RECT 46.905 0.515 47.075 0.595 ;
        RECT 48.340 0.505 48.510 1.635 ;
        RECT 49.310 0.755 49.480 1.635 ;
        RECT 49.795 1.710 50.405 1.880 ;
        RECT 51.670 1.805 51.840 1.885 ;
        RECT 52.640 1.805 52.810 1.885 ;
        RECT 53.565 1.880 53.735 5.345 ;
        RECT 55.415 2.055 55.585 5.095 ;
        RECT 49.795 0.975 49.965 1.710 ;
        RECT 51.670 1.635 52.810 1.805 ;
        RECT 50.280 0.755 50.450 1.525 ;
        RECT 49.310 0.585 50.450 0.755 ;
        RECT 49.310 0.505 49.480 0.585 ;
        RECT 50.280 0.505 50.450 0.585 ;
        RECT 51.670 0.505 51.840 1.635 ;
        RECT 52.640 0.755 52.810 1.635 ;
        RECT 53.125 1.710 53.735 1.880 ;
        RECT 55.000 1.805 55.170 1.885 ;
        RECT 55.970 1.805 56.140 1.885 ;
        RECT 56.895 1.880 57.065 5.345 ;
        RECT 58.745 2.055 58.915 5.095 ;
        RECT 59.515 4.940 59.685 5.095 ;
        RECT 59.485 4.765 59.685 4.940 ;
        RECT 59.485 2.055 59.655 4.765 ;
        RECT 53.125 0.975 53.295 1.710 ;
        RECT 55.000 1.635 56.140 1.805 ;
        RECT 53.610 0.755 53.780 1.525 ;
        RECT 52.640 0.585 53.780 0.755 ;
        RECT 52.640 0.505 52.810 0.585 ;
        RECT 53.610 0.505 53.780 0.585 ;
        RECT 55.000 0.505 55.170 1.635 ;
        RECT 55.970 0.755 56.140 1.635 ;
        RECT 56.455 1.710 57.065 1.880 ;
        RECT 58.330 1.805 58.500 1.885 ;
        RECT 59.300 1.805 59.470 1.885 ;
        RECT 60.225 1.880 60.395 5.345 ;
        RECT 62.075 2.055 62.245 5.095 ;
        RECT 62.845 4.940 63.015 5.095 ;
        RECT 62.815 4.765 63.015 4.940 ;
        RECT 62.815 2.055 62.985 4.765 ;
        RECT 56.455 0.975 56.625 1.710 ;
        RECT 58.330 1.635 59.470 1.805 ;
        RECT 56.940 0.755 57.110 1.525 ;
        RECT 55.970 0.585 57.110 0.755 ;
        RECT 55.970 0.505 56.140 0.585 ;
        RECT 56.940 0.505 57.110 0.585 ;
        RECT 58.330 0.505 58.500 1.635 ;
        RECT 59.300 0.755 59.470 1.635 ;
        RECT 59.785 1.710 60.395 1.880 ;
        RECT 61.660 1.805 61.830 1.885 ;
        RECT 62.630 1.805 62.800 1.885 ;
        RECT 63.555 1.880 63.725 5.345 ;
        RECT 66.405 5.275 66.575 5.355 ;
        RECT 68.405 7.055 70.335 7.225 ;
        RECT 68.405 5.275 68.575 7.055 ;
        RECT 68.845 5.525 69.015 6.795 ;
        RECT 69.285 5.785 69.455 7.055 ;
        RECT 69.725 5.525 69.895 6.795 ;
        RECT 70.165 5.605 70.335 7.055 ;
        RECT 71.745 7.055 73.675 7.225 ;
        RECT 68.845 5.355 69.895 5.525 ;
        RECT 69.725 5.275 69.895 5.355 ;
        RECT 71.745 5.275 71.915 7.055 ;
        RECT 72.625 5.785 72.795 7.055 ;
        RECT 73.505 5.785 73.675 7.055 ;
        RECT 65.035 2.055 65.205 5.100 ;
        RECT 66.185 4.940 66.355 5.100 ;
        RECT 66.145 4.770 66.355 4.940 ;
        RECT 66.145 2.055 66.315 4.770 ;
        RECT 68.735 2.055 68.905 5.100 ;
        RECT 70.215 2.055 70.385 5.100 ;
        RECT 71.695 2.055 71.865 5.100 ;
        RECT 72.805 4.770 72.995 5.100 ;
        RECT 72.805 2.055 72.975 4.770 ;
        RECT 59.785 0.975 59.955 1.710 ;
        RECT 61.660 1.635 62.800 1.805 ;
        RECT 60.270 0.755 60.440 1.525 ;
        RECT 59.300 0.585 60.440 0.755 ;
        RECT 59.300 0.505 59.470 0.585 ;
        RECT 60.270 0.505 60.440 0.585 ;
        RECT 61.660 0.505 61.830 1.635 ;
        RECT 62.630 0.755 62.800 1.635 ;
        RECT 63.115 1.710 63.725 1.880 ;
        RECT 64.990 1.805 65.160 1.885 ;
        RECT 65.960 1.805 66.130 1.885 ;
        RECT 63.115 0.975 63.285 1.710 ;
        RECT 64.990 1.635 66.130 1.805 ;
        RECT 63.600 0.755 63.770 1.525 ;
        RECT 62.630 0.585 63.770 0.755 ;
        RECT 62.630 0.505 62.800 0.585 ;
        RECT 63.600 0.505 63.770 0.585 ;
        RECT 64.990 0.505 65.160 1.635 ;
        RECT 65.960 0.755 66.130 1.635 ;
        RECT 66.930 0.755 67.100 1.885 ;
        RECT 65.960 0.585 67.100 0.755 ;
        RECT 65.960 0.505 66.130 0.585 ;
        RECT 66.930 0.505 67.100 0.585 ;
        RECT 68.320 1.805 68.490 1.885 ;
        RECT 69.290 1.805 69.460 1.885 ;
        RECT 68.320 1.635 69.460 1.805 ;
        RECT 68.320 0.505 68.490 1.635 ;
        RECT 69.290 0.755 69.460 1.635 ;
        RECT 70.260 0.755 70.430 1.885 ;
        RECT 69.290 0.585 70.430 0.755 ;
        RECT 69.290 0.505 69.460 0.585 ;
        RECT 70.260 0.505 70.430 0.585 ;
        RECT 71.650 1.805 71.820 1.885 ;
        RECT 72.620 1.805 72.790 1.885 ;
        RECT 71.650 1.635 72.790 1.805 ;
        RECT 71.650 0.505 71.820 1.635 ;
        RECT 72.620 0.755 72.790 1.635 ;
        RECT 73.590 0.755 73.760 1.530 ;
        RECT 72.620 0.585 73.760 0.755 ;
        RECT 72.620 0.505 72.790 0.585 ;
        RECT 73.590 0.505 73.760 0.585 ;
      LAYER mcon ;
        RECT 1.025 4.355 1.195 4.525 ;
        RECT 3.245 3.615 3.415 3.785 ;
        RECT 3.985 3.985 4.155 4.155 ;
        RECT 5.835 3.985 6.005 4.155 ;
        RECT 7.315 3.615 7.485 3.785 ;
        RECT 9.165 3.615 9.335 3.785 ;
        RECT 9.905 4.355 10.075 4.525 ;
        RECT 10.645 3.615 10.815 3.785 ;
        RECT 12.495 3.615 12.665 3.785 ;
        RECT 13.975 4.355 14.145 4.525 ;
        RECT 15.825 3.985 15.995 4.155 ;
        RECT 16.565 3.245 16.735 3.415 ;
        RECT 17.305 3.985 17.475 4.155 ;
        RECT 19.155 3.985 19.325 4.155 ;
        RECT 19.895 4.355 20.065 4.525 ;
        RECT 20.635 3.245 20.805 3.415 ;
        RECT 22.485 4.355 22.655 4.525 ;
        RECT 24.705 3.615 24.875 3.785 ;
        RECT 25.445 3.985 25.615 4.155 ;
        RECT 27.295 3.985 27.465 4.155 ;
        RECT 28.775 3.615 28.945 3.785 ;
        RECT 30.625 3.615 30.795 3.785 ;
        RECT 31.365 4.355 31.535 4.525 ;
        RECT 32.105 3.615 32.275 3.785 ;
        RECT 33.955 3.615 34.125 3.785 ;
        RECT 35.435 4.355 35.605 4.525 ;
        RECT 37.285 3.985 37.455 4.155 ;
        RECT 38.025 2.505 38.195 2.675 ;
        RECT 38.765 3.985 38.935 4.155 ;
        RECT 40.615 3.985 40.785 4.155 ;
        RECT 41.355 4.355 41.525 4.525 ;
        RECT 66.405 5.355 66.575 5.525 ;
        RECT 42.095 2.505 42.265 2.675 ;
        RECT 43.945 4.355 44.115 4.525 ;
        RECT 46.165 3.615 46.335 3.785 ;
        RECT 46.905 3.985 47.075 4.155 ;
        RECT 48.755 3.985 48.925 4.155 ;
        RECT 50.235 3.615 50.405 3.785 ;
        RECT 52.085 3.615 52.255 3.785 ;
        RECT 52.825 4.355 52.995 4.525 ;
        RECT 53.565 3.615 53.735 3.785 ;
        RECT 55.415 3.615 55.585 3.785 ;
        RECT 56.895 4.355 57.065 4.525 ;
        RECT 58.745 3.985 58.915 4.155 ;
        RECT 59.485 3.985 59.655 4.155 ;
        RECT 60.225 4.725 60.395 4.895 ;
        RECT 62.075 4.725 62.245 4.895 ;
        RECT 62.815 4.355 62.985 4.525 ;
        RECT 68.405 5.355 68.575 5.525 ;
        RECT 69.725 5.355 69.895 5.525 ;
        RECT 71.745 5.355 71.915 5.525 ;
        RECT 63.555 3.985 63.725 4.155 ;
        RECT 65.035 4.725 65.205 4.895 ;
        RECT 65.035 3.985 65.205 4.155 ;
        RECT 66.145 4.355 66.315 4.525 ;
        RECT 66.145 2.505 66.315 2.675 ;
        RECT 68.735 4.725 68.905 4.895 ;
        RECT 70.215 3.245 70.385 3.415 ;
        RECT 70.215 2.135 70.385 2.305 ;
        RECT 71.695 2.135 71.865 2.305 ;
        RECT 72.805 4.355 72.975 4.525 ;
      LAYER met1 ;
        RECT 66.375 5.525 66.605 5.555 ;
        RECT 68.375 5.525 68.605 5.555 ;
        RECT 69.695 5.525 69.925 5.555 ;
        RECT 71.715 5.525 71.945 5.555 ;
        RECT 66.345 5.355 68.635 5.525 ;
        RECT 69.665 5.355 71.975 5.525 ;
        RECT 66.375 5.325 66.605 5.355 ;
        RECT 68.375 5.325 68.605 5.355 ;
        RECT 69.695 5.325 69.925 5.355 ;
        RECT 71.715 5.325 71.945 5.355 ;
        RECT 60.195 4.895 60.425 4.925 ;
        RECT 62.045 4.895 62.275 4.925 ;
        RECT 65.005 4.895 65.235 4.925 ;
        RECT 68.705 4.895 68.935 4.925 ;
        RECT 60.165 4.725 62.305 4.895 ;
        RECT 64.975 4.725 68.965 4.895 ;
        RECT 60.195 4.695 60.425 4.725 ;
        RECT 62.045 4.695 62.275 4.725 ;
        RECT 65.005 4.695 65.235 4.725 ;
        RECT 68.705 4.695 68.935 4.725 ;
        RECT 0.995 4.525 1.225 4.555 ;
        RECT 9.875 4.525 10.105 4.555 ;
        RECT 13.945 4.525 14.175 4.555 ;
        RECT 19.865 4.525 20.095 4.555 ;
        RECT 22.455 4.525 22.685 4.555 ;
        RECT 31.335 4.525 31.565 4.555 ;
        RECT 35.405 4.525 35.635 4.555 ;
        RECT 41.325 4.525 41.555 4.555 ;
        RECT 43.915 4.525 44.145 4.555 ;
        RECT 52.795 4.525 53.025 4.555 ;
        RECT 56.865 4.525 57.095 4.555 ;
        RECT 62.785 4.525 63.015 4.555 ;
        RECT 66.115 4.525 66.345 4.555 ;
        RECT 72.775 4.525 73.005 4.555 ;
        RECT 0.965 4.355 20.125 4.525 ;
        RECT 22.425 4.355 41.585 4.525 ;
        RECT 43.885 4.355 63.045 4.525 ;
        RECT 66.085 4.355 73.035 4.525 ;
        RECT 0.995 4.325 1.225 4.355 ;
        RECT 9.875 4.325 10.105 4.355 ;
        RECT 13.945 4.325 14.175 4.355 ;
        RECT 19.865 4.325 20.095 4.355 ;
        RECT 22.455 4.325 22.685 4.355 ;
        RECT 31.335 4.325 31.565 4.355 ;
        RECT 35.405 4.325 35.635 4.355 ;
        RECT 41.325 4.325 41.555 4.355 ;
        RECT 43.915 4.325 44.145 4.355 ;
        RECT 52.795 4.325 53.025 4.355 ;
        RECT 56.865 4.325 57.095 4.355 ;
        RECT 62.785 4.325 63.015 4.355 ;
        RECT 66.115 4.325 66.345 4.355 ;
        RECT 72.775 4.325 73.005 4.355 ;
        RECT 3.955 4.155 4.185 4.185 ;
        RECT 5.805 4.155 6.035 4.185 ;
        RECT 15.795 4.155 16.025 4.185 ;
        RECT 17.275 4.155 17.505 4.185 ;
        RECT 19.125 4.155 19.355 4.185 ;
        RECT 25.415 4.155 25.645 4.185 ;
        RECT 27.265 4.155 27.495 4.185 ;
        RECT 37.255 4.155 37.485 4.185 ;
        RECT 38.735 4.155 38.965 4.185 ;
        RECT 40.585 4.155 40.815 4.185 ;
        RECT 46.875 4.155 47.105 4.185 ;
        RECT 48.725 4.155 48.955 4.185 ;
        RECT 58.715 4.155 58.945 4.185 ;
        RECT 59.455 4.155 59.685 4.185 ;
        RECT 63.525 4.155 63.755 4.185 ;
        RECT 65.005 4.155 65.235 4.185 ;
        RECT 3.925 3.985 16.055 4.155 ;
        RECT 17.245 3.985 19.385 4.155 ;
        RECT 25.385 3.985 37.515 4.155 ;
        RECT 38.705 3.985 40.845 4.155 ;
        RECT 46.845 3.985 58.975 4.155 ;
        RECT 59.425 3.985 65.265 4.155 ;
        RECT 3.955 3.955 4.185 3.985 ;
        RECT 5.805 3.955 6.035 3.985 ;
        RECT 15.795 3.955 16.025 3.985 ;
        RECT 17.275 3.955 17.505 3.985 ;
        RECT 19.125 3.955 19.355 3.985 ;
        RECT 25.415 3.955 25.645 3.985 ;
        RECT 27.265 3.955 27.495 3.985 ;
        RECT 37.255 3.955 37.485 3.985 ;
        RECT 38.735 3.955 38.965 3.985 ;
        RECT 40.585 3.955 40.815 3.985 ;
        RECT 46.875 3.955 47.105 3.985 ;
        RECT 48.725 3.955 48.955 3.985 ;
        RECT 58.715 3.955 58.945 3.985 ;
        RECT 59.455 3.955 59.685 3.985 ;
        RECT 63.525 3.955 63.755 3.985 ;
        RECT 65.005 3.955 65.235 3.985 ;
        RECT 3.215 3.785 3.445 3.815 ;
        RECT 7.285 3.785 7.515 3.815 ;
        RECT 9.135 3.785 9.365 3.815 ;
        RECT 10.615 3.785 10.845 3.815 ;
        RECT 12.465 3.785 12.695 3.815 ;
        RECT 24.675 3.785 24.905 3.815 ;
        RECT 28.745 3.785 28.975 3.815 ;
        RECT 30.595 3.785 30.825 3.815 ;
        RECT 32.075 3.785 32.305 3.815 ;
        RECT 33.925 3.785 34.155 3.815 ;
        RECT 46.135 3.785 46.365 3.815 ;
        RECT 50.205 3.785 50.435 3.815 ;
        RECT 52.055 3.785 52.285 3.815 ;
        RECT 53.535 3.785 53.765 3.815 ;
        RECT 55.385 3.785 55.615 3.815 ;
        RECT 3.185 3.615 9.395 3.785 ;
        RECT 10.585 3.615 12.725 3.785 ;
        RECT 24.645 3.615 30.855 3.785 ;
        RECT 32.045 3.615 34.185 3.785 ;
        RECT 46.105 3.615 52.315 3.785 ;
        RECT 53.505 3.615 55.645 3.785 ;
        RECT 3.215 3.585 3.445 3.615 ;
        RECT 7.285 3.585 7.515 3.615 ;
        RECT 9.135 3.585 9.365 3.615 ;
        RECT 10.615 3.585 10.845 3.615 ;
        RECT 12.465 3.585 12.695 3.615 ;
        RECT 24.675 3.585 24.905 3.615 ;
        RECT 28.745 3.585 28.975 3.615 ;
        RECT 30.595 3.585 30.825 3.615 ;
        RECT 32.075 3.585 32.305 3.615 ;
        RECT 33.925 3.585 34.155 3.615 ;
        RECT 46.135 3.585 46.365 3.615 ;
        RECT 50.205 3.585 50.435 3.615 ;
        RECT 52.055 3.585 52.285 3.615 ;
        RECT 53.535 3.585 53.765 3.615 ;
        RECT 55.385 3.585 55.615 3.615 ;
        RECT 16.535 3.415 16.765 3.445 ;
        RECT 20.605 3.415 20.835 3.445 ;
        RECT 70.185 3.415 70.415 3.445 ;
        RECT 16.505 3.245 70.445 3.415 ;
        RECT 16.535 3.215 16.765 3.245 ;
        RECT 20.605 3.215 20.835 3.245 ;
        RECT 70.185 3.215 70.415 3.245 ;
        RECT 37.995 2.675 38.225 2.705 ;
        RECT 42.065 2.675 42.295 2.705 ;
        RECT 66.115 2.675 66.345 2.705 ;
        RECT 37.965 2.505 66.375 2.675 ;
        RECT 37.995 2.475 38.225 2.505 ;
        RECT 42.065 2.475 42.295 2.505 ;
        RECT 66.115 2.475 66.345 2.505 ;
        RECT 70.185 2.305 70.415 2.335 ;
        RECT 71.665 2.305 71.895 2.335 ;
        RECT 70.155 2.135 71.925 2.305 ;
        RECT 70.185 2.105 70.415 2.135 ;
        RECT 71.665 2.105 71.895 2.135 ;
  END
END TMRDFFQNX1






MACRO TMRDFFQX1
  CLASS BLOCK ;
  FOREIGN TMRDFFQX1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 77.430 BY 7.950 ;
  PIN D
    ANTENNAGATEAREA 3.081750 ;
    PORT
      LAYER li1 ;
        RECT 6.605 4.940 6.775 5.095 ;
        RECT 28.065 4.940 28.235 5.095 ;
        RECT 49.525 4.940 49.695 5.095 ;
        RECT 6.575 4.765 6.775 4.940 ;
        RECT 28.035 4.765 28.235 4.940 ;
        RECT 49.495 4.765 49.695 4.940 ;
        RECT 6.575 2.055 6.745 4.765 ;
        RECT 28.035 2.055 28.205 4.765 ;
        RECT 49.495 2.055 49.665 4.765 ;
      LAYER mcon ;
        RECT 6.575 2.135 6.745 2.305 ;
        RECT 28.035 2.135 28.205 2.305 ;
        RECT 49.495 2.135 49.665 2.305 ;
      LAYER met1 ;
        RECT 6.545 2.305 6.775 2.335 ;
        RECT 28.005 2.305 28.235 2.335 ;
        RECT 49.465 2.305 49.695 2.335 ;
        RECT 6.395 2.135 49.725 2.305 ;
        RECT 6.545 2.105 6.775 2.135 ;
        RECT 28.005 2.105 28.235 2.135 ;
        RECT 49.465 2.105 49.695 2.135 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 6.126300 ;
    PORT
      LAYER li1 ;
        RECT 2.135 2.055 2.305 5.095 ;
        RECT 13.265 4.975 13.435 5.095 ;
        RECT 13.235 4.765 13.435 4.975 ;
        RECT 13.235 2.055 13.405 4.765 ;
        RECT 23.595 2.055 23.765 5.095 ;
        RECT 34.725 4.975 34.895 5.095 ;
        RECT 34.695 4.765 34.895 4.975 ;
        RECT 34.695 2.055 34.865 4.765 ;
        RECT 45.055 2.055 45.225 5.095 ;
        RECT 56.185 4.975 56.355 5.095 ;
        RECT 56.155 4.765 56.355 4.975 ;
        RECT 56.155 2.055 56.325 4.765 ;
      LAYER mcon ;
        RECT 2.135 4.725 2.305 4.895 ;
        RECT 13.235 4.725 13.405 4.895 ;
        RECT 23.595 4.725 23.765 4.895 ;
        RECT 34.695 4.725 34.865 4.895 ;
        RECT 45.055 4.725 45.225 4.895 ;
        RECT 56.155 4.725 56.325 4.895 ;
      LAYER met1 ;
        RECT 2.105 4.895 2.335 4.925 ;
        RECT 13.205 4.895 13.435 4.925 ;
        RECT 23.565 4.895 23.795 4.925 ;
        RECT 34.665 4.895 34.895 4.925 ;
        RECT 45.025 4.895 45.255 4.925 ;
        RECT 56.125 4.895 56.355 4.925 ;
        RECT 2.075 4.890 13.465 4.895 ;
        RECT 16.745 4.890 56.385 4.895 ;
        RECT 2.075 4.735 56.385 4.890 ;
        RECT 2.075 4.725 13.465 4.735 ;
        RECT 16.745 4.725 56.385 4.735 ;
        RECT 2.105 4.695 2.335 4.725 ;
        RECT 13.205 4.695 13.435 4.725 ;
        RECT 23.565 4.695 23.795 4.725 ;
        RECT 34.665 4.695 34.895 4.725 ;
        RECT 45.025 4.695 45.255 4.725 ;
        RECT 56.125 4.695 56.355 4.725 ;
    END
  END CLK
  PIN VDD
    ANTENNADIFFAREA 92.170746 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 77.010 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 76.745 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 1.005 5.445 1.175 7.460 ;
        RECT 1.885 5.785 2.055 7.460 ;
        RECT 2.765 5.785 2.935 7.460 ;
        RECT 3.645 5.785 3.815 7.460 ;
        RECT 4.655 4.340 4.965 7.460 ;
        RECT 5.515 5.365 5.685 7.460 ;
        RECT 6.395 5.785 6.565 7.460 ;
        RECT 7.275 5.785 7.445 7.460 ;
        RECT 7.985 4.340 8.295 7.460 ;
        RECT 8.845 5.365 9.015 7.460 ;
        RECT 9.725 5.785 9.895 7.460 ;
        RECT 10.605 5.785 10.775 7.460 ;
        RECT 11.315 4.340 11.625 7.460 ;
        RECT 12.175 5.365 12.345 7.460 ;
        RECT 13.055 5.785 13.225 7.460 ;
        RECT 13.935 5.785 14.105 7.460 ;
        RECT 14.645 4.340 14.955 7.460 ;
        RECT 15.505 5.365 15.675 7.460 ;
        RECT 16.385 5.785 16.555 7.460 ;
        RECT 17.265 5.785 17.435 7.460 ;
        RECT 17.975 4.340 18.285 7.460 ;
        RECT 18.835 5.365 19.005 7.460 ;
        RECT 19.715 5.785 19.885 7.460 ;
        RECT 20.595 5.785 20.765 7.460 ;
        RECT 21.305 4.340 21.615 7.460 ;
        RECT 22.465 5.445 22.635 7.460 ;
        RECT 23.345 5.785 23.515 7.460 ;
        RECT 24.225 5.785 24.395 7.460 ;
        RECT 25.105 5.785 25.275 7.460 ;
        RECT 26.115 4.340 26.425 7.460 ;
        RECT 26.975 5.365 27.145 7.460 ;
        RECT 27.855 5.785 28.025 7.460 ;
        RECT 28.735 5.785 28.905 7.460 ;
        RECT 29.445 4.340 29.755 7.460 ;
        RECT 30.305 5.365 30.475 7.460 ;
        RECT 31.185 5.785 31.355 7.460 ;
        RECT 32.065 5.785 32.235 7.460 ;
        RECT 32.775 4.340 33.085 7.460 ;
        RECT 33.635 5.365 33.805 7.460 ;
        RECT 34.515 5.785 34.685 7.460 ;
        RECT 35.395 5.785 35.565 7.460 ;
        RECT 36.105 4.340 36.415 7.460 ;
        RECT 36.965 5.365 37.135 7.460 ;
        RECT 37.845 5.785 38.015 7.460 ;
        RECT 38.725 5.785 38.895 7.460 ;
        RECT 39.435 4.340 39.745 7.460 ;
        RECT 40.295 5.365 40.465 7.460 ;
        RECT 41.175 5.785 41.345 7.460 ;
        RECT 42.055 5.785 42.225 7.460 ;
        RECT 42.765 4.340 43.075 7.460 ;
        RECT 43.925 5.445 44.095 7.460 ;
        RECT 44.805 5.785 44.975 7.460 ;
        RECT 45.685 5.785 45.855 7.460 ;
        RECT 46.565 5.785 46.735 7.460 ;
        RECT 47.575 4.340 47.885 7.460 ;
        RECT 48.435 5.365 48.605 7.460 ;
        RECT 49.315 5.785 49.485 7.460 ;
        RECT 50.195 5.785 50.365 7.460 ;
        RECT 50.905 4.340 51.215 7.460 ;
        RECT 51.765 5.365 51.935 7.460 ;
        RECT 52.645 5.785 52.815 7.460 ;
        RECT 53.525 5.785 53.695 7.460 ;
        RECT 54.235 4.340 54.545 7.460 ;
        RECT 55.095 5.365 55.265 7.460 ;
        RECT 55.975 5.785 56.145 7.460 ;
        RECT 56.855 5.785 57.025 7.460 ;
        RECT 57.565 4.340 57.875 7.460 ;
        RECT 58.425 5.365 58.595 7.460 ;
        RECT 59.305 5.785 59.475 7.460 ;
        RECT 60.185 5.785 60.355 7.460 ;
        RECT 60.895 4.340 61.205 7.460 ;
        RECT 61.755 5.365 61.925 7.460 ;
        RECT 62.635 5.785 62.805 7.460 ;
        RECT 63.515 5.785 63.685 7.460 ;
        RECT 64.225 4.340 64.535 7.460 ;
        RECT 65.085 5.355 65.255 7.460 ;
        RECT 65.965 5.785 66.135 7.460 ;
        RECT 66.845 5.355 67.015 7.460 ;
        RECT 67.555 4.340 67.865 7.460 ;
        RECT 70.885 4.340 71.195 7.460 ;
        RECT 74.215 4.340 74.525 7.460 ;
        RECT 74.955 5.415 75.125 7.460 ;
        RECT 75.835 5.415 76.005 7.460 ;
        RECT 76.435 4.340 76.745 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 0.995 7.525 1.165 7.695 ;
        RECT 1.355 7.525 1.525 7.695 ;
        RECT 1.715 7.525 1.885 7.695 ;
        RECT 2.075 7.525 2.245 7.695 ;
        RECT 2.565 7.525 2.735 7.695 ;
        RECT 2.925 7.525 3.095 7.695 ;
        RECT 3.285 7.525 3.455 7.695 ;
        RECT 3.645 7.525 3.815 7.695 ;
        RECT 4.005 7.525 4.175 7.695 ;
        RECT 4.365 7.525 4.535 7.695 ;
        RECT 5.085 7.525 5.255 7.695 ;
        RECT 5.445 7.525 5.615 7.695 ;
        RECT 5.805 7.525 5.975 7.695 ;
        RECT 6.165 7.525 6.335 7.695 ;
        RECT 6.615 7.525 6.785 7.695 ;
        RECT 6.975 7.525 7.145 7.695 ;
        RECT 7.335 7.525 7.505 7.695 ;
        RECT 7.695 7.525 7.865 7.695 ;
        RECT 8.415 7.525 8.585 7.695 ;
        RECT 8.775 7.525 8.945 7.695 ;
        RECT 9.135 7.525 9.305 7.695 ;
        RECT 9.495 7.525 9.665 7.695 ;
        RECT 9.945 7.525 10.115 7.695 ;
        RECT 10.305 7.525 10.475 7.695 ;
        RECT 10.665 7.525 10.835 7.695 ;
        RECT 11.025 7.525 11.195 7.695 ;
        RECT 11.745 7.525 11.915 7.695 ;
        RECT 12.105 7.525 12.275 7.695 ;
        RECT 12.465 7.525 12.635 7.695 ;
        RECT 12.825 7.525 12.995 7.695 ;
        RECT 13.275 7.525 13.445 7.695 ;
        RECT 13.635 7.525 13.805 7.695 ;
        RECT 13.995 7.525 14.165 7.695 ;
        RECT 14.355 7.525 14.525 7.695 ;
        RECT 15.075 7.525 15.245 7.695 ;
        RECT 15.435 7.525 15.605 7.695 ;
        RECT 15.795 7.525 15.965 7.695 ;
        RECT 16.155 7.525 16.325 7.695 ;
        RECT 16.605 7.525 16.775 7.695 ;
        RECT 16.965 7.525 17.135 7.695 ;
        RECT 17.325 7.525 17.495 7.695 ;
        RECT 17.685 7.525 17.855 7.695 ;
        RECT 18.405 7.525 18.575 7.695 ;
        RECT 18.765 7.525 18.935 7.695 ;
        RECT 19.125 7.525 19.295 7.695 ;
        RECT 19.485 7.525 19.655 7.695 ;
        RECT 19.935 7.525 20.105 7.695 ;
        RECT 20.295 7.525 20.465 7.695 ;
        RECT 20.655 7.525 20.825 7.695 ;
        RECT 21.015 7.525 21.185 7.695 ;
        RECT 21.735 7.525 21.905 7.695 ;
        RECT 22.095 7.525 22.265 7.695 ;
        RECT 22.455 7.525 22.625 7.695 ;
        RECT 22.815 7.525 22.985 7.695 ;
        RECT 23.175 7.525 23.345 7.695 ;
        RECT 23.535 7.525 23.705 7.695 ;
        RECT 24.025 7.525 24.195 7.695 ;
        RECT 24.385 7.525 24.555 7.695 ;
        RECT 24.745 7.525 24.915 7.695 ;
        RECT 25.105 7.525 25.275 7.695 ;
        RECT 25.465 7.525 25.635 7.695 ;
        RECT 25.825 7.525 25.995 7.695 ;
        RECT 26.545 7.525 26.715 7.695 ;
        RECT 26.905 7.525 27.075 7.695 ;
        RECT 27.265 7.525 27.435 7.695 ;
        RECT 27.625 7.525 27.795 7.695 ;
        RECT 28.075 7.525 28.245 7.695 ;
        RECT 28.435 7.525 28.605 7.695 ;
        RECT 28.795 7.525 28.965 7.695 ;
        RECT 29.155 7.525 29.325 7.695 ;
        RECT 29.875 7.525 30.045 7.695 ;
        RECT 30.235 7.525 30.405 7.695 ;
        RECT 30.595 7.525 30.765 7.695 ;
        RECT 30.955 7.525 31.125 7.695 ;
        RECT 31.405 7.525 31.575 7.695 ;
        RECT 31.765 7.525 31.935 7.695 ;
        RECT 32.125 7.525 32.295 7.695 ;
        RECT 32.485 7.525 32.655 7.695 ;
        RECT 33.205 7.525 33.375 7.695 ;
        RECT 33.565 7.525 33.735 7.695 ;
        RECT 33.925 7.525 34.095 7.695 ;
        RECT 34.285 7.525 34.455 7.695 ;
        RECT 34.735 7.525 34.905 7.695 ;
        RECT 35.095 7.525 35.265 7.695 ;
        RECT 35.455 7.525 35.625 7.695 ;
        RECT 35.815 7.525 35.985 7.695 ;
        RECT 36.535 7.525 36.705 7.695 ;
        RECT 36.895 7.525 37.065 7.695 ;
        RECT 37.255 7.525 37.425 7.695 ;
        RECT 37.615 7.525 37.785 7.695 ;
        RECT 38.065 7.525 38.235 7.695 ;
        RECT 38.425 7.525 38.595 7.695 ;
        RECT 38.785 7.525 38.955 7.695 ;
        RECT 39.145 7.525 39.315 7.695 ;
        RECT 39.865 7.525 40.035 7.695 ;
        RECT 40.225 7.525 40.395 7.695 ;
        RECT 40.585 7.525 40.755 7.695 ;
        RECT 40.945 7.525 41.115 7.695 ;
        RECT 41.395 7.525 41.565 7.695 ;
        RECT 41.755 7.525 41.925 7.695 ;
        RECT 42.115 7.525 42.285 7.695 ;
        RECT 42.475 7.525 42.645 7.695 ;
        RECT 43.195 7.525 43.365 7.695 ;
        RECT 43.555 7.525 43.725 7.695 ;
        RECT 43.915 7.525 44.085 7.695 ;
        RECT 44.275 7.525 44.445 7.695 ;
        RECT 44.635 7.525 44.805 7.695 ;
        RECT 44.995 7.525 45.165 7.695 ;
        RECT 45.485 7.525 45.655 7.695 ;
        RECT 45.845 7.525 46.015 7.695 ;
        RECT 46.205 7.525 46.375 7.695 ;
        RECT 46.565 7.525 46.735 7.695 ;
        RECT 46.925 7.525 47.095 7.695 ;
        RECT 47.285 7.525 47.455 7.695 ;
        RECT 48.005 7.525 48.175 7.695 ;
        RECT 48.365 7.525 48.535 7.695 ;
        RECT 48.725 7.525 48.895 7.695 ;
        RECT 49.085 7.525 49.255 7.695 ;
        RECT 49.535 7.525 49.705 7.695 ;
        RECT 49.895 7.525 50.065 7.695 ;
        RECT 50.255 7.525 50.425 7.695 ;
        RECT 50.615 7.525 50.785 7.695 ;
        RECT 51.335 7.525 51.505 7.695 ;
        RECT 51.695 7.525 51.865 7.695 ;
        RECT 52.055 7.525 52.225 7.695 ;
        RECT 52.415 7.525 52.585 7.695 ;
        RECT 52.865 7.525 53.035 7.695 ;
        RECT 53.225 7.525 53.395 7.695 ;
        RECT 53.585 7.525 53.755 7.695 ;
        RECT 53.945 7.525 54.115 7.695 ;
        RECT 54.665 7.525 54.835 7.695 ;
        RECT 55.025 7.525 55.195 7.695 ;
        RECT 55.385 7.525 55.555 7.695 ;
        RECT 55.745 7.525 55.915 7.695 ;
        RECT 56.195 7.525 56.365 7.695 ;
        RECT 56.555 7.525 56.725 7.695 ;
        RECT 56.915 7.525 57.085 7.695 ;
        RECT 57.275 7.525 57.445 7.695 ;
        RECT 57.995 7.525 58.165 7.695 ;
        RECT 58.355 7.525 58.525 7.695 ;
        RECT 58.715 7.525 58.885 7.695 ;
        RECT 59.075 7.525 59.245 7.695 ;
        RECT 59.525 7.525 59.695 7.695 ;
        RECT 59.885 7.525 60.055 7.695 ;
        RECT 60.245 7.525 60.415 7.695 ;
        RECT 60.605 7.525 60.775 7.695 ;
        RECT 61.325 7.525 61.495 7.695 ;
        RECT 61.685 7.525 61.855 7.695 ;
        RECT 62.045 7.525 62.215 7.695 ;
        RECT 62.405 7.525 62.575 7.695 ;
        RECT 62.855 7.525 63.025 7.695 ;
        RECT 63.215 7.525 63.385 7.695 ;
        RECT 63.575 7.525 63.745 7.695 ;
        RECT 63.935 7.525 64.105 7.695 ;
        RECT 64.655 7.525 64.825 7.695 ;
        RECT 65.015 7.525 65.185 7.695 ;
        RECT 65.375 7.525 65.545 7.695 ;
        RECT 65.735 7.525 65.905 7.695 ;
        RECT 66.185 7.525 66.355 7.695 ;
        RECT 66.545 7.525 66.715 7.695 ;
        RECT 66.905 7.525 67.075 7.695 ;
        RECT 67.265 7.525 67.435 7.695 ;
        RECT 67.985 7.525 68.155 7.695 ;
        RECT 68.345 7.525 68.515 7.695 ;
        RECT 68.705 7.525 68.875 7.695 ;
        RECT 69.065 7.525 69.235 7.695 ;
        RECT 69.515 7.525 69.685 7.695 ;
        RECT 69.875 7.525 70.045 7.695 ;
        RECT 70.235 7.525 70.405 7.695 ;
        RECT 70.595 7.525 70.765 7.695 ;
        RECT 71.315 7.525 71.485 7.695 ;
        RECT 71.675 7.525 71.845 7.695 ;
        RECT 72.035 7.525 72.205 7.695 ;
        RECT 72.395 7.525 72.565 7.695 ;
        RECT 72.845 7.525 73.015 7.695 ;
        RECT 73.205 7.525 73.375 7.695 ;
        RECT 73.565 7.525 73.735 7.695 ;
        RECT 73.925 7.525 74.095 7.695 ;
        RECT 74.645 7.525 74.815 7.695 ;
        RECT 75.005 7.525 75.175 7.695 ;
        RECT 75.395 7.525 75.565 7.695 ;
        RECT 75.785 7.525 75.955 7.695 ;
        RECT 76.145 7.525 76.315 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 76.745 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 58.696899 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 76.875 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 4.525 -0.075 5.095 -0.065 ;
        RECT 7.855 -0.075 8.425 -0.065 ;
        RECT 11.185 -0.075 11.755 -0.065 ;
        RECT 14.515 -0.075 15.085 -0.065 ;
        RECT 17.845 -0.075 18.415 -0.065 ;
        RECT 21.175 -0.075 21.745 -0.065 ;
        RECT 25.985 -0.075 26.555 -0.065 ;
        RECT 29.315 -0.075 29.885 -0.065 ;
        RECT 32.645 -0.075 33.215 -0.065 ;
        RECT 35.975 -0.075 36.545 -0.065 ;
        RECT 39.305 -0.075 39.875 -0.065 ;
        RECT 42.635 -0.075 43.205 -0.065 ;
        RECT 47.445 -0.075 48.015 -0.065 ;
        RECT 50.775 -0.075 51.345 -0.065 ;
        RECT 54.105 -0.075 54.675 -0.065 ;
        RECT 57.435 -0.075 58.005 -0.065 ;
        RECT 60.765 -0.075 61.335 -0.065 ;
        RECT 64.095 -0.075 64.665 -0.065 ;
        RECT 67.425 -0.075 67.995 -0.065 ;
        RECT 70.755 -0.075 71.325 -0.065 ;
        RECT 74.085 -0.075 74.655 -0.065 ;
        RECT 76.305 -0.075 76.875 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 0.990 0.310 1.160 1.270 ;
        RECT 4.655 0.310 4.965 2.860 ;
        RECT 5.905 0.310 6.075 1.260 ;
        RECT 7.985 0.310 8.295 2.860 ;
        RECT 9.235 0.310 9.405 1.260 ;
        RECT 11.315 0.310 11.625 2.860 ;
        RECT 12.565 0.310 12.735 1.260 ;
        RECT 14.645 0.310 14.955 2.860 ;
        RECT 15.895 0.310 16.065 1.260 ;
        RECT 17.975 0.310 18.285 2.860 ;
        RECT 19.225 0.310 19.395 1.260 ;
        RECT 21.305 0.310 21.615 2.860 ;
        RECT 22.450 0.310 22.620 1.270 ;
        RECT 26.115 0.310 26.425 2.860 ;
        RECT 27.365 0.310 27.535 1.260 ;
        RECT 29.445 0.310 29.755 2.860 ;
        RECT 30.695 0.310 30.865 1.260 ;
        RECT 32.775 0.310 33.085 2.860 ;
        RECT 34.025 0.310 34.195 1.260 ;
        RECT 36.105 0.310 36.415 2.860 ;
        RECT 37.355 0.310 37.525 1.260 ;
        RECT 39.435 0.310 39.745 2.860 ;
        RECT 40.685 0.310 40.855 1.260 ;
        RECT 42.765 0.310 43.075 2.860 ;
        RECT 43.910 0.310 44.080 1.270 ;
        RECT 47.575 0.310 47.885 2.860 ;
        RECT 48.825 0.310 48.995 1.260 ;
        RECT 50.905 0.310 51.215 2.860 ;
        RECT 52.155 0.310 52.325 1.260 ;
        RECT 54.235 0.310 54.545 2.860 ;
        RECT 55.485 0.310 55.655 1.260 ;
        RECT 57.565 0.310 57.875 2.860 ;
        RECT 58.815 0.310 58.985 1.260 ;
        RECT 60.895 0.310 61.205 2.860 ;
        RECT 62.145 0.310 62.315 1.260 ;
        RECT 64.225 0.310 64.535 2.860 ;
        RECT 65.475 0.310 65.645 1.260 ;
        RECT 67.555 0.310 67.865 2.860 ;
        RECT 68.805 0.310 68.975 1.260 ;
        RECT 70.885 0.310 71.195 2.860 ;
        RECT 72.135 0.310 72.305 1.260 ;
        RECT 74.215 0.310 74.525 2.860 ;
        RECT 74.915 0.755 75.085 1.885 ;
        RECT 75.885 0.755 76.055 1.885 ;
        RECT 74.915 0.585 76.055 0.755 ;
        RECT 74.915 0.310 75.085 0.585 ;
        RECT 75.400 0.310 75.570 0.585 ;
        RECT 75.885 0.310 76.055 0.585 ;
        RECT 76.435 0.310 76.745 2.860 ;
        RECT -0.155 0.235 69.775 0.310 ;
        RECT 69.945 0.235 76.745 0.310 ;
        RECT -0.155 0.000 76.745 0.235 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 0.995 0.065 1.165 0.235 ;
        RECT 1.355 0.065 1.525 0.235 ;
        RECT 1.715 0.065 1.885 0.235 ;
        RECT 2.075 0.065 2.245 0.235 ;
        RECT 2.565 0.065 2.735 0.235 ;
        RECT 2.925 0.065 3.095 0.235 ;
        RECT 3.285 0.065 3.455 0.235 ;
        RECT 3.645 0.065 3.815 0.235 ;
        RECT 4.005 0.065 4.175 0.235 ;
        RECT 4.365 0.065 4.535 0.235 ;
        RECT 5.085 0.065 5.255 0.235 ;
        RECT 5.445 0.065 5.615 0.235 ;
        RECT 5.805 0.065 5.975 0.235 ;
        RECT 6.165 0.065 6.335 0.235 ;
        RECT 6.615 0.065 6.785 0.235 ;
        RECT 6.975 0.065 7.145 0.235 ;
        RECT 7.335 0.065 7.505 0.235 ;
        RECT 7.695 0.065 7.865 0.235 ;
        RECT 8.415 0.065 8.585 0.235 ;
        RECT 8.775 0.065 8.945 0.235 ;
        RECT 9.135 0.065 9.305 0.235 ;
        RECT 9.495 0.065 9.665 0.235 ;
        RECT 9.945 0.065 10.115 0.235 ;
        RECT 10.305 0.065 10.475 0.235 ;
        RECT 10.665 0.065 10.835 0.235 ;
        RECT 11.025 0.065 11.195 0.235 ;
        RECT 11.745 0.065 11.915 0.235 ;
        RECT 12.105 0.065 12.275 0.235 ;
        RECT 12.465 0.065 12.635 0.235 ;
        RECT 12.825 0.065 12.995 0.235 ;
        RECT 13.275 0.065 13.445 0.235 ;
        RECT 13.635 0.065 13.805 0.235 ;
        RECT 13.995 0.065 14.165 0.235 ;
        RECT 14.355 0.065 14.525 0.235 ;
        RECT 15.075 0.065 15.245 0.235 ;
        RECT 15.435 0.065 15.605 0.235 ;
        RECT 15.795 0.065 15.965 0.235 ;
        RECT 16.155 0.065 16.325 0.235 ;
        RECT 16.605 0.065 16.775 0.235 ;
        RECT 16.965 0.065 17.135 0.235 ;
        RECT 17.325 0.065 17.495 0.235 ;
        RECT 17.685 0.065 17.855 0.235 ;
        RECT 18.405 0.065 18.575 0.235 ;
        RECT 18.765 0.065 18.935 0.235 ;
        RECT 19.125 0.065 19.295 0.235 ;
        RECT 19.485 0.065 19.655 0.235 ;
        RECT 19.935 0.065 20.105 0.235 ;
        RECT 20.295 0.065 20.465 0.235 ;
        RECT 20.655 0.065 20.825 0.235 ;
        RECT 21.015 0.065 21.185 0.235 ;
        RECT 21.735 0.065 21.905 0.235 ;
        RECT 22.095 0.065 22.265 0.235 ;
        RECT 22.455 0.065 22.625 0.235 ;
        RECT 22.815 0.065 22.985 0.235 ;
        RECT 23.175 0.065 23.345 0.235 ;
        RECT 23.535 0.065 23.705 0.235 ;
        RECT 24.025 0.065 24.195 0.235 ;
        RECT 24.385 0.065 24.555 0.235 ;
        RECT 24.745 0.065 24.915 0.235 ;
        RECT 25.105 0.065 25.275 0.235 ;
        RECT 25.465 0.065 25.635 0.235 ;
        RECT 25.825 0.065 25.995 0.235 ;
        RECT 26.545 0.065 26.715 0.235 ;
        RECT 26.905 0.065 27.075 0.235 ;
        RECT 27.265 0.065 27.435 0.235 ;
        RECT 27.625 0.065 27.795 0.235 ;
        RECT 28.075 0.065 28.245 0.235 ;
        RECT 28.435 0.065 28.605 0.235 ;
        RECT 28.795 0.065 28.965 0.235 ;
        RECT 29.155 0.065 29.325 0.235 ;
        RECT 29.875 0.065 30.045 0.235 ;
        RECT 30.235 0.065 30.405 0.235 ;
        RECT 30.595 0.065 30.765 0.235 ;
        RECT 30.955 0.065 31.125 0.235 ;
        RECT 31.405 0.065 31.575 0.235 ;
        RECT 31.765 0.065 31.935 0.235 ;
        RECT 32.125 0.065 32.295 0.235 ;
        RECT 32.485 0.065 32.655 0.235 ;
        RECT 33.205 0.065 33.375 0.235 ;
        RECT 33.565 0.065 33.735 0.235 ;
        RECT 33.925 0.065 34.095 0.235 ;
        RECT 34.285 0.065 34.455 0.235 ;
        RECT 34.735 0.065 34.905 0.235 ;
        RECT 35.095 0.065 35.265 0.235 ;
        RECT 35.455 0.065 35.625 0.235 ;
        RECT 35.815 0.065 35.985 0.235 ;
        RECT 36.535 0.065 36.705 0.235 ;
        RECT 36.895 0.065 37.065 0.235 ;
        RECT 37.255 0.065 37.425 0.235 ;
        RECT 37.615 0.065 37.785 0.235 ;
        RECT 38.065 0.065 38.235 0.235 ;
        RECT 38.425 0.065 38.595 0.235 ;
        RECT 38.785 0.065 38.955 0.235 ;
        RECT 39.145 0.065 39.315 0.235 ;
        RECT 39.865 0.065 40.035 0.235 ;
        RECT 40.225 0.065 40.395 0.235 ;
        RECT 40.585 0.065 40.755 0.235 ;
        RECT 40.945 0.065 41.115 0.235 ;
        RECT 41.395 0.065 41.565 0.235 ;
        RECT 41.755 0.065 41.925 0.235 ;
        RECT 42.115 0.065 42.285 0.235 ;
        RECT 42.475 0.065 42.645 0.235 ;
        RECT 43.195 0.065 43.365 0.235 ;
        RECT 43.555 0.065 43.725 0.235 ;
        RECT 43.915 0.065 44.085 0.235 ;
        RECT 44.275 0.065 44.445 0.235 ;
        RECT 44.635 0.065 44.805 0.235 ;
        RECT 44.995 0.065 45.165 0.235 ;
        RECT 45.485 0.065 45.655 0.235 ;
        RECT 45.845 0.065 46.015 0.235 ;
        RECT 46.205 0.065 46.375 0.235 ;
        RECT 46.565 0.065 46.735 0.235 ;
        RECT 46.925 0.065 47.095 0.235 ;
        RECT 47.285 0.065 47.455 0.235 ;
        RECT 48.005 0.065 48.175 0.235 ;
        RECT 48.365 0.065 48.535 0.235 ;
        RECT 48.725 0.065 48.895 0.235 ;
        RECT 49.085 0.065 49.255 0.235 ;
        RECT 49.535 0.065 49.705 0.235 ;
        RECT 49.895 0.065 50.065 0.235 ;
        RECT 50.255 0.065 50.425 0.235 ;
        RECT 50.615 0.065 50.785 0.235 ;
        RECT 51.335 0.065 51.505 0.235 ;
        RECT 51.695 0.065 51.865 0.235 ;
        RECT 52.055 0.065 52.225 0.235 ;
        RECT 52.415 0.065 52.585 0.235 ;
        RECT 52.865 0.065 53.035 0.235 ;
        RECT 53.225 0.065 53.395 0.235 ;
        RECT 53.585 0.065 53.755 0.235 ;
        RECT 53.945 0.065 54.115 0.235 ;
        RECT 54.665 0.065 54.835 0.235 ;
        RECT 55.025 0.065 55.195 0.235 ;
        RECT 55.385 0.065 55.555 0.235 ;
        RECT 55.745 0.065 55.915 0.235 ;
        RECT 56.195 0.065 56.365 0.235 ;
        RECT 56.555 0.065 56.725 0.235 ;
        RECT 56.915 0.065 57.085 0.235 ;
        RECT 57.275 0.065 57.445 0.235 ;
        RECT 57.995 0.065 58.165 0.235 ;
        RECT 58.355 0.065 58.525 0.235 ;
        RECT 58.715 0.065 58.885 0.235 ;
        RECT 59.075 0.065 59.245 0.235 ;
        RECT 59.525 0.065 59.695 0.235 ;
        RECT 59.885 0.065 60.055 0.235 ;
        RECT 60.245 0.065 60.415 0.235 ;
        RECT 60.605 0.065 60.775 0.235 ;
        RECT 61.325 0.065 61.495 0.235 ;
        RECT 61.685 0.065 61.855 0.235 ;
        RECT 62.045 0.065 62.215 0.235 ;
        RECT 62.405 0.065 62.575 0.235 ;
        RECT 62.855 0.065 63.025 0.235 ;
        RECT 63.215 0.065 63.385 0.235 ;
        RECT 63.575 0.065 63.745 0.235 ;
        RECT 63.935 0.065 64.105 0.235 ;
        RECT 64.655 0.065 64.825 0.235 ;
        RECT 65.015 0.065 65.185 0.235 ;
        RECT 65.375 0.065 65.545 0.235 ;
        RECT 65.735 0.065 65.905 0.235 ;
        RECT 66.185 0.065 66.355 0.235 ;
        RECT 66.545 0.065 66.715 0.235 ;
        RECT 66.905 0.065 67.075 0.235 ;
        RECT 67.265 0.065 67.435 0.235 ;
        RECT 67.985 0.065 68.155 0.235 ;
        RECT 68.345 0.065 68.515 0.235 ;
        RECT 68.705 0.065 68.875 0.235 ;
        RECT 69.065 0.065 69.235 0.235 ;
        RECT 69.515 0.065 69.685 0.235 ;
        RECT 69.875 0.065 70.045 0.235 ;
        RECT 70.235 0.065 70.405 0.235 ;
        RECT 70.595 0.065 70.765 0.235 ;
        RECT 71.315 0.065 71.485 0.235 ;
        RECT 71.675 0.065 71.845 0.235 ;
        RECT 72.035 0.065 72.205 0.235 ;
        RECT 72.395 0.065 72.565 0.235 ;
        RECT 72.845 0.065 73.015 0.235 ;
        RECT 73.205 0.065 73.375 0.235 ;
        RECT 73.565 0.065 73.735 0.235 ;
        RECT 73.925 0.065 74.095 0.235 ;
        RECT 74.645 0.065 74.815 0.235 ;
        RECT 75.005 0.065 75.175 0.235 ;
        RECT 75.395 0.065 75.565 0.235 ;
        RECT 75.785 0.065 75.955 0.235 ;
        RECT 76.145 0.065 76.315 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 76.745 0.310 ;
    END
  END VSS
  PIN Q
    ANTENNADIFFAREA 0.771900 ;
    PORT
      LAYER li1 ;
        RECT 75.395 4.895 75.565 7.250 ;
        RECT 75.395 4.725 75.935 4.895 ;
        RECT 75.765 2.305 75.935 4.725 ;
        RECT 75.395 2.135 75.935 2.305 ;
        RECT 75.395 0.975 75.565 2.135 ;
      LAYER mcon ;
        RECT 75.765 3.985 75.935 4.155 ;
      LAYER met1 ;
        RECT 75.735 4.155 75.965 4.185 ;
        RECT 75.705 3.985 76.115 4.155 ;
        RECT 75.735 3.955 75.965 3.985 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 1.445 5.470 1.615 7.250 ;
        RECT 2.325 5.470 2.495 7.250 ;
        RECT 3.205 5.470 3.375 7.250 ;
        RECT 5.955 5.515 6.125 7.250 ;
        RECT 6.835 5.515 7.005 7.250 ;
        RECT 9.285 5.515 9.455 7.250 ;
        RECT 10.165 5.515 10.335 7.250 ;
        RECT 12.615 5.515 12.785 7.250 ;
        RECT 13.495 5.515 13.665 7.250 ;
        RECT 15.945 5.515 16.115 7.250 ;
        RECT 16.825 5.515 16.995 7.250 ;
        RECT 19.275 5.515 19.445 7.250 ;
        RECT 20.155 5.515 20.325 7.250 ;
        RECT 1.445 5.300 4.155 5.470 ;
        RECT 5.955 5.345 7.485 5.515 ;
        RECT 9.285 5.345 10.815 5.515 ;
        RECT 12.615 5.345 14.145 5.515 ;
        RECT 15.945 5.345 17.475 5.515 ;
        RECT 19.275 5.345 20.805 5.515 ;
        RECT 1.025 2.055 1.195 5.095 ;
        RECT 3.245 2.055 3.415 5.095 ;
        RECT 0.505 1.815 0.675 1.895 ;
        RECT 1.475 1.815 1.645 1.895 ;
        RECT 2.445 1.815 2.615 1.895 ;
        RECT 0.505 1.645 2.615 1.815 ;
        RECT 0.505 0.515 0.675 1.645 ;
        RECT 1.475 0.765 1.645 1.645 ;
        RECT 2.445 1.565 2.615 1.645 ;
        RECT 1.965 1.220 2.135 1.300 ;
        RECT 3.015 1.220 3.185 1.895 ;
        RECT 3.985 1.890 4.155 5.300 ;
        RECT 5.835 2.055 6.005 5.095 ;
        RECT 1.965 1.050 3.185 1.220 ;
        RECT 1.965 0.970 2.135 1.050 ;
        RECT 2.445 0.765 2.615 0.845 ;
        RECT 1.475 0.595 2.615 0.765 ;
        RECT 1.475 0.515 1.645 0.595 ;
        RECT 2.445 0.515 2.615 0.595 ;
        RECT 3.015 0.765 3.185 1.050 ;
        RECT 3.500 1.720 4.155 1.890 ;
        RECT 5.420 1.805 5.590 1.885 ;
        RECT 6.390 1.805 6.560 1.885 ;
        RECT 7.315 1.880 7.485 5.345 ;
        RECT 9.165 2.055 9.335 5.095 ;
        RECT 9.935 4.940 10.105 5.095 ;
        RECT 9.905 4.765 10.105 4.940 ;
        RECT 9.905 2.055 10.075 4.765 ;
        RECT 3.500 0.985 3.670 1.720 ;
        RECT 5.420 1.635 6.560 1.805 ;
        RECT 3.985 0.765 4.155 1.535 ;
        RECT 3.015 0.595 4.155 0.765 ;
        RECT 3.015 0.515 3.185 0.595 ;
        RECT 3.985 0.515 4.155 0.595 ;
        RECT 5.420 0.505 5.590 1.635 ;
        RECT 6.390 0.755 6.560 1.635 ;
        RECT 6.875 1.710 7.485 1.880 ;
        RECT 8.750 1.805 8.920 1.885 ;
        RECT 9.720 1.805 9.890 1.885 ;
        RECT 10.645 1.880 10.815 5.345 ;
        RECT 12.495 2.055 12.665 5.095 ;
        RECT 6.875 0.975 7.045 1.710 ;
        RECT 8.750 1.635 9.890 1.805 ;
        RECT 7.360 0.755 7.530 1.525 ;
        RECT 6.390 0.585 7.530 0.755 ;
        RECT 6.390 0.505 6.560 0.585 ;
        RECT 7.360 0.505 7.530 0.585 ;
        RECT 8.750 0.505 8.920 1.635 ;
        RECT 9.720 0.755 9.890 1.635 ;
        RECT 10.205 1.710 10.815 1.880 ;
        RECT 12.080 1.805 12.250 1.885 ;
        RECT 13.050 1.805 13.220 1.885 ;
        RECT 13.975 1.880 14.145 5.345 ;
        RECT 15.825 2.055 15.995 5.095 ;
        RECT 16.595 4.940 16.765 5.095 ;
        RECT 16.565 4.765 16.765 4.940 ;
        RECT 16.565 2.055 16.735 4.765 ;
        RECT 10.205 0.975 10.375 1.710 ;
        RECT 12.080 1.635 13.220 1.805 ;
        RECT 10.690 0.755 10.860 1.525 ;
        RECT 9.720 0.585 10.860 0.755 ;
        RECT 9.720 0.505 9.890 0.585 ;
        RECT 10.690 0.505 10.860 0.585 ;
        RECT 12.080 0.505 12.250 1.635 ;
        RECT 13.050 0.755 13.220 1.635 ;
        RECT 13.535 1.710 14.145 1.880 ;
        RECT 15.410 1.805 15.580 1.885 ;
        RECT 16.380 1.805 16.550 1.885 ;
        RECT 17.305 1.880 17.475 5.345 ;
        RECT 19.155 2.055 19.325 5.095 ;
        RECT 19.925 4.940 20.095 5.095 ;
        RECT 19.895 4.765 20.095 4.940 ;
        RECT 19.895 2.055 20.065 4.765 ;
        RECT 13.535 0.975 13.705 1.710 ;
        RECT 15.410 1.635 16.550 1.805 ;
        RECT 14.020 0.755 14.190 1.525 ;
        RECT 13.050 0.585 14.190 0.755 ;
        RECT 13.050 0.505 13.220 0.585 ;
        RECT 14.020 0.505 14.190 0.585 ;
        RECT 15.410 0.505 15.580 1.635 ;
        RECT 16.380 0.755 16.550 1.635 ;
        RECT 16.865 1.710 17.475 1.880 ;
        RECT 18.740 1.805 18.910 1.885 ;
        RECT 19.710 1.805 19.880 1.885 ;
        RECT 20.635 1.880 20.805 5.345 ;
        RECT 22.905 5.470 23.075 7.250 ;
        RECT 23.785 5.470 23.955 7.250 ;
        RECT 24.665 5.470 24.835 7.250 ;
        RECT 27.415 5.515 27.585 7.250 ;
        RECT 28.295 5.515 28.465 7.250 ;
        RECT 30.745 5.515 30.915 7.250 ;
        RECT 31.625 5.515 31.795 7.250 ;
        RECT 34.075 5.515 34.245 7.250 ;
        RECT 34.955 5.515 35.125 7.250 ;
        RECT 37.405 5.515 37.575 7.250 ;
        RECT 38.285 5.515 38.455 7.250 ;
        RECT 40.735 5.515 40.905 7.250 ;
        RECT 41.615 5.515 41.785 7.250 ;
        RECT 22.905 5.300 25.615 5.470 ;
        RECT 27.415 5.345 28.945 5.515 ;
        RECT 30.745 5.345 32.275 5.515 ;
        RECT 34.075 5.345 35.605 5.515 ;
        RECT 37.405 5.345 38.935 5.515 ;
        RECT 40.735 5.345 42.265 5.515 ;
        RECT 22.485 2.055 22.655 5.095 ;
        RECT 24.705 2.055 24.875 5.095 ;
        RECT 16.865 0.975 17.035 1.710 ;
        RECT 18.740 1.635 19.880 1.805 ;
        RECT 17.350 0.755 17.520 1.525 ;
        RECT 16.380 0.585 17.520 0.755 ;
        RECT 16.380 0.505 16.550 0.585 ;
        RECT 17.350 0.505 17.520 0.585 ;
        RECT 18.740 0.505 18.910 1.635 ;
        RECT 19.710 0.755 19.880 1.635 ;
        RECT 20.195 1.710 20.805 1.880 ;
        RECT 21.965 1.815 22.135 1.895 ;
        RECT 22.935 1.815 23.105 1.895 ;
        RECT 23.905 1.815 24.075 1.895 ;
        RECT 20.195 0.975 20.365 1.710 ;
        RECT 21.965 1.645 24.075 1.815 ;
        RECT 20.680 0.755 20.850 1.525 ;
        RECT 19.710 0.585 20.850 0.755 ;
        RECT 19.710 0.505 19.880 0.585 ;
        RECT 20.680 0.505 20.850 0.585 ;
        RECT 21.965 0.515 22.135 1.645 ;
        RECT 22.935 0.765 23.105 1.645 ;
        RECT 23.905 1.565 24.075 1.645 ;
        RECT 23.425 1.220 23.595 1.300 ;
        RECT 24.475 1.220 24.645 1.895 ;
        RECT 25.445 1.890 25.615 5.300 ;
        RECT 27.295 2.055 27.465 5.095 ;
        RECT 23.425 1.050 24.645 1.220 ;
        RECT 23.425 0.970 23.595 1.050 ;
        RECT 23.905 0.765 24.075 0.845 ;
        RECT 22.935 0.595 24.075 0.765 ;
        RECT 22.935 0.515 23.105 0.595 ;
        RECT 23.905 0.515 24.075 0.595 ;
        RECT 24.475 0.765 24.645 1.050 ;
        RECT 24.960 1.720 25.615 1.890 ;
        RECT 26.880 1.805 27.050 1.885 ;
        RECT 27.850 1.805 28.020 1.885 ;
        RECT 28.775 1.880 28.945 5.345 ;
        RECT 30.625 2.055 30.795 5.095 ;
        RECT 31.395 4.940 31.565 5.095 ;
        RECT 31.365 4.765 31.565 4.940 ;
        RECT 31.365 2.055 31.535 4.765 ;
        RECT 24.960 0.985 25.130 1.720 ;
        RECT 26.880 1.635 28.020 1.805 ;
        RECT 25.445 0.765 25.615 1.535 ;
        RECT 24.475 0.595 25.615 0.765 ;
        RECT 24.475 0.515 24.645 0.595 ;
        RECT 25.445 0.515 25.615 0.595 ;
        RECT 26.880 0.505 27.050 1.635 ;
        RECT 27.850 0.755 28.020 1.635 ;
        RECT 28.335 1.710 28.945 1.880 ;
        RECT 30.210 1.805 30.380 1.885 ;
        RECT 31.180 1.805 31.350 1.885 ;
        RECT 32.105 1.880 32.275 5.345 ;
        RECT 33.955 2.055 34.125 5.095 ;
        RECT 28.335 0.975 28.505 1.710 ;
        RECT 30.210 1.635 31.350 1.805 ;
        RECT 28.820 0.755 28.990 1.525 ;
        RECT 27.850 0.585 28.990 0.755 ;
        RECT 27.850 0.505 28.020 0.585 ;
        RECT 28.820 0.505 28.990 0.585 ;
        RECT 30.210 0.505 30.380 1.635 ;
        RECT 31.180 0.755 31.350 1.635 ;
        RECT 31.665 1.710 32.275 1.880 ;
        RECT 33.540 1.805 33.710 1.885 ;
        RECT 34.510 1.805 34.680 1.885 ;
        RECT 35.435 1.880 35.605 5.345 ;
        RECT 37.285 2.055 37.455 5.095 ;
        RECT 38.055 4.940 38.225 5.095 ;
        RECT 38.025 4.765 38.225 4.940 ;
        RECT 38.025 2.055 38.195 4.765 ;
        RECT 31.665 0.975 31.835 1.710 ;
        RECT 33.540 1.635 34.680 1.805 ;
        RECT 32.150 0.755 32.320 1.525 ;
        RECT 31.180 0.585 32.320 0.755 ;
        RECT 31.180 0.505 31.350 0.585 ;
        RECT 32.150 0.505 32.320 0.585 ;
        RECT 33.540 0.505 33.710 1.635 ;
        RECT 34.510 0.755 34.680 1.635 ;
        RECT 34.995 1.710 35.605 1.880 ;
        RECT 36.870 1.805 37.040 1.885 ;
        RECT 37.840 1.805 38.010 1.885 ;
        RECT 38.765 1.880 38.935 5.345 ;
        RECT 40.615 2.055 40.785 5.095 ;
        RECT 41.385 4.940 41.555 5.095 ;
        RECT 41.355 4.765 41.555 4.940 ;
        RECT 41.355 2.055 41.525 4.765 ;
        RECT 34.995 0.975 35.165 1.710 ;
        RECT 36.870 1.635 38.010 1.805 ;
        RECT 35.480 0.755 35.650 1.525 ;
        RECT 34.510 0.585 35.650 0.755 ;
        RECT 34.510 0.505 34.680 0.585 ;
        RECT 35.480 0.505 35.650 0.585 ;
        RECT 36.870 0.505 37.040 1.635 ;
        RECT 37.840 0.755 38.010 1.635 ;
        RECT 38.325 1.710 38.935 1.880 ;
        RECT 40.200 1.805 40.370 1.885 ;
        RECT 41.170 1.805 41.340 1.885 ;
        RECT 42.095 1.880 42.265 5.345 ;
        RECT 44.365 5.470 44.535 7.250 ;
        RECT 45.245 5.470 45.415 7.250 ;
        RECT 46.125 5.470 46.295 7.250 ;
        RECT 48.875 5.515 49.045 7.250 ;
        RECT 49.755 5.515 49.925 7.250 ;
        RECT 52.205 5.515 52.375 7.250 ;
        RECT 53.085 5.515 53.255 7.250 ;
        RECT 55.535 5.515 55.705 7.250 ;
        RECT 56.415 5.515 56.585 7.250 ;
        RECT 58.865 5.515 59.035 7.250 ;
        RECT 59.745 5.515 59.915 7.250 ;
        RECT 62.195 5.515 62.365 7.250 ;
        RECT 63.075 5.515 63.245 7.250 ;
        RECT 65.525 7.055 65.705 7.225 ;
        RECT 65.525 5.525 65.695 7.055 ;
        RECT 66.405 5.525 66.575 7.225 ;
        RECT 44.365 5.300 47.075 5.470 ;
        RECT 48.875 5.345 50.405 5.515 ;
        RECT 52.205 5.345 53.735 5.515 ;
        RECT 55.535 5.345 57.065 5.515 ;
        RECT 58.865 5.345 60.395 5.515 ;
        RECT 62.195 5.345 63.725 5.515 ;
        RECT 65.525 5.355 66.575 5.525 ;
        RECT 43.945 2.055 44.115 5.095 ;
        RECT 46.165 2.055 46.335 5.095 ;
        RECT 38.325 0.975 38.495 1.710 ;
        RECT 40.200 1.635 41.340 1.805 ;
        RECT 38.810 0.755 38.980 1.525 ;
        RECT 37.840 0.585 38.980 0.755 ;
        RECT 37.840 0.505 38.010 0.585 ;
        RECT 38.810 0.505 38.980 0.585 ;
        RECT 40.200 0.505 40.370 1.635 ;
        RECT 41.170 0.755 41.340 1.635 ;
        RECT 41.655 1.710 42.265 1.880 ;
        RECT 43.425 1.815 43.595 1.895 ;
        RECT 44.395 1.815 44.565 1.895 ;
        RECT 45.365 1.815 45.535 1.895 ;
        RECT 41.655 0.975 41.825 1.710 ;
        RECT 43.425 1.645 45.535 1.815 ;
        RECT 42.140 0.755 42.310 1.525 ;
        RECT 41.170 0.585 42.310 0.755 ;
        RECT 41.170 0.505 41.340 0.585 ;
        RECT 42.140 0.505 42.310 0.585 ;
        RECT 43.425 0.515 43.595 1.645 ;
        RECT 44.395 0.765 44.565 1.645 ;
        RECT 45.365 1.565 45.535 1.645 ;
        RECT 44.885 1.220 45.055 1.300 ;
        RECT 45.935 1.220 46.105 1.895 ;
        RECT 46.905 1.890 47.075 5.300 ;
        RECT 48.755 2.055 48.925 5.095 ;
        RECT 44.885 1.050 46.105 1.220 ;
        RECT 44.885 0.970 45.055 1.050 ;
        RECT 45.365 0.765 45.535 0.845 ;
        RECT 44.395 0.595 45.535 0.765 ;
        RECT 44.395 0.515 44.565 0.595 ;
        RECT 45.365 0.515 45.535 0.595 ;
        RECT 45.935 0.765 46.105 1.050 ;
        RECT 46.420 1.720 47.075 1.890 ;
        RECT 48.340 1.805 48.510 1.885 ;
        RECT 49.310 1.805 49.480 1.885 ;
        RECT 50.235 1.880 50.405 5.345 ;
        RECT 52.085 2.055 52.255 5.095 ;
        RECT 52.855 4.940 53.025 5.095 ;
        RECT 52.825 4.765 53.025 4.940 ;
        RECT 52.825 2.055 52.995 4.765 ;
        RECT 46.420 0.985 46.590 1.720 ;
        RECT 48.340 1.635 49.480 1.805 ;
        RECT 46.905 0.765 47.075 1.535 ;
        RECT 45.935 0.595 47.075 0.765 ;
        RECT 45.935 0.515 46.105 0.595 ;
        RECT 46.905 0.515 47.075 0.595 ;
        RECT 48.340 0.505 48.510 1.635 ;
        RECT 49.310 0.755 49.480 1.635 ;
        RECT 49.795 1.710 50.405 1.880 ;
        RECT 51.670 1.805 51.840 1.885 ;
        RECT 52.640 1.805 52.810 1.885 ;
        RECT 53.565 1.880 53.735 5.345 ;
        RECT 55.415 2.055 55.585 5.095 ;
        RECT 49.795 0.975 49.965 1.710 ;
        RECT 51.670 1.635 52.810 1.805 ;
        RECT 50.280 0.755 50.450 1.525 ;
        RECT 49.310 0.585 50.450 0.755 ;
        RECT 49.310 0.505 49.480 0.585 ;
        RECT 50.280 0.505 50.450 0.585 ;
        RECT 51.670 0.505 51.840 1.635 ;
        RECT 52.640 0.755 52.810 1.635 ;
        RECT 53.125 1.710 53.735 1.880 ;
        RECT 55.000 1.805 55.170 1.885 ;
        RECT 55.970 1.805 56.140 1.885 ;
        RECT 56.895 1.880 57.065 5.345 ;
        RECT 58.745 2.055 58.915 5.095 ;
        RECT 59.515 4.940 59.685 5.095 ;
        RECT 59.485 4.765 59.685 4.940 ;
        RECT 59.485 2.055 59.655 4.765 ;
        RECT 53.125 0.975 53.295 1.710 ;
        RECT 55.000 1.635 56.140 1.805 ;
        RECT 53.610 0.755 53.780 1.525 ;
        RECT 52.640 0.585 53.780 0.755 ;
        RECT 52.640 0.505 52.810 0.585 ;
        RECT 53.610 0.505 53.780 0.585 ;
        RECT 55.000 0.505 55.170 1.635 ;
        RECT 55.970 0.755 56.140 1.635 ;
        RECT 56.455 1.710 57.065 1.880 ;
        RECT 58.330 1.805 58.500 1.885 ;
        RECT 59.300 1.805 59.470 1.885 ;
        RECT 60.225 1.880 60.395 5.345 ;
        RECT 62.075 2.055 62.245 5.095 ;
        RECT 62.845 4.940 63.015 5.095 ;
        RECT 62.815 4.765 63.015 4.940 ;
        RECT 62.815 2.055 62.985 4.765 ;
        RECT 56.455 0.975 56.625 1.710 ;
        RECT 58.330 1.635 59.470 1.805 ;
        RECT 56.940 0.755 57.110 1.525 ;
        RECT 55.970 0.585 57.110 0.755 ;
        RECT 55.970 0.505 56.140 0.585 ;
        RECT 56.940 0.505 57.110 0.585 ;
        RECT 58.330 0.505 58.500 1.635 ;
        RECT 59.300 0.755 59.470 1.635 ;
        RECT 59.785 1.710 60.395 1.880 ;
        RECT 61.660 1.805 61.830 1.885 ;
        RECT 62.630 1.805 62.800 1.885 ;
        RECT 63.555 1.880 63.725 5.345 ;
        RECT 66.405 5.275 66.575 5.355 ;
        RECT 68.405 7.055 70.335 7.225 ;
        RECT 68.405 5.275 68.575 7.055 ;
        RECT 68.845 5.525 69.015 6.795 ;
        RECT 69.285 5.785 69.455 7.055 ;
        RECT 69.725 5.525 69.895 6.795 ;
        RECT 70.165 5.605 70.335 7.055 ;
        RECT 71.745 7.055 73.675 7.225 ;
        RECT 68.845 5.355 69.895 5.525 ;
        RECT 69.725 5.275 69.895 5.355 ;
        RECT 71.745 5.275 71.915 7.055 ;
        RECT 72.185 5.525 72.355 6.795 ;
        RECT 72.625 5.785 72.795 7.055 ;
        RECT 73.065 5.525 73.235 6.795 ;
        RECT 73.505 5.785 73.675 7.055 ;
        RECT 72.185 5.355 73.715 5.525 ;
        RECT 65.035 2.055 65.205 5.100 ;
        RECT 66.185 4.940 66.355 5.100 ;
        RECT 66.145 4.770 66.355 4.940 ;
        RECT 66.145 2.055 66.315 4.770 ;
        RECT 68.735 2.055 68.905 5.100 ;
        RECT 70.215 2.055 70.385 5.100 ;
        RECT 71.695 2.055 71.865 5.100 ;
        RECT 72.805 4.770 72.995 5.100 ;
        RECT 72.805 2.055 72.975 4.770 ;
        RECT 59.785 0.975 59.955 1.710 ;
        RECT 61.660 1.635 62.800 1.805 ;
        RECT 60.270 0.755 60.440 1.525 ;
        RECT 59.300 0.585 60.440 0.755 ;
        RECT 59.300 0.505 59.470 0.585 ;
        RECT 60.270 0.505 60.440 0.585 ;
        RECT 61.660 0.505 61.830 1.635 ;
        RECT 62.630 0.755 62.800 1.635 ;
        RECT 63.115 1.710 63.725 1.880 ;
        RECT 64.990 1.805 65.160 1.885 ;
        RECT 65.960 1.805 66.130 1.885 ;
        RECT 63.115 0.975 63.285 1.710 ;
        RECT 64.990 1.635 66.130 1.805 ;
        RECT 63.600 0.755 63.770 1.525 ;
        RECT 62.630 0.585 63.770 0.755 ;
        RECT 62.630 0.505 62.800 0.585 ;
        RECT 63.600 0.505 63.770 0.585 ;
        RECT 64.990 0.505 65.160 1.635 ;
        RECT 65.960 0.755 66.130 1.635 ;
        RECT 66.445 1.310 66.615 1.485 ;
        RECT 66.440 1.155 66.615 1.310 ;
        RECT 66.440 0.975 66.610 1.155 ;
        RECT 66.930 0.755 67.100 1.885 ;
        RECT 65.960 0.585 67.100 0.755 ;
        RECT 65.960 0.505 66.130 0.585 ;
        RECT 66.930 0.505 67.100 0.585 ;
        RECT 68.320 1.805 68.490 1.885 ;
        RECT 69.290 1.805 69.460 1.885 ;
        RECT 68.320 1.635 69.460 1.805 ;
        RECT 68.320 0.505 68.490 1.635 ;
        RECT 69.290 0.755 69.460 1.635 ;
        RECT 69.775 0.975 69.945 1.485 ;
        RECT 70.260 0.755 70.430 1.885 ;
        RECT 69.290 0.585 70.430 0.755 ;
        RECT 69.290 0.505 69.460 0.585 ;
        RECT 70.260 0.505 70.430 0.585 ;
        RECT 71.650 1.805 71.820 1.885 ;
        RECT 72.620 1.805 72.790 1.885 ;
        RECT 73.545 1.870 73.715 5.355 ;
        RECT 75.025 2.055 75.195 5.095 ;
        RECT 71.650 1.635 72.790 1.805 ;
        RECT 71.650 0.505 71.820 1.635 ;
        RECT 72.620 0.755 72.790 1.635 ;
        RECT 73.105 1.700 73.715 1.870 ;
        RECT 73.105 0.975 73.275 1.700 ;
        RECT 73.590 0.755 73.760 1.530 ;
        RECT 72.620 0.585 73.760 0.755 ;
        RECT 72.620 0.505 72.790 0.585 ;
        RECT 73.590 0.505 73.760 0.585 ;
      LAYER mcon ;
        RECT 1.025 4.355 1.195 4.525 ;
        RECT 3.245 3.615 3.415 3.785 ;
        RECT 3.985 3.985 4.155 4.155 ;
        RECT 5.835 3.985 6.005 4.155 ;
        RECT 7.315 3.615 7.485 3.785 ;
        RECT 9.165 3.615 9.335 3.785 ;
        RECT 9.905 4.355 10.075 4.525 ;
        RECT 10.645 3.615 10.815 3.785 ;
        RECT 12.495 3.615 12.665 3.785 ;
        RECT 13.975 4.355 14.145 4.525 ;
        RECT 15.825 3.985 15.995 4.155 ;
        RECT 16.565 3.245 16.735 3.415 ;
        RECT 17.305 3.985 17.475 4.155 ;
        RECT 19.155 3.985 19.325 4.155 ;
        RECT 19.895 4.355 20.065 4.525 ;
        RECT 20.635 3.245 20.805 3.415 ;
        RECT 22.485 4.355 22.655 4.525 ;
        RECT 24.705 3.615 24.875 3.785 ;
        RECT 25.445 3.985 25.615 4.155 ;
        RECT 27.295 3.985 27.465 4.155 ;
        RECT 28.775 3.615 28.945 3.785 ;
        RECT 30.625 3.615 30.795 3.785 ;
        RECT 31.365 4.355 31.535 4.525 ;
        RECT 32.105 3.615 32.275 3.785 ;
        RECT 33.955 3.615 34.125 3.785 ;
        RECT 35.435 4.355 35.605 4.525 ;
        RECT 37.285 3.985 37.455 4.155 ;
        RECT 38.025 2.505 38.195 2.675 ;
        RECT 38.765 3.985 38.935 4.155 ;
        RECT 40.615 3.985 40.785 4.155 ;
        RECT 41.355 4.355 41.525 4.525 ;
        RECT 66.405 5.355 66.575 5.525 ;
        RECT 42.095 2.505 42.265 2.675 ;
        RECT 43.945 4.355 44.115 4.525 ;
        RECT 46.165 3.615 46.335 3.785 ;
        RECT 46.905 3.985 47.075 4.155 ;
        RECT 48.755 3.985 48.925 4.155 ;
        RECT 50.235 3.615 50.405 3.785 ;
        RECT 52.085 3.615 52.255 3.785 ;
        RECT 52.825 4.355 52.995 4.525 ;
        RECT 53.565 3.615 53.735 3.785 ;
        RECT 55.415 3.615 55.585 3.785 ;
        RECT 56.895 4.355 57.065 4.525 ;
        RECT 58.745 3.985 58.915 4.155 ;
        RECT 59.485 3.985 59.655 4.155 ;
        RECT 60.225 4.725 60.395 4.895 ;
        RECT 62.075 4.725 62.245 4.895 ;
        RECT 62.815 4.355 62.985 4.525 ;
        RECT 68.405 5.355 68.575 5.525 ;
        RECT 69.725 5.355 69.895 5.525 ;
        RECT 71.745 5.355 71.915 5.525 ;
        RECT 63.555 3.985 63.725 4.155 ;
        RECT 65.035 4.725 65.205 4.895 ;
        RECT 65.035 3.985 65.205 4.155 ;
        RECT 66.145 4.355 66.315 4.525 ;
        RECT 66.145 2.505 66.315 2.675 ;
        RECT 68.735 4.725 68.905 4.895 ;
        RECT 70.215 3.245 70.385 3.415 ;
        RECT 70.215 2.135 70.385 2.305 ;
        RECT 71.695 2.135 71.865 2.305 ;
        RECT 72.805 4.355 72.975 4.525 ;
        RECT 73.545 3.985 73.715 4.155 ;
        RECT 66.445 1.235 66.615 1.405 ;
        RECT 69.775 1.235 69.945 1.405 ;
        RECT 75.025 3.985 75.195 4.155 ;
        RECT 73.105 1.235 73.275 1.405 ;
      LAYER met1 ;
        RECT 66.375 5.525 66.605 5.555 ;
        RECT 68.375 5.525 68.605 5.555 ;
        RECT 69.695 5.525 69.925 5.555 ;
        RECT 71.715 5.525 71.945 5.555 ;
        RECT 66.345 5.355 68.635 5.525 ;
        RECT 69.665 5.355 71.975 5.525 ;
        RECT 66.375 5.325 66.605 5.355 ;
        RECT 68.375 5.325 68.605 5.355 ;
        RECT 69.695 5.325 69.925 5.355 ;
        RECT 71.715 5.325 71.945 5.355 ;
        RECT 60.195 4.895 60.425 4.925 ;
        RECT 62.045 4.895 62.275 4.925 ;
        RECT 65.005 4.895 65.235 4.925 ;
        RECT 68.705 4.895 68.935 4.925 ;
        RECT 60.165 4.725 62.305 4.895 ;
        RECT 64.975 4.725 68.965 4.895 ;
        RECT 60.195 4.695 60.425 4.725 ;
        RECT 62.045 4.695 62.275 4.725 ;
        RECT 65.005 4.695 65.235 4.725 ;
        RECT 68.705 4.695 68.935 4.725 ;
        RECT 0.995 4.525 1.225 4.555 ;
        RECT 9.875 4.525 10.105 4.555 ;
        RECT 13.945 4.525 14.175 4.555 ;
        RECT 19.865 4.525 20.095 4.555 ;
        RECT 22.455 4.525 22.685 4.555 ;
        RECT 31.335 4.525 31.565 4.555 ;
        RECT 35.405 4.525 35.635 4.555 ;
        RECT 41.325 4.525 41.555 4.555 ;
        RECT 43.915 4.525 44.145 4.555 ;
        RECT 52.795 4.525 53.025 4.555 ;
        RECT 56.865 4.525 57.095 4.555 ;
        RECT 62.785 4.525 63.015 4.555 ;
        RECT 66.115 4.525 66.345 4.555 ;
        RECT 72.775 4.525 73.005 4.555 ;
        RECT 0.965 4.355 20.125 4.525 ;
        RECT 22.425 4.355 41.585 4.525 ;
        RECT 43.885 4.355 63.045 4.525 ;
        RECT 66.085 4.355 73.035 4.525 ;
        RECT 0.995 4.325 1.225 4.355 ;
        RECT 9.875 4.325 10.105 4.355 ;
        RECT 13.945 4.325 14.175 4.355 ;
        RECT 19.865 4.325 20.095 4.355 ;
        RECT 22.455 4.325 22.685 4.355 ;
        RECT 31.335 4.325 31.565 4.355 ;
        RECT 35.405 4.325 35.635 4.355 ;
        RECT 41.325 4.325 41.555 4.355 ;
        RECT 43.915 4.325 44.145 4.355 ;
        RECT 52.795 4.325 53.025 4.355 ;
        RECT 56.865 4.325 57.095 4.355 ;
        RECT 62.785 4.325 63.015 4.355 ;
        RECT 66.115 4.325 66.345 4.355 ;
        RECT 72.775 4.325 73.005 4.355 ;
        RECT 3.955 4.155 4.185 4.185 ;
        RECT 5.805 4.155 6.035 4.185 ;
        RECT 15.795 4.155 16.025 4.185 ;
        RECT 17.275 4.155 17.505 4.185 ;
        RECT 19.125 4.155 19.355 4.185 ;
        RECT 25.415 4.155 25.645 4.185 ;
        RECT 27.265 4.155 27.495 4.185 ;
        RECT 37.255 4.155 37.485 4.185 ;
        RECT 38.735 4.155 38.965 4.185 ;
        RECT 40.585 4.155 40.815 4.185 ;
        RECT 46.875 4.155 47.105 4.185 ;
        RECT 48.725 4.155 48.955 4.185 ;
        RECT 58.715 4.155 58.945 4.185 ;
        RECT 59.455 4.155 59.685 4.185 ;
        RECT 63.525 4.155 63.755 4.185 ;
        RECT 65.005 4.155 65.235 4.185 ;
        RECT 73.515 4.155 73.745 4.185 ;
        RECT 74.995 4.155 75.225 4.185 ;
        RECT 3.925 3.985 16.055 4.155 ;
        RECT 17.245 3.985 19.385 4.155 ;
        RECT 25.385 3.985 37.515 4.155 ;
        RECT 38.705 3.985 40.845 4.155 ;
        RECT 46.845 3.985 58.975 4.155 ;
        RECT 59.425 3.985 65.265 4.155 ;
        RECT 73.485 3.985 75.255 4.155 ;
        RECT 3.955 3.955 4.185 3.985 ;
        RECT 5.805 3.955 6.035 3.985 ;
        RECT 15.795 3.955 16.025 3.985 ;
        RECT 17.275 3.955 17.505 3.985 ;
        RECT 19.125 3.955 19.355 3.985 ;
        RECT 25.415 3.955 25.645 3.985 ;
        RECT 27.265 3.955 27.495 3.985 ;
        RECT 37.255 3.955 37.485 3.985 ;
        RECT 38.735 3.955 38.965 3.985 ;
        RECT 40.585 3.955 40.815 3.985 ;
        RECT 46.875 3.955 47.105 3.985 ;
        RECT 48.725 3.955 48.955 3.985 ;
        RECT 58.715 3.955 58.945 3.985 ;
        RECT 59.455 3.955 59.685 3.985 ;
        RECT 63.525 3.955 63.755 3.985 ;
        RECT 65.005 3.955 65.235 3.985 ;
        RECT 73.515 3.955 73.745 3.985 ;
        RECT 74.995 3.955 75.225 3.985 ;
        RECT 3.215 3.785 3.445 3.815 ;
        RECT 7.285 3.785 7.515 3.815 ;
        RECT 9.135 3.785 9.365 3.815 ;
        RECT 10.615 3.785 10.845 3.815 ;
        RECT 12.465 3.785 12.695 3.815 ;
        RECT 24.675 3.785 24.905 3.815 ;
        RECT 28.745 3.785 28.975 3.815 ;
        RECT 30.595 3.785 30.825 3.815 ;
        RECT 32.075 3.785 32.305 3.815 ;
        RECT 33.925 3.785 34.155 3.815 ;
        RECT 46.135 3.785 46.365 3.815 ;
        RECT 50.205 3.785 50.435 3.815 ;
        RECT 52.055 3.785 52.285 3.815 ;
        RECT 53.535 3.785 53.765 3.815 ;
        RECT 55.385 3.785 55.615 3.815 ;
        RECT 3.185 3.615 9.395 3.785 ;
        RECT 10.585 3.615 12.725 3.785 ;
        RECT 24.645 3.615 30.855 3.785 ;
        RECT 32.045 3.615 34.185 3.785 ;
        RECT 46.105 3.615 52.315 3.785 ;
        RECT 53.505 3.615 55.645 3.785 ;
        RECT 3.215 3.585 3.445 3.615 ;
        RECT 7.285 3.585 7.515 3.615 ;
        RECT 9.135 3.585 9.365 3.615 ;
        RECT 10.615 3.585 10.845 3.615 ;
        RECT 12.465 3.585 12.695 3.615 ;
        RECT 24.675 3.585 24.905 3.615 ;
        RECT 28.745 3.585 28.975 3.615 ;
        RECT 30.595 3.585 30.825 3.615 ;
        RECT 32.075 3.585 32.305 3.615 ;
        RECT 33.925 3.585 34.155 3.615 ;
        RECT 46.135 3.585 46.365 3.615 ;
        RECT 50.205 3.585 50.435 3.615 ;
        RECT 52.055 3.585 52.285 3.615 ;
        RECT 53.535 3.585 53.765 3.615 ;
        RECT 55.385 3.585 55.615 3.615 ;
        RECT 16.535 3.415 16.765 3.445 ;
        RECT 20.605 3.415 20.835 3.445 ;
        RECT 70.185 3.415 70.415 3.445 ;
        RECT 16.505 3.245 70.445 3.415 ;
        RECT 16.535 3.215 16.765 3.245 ;
        RECT 20.605 3.215 20.835 3.245 ;
        RECT 70.185 3.215 70.415 3.245 ;
        RECT 37.995 2.675 38.225 2.705 ;
        RECT 42.065 2.675 42.295 2.705 ;
        RECT 66.115 2.675 66.345 2.705 ;
        RECT 37.965 2.505 66.375 2.675 ;
        RECT 37.995 2.475 38.225 2.505 ;
        RECT 42.065 2.475 42.295 2.505 ;
        RECT 66.115 2.475 66.345 2.505 ;
        RECT 70.185 2.305 70.415 2.335 ;
        RECT 71.665 2.305 71.895 2.335 ;
        RECT 70.155 2.135 71.925 2.305 ;
        RECT 70.185 2.105 70.415 2.135 ;
        RECT 71.665 2.105 71.895 2.135 ;
        RECT 66.415 1.405 66.645 1.435 ;
        RECT 69.745 1.405 69.975 1.435 ;
        RECT 73.075 1.405 73.305 1.435 ;
        RECT 66.385 1.235 73.335 1.405 ;
        RECT 66.415 1.205 66.645 1.235 ;
        RECT 69.745 1.205 69.975 1.235 ;
        RECT 73.075 1.205 73.305 1.235 ;
  END
END TMRDFFQX1






MACRO TMRDFFRNQNX1
  CLASS BLOCK ;
  FOREIGN TMRDFFRNQNX1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 88.530 BY 7.950 ;
  PIN QN
    ANTENNADIFFAREA 1.734950 ;
    PORT
      LAYER li1 ;
        RECT 85.505 5.525 85.675 6.795 ;
        RECT 86.385 5.525 86.555 6.795 ;
        RECT 85.505 5.355 87.035 5.525 ;
        RECT 86.865 1.870 87.035 5.355 ;
        RECT 86.425 1.700 87.035 1.870 ;
        RECT 79.765 1.310 79.935 1.485 ;
        RECT 79.760 1.155 79.935 1.310 ;
        RECT 79.760 0.975 79.930 1.155 ;
        RECT 83.095 0.975 83.265 1.485 ;
        RECT 86.425 0.975 86.595 1.700 ;
      LAYER mcon ;
        RECT 86.865 3.985 87.035 4.155 ;
        RECT 79.765 1.235 79.935 1.405 ;
        RECT 83.095 1.235 83.265 1.405 ;
        RECT 86.425 1.235 86.595 1.405 ;
      LAYER met1 ;
        RECT 86.835 4.155 87.065 4.185 ;
        RECT 86.805 3.985 87.215 4.155 ;
        RECT 86.835 3.955 87.065 3.985 ;
        RECT 79.735 1.405 79.965 1.435 ;
        RECT 83.065 1.405 83.295 1.435 ;
        RECT 86.395 1.405 86.625 1.435 ;
        RECT 79.705 1.235 86.655 1.405 ;
        RECT 79.735 1.205 79.965 1.235 ;
        RECT 83.065 1.205 83.295 1.235 ;
        RECT 86.395 1.205 86.625 1.235 ;
    END
  END QN
  PIN D
    ANTENNAGATEAREA 3.044550 ;
    PORT
      LAYER li1 ;
        RECT 6.945 2.055 7.115 5.095 ;
        RECT 32.845 2.055 33.015 5.095 ;
        RECT 58.745 2.055 58.915 5.095 ;
      LAYER mcon ;
        RECT 6.945 2.135 7.115 2.305 ;
        RECT 32.845 2.135 33.015 2.305 ;
        RECT 58.745 2.135 58.915 2.305 ;
      LAYER met1 ;
        RECT 6.915 2.305 7.145 2.335 ;
        RECT 32.815 2.305 33.045 2.335 ;
        RECT 58.715 2.305 58.945 2.335 ;
        RECT 6.885 2.135 59.095 2.305 ;
        RECT 6.915 2.105 7.145 2.135 ;
        RECT 32.815 2.105 33.045 2.135 ;
        RECT 58.715 2.105 58.945 2.135 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 6.089100 ;
    PORT
      LAYER li1 ;
        RECT 2.135 2.055 2.305 5.095 ;
        RECT 15.085 2.055 15.255 5.095 ;
        RECT 28.035 2.055 28.205 5.095 ;
        RECT 40.985 2.055 41.155 5.095 ;
        RECT 53.935 2.055 54.105 5.095 ;
        RECT 66.885 2.055 67.055 5.095 ;
      LAYER mcon ;
        RECT 2.135 4.725 2.305 4.895 ;
        RECT 15.085 4.725 15.255 4.895 ;
        RECT 28.035 4.725 28.205 4.895 ;
        RECT 40.985 4.725 41.155 4.895 ;
        RECT 53.935 4.725 54.105 4.895 ;
        RECT 66.885 4.725 67.055 4.895 ;
      LAYER met1 ;
        RECT 2.105 4.895 2.335 4.925 ;
        RECT 15.055 4.895 15.285 4.925 ;
        RECT 28.005 4.895 28.235 4.925 ;
        RECT 40.955 4.895 41.185 4.925 ;
        RECT 53.905 4.895 54.135 4.925 ;
        RECT 66.855 4.895 67.085 4.925 ;
        RECT 2.075 4.725 67.115 4.895 ;
        RECT 2.105 4.695 2.335 4.725 ;
        RECT 15.055 4.695 15.285 4.725 ;
        RECT 28.005 4.695 28.235 4.725 ;
        RECT 40.955 4.695 41.185 4.725 ;
        RECT 53.905 4.695 54.135 4.725 ;
        RECT 66.855 4.695 67.085 4.725 ;
    END
  END CLK
  PIN RN
    ANTENNAGATEAREA 9.208050 ;
    PORT
      LAYER li1 ;
        RECT 8.055 2.055 8.225 5.095 ;
        RECT 16.195 2.055 16.365 5.095 ;
        RECT 19.895 2.055 20.065 5.095 ;
        RECT 33.955 2.055 34.125 5.095 ;
        RECT 42.095 2.055 42.265 5.095 ;
        RECT 45.795 2.055 45.965 5.095 ;
        RECT 59.855 2.055 60.025 5.095 ;
        RECT 67.995 2.055 68.165 5.095 ;
        RECT 71.695 2.055 71.865 5.095 ;
      LAYER mcon ;
        RECT 8.055 2.505 8.225 2.675 ;
        RECT 16.195 2.505 16.365 2.675 ;
        RECT 19.895 2.505 20.065 2.675 ;
        RECT 33.955 2.505 34.125 2.675 ;
        RECT 42.095 2.505 42.265 2.675 ;
        RECT 45.795 2.505 45.965 2.675 ;
        RECT 59.855 2.505 60.025 2.675 ;
        RECT 67.995 2.505 68.165 2.675 ;
        RECT 71.695 2.505 71.865 2.675 ;
      LAYER met1 ;
        RECT 8.025 2.675 8.255 2.705 ;
        RECT 16.165 2.675 16.395 2.705 ;
        RECT 19.865 2.675 20.095 2.705 ;
        RECT 33.925 2.675 34.155 2.705 ;
        RECT 42.065 2.675 42.295 2.705 ;
        RECT 45.765 2.675 45.995 2.705 ;
        RECT 59.825 2.675 60.055 2.705 ;
        RECT 67.965 2.675 68.195 2.705 ;
        RECT 71.665 2.675 71.895 2.705 ;
        RECT 7.995 2.505 71.925 2.675 ;
        RECT 8.025 2.475 8.255 2.505 ;
        RECT 16.165 2.475 16.395 2.505 ;
        RECT 19.865 2.475 20.095 2.505 ;
        RECT 33.925 2.475 34.155 2.505 ;
        RECT 42.065 2.475 42.295 2.505 ;
        RECT 45.765 2.475 45.995 2.505 ;
        RECT 59.825 2.475 60.055 2.505 ;
        RECT 67.965 2.475 68.195 2.505 ;
        RECT 71.665 2.475 71.895 2.505 ;
    END
  END RN
  PIN VDD
    ANTENNADIFFAREA 100.727501 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 88.110 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 87.845 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 1.005 5.445 1.175 7.460 ;
        RECT 1.885 5.785 2.055 7.460 ;
        RECT 2.765 5.785 2.935 7.460 ;
        RECT 3.645 5.785 3.815 7.460 ;
        RECT 4.655 4.340 4.965 7.460 ;
        RECT 5.815 5.445 5.985 7.460 ;
        RECT 6.695 5.785 6.865 7.460 ;
        RECT 7.575 5.785 7.745 7.460 ;
        RECT 8.455 5.785 8.625 7.460 ;
        RECT 9.465 4.340 9.775 7.460 ;
        RECT 10.325 5.365 10.495 7.460 ;
        RECT 11.205 5.785 11.375 7.460 ;
        RECT 12.085 5.785 12.255 7.460 ;
        RECT 12.795 4.340 13.105 7.460 ;
        RECT 13.955 5.445 14.125 7.460 ;
        RECT 14.835 5.785 15.005 7.460 ;
        RECT 15.715 5.785 15.885 7.460 ;
        RECT 16.595 5.785 16.765 7.460 ;
        RECT 17.605 4.340 17.915 7.460 ;
        RECT 18.765 5.445 18.935 7.460 ;
        RECT 19.645 5.785 19.815 7.460 ;
        RECT 20.525 5.785 20.695 7.460 ;
        RECT 21.405 5.785 21.575 7.460 ;
        RECT 22.415 4.340 22.725 7.460 ;
        RECT 23.275 5.365 23.445 7.460 ;
        RECT 24.155 5.785 24.325 7.460 ;
        RECT 25.035 5.785 25.205 7.460 ;
        RECT 25.745 4.340 26.055 7.460 ;
        RECT 26.905 5.445 27.075 7.460 ;
        RECT 27.785 5.785 27.955 7.460 ;
        RECT 28.665 5.785 28.835 7.460 ;
        RECT 29.545 5.785 29.715 7.460 ;
        RECT 30.555 4.340 30.865 7.460 ;
        RECT 31.715 5.445 31.885 7.460 ;
        RECT 32.595 5.785 32.765 7.460 ;
        RECT 33.475 5.785 33.645 7.460 ;
        RECT 34.355 5.785 34.525 7.460 ;
        RECT 35.365 4.340 35.675 7.460 ;
        RECT 36.225 5.365 36.395 7.460 ;
        RECT 37.105 5.785 37.275 7.460 ;
        RECT 37.985 5.785 38.155 7.460 ;
        RECT 38.695 4.340 39.005 7.460 ;
        RECT 39.855 5.445 40.025 7.460 ;
        RECT 40.735 5.785 40.905 7.460 ;
        RECT 41.615 5.785 41.785 7.460 ;
        RECT 42.495 5.785 42.665 7.460 ;
        RECT 43.505 4.340 43.815 7.460 ;
        RECT 44.665 5.445 44.835 7.460 ;
        RECT 45.545 5.785 45.715 7.460 ;
        RECT 46.425 5.785 46.595 7.460 ;
        RECT 47.305 5.785 47.475 7.460 ;
        RECT 48.315 4.340 48.625 7.460 ;
        RECT 49.175 5.365 49.345 7.460 ;
        RECT 50.055 5.785 50.225 7.460 ;
        RECT 50.935 5.785 51.105 7.460 ;
        RECT 51.645 4.340 51.955 7.460 ;
        RECT 52.805 5.445 52.975 7.460 ;
        RECT 53.685 5.785 53.855 7.460 ;
        RECT 54.565 5.785 54.735 7.460 ;
        RECT 55.445 5.785 55.615 7.460 ;
        RECT 56.455 4.340 56.765 7.460 ;
        RECT 57.615 5.445 57.785 7.460 ;
        RECT 58.495 5.785 58.665 7.460 ;
        RECT 59.375 5.785 59.545 7.460 ;
        RECT 60.255 5.785 60.425 7.460 ;
        RECT 61.265 4.340 61.575 7.460 ;
        RECT 62.125 5.365 62.295 7.460 ;
        RECT 63.005 5.785 63.175 7.460 ;
        RECT 63.885 5.785 64.055 7.460 ;
        RECT 64.595 4.340 64.905 7.460 ;
        RECT 65.755 5.445 65.925 7.460 ;
        RECT 66.635 5.785 66.805 7.460 ;
        RECT 67.515 5.785 67.685 7.460 ;
        RECT 68.395 5.785 68.565 7.460 ;
        RECT 69.405 4.340 69.715 7.460 ;
        RECT 70.565 5.445 70.735 7.460 ;
        RECT 71.445 5.785 71.615 7.460 ;
        RECT 72.325 5.785 72.495 7.460 ;
        RECT 73.205 5.785 73.375 7.460 ;
        RECT 74.215 4.340 74.525 7.460 ;
        RECT 75.075 5.365 75.245 7.460 ;
        RECT 75.955 5.785 76.125 7.460 ;
        RECT 76.835 5.785 77.005 7.460 ;
        RECT 77.545 4.340 77.855 7.460 ;
        RECT 78.405 5.355 78.575 7.460 ;
        RECT 79.285 5.785 79.455 7.460 ;
        RECT 80.165 5.355 80.335 7.460 ;
        RECT 80.875 4.340 81.185 7.460 ;
        RECT 84.205 4.340 84.515 7.460 ;
        RECT 87.535 4.340 87.845 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 0.995 7.525 1.165 7.695 ;
        RECT 1.355 7.525 1.525 7.695 ;
        RECT 1.715 7.525 1.885 7.695 ;
        RECT 2.075 7.525 2.245 7.695 ;
        RECT 2.565 7.525 2.735 7.695 ;
        RECT 2.925 7.525 3.095 7.695 ;
        RECT 3.285 7.525 3.455 7.695 ;
        RECT 3.645 7.525 3.815 7.695 ;
        RECT 4.005 7.525 4.175 7.695 ;
        RECT 4.365 7.525 4.535 7.695 ;
        RECT 5.085 7.525 5.255 7.695 ;
        RECT 5.445 7.525 5.615 7.695 ;
        RECT 5.805 7.525 5.975 7.695 ;
        RECT 6.165 7.525 6.335 7.695 ;
        RECT 6.525 7.525 6.695 7.695 ;
        RECT 6.885 7.525 7.055 7.695 ;
        RECT 7.375 7.525 7.545 7.695 ;
        RECT 7.735 7.525 7.905 7.695 ;
        RECT 8.095 7.525 8.265 7.695 ;
        RECT 8.455 7.525 8.625 7.695 ;
        RECT 8.815 7.525 8.985 7.695 ;
        RECT 9.175 7.525 9.345 7.695 ;
        RECT 9.895 7.525 10.065 7.695 ;
        RECT 10.255 7.525 10.425 7.695 ;
        RECT 10.615 7.525 10.785 7.695 ;
        RECT 10.975 7.525 11.145 7.695 ;
        RECT 11.425 7.525 11.595 7.695 ;
        RECT 11.785 7.525 11.955 7.695 ;
        RECT 12.145 7.525 12.315 7.695 ;
        RECT 12.505 7.525 12.675 7.695 ;
        RECT 13.225 7.525 13.395 7.695 ;
        RECT 13.585 7.525 13.755 7.695 ;
        RECT 13.945 7.525 14.115 7.695 ;
        RECT 14.305 7.525 14.475 7.695 ;
        RECT 14.665 7.525 14.835 7.695 ;
        RECT 15.025 7.525 15.195 7.695 ;
        RECT 15.515 7.525 15.685 7.695 ;
        RECT 15.875 7.525 16.045 7.695 ;
        RECT 16.235 7.525 16.405 7.695 ;
        RECT 16.595 7.525 16.765 7.695 ;
        RECT 16.955 7.525 17.125 7.695 ;
        RECT 17.315 7.525 17.485 7.695 ;
        RECT 18.035 7.525 18.205 7.695 ;
        RECT 18.395 7.525 18.565 7.695 ;
        RECT 18.755 7.525 18.925 7.695 ;
        RECT 19.115 7.525 19.285 7.695 ;
        RECT 19.475 7.525 19.645 7.695 ;
        RECT 19.835 7.525 20.005 7.695 ;
        RECT 20.325 7.525 20.495 7.695 ;
        RECT 20.685 7.525 20.855 7.695 ;
        RECT 21.045 7.525 21.215 7.695 ;
        RECT 21.405 7.525 21.575 7.695 ;
        RECT 21.765 7.525 21.935 7.695 ;
        RECT 22.125 7.525 22.295 7.695 ;
        RECT 22.845 7.525 23.015 7.695 ;
        RECT 23.205 7.525 23.375 7.695 ;
        RECT 23.565 7.525 23.735 7.695 ;
        RECT 23.925 7.525 24.095 7.695 ;
        RECT 24.375 7.525 24.545 7.695 ;
        RECT 24.735 7.525 24.905 7.695 ;
        RECT 25.095 7.525 25.265 7.695 ;
        RECT 25.455 7.525 25.625 7.695 ;
        RECT 26.175 7.525 26.345 7.695 ;
        RECT 26.535 7.525 26.705 7.695 ;
        RECT 26.895 7.525 27.065 7.695 ;
        RECT 27.255 7.525 27.425 7.695 ;
        RECT 27.615 7.525 27.785 7.695 ;
        RECT 27.975 7.525 28.145 7.695 ;
        RECT 28.465 7.525 28.635 7.695 ;
        RECT 28.825 7.525 28.995 7.695 ;
        RECT 29.185 7.525 29.355 7.695 ;
        RECT 29.545 7.525 29.715 7.695 ;
        RECT 29.905 7.525 30.075 7.695 ;
        RECT 30.265 7.525 30.435 7.695 ;
        RECT 30.985 7.525 31.155 7.695 ;
        RECT 31.345 7.525 31.515 7.695 ;
        RECT 31.705 7.525 31.875 7.695 ;
        RECT 32.065 7.525 32.235 7.695 ;
        RECT 32.425 7.525 32.595 7.695 ;
        RECT 32.785 7.525 32.955 7.695 ;
        RECT 33.275 7.525 33.445 7.695 ;
        RECT 33.635 7.525 33.805 7.695 ;
        RECT 33.995 7.525 34.165 7.695 ;
        RECT 34.355 7.525 34.525 7.695 ;
        RECT 34.715 7.525 34.885 7.695 ;
        RECT 35.075 7.525 35.245 7.695 ;
        RECT 35.795 7.525 35.965 7.695 ;
        RECT 36.155 7.525 36.325 7.695 ;
        RECT 36.515 7.525 36.685 7.695 ;
        RECT 36.875 7.525 37.045 7.695 ;
        RECT 37.325 7.525 37.495 7.695 ;
        RECT 37.685 7.525 37.855 7.695 ;
        RECT 38.045 7.525 38.215 7.695 ;
        RECT 38.405 7.525 38.575 7.695 ;
        RECT 39.125 7.525 39.295 7.695 ;
        RECT 39.485 7.525 39.655 7.695 ;
        RECT 39.845 7.525 40.015 7.695 ;
        RECT 40.205 7.525 40.375 7.695 ;
        RECT 40.565 7.525 40.735 7.695 ;
        RECT 40.925 7.525 41.095 7.695 ;
        RECT 41.415 7.525 41.585 7.695 ;
        RECT 41.775 7.525 41.945 7.695 ;
        RECT 42.135 7.525 42.305 7.695 ;
        RECT 42.495 7.525 42.665 7.695 ;
        RECT 42.855 7.525 43.025 7.695 ;
        RECT 43.215 7.525 43.385 7.695 ;
        RECT 43.935 7.525 44.105 7.695 ;
        RECT 44.295 7.525 44.465 7.695 ;
        RECT 44.655 7.525 44.825 7.695 ;
        RECT 45.015 7.525 45.185 7.695 ;
        RECT 45.375 7.525 45.545 7.695 ;
        RECT 45.735 7.525 45.905 7.695 ;
        RECT 46.225 7.525 46.395 7.695 ;
        RECT 46.585 7.525 46.755 7.695 ;
        RECT 46.945 7.525 47.115 7.695 ;
        RECT 47.305 7.525 47.475 7.695 ;
        RECT 47.665 7.525 47.835 7.695 ;
        RECT 48.025 7.525 48.195 7.695 ;
        RECT 48.745 7.525 48.915 7.695 ;
        RECT 49.105 7.525 49.275 7.695 ;
        RECT 49.465 7.525 49.635 7.695 ;
        RECT 49.825 7.525 49.995 7.695 ;
        RECT 50.275 7.525 50.445 7.695 ;
        RECT 50.635 7.525 50.805 7.695 ;
        RECT 50.995 7.525 51.165 7.695 ;
        RECT 51.355 7.525 51.525 7.695 ;
        RECT 52.075 7.525 52.245 7.695 ;
        RECT 52.435 7.525 52.605 7.695 ;
        RECT 52.795 7.525 52.965 7.695 ;
        RECT 53.155 7.525 53.325 7.695 ;
        RECT 53.515 7.525 53.685 7.695 ;
        RECT 53.875 7.525 54.045 7.695 ;
        RECT 54.365 7.525 54.535 7.695 ;
        RECT 54.725 7.525 54.895 7.695 ;
        RECT 55.085 7.525 55.255 7.695 ;
        RECT 55.445 7.525 55.615 7.695 ;
        RECT 55.805 7.525 55.975 7.695 ;
        RECT 56.165 7.525 56.335 7.695 ;
        RECT 56.885 7.525 57.055 7.695 ;
        RECT 57.245 7.525 57.415 7.695 ;
        RECT 57.605 7.525 57.775 7.695 ;
        RECT 57.965 7.525 58.135 7.695 ;
        RECT 58.325 7.525 58.495 7.695 ;
        RECT 58.685 7.525 58.855 7.695 ;
        RECT 59.175 7.525 59.345 7.695 ;
        RECT 59.535 7.525 59.705 7.695 ;
        RECT 59.895 7.525 60.065 7.695 ;
        RECT 60.255 7.525 60.425 7.695 ;
        RECT 60.615 7.525 60.785 7.695 ;
        RECT 60.975 7.525 61.145 7.695 ;
        RECT 61.695 7.525 61.865 7.695 ;
        RECT 62.055 7.525 62.225 7.695 ;
        RECT 62.415 7.525 62.585 7.695 ;
        RECT 62.775 7.525 62.945 7.695 ;
        RECT 63.225 7.525 63.395 7.695 ;
        RECT 63.585 7.525 63.755 7.695 ;
        RECT 63.945 7.525 64.115 7.695 ;
        RECT 64.305 7.525 64.475 7.695 ;
        RECT 65.025 7.525 65.195 7.695 ;
        RECT 65.385 7.525 65.555 7.695 ;
        RECT 65.745 7.525 65.915 7.695 ;
        RECT 66.105 7.525 66.275 7.695 ;
        RECT 66.465 7.525 66.635 7.695 ;
        RECT 66.825 7.525 66.995 7.695 ;
        RECT 67.315 7.525 67.485 7.695 ;
        RECT 67.675 7.525 67.845 7.695 ;
        RECT 68.035 7.525 68.205 7.695 ;
        RECT 68.395 7.525 68.565 7.695 ;
        RECT 68.755 7.525 68.925 7.695 ;
        RECT 69.115 7.525 69.285 7.695 ;
        RECT 69.835 7.525 70.005 7.695 ;
        RECT 70.195 7.525 70.365 7.695 ;
        RECT 70.555 7.525 70.725 7.695 ;
        RECT 70.915 7.525 71.085 7.695 ;
        RECT 71.275 7.525 71.445 7.695 ;
        RECT 71.635 7.525 71.805 7.695 ;
        RECT 72.125 7.525 72.295 7.695 ;
        RECT 72.485 7.525 72.655 7.695 ;
        RECT 72.845 7.525 73.015 7.695 ;
        RECT 73.205 7.525 73.375 7.695 ;
        RECT 73.565 7.525 73.735 7.695 ;
        RECT 73.925 7.525 74.095 7.695 ;
        RECT 74.645 7.525 74.815 7.695 ;
        RECT 75.005 7.525 75.175 7.695 ;
        RECT 75.365 7.525 75.535 7.695 ;
        RECT 75.725 7.525 75.895 7.695 ;
        RECT 76.175 7.525 76.345 7.695 ;
        RECT 76.535 7.525 76.705 7.695 ;
        RECT 76.895 7.525 77.065 7.695 ;
        RECT 77.255 7.525 77.425 7.695 ;
        RECT 77.975 7.525 78.145 7.695 ;
        RECT 78.335 7.525 78.505 7.695 ;
        RECT 78.695 7.525 78.865 7.695 ;
        RECT 79.055 7.525 79.225 7.695 ;
        RECT 79.505 7.525 79.675 7.695 ;
        RECT 79.865 7.525 80.035 7.695 ;
        RECT 80.225 7.525 80.395 7.695 ;
        RECT 80.585 7.525 80.755 7.695 ;
        RECT 81.305 7.525 81.475 7.695 ;
        RECT 81.665 7.525 81.835 7.695 ;
        RECT 82.025 7.525 82.195 7.695 ;
        RECT 82.385 7.525 82.555 7.695 ;
        RECT 82.835 7.525 83.005 7.695 ;
        RECT 83.195 7.525 83.365 7.695 ;
        RECT 83.555 7.525 83.725 7.695 ;
        RECT 83.915 7.525 84.085 7.695 ;
        RECT 84.635 7.525 84.805 7.695 ;
        RECT 84.995 7.525 85.165 7.695 ;
        RECT 85.355 7.525 85.525 7.695 ;
        RECT 85.715 7.525 85.885 7.695 ;
        RECT 86.165 7.525 86.335 7.695 ;
        RECT 86.525 7.525 86.695 7.695 ;
        RECT 86.885 7.525 87.055 7.695 ;
        RECT 87.245 7.525 87.415 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 87.845 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 62.126400 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 87.975 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 4.525 -0.075 5.095 -0.065 ;
        RECT 9.335 -0.075 9.905 -0.065 ;
        RECT 12.665 -0.075 13.235 -0.065 ;
        RECT 17.475 -0.075 18.045 -0.065 ;
        RECT 22.285 -0.075 22.855 -0.065 ;
        RECT 25.615 -0.075 26.185 -0.065 ;
        RECT 30.425 -0.075 30.995 -0.065 ;
        RECT 35.235 -0.075 35.805 -0.065 ;
        RECT 38.565 -0.075 39.135 -0.065 ;
        RECT 43.375 -0.075 43.945 -0.065 ;
        RECT 48.185 -0.075 48.755 -0.065 ;
        RECT 51.515 -0.075 52.085 -0.065 ;
        RECT 56.325 -0.075 56.895 -0.065 ;
        RECT 61.135 -0.075 61.705 -0.065 ;
        RECT 64.465 -0.075 65.035 -0.065 ;
        RECT 69.275 -0.075 69.845 -0.065 ;
        RECT 74.085 -0.075 74.655 -0.065 ;
        RECT 77.415 -0.075 77.985 -0.065 ;
        RECT 80.745 -0.075 81.315 -0.065 ;
        RECT 84.075 -0.075 84.645 -0.065 ;
        RECT 87.405 -0.075 87.975 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 0.990 0.310 1.160 1.270 ;
        RECT 4.655 0.310 4.965 2.860 ;
        RECT 5.800 0.310 5.970 1.270 ;
        RECT 9.465 0.310 9.775 2.860 ;
        RECT 10.715 0.310 10.885 1.260 ;
        RECT 12.795 0.310 13.105 2.860 ;
        RECT 13.940 0.310 14.110 1.270 ;
        RECT 17.605 0.310 17.915 2.860 ;
        RECT 18.750 0.310 18.920 1.270 ;
        RECT 22.415 0.310 22.725 2.860 ;
        RECT 23.665 0.310 23.835 1.260 ;
        RECT 25.745 0.310 26.055 2.860 ;
        RECT 26.890 0.310 27.060 1.270 ;
        RECT 30.555 0.310 30.865 2.860 ;
        RECT 31.700 0.310 31.870 1.270 ;
        RECT 35.365 0.310 35.675 2.860 ;
        RECT 36.615 0.310 36.785 1.260 ;
        RECT 38.695 0.310 39.005 2.860 ;
        RECT 39.840 0.310 40.010 1.270 ;
        RECT 43.505 0.310 43.815 2.860 ;
        RECT 44.650 0.310 44.820 1.270 ;
        RECT 48.315 0.310 48.625 2.860 ;
        RECT 49.565 0.310 49.735 1.260 ;
        RECT 51.645 0.310 51.955 2.860 ;
        RECT 52.790 0.310 52.960 1.270 ;
        RECT 56.455 0.310 56.765 2.860 ;
        RECT 57.600 0.310 57.770 1.270 ;
        RECT 61.265 0.310 61.575 2.860 ;
        RECT 62.515 0.310 62.685 1.260 ;
        RECT 64.595 0.310 64.905 2.860 ;
        RECT 65.740 0.310 65.910 1.270 ;
        RECT 69.405 0.310 69.715 2.860 ;
        RECT 70.550 0.310 70.720 1.270 ;
        RECT 74.215 0.310 74.525 2.860 ;
        RECT 75.465 0.310 75.635 1.260 ;
        RECT 77.545 0.310 77.855 2.860 ;
        RECT 78.795 0.310 78.965 1.260 ;
        RECT 80.875 0.310 81.185 2.860 ;
        RECT 82.125 0.310 82.295 1.260 ;
        RECT 84.205 0.310 84.515 2.860 ;
        RECT 85.455 0.310 85.625 1.260 ;
        RECT 87.535 0.310 87.845 2.860 ;
        RECT -0.155 0.235 83.095 0.310 ;
        RECT 83.265 0.235 87.845 0.310 ;
        RECT -0.155 0.000 87.845 0.235 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 0.995 0.065 1.165 0.235 ;
        RECT 1.355 0.065 1.525 0.235 ;
        RECT 1.715 0.065 1.885 0.235 ;
        RECT 2.075 0.065 2.245 0.235 ;
        RECT 2.565 0.065 2.735 0.235 ;
        RECT 2.925 0.065 3.095 0.235 ;
        RECT 3.285 0.065 3.455 0.235 ;
        RECT 3.645 0.065 3.815 0.235 ;
        RECT 4.005 0.065 4.175 0.235 ;
        RECT 4.365 0.065 4.535 0.235 ;
        RECT 5.085 0.065 5.255 0.235 ;
        RECT 5.445 0.065 5.615 0.235 ;
        RECT 5.805 0.065 5.975 0.235 ;
        RECT 6.165 0.065 6.335 0.235 ;
        RECT 6.525 0.065 6.695 0.235 ;
        RECT 6.885 0.065 7.055 0.235 ;
        RECT 7.375 0.065 7.545 0.235 ;
        RECT 7.735 0.065 7.905 0.235 ;
        RECT 8.095 0.065 8.265 0.235 ;
        RECT 8.455 0.065 8.625 0.235 ;
        RECT 8.815 0.065 8.985 0.235 ;
        RECT 9.175 0.065 9.345 0.235 ;
        RECT 9.895 0.065 10.065 0.235 ;
        RECT 10.255 0.065 10.425 0.235 ;
        RECT 10.615 0.065 10.785 0.235 ;
        RECT 10.975 0.065 11.145 0.235 ;
        RECT 11.425 0.065 11.595 0.235 ;
        RECT 11.785 0.065 11.955 0.235 ;
        RECT 12.145 0.065 12.315 0.235 ;
        RECT 12.505 0.065 12.675 0.235 ;
        RECT 13.225 0.065 13.395 0.235 ;
        RECT 13.585 0.065 13.755 0.235 ;
        RECT 13.945 0.065 14.115 0.235 ;
        RECT 14.305 0.065 14.475 0.235 ;
        RECT 14.665 0.065 14.835 0.235 ;
        RECT 15.025 0.065 15.195 0.235 ;
        RECT 15.515 0.065 15.685 0.235 ;
        RECT 15.875 0.065 16.045 0.235 ;
        RECT 16.235 0.065 16.405 0.235 ;
        RECT 16.595 0.065 16.765 0.235 ;
        RECT 16.955 0.065 17.125 0.235 ;
        RECT 17.315 0.065 17.485 0.235 ;
        RECT 18.035 0.065 18.205 0.235 ;
        RECT 18.395 0.065 18.565 0.235 ;
        RECT 18.755 0.065 18.925 0.235 ;
        RECT 19.115 0.065 19.285 0.235 ;
        RECT 19.475 0.065 19.645 0.235 ;
        RECT 19.835 0.065 20.005 0.235 ;
        RECT 20.325 0.065 20.495 0.235 ;
        RECT 20.685 0.065 20.855 0.235 ;
        RECT 21.045 0.065 21.215 0.235 ;
        RECT 21.405 0.065 21.575 0.235 ;
        RECT 21.765 0.065 21.935 0.235 ;
        RECT 22.125 0.065 22.295 0.235 ;
        RECT 22.845 0.065 23.015 0.235 ;
        RECT 23.205 0.065 23.375 0.235 ;
        RECT 23.565 0.065 23.735 0.235 ;
        RECT 23.925 0.065 24.095 0.235 ;
        RECT 24.375 0.065 24.545 0.235 ;
        RECT 24.735 0.065 24.905 0.235 ;
        RECT 25.095 0.065 25.265 0.235 ;
        RECT 25.455 0.065 25.625 0.235 ;
        RECT 26.175 0.065 26.345 0.235 ;
        RECT 26.535 0.065 26.705 0.235 ;
        RECT 26.895 0.065 27.065 0.235 ;
        RECT 27.255 0.065 27.425 0.235 ;
        RECT 27.615 0.065 27.785 0.235 ;
        RECT 27.975 0.065 28.145 0.235 ;
        RECT 28.465 0.065 28.635 0.235 ;
        RECT 28.825 0.065 28.995 0.235 ;
        RECT 29.185 0.065 29.355 0.235 ;
        RECT 29.545 0.065 29.715 0.235 ;
        RECT 29.905 0.065 30.075 0.235 ;
        RECT 30.265 0.065 30.435 0.235 ;
        RECT 30.985 0.065 31.155 0.235 ;
        RECT 31.345 0.065 31.515 0.235 ;
        RECT 31.705 0.065 31.875 0.235 ;
        RECT 32.065 0.065 32.235 0.235 ;
        RECT 32.425 0.065 32.595 0.235 ;
        RECT 32.785 0.065 32.955 0.235 ;
        RECT 33.275 0.065 33.445 0.235 ;
        RECT 33.635 0.065 33.805 0.235 ;
        RECT 33.995 0.065 34.165 0.235 ;
        RECT 34.355 0.065 34.525 0.235 ;
        RECT 34.715 0.065 34.885 0.235 ;
        RECT 35.075 0.065 35.245 0.235 ;
        RECT 35.795 0.065 35.965 0.235 ;
        RECT 36.155 0.065 36.325 0.235 ;
        RECT 36.515 0.065 36.685 0.235 ;
        RECT 36.875 0.065 37.045 0.235 ;
        RECT 37.325 0.065 37.495 0.235 ;
        RECT 37.685 0.065 37.855 0.235 ;
        RECT 38.045 0.065 38.215 0.235 ;
        RECT 38.405 0.065 38.575 0.235 ;
        RECT 39.125 0.065 39.295 0.235 ;
        RECT 39.485 0.065 39.655 0.235 ;
        RECT 39.845 0.065 40.015 0.235 ;
        RECT 40.205 0.065 40.375 0.235 ;
        RECT 40.565 0.065 40.735 0.235 ;
        RECT 40.925 0.065 41.095 0.235 ;
        RECT 41.415 0.065 41.585 0.235 ;
        RECT 41.775 0.065 41.945 0.235 ;
        RECT 42.135 0.065 42.305 0.235 ;
        RECT 42.495 0.065 42.665 0.235 ;
        RECT 42.855 0.065 43.025 0.235 ;
        RECT 43.215 0.065 43.385 0.235 ;
        RECT 43.935 0.065 44.105 0.235 ;
        RECT 44.295 0.065 44.465 0.235 ;
        RECT 44.655 0.065 44.825 0.235 ;
        RECT 45.015 0.065 45.185 0.235 ;
        RECT 45.375 0.065 45.545 0.235 ;
        RECT 45.735 0.065 45.905 0.235 ;
        RECT 46.225 0.065 46.395 0.235 ;
        RECT 46.585 0.065 46.755 0.235 ;
        RECT 46.945 0.065 47.115 0.235 ;
        RECT 47.305 0.065 47.475 0.235 ;
        RECT 47.665 0.065 47.835 0.235 ;
        RECT 48.025 0.065 48.195 0.235 ;
        RECT 48.745 0.065 48.915 0.235 ;
        RECT 49.105 0.065 49.275 0.235 ;
        RECT 49.465 0.065 49.635 0.235 ;
        RECT 49.825 0.065 49.995 0.235 ;
        RECT 50.275 0.065 50.445 0.235 ;
        RECT 50.635 0.065 50.805 0.235 ;
        RECT 50.995 0.065 51.165 0.235 ;
        RECT 51.355 0.065 51.525 0.235 ;
        RECT 52.075 0.065 52.245 0.235 ;
        RECT 52.435 0.065 52.605 0.235 ;
        RECT 52.795 0.065 52.965 0.235 ;
        RECT 53.155 0.065 53.325 0.235 ;
        RECT 53.515 0.065 53.685 0.235 ;
        RECT 53.875 0.065 54.045 0.235 ;
        RECT 54.365 0.065 54.535 0.235 ;
        RECT 54.725 0.065 54.895 0.235 ;
        RECT 55.085 0.065 55.255 0.235 ;
        RECT 55.445 0.065 55.615 0.235 ;
        RECT 55.805 0.065 55.975 0.235 ;
        RECT 56.165 0.065 56.335 0.235 ;
        RECT 56.885 0.065 57.055 0.235 ;
        RECT 57.245 0.065 57.415 0.235 ;
        RECT 57.605 0.065 57.775 0.235 ;
        RECT 57.965 0.065 58.135 0.235 ;
        RECT 58.325 0.065 58.495 0.235 ;
        RECT 58.685 0.065 58.855 0.235 ;
        RECT 59.175 0.065 59.345 0.235 ;
        RECT 59.535 0.065 59.705 0.235 ;
        RECT 59.895 0.065 60.065 0.235 ;
        RECT 60.255 0.065 60.425 0.235 ;
        RECT 60.615 0.065 60.785 0.235 ;
        RECT 60.975 0.065 61.145 0.235 ;
        RECT 61.695 0.065 61.865 0.235 ;
        RECT 62.055 0.065 62.225 0.235 ;
        RECT 62.415 0.065 62.585 0.235 ;
        RECT 62.775 0.065 62.945 0.235 ;
        RECT 63.225 0.065 63.395 0.235 ;
        RECT 63.585 0.065 63.755 0.235 ;
        RECT 63.945 0.065 64.115 0.235 ;
        RECT 64.305 0.065 64.475 0.235 ;
        RECT 65.025 0.065 65.195 0.235 ;
        RECT 65.385 0.065 65.555 0.235 ;
        RECT 65.745 0.065 65.915 0.235 ;
        RECT 66.105 0.065 66.275 0.235 ;
        RECT 66.465 0.065 66.635 0.235 ;
        RECT 66.825 0.065 66.995 0.235 ;
        RECT 67.315 0.065 67.485 0.235 ;
        RECT 67.675 0.065 67.845 0.235 ;
        RECT 68.035 0.065 68.205 0.235 ;
        RECT 68.395 0.065 68.565 0.235 ;
        RECT 68.755 0.065 68.925 0.235 ;
        RECT 69.115 0.065 69.285 0.235 ;
        RECT 69.835 0.065 70.005 0.235 ;
        RECT 70.195 0.065 70.365 0.235 ;
        RECT 70.555 0.065 70.725 0.235 ;
        RECT 70.915 0.065 71.085 0.235 ;
        RECT 71.275 0.065 71.445 0.235 ;
        RECT 71.635 0.065 71.805 0.235 ;
        RECT 72.125 0.065 72.295 0.235 ;
        RECT 72.485 0.065 72.655 0.235 ;
        RECT 72.845 0.065 73.015 0.235 ;
        RECT 73.205 0.065 73.375 0.235 ;
        RECT 73.565 0.065 73.735 0.235 ;
        RECT 73.925 0.065 74.095 0.235 ;
        RECT 74.645 0.065 74.815 0.235 ;
        RECT 75.005 0.065 75.175 0.235 ;
        RECT 75.365 0.065 75.535 0.235 ;
        RECT 75.725 0.065 75.895 0.235 ;
        RECT 76.175 0.065 76.345 0.235 ;
        RECT 76.535 0.065 76.705 0.235 ;
        RECT 76.895 0.065 77.065 0.235 ;
        RECT 77.255 0.065 77.425 0.235 ;
        RECT 77.975 0.065 78.145 0.235 ;
        RECT 78.335 0.065 78.505 0.235 ;
        RECT 78.695 0.065 78.865 0.235 ;
        RECT 79.055 0.065 79.225 0.235 ;
        RECT 79.505 0.065 79.675 0.235 ;
        RECT 79.865 0.065 80.035 0.235 ;
        RECT 80.225 0.065 80.395 0.235 ;
        RECT 80.585 0.065 80.755 0.235 ;
        RECT 81.305 0.065 81.475 0.235 ;
        RECT 81.665 0.065 81.835 0.235 ;
        RECT 82.025 0.065 82.195 0.235 ;
        RECT 82.385 0.065 82.555 0.235 ;
        RECT 82.835 0.065 83.005 0.235 ;
        RECT 83.195 0.065 83.365 0.235 ;
        RECT 83.555 0.065 83.725 0.235 ;
        RECT 83.915 0.065 84.085 0.235 ;
        RECT 84.635 0.065 84.805 0.235 ;
        RECT 84.995 0.065 85.165 0.235 ;
        RECT 85.355 0.065 85.525 0.235 ;
        RECT 85.715 0.065 85.885 0.235 ;
        RECT 86.165 0.065 86.335 0.235 ;
        RECT 86.525 0.065 86.695 0.235 ;
        RECT 86.885 0.065 87.055 0.235 ;
        RECT 87.245 0.065 87.415 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 87.845 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 1.445 5.470 1.615 7.250 ;
        RECT 2.325 5.470 2.495 7.250 ;
        RECT 3.205 5.470 3.375 7.250 ;
        RECT 6.255 5.470 6.425 7.250 ;
        RECT 7.135 5.470 7.305 7.250 ;
        RECT 8.015 5.470 8.185 7.250 ;
        RECT 10.765 5.515 10.935 7.250 ;
        RECT 11.645 5.515 11.815 7.250 ;
        RECT 1.445 5.300 4.155 5.470 ;
        RECT 6.255 5.300 8.965 5.470 ;
        RECT 10.765 5.345 12.295 5.515 ;
        RECT 1.025 2.055 1.195 5.095 ;
        RECT 3.245 2.055 3.415 5.095 ;
        RECT 0.505 1.815 0.675 1.895 ;
        RECT 1.475 1.815 1.645 1.895 ;
        RECT 2.445 1.815 2.615 1.895 ;
        RECT 0.505 1.645 2.615 1.815 ;
        RECT 0.505 0.515 0.675 1.645 ;
        RECT 1.475 0.765 1.645 1.645 ;
        RECT 2.445 1.565 2.615 1.645 ;
        RECT 1.965 1.220 2.135 1.300 ;
        RECT 3.015 1.220 3.185 1.895 ;
        RECT 3.985 1.890 4.155 5.300 ;
        RECT 5.835 2.055 6.005 5.095 ;
        RECT 1.965 1.050 3.185 1.220 ;
        RECT 1.965 0.970 2.135 1.050 ;
        RECT 2.445 0.765 2.615 0.845 ;
        RECT 1.475 0.595 2.615 0.765 ;
        RECT 1.475 0.515 1.645 0.595 ;
        RECT 2.445 0.515 2.615 0.595 ;
        RECT 3.015 0.765 3.185 1.050 ;
        RECT 3.500 1.720 4.155 1.890 ;
        RECT 5.315 1.815 5.485 1.895 ;
        RECT 6.285 1.815 6.455 1.895 ;
        RECT 7.255 1.815 7.425 1.895 ;
        RECT 3.500 0.985 3.670 1.720 ;
        RECT 5.315 1.645 7.425 1.815 ;
        RECT 3.985 0.765 4.155 1.535 ;
        RECT 3.015 0.595 4.155 0.765 ;
        RECT 3.015 0.515 3.185 0.595 ;
        RECT 3.985 0.515 4.155 0.595 ;
        RECT 5.315 0.515 5.485 1.645 ;
        RECT 6.285 0.765 6.455 1.645 ;
        RECT 7.255 1.565 7.425 1.645 ;
        RECT 6.775 1.220 6.945 1.300 ;
        RECT 7.825 1.220 7.995 1.895 ;
        RECT 8.795 1.890 8.965 5.300 ;
        RECT 10.645 2.055 10.815 5.095 ;
        RECT 11.415 4.940 11.585 5.095 ;
        RECT 11.385 4.765 11.585 4.940 ;
        RECT 11.385 2.055 11.555 4.765 ;
        RECT 6.775 1.050 7.995 1.220 ;
        RECT 6.775 0.970 6.945 1.050 ;
        RECT 7.255 0.765 7.425 0.845 ;
        RECT 6.285 0.595 7.425 0.765 ;
        RECT 6.285 0.515 6.455 0.595 ;
        RECT 7.255 0.515 7.425 0.595 ;
        RECT 7.825 0.765 7.995 1.050 ;
        RECT 8.310 1.720 8.965 1.890 ;
        RECT 10.230 1.805 10.400 1.885 ;
        RECT 11.200 1.805 11.370 1.885 ;
        RECT 12.125 1.880 12.295 5.345 ;
        RECT 14.395 5.470 14.565 7.250 ;
        RECT 15.275 5.470 15.445 7.250 ;
        RECT 16.155 5.470 16.325 7.250 ;
        RECT 19.205 5.470 19.375 7.250 ;
        RECT 20.085 5.470 20.255 7.250 ;
        RECT 20.965 5.470 21.135 7.250 ;
        RECT 23.715 5.515 23.885 7.250 ;
        RECT 24.595 5.515 24.765 7.250 ;
        RECT 14.395 5.300 17.105 5.470 ;
        RECT 19.205 5.300 21.915 5.470 ;
        RECT 23.715 5.345 25.245 5.515 ;
        RECT 13.975 2.055 14.145 5.095 ;
        RECT 8.310 0.985 8.480 1.720 ;
        RECT 10.230 1.635 11.370 1.805 ;
        RECT 8.795 0.765 8.965 1.535 ;
        RECT 7.825 0.595 8.965 0.765 ;
        RECT 7.825 0.515 7.995 0.595 ;
        RECT 8.795 0.515 8.965 0.595 ;
        RECT 10.230 0.505 10.400 1.635 ;
        RECT 11.200 0.755 11.370 1.635 ;
        RECT 11.685 1.710 12.295 1.880 ;
        RECT 13.455 1.815 13.625 1.895 ;
        RECT 14.425 1.815 14.595 1.895 ;
        RECT 15.395 1.815 15.565 1.895 ;
        RECT 11.685 0.975 11.855 1.710 ;
        RECT 13.455 1.645 15.565 1.815 ;
        RECT 12.170 0.755 12.340 1.525 ;
        RECT 11.200 0.585 12.340 0.755 ;
        RECT 11.200 0.505 11.370 0.585 ;
        RECT 12.170 0.505 12.340 0.585 ;
        RECT 13.455 0.515 13.625 1.645 ;
        RECT 14.425 0.765 14.595 1.645 ;
        RECT 15.395 1.565 15.565 1.645 ;
        RECT 14.915 1.220 15.085 1.300 ;
        RECT 15.965 1.220 16.135 1.895 ;
        RECT 16.935 1.890 17.105 5.300 ;
        RECT 18.785 2.055 18.955 5.095 ;
        RECT 21.005 2.055 21.175 5.095 ;
        RECT 14.915 1.050 16.135 1.220 ;
        RECT 14.915 0.970 15.085 1.050 ;
        RECT 15.395 0.765 15.565 0.845 ;
        RECT 14.425 0.595 15.565 0.765 ;
        RECT 14.425 0.515 14.595 0.595 ;
        RECT 15.395 0.515 15.565 0.595 ;
        RECT 15.965 0.765 16.135 1.050 ;
        RECT 16.450 1.720 17.105 1.890 ;
        RECT 18.265 1.815 18.435 1.895 ;
        RECT 19.235 1.815 19.405 1.895 ;
        RECT 20.205 1.815 20.375 1.895 ;
        RECT 16.450 0.985 16.620 1.720 ;
        RECT 18.265 1.645 20.375 1.815 ;
        RECT 16.935 0.765 17.105 1.535 ;
        RECT 15.965 0.595 17.105 0.765 ;
        RECT 15.965 0.515 16.135 0.595 ;
        RECT 16.935 0.515 17.105 0.595 ;
        RECT 18.265 0.515 18.435 1.645 ;
        RECT 19.235 0.765 19.405 1.645 ;
        RECT 20.205 1.565 20.375 1.645 ;
        RECT 19.725 1.220 19.895 1.300 ;
        RECT 20.775 1.220 20.945 1.895 ;
        RECT 21.745 1.890 21.915 5.300 ;
        RECT 23.595 2.055 23.765 5.095 ;
        RECT 24.365 4.940 24.535 5.095 ;
        RECT 24.335 4.765 24.535 4.940 ;
        RECT 24.335 2.055 24.505 4.765 ;
        RECT 19.725 1.050 20.945 1.220 ;
        RECT 19.725 0.970 19.895 1.050 ;
        RECT 20.205 0.765 20.375 0.845 ;
        RECT 19.235 0.595 20.375 0.765 ;
        RECT 19.235 0.515 19.405 0.595 ;
        RECT 20.205 0.515 20.375 0.595 ;
        RECT 20.775 0.765 20.945 1.050 ;
        RECT 21.260 1.720 21.915 1.890 ;
        RECT 23.180 1.805 23.350 1.885 ;
        RECT 24.150 1.805 24.320 1.885 ;
        RECT 25.075 1.880 25.245 5.345 ;
        RECT 27.345 5.470 27.515 7.250 ;
        RECT 28.225 5.470 28.395 7.250 ;
        RECT 29.105 5.470 29.275 7.250 ;
        RECT 32.155 5.470 32.325 7.250 ;
        RECT 33.035 5.470 33.205 7.250 ;
        RECT 33.915 5.470 34.085 7.250 ;
        RECT 36.665 5.515 36.835 7.250 ;
        RECT 37.545 5.515 37.715 7.250 ;
        RECT 27.345 5.300 30.055 5.470 ;
        RECT 32.155 5.300 34.865 5.470 ;
        RECT 36.665 5.345 38.195 5.515 ;
        RECT 26.925 2.055 27.095 5.095 ;
        RECT 29.145 2.055 29.315 5.095 ;
        RECT 21.260 0.985 21.430 1.720 ;
        RECT 23.180 1.635 24.320 1.805 ;
        RECT 21.745 0.765 21.915 1.535 ;
        RECT 20.775 0.595 21.915 0.765 ;
        RECT 20.775 0.515 20.945 0.595 ;
        RECT 21.745 0.515 21.915 0.595 ;
        RECT 23.180 0.505 23.350 1.635 ;
        RECT 24.150 0.755 24.320 1.635 ;
        RECT 24.635 1.710 25.245 1.880 ;
        RECT 26.405 1.815 26.575 1.895 ;
        RECT 27.375 1.815 27.545 1.895 ;
        RECT 28.345 1.815 28.515 1.895 ;
        RECT 24.635 0.975 24.805 1.710 ;
        RECT 26.405 1.645 28.515 1.815 ;
        RECT 25.120 0.755 25.290 1.525 ;
        RECT 24.150 0.585 25.290 0.755 ;
        RECT 24.150 0.505 24.320 0.585 ;
        RECT 25.120 0.505 25.290 0.585 ;
        RECT 26.405 0.515 26.575 1.645 ;
        RECT 27.375 0.765 27.545 1.645 ;
        RECT 28.345 1.565 28.515 1.645 ;
        RECT 27.865 1.220 28.035 1.300 ;
        RECT 28.915 1.220 29.085 1.895 ;
        RECT 29.885 1.890 30.055 5.300 ;
        RECT 31.735 2.055 31.905 5.095 ;
        RECT 27.865 1.050 29.085 1.220 ;
        RECT 27.865 0.970 28.035 1.050 ;
        RECT 28.345 0.765 28.515 0.845 ;
        RECT 27.375 0.595 28.515 0.765 ;
        RECT 27.375 0.515 27.545 0.595 ;
        RECT 28.345 0.515 28.515 0.595 ;
        RECT 28.915 0.765 29.085 1.050 ;
        RECT 29.400 1.720 30.055 1.890 ;
        RECT 31.215 1.815 31.385 1.895 ;
        RECT 32.185 1.815 32.355 1.895 ;
        RECT 33.155 1.815 33.325 1.895 ;
        RECT 29.400 0.985 29.570 1.720 ;
        RECT 31.215 1.645 33.325 1.815 ;
        RECT 29.885 0.765 30.055 1.535 ;
        RECT 28.915 0.595 30.055 0.765 ;
        RECT 28.915 0.515 29.085 0.595 ;
        RECT 29.885 0.515 30.055 0.595 ;
        RECT 31.215 0.515 31.385 1.645 ;
        RECT 32.185 0.765 32.355 1.645 ;
        RECT 33.155 1.565 33.325 1.645 ;
        RECT 32.675 1.220 32.845 1.300 ;
        RECT 33.725 1.220 33.895 1.895 ;
        RECT 34.695 1.890 34.865 5.300 ;
        RECT 36.545 2.055 36.715 5.095 ;
        RECT 37.315 4.940 37.485 5.095 ;
        RECT 37.285 4.765 37.485 4.940 ;
        RECT 37.285 2.055 37.455 4.765 ;
        RECT 32.675 1.050 33.895 1.220 ;
        RECT 32.675 0.970 32.845 1.050 ;
        RECT 33.155 0.765 33.325 0.845 ;
        RECT 32.185 0.595 33.325 0.765 ;
        RECT 32.185 0.515 32.355 0.595 ;
        RECT 33.155 0.515 33.325 0.595 ;
        RECT 33.725 0.765 33.895 1.050 ;
        RECT 34.210 1.720 34.865 1.890 ;
        RECT 36.130 1.805 36.300 1.885 ;
        RECT 37.100 1.805 37.270 1.885 ;
        RECT 38.025 1.880 38.195 5.345 ;
        RECT 40.295 5.470 40.465 7.250 ;
        RECT 41.175 5.470 41.345 7.250 ;
        RECT 42.055 5.470 42.225 7.250 ;
        RECT 45.105 5.470 45.275 7.250 ;
        RECT 45.985 5.470 46.155 7.250 ;
        RECT 46.865 5.470 47.035 7.250 ;
        RECT 49.615 5.515 49.785 7.250 ;
        RECT 50.495 5.515 50.665 7.250 ;
        RECT 40.295 5.300 43.005 5.470 ;
        RECT 45.105 5.300 47.815 5.470 ;
        RECT 49.615 5.345 51.145 5.515 ;
        RECT 39.875 2.055 40.045 5.095 ;
        RECT 34.210 0.985 34.380 1.720 ;
        RECT 36.130 1.635 37.270 1.805 ;
        RECT 34.695 0.765 34.865 1.535 ;
        RECT 33.725 0.595 34.865 0.765 ;
        RECT 33.725 0.515 33.895 0.595 ;
        RECT 34.695 0.515 34.865 0.595 ;
        RECT 36.130 0.505 36.300 1.635 ;
        RECT 37.100 0.755 37.270 1.635 ;
        RECT 37.585 1.710 38.195 1.880 ;
        RECT 39.355 1.815 39.525 1.895 ;
        RECT 40.325 1.815 40.495 1.895 ;
        RECT 41.295 1.815 41.465 1.895 ;
        RECT 37.585 0.975 37.755 1.710 ;
        RECT 39.355 1.645 41.465 1.815 ;
        RECT 38.070 0.755 38.240 1.525 ;
        RECT 37.100 0.585 38.240 0.755 ;
        RECT 37.100 0.505 37.270 0.585 ;
        RECT 38.070 0.505 38.240 0.585 ;
        RECT 39.355 0.515 39.525 1.645 ;
        RECT 40.325 0.765 40.495 1.645 ;
        RECT 41.295 1.565 41.465 1.645 ;
        RECT 40.815 1.220 40.985 1.300 ;
        RECT 41.865 1.220 42.035 1.895 ;
        RECT 42.835 1.890 43.005 5.300 ;
        RECT 44.685 2.055 44.855 5.095 ;
        RECT 46.905 2.055 47.075 5.095 ;
        RECT 40.815 1.050 42.035 1.220 ;
        RECT 40.815 0.970 40.985 1.050 ;
        RECT 41.295 0.765 41.465 0.845 ;
        RECT 40.325 0.595 41.465 0.765 ;
        RECT 40.325 0.515 40.495 0.595 ;
        RECT 41.295 0.515 41.465 0.595 ;
        RECT 41.865 0.765 42.035 1.050 ;
        RECT 42.350 1.720 43.005 1.890 ;
        RECT 44.165 1.815 44.335 1.895 ;
        RECT 45.135 1.815 45.305 1.895 ;
        RECT 46.105 1.815 46.275 1.895 ;
        RECT 42.350 0.985 42.520 1.720 ;
        RECT 44.165 1.645 46.275 1.815 ;
        RECT 42.835 0.765 43.005 1.535 ;
        RECT 41.865 0.595 43.005 0.765 ;
        RECT 41.865 0.515 42.035 0.595 ;
        RECT 42.835 0.515 43.005 0.595 ;
        RECT 44.165 0.515 44.335 1.645 ;
        RECT 45.135 0.765 45.305 1.645 ;
        RECT 46.105 1.565 46.275 1.645 ;
        RECT 45.625 1.220 45.795 1.300 ;
        RECT 46.675 1.220 46.845 1.895 ;
        RECT 47.645 1.890 47.815 5.300 ;
        RECT 49.495 2.055 49.665 5.095 ;
        RECT 50.265 4.940 50.435 5.095 ;
        RECT 50.235 4.765 50.435 4.940 ;
        RECT 50.235 2.055 50.405 4.765 ;
        RECT 45.625 1.050 46.845 1.220 ;
        RECT 45.625 0.970 45.795 1.050 ;
        RECT 46.105 0.765 46.275 0.845 ;
        RECT 45.135 0.595 46.275 0.765 ;
        RECT 45.135 0.515 45.305 0.595 ;
        RECT 46.105 0.515 46.275 0.595 ;
        RECT 46.675 0.765 46.845 1.050 ;
        RECT 47.160 1.720 47.815 1.890 ;
        RECT 49.080 1.805 49.250 1.885 ;
        RECT 50.050 1.805 50.220 1.885 ;
        RECT 50.975 1.880 51.145 5.345 ;
        RECT 53.245 5.470 53.415 7.250 ;
        RECT 54.125 5.470 54.295 7.250 ;
        RECT 55.005 5.470 55.175 7.250 ;
        RECT 58.055 5.470 58.225 7.250 ;
        RECT 58.935 5.470 59.105 7.250 ;
        RECT 59.815 5.470 59.985 7.250 ;
        RECT 62.565 5.515 62.735 7.250 ;
        RECT 63.445 5.515 63.615 7.250 ;
        RECT 53.245 5.300 55.955 5.470 ;
        RECT 58.055 5.300 60.765 5.470 ;
        RECT 62.565 5.345 64.095 5.515 ;
        RECT 52.825 2.055 52.995 5.095 ;
        RECT 55.045 2.055 55.215 5.095 ;
        RECT 47.160 0.985 47.330 1.720 ;
        RECT 49.080 1.635 50.220 1.805 ;
        RECT 47.645 0.765 47.815 1.535 ;
        RECT 46.675 0.595 47.815 0.765 ;
        RECT 46.675 0.515 46.845 0.595 ;
        RECT 47.645 0.515 47.815 0.595 ;
        RECT 49.080 0.505 49.250 1.635 ;
        RECT 50.050 0.755 50.220 1.635 ;
        RECT 50.535 1.710 51.145 1.880 ;
        RECT 52.305 1.815 52.475 1.895 ;
        RECT 53.275 1.815 53.445 1.895 ;
        RECT 54.245 1.815 54.415 1.895 ;
        RECT 50.535 0.975 50.705 1.710 ;
        RECT 52.305 1.645 54.415 1.815 ;
        RECT 51.020 0.755 51.190 1.525 ;
        RECT 50.050 0.585 51.190 0.755 ;
        RECT 50.050 0.505 50.220 0.585 ;
        RECT 51.020 0.505 51.190 0.585 ;
        RECT 52.305 0.515 52.475 1.645 ;
        RECT 53.275 0.765 53.445 1.645 ;
        RECT 54.245 1.565 54.415 1.645 ;
        RECT 53.765 1.220 53.935 1.300 ;
        RECT 54.815 1.220 54.985 1.895 ;
        RECT 55.785 1.890 55.955 5.300 ;
        RECT 57.635 2.055 57.805 5.095 ;
        RECT 53.765 1.050 54.985 1.220 ;
        RECT 53.765 0.970 53.935 1.050 ;
        RECT 54.245 0.765 54.415 0.845 ;
        RECT 53.275 0.595 54.415 0.765 ;
        RECT 53.275 0.515 53.445 0.595 ;
        RECT 54.245 0.515 54.415 0.595 ;
        RECT 54.815 0.765 54.985 1.050 ;
        RECT 55.300 1.720 55.955 1.890 ;
        RECT 57.115 1.815 57.285 1.895 ;
        RECT 58.085 1.815 58.255 1.895 ;
        RECT 59.055 1.815 59.225 1.895 ;
        RECT 55.300 0.985 55.470 1.720 ;
        RECT 57.115 1.645 59.225 1.815 ;
        RECT 55.785 0.765 55.955 1.535 ;
        RECT 54.815 0.595 55.955 0.765 ;
        RECT 54.815 0.515 54.985 0.595 ;
        RECT 55.785 0.515 55.955 0.595 ;
        RECT 57.115 0.515 57.285 1.645 ;
        RECT 58.085 0.765 58.255 1.645 ;
        RECT 59.055 1.565 59.225 1.645 ;
        RECT 58.575 1.220 58.745 1.300 ;
        RECT 59.625 1.220 59.795 1.895 ;
        RECT 60.595 1.890 60.765 5.300 ;
        RECT 62.445 2.055 62.615 5.095 ;
        RECT 63.215 4.940 63.385 5.095 ;
        RECT 63.185 4.765 63.385 4.940 ;
        RECT 63.185 2.055 63.355 4.765 ;
        RECT 58.575 1.050 59.795 1.220 ;
        RECT 58.575 0.970 58.745 1.050 ;
        RECT 59.055 0.765 59.225 0.845 ;
        RECT 58.085 0.595 59.225 0.765 ;
        RECT 58.085 0.515 58.255 0.595 ;
        RECT 59.055 0.515 59.225 0.595 ;
        RECT 59.625 0.765 59.795 1.050 ;
        RECT 60.110 1.720 60.765 1.890 ;
        RECT 62.030 1.805 62.200 1.885 ;
        RECT 63.000 1.805 63.170 1.885 ;
        RECT 63.925 1.880 64.095 5.345 ;
        RECT 66.195 5.470 66.365 7.250 ;
        RECT 67.075 5.470 67.245 7.250 ;
        RECT 67.955 5.470 68.125 7.250 ;
        RECT 71.005 5.470 71.175 7.250 ;
        RECT 71.885 5.470 72.055 7.250 ;
        RECT 72.765 5.470 72.935 7.250 ;
        RECT 75.515 5.515 75.685 7.250 ;
        RECT 76.395 5.515 76.565 7.250 ;
        RECT 78.845 7.055 79.025 7.225 ;
        RECT 78.845 5.525 79.015 7.055 ;
        RECT 79.725 5.525 79.895 7.225 ;
        RECT 66.195 5.300 68.905 5.470 ;
        RECT 71.005 5.300 73.715 5.470 ;
        RECT 75.515 5.345 77.045 5.515 ;
        RECT 78.845 5.355 79.895 5.525 ;
        RECT 65.775 2.055 65.945 5.095 ;
        RECT 60.110 0.985 60.280 1.720 ;
        RECT 62.030 1.635 63.170 1.805 ;
        RECT 60.595 0.765 60.765 1.535 ;
        RECT 59.625 0.595 60.765 0.765 ;
        RECT 59.625 0.515 59.795 0.595 ;
        RECT 60.595 0.515 60.765 0.595 ;
        RECT 62.030 0.505 62.200 1.635 ;
        RECT 63.000 0.755 63.170 1.635 ;
        RECT 63.485 1.710 64.095 1.880 ;
        RECT 65.255 1.815 65.425 1.895 ;
        RECT 66.225 1.815 66.395 1.895 ;
        RECT 67.195 1.815 67.365 1.895 ;
        RECT 63.485 0.975 63.655 1.710 ;
        RECT 65.255 1.645 67.365 1.815 ;
        RECT 63.970 0.755 64.140 1.525 ;
        RECT 63.000 0.585 64.140 0.755 ;
        RECT 63.000 0.505 63.170 0.585 ;
        RECT 63.970 0.505 64.140 0.585 ;
        RECT 65.255 0.515 65.425 1.645 ;
        RECT 66.225 0.765 66.395 1.645 ;
        RECT 67.195 1.565 67.365 1.645 ;
        RECT 66.715 1.220 66.885 1.300 ;
        RECT 67.765 1.220 67.935 1.895 ;
        RECT 68.735 1.890 68.905 5.300 ;
        RECT 70.585 2.055 70.755 5.095 ;
        RECT 72.805 2.055 72.975 5.095 ;
        RECT 66.715 1.050 67.935 1.220 ;
        RECT 66.715 0.970 66.885 1.050 ;
        RECT 67.195 0.765 67.365 0.845 ;
        RECT 66.225 0.595 67.365 0.765 ;
        RECT 66.225 0.515 66.395 0.595 ;
        RECT 67.195 0.515 67.365 0.595 ;
        RECT 67.765 0.765 67.935 1.050 ;
        RECT 68.250 1.720 68.905 1.890 ;
        RECT 70.065 1.815 70.235 1.895 ;
        RECT 71.035 1.815 71.205 1.895 ;
        RECT 72.005 1.815 72.175 1.895 ;
        RECT 68.250 0.985 68.420 1.720 ;
        RECT 70.065 1.645 72.175 1.815 ;
        RECT 68.735 0.765 68.905 1.535 ;
        RECT 67.765 0.595 68.905 0.765 ;
        RECT 67.765 0.515 67.935 0.595 ;
        RECT 68.735 0.515 68.905 0.595 ;
        RECT 70.065 0.515 70.235 1.645 ;
        RECT 71.035 0.765 71.205 1.645 ;
        RECT 72.005 1.565 72.175 1.645 ;
        RECT 71.525 1.220 71.695 1.300 ;
        RECT 72.575 1.220 72.745 1.895 ;
        RECT 73.545 1.890 73.715 5.300 ;
        RECT 75.395 2.055 75.565 5.095 ;
        RECT 76.165 4.940 76.335 5.095 ;
        RECT 76.135 4.765 76.335 4.940 ;
        RECT 76.135 2.055 76.305 4.765 ;
        RECT 71.525 1.050 72.745 1.220 ;
        RECT 71.525 0.970 71.695 1.050 ;
        RECT 72.005 0.765 72.175 0.845 ;
        RECT 71.035 0.595 72.175 0.765 ;
        RECT 71.035 0.515 71.205 0.595 ;
        RECT 72.005 0.515 72.175 0.595 ;
        RECT 72.575 0.765 72.745 1.050 ;
        RECT 73.060 1.720 73.715 1.890 ;
        RECT 74.980 1.805 75.150 1.885 ;
        RECT 75.950 1.805 76.120 1.885 ;
        RECT 76.875 1.880 77.045 5.345 ;
        RECT 79.725 5.275 79.895 5.355 ;
        RECT 81.725 7.055 83.655 7.225 ;
        RECT 81.725 5.275 81.895 7.055 ;
        RECT 82.165 5.525 82.335 6.795 ;
        RECT 82.605 5.785 82.775 7.055 ;
        RECT 83.045 5.525 83.215 6.795 ;
        RECT 83.485 5.605 83.655 7.055 ;
        RECT 85.065 7.055 86.995 7.225 ;
        RECT 82.165 5.355 83.215 5.525 ;
        RECT 83.045 5.275 83.215 5.355 ;
        RECT 85.065 5.275 85.235 7.055 ;
        RECT 85.945 5.785 86.115 7.055 ;
        RECT 86.825 5.785 86.995 7.055 ;
        RECT 78.355 2.055 78.525 5.100 ;
        RECT 79.505 4.940 79.675 5.100 ;
        RECT 79.465 4.770 79.675 4.940 ;
        RECT 79.465 2.055 79.635 4.770 ;
        RECT 82.055 2.055 82.225 5.100 ;
        RECT 83.535 2.055 83.705 5.100 ;
        RECT 85.015 2.055 85.185 5.100 ;
        RECT 86.125 4.770 86.315 5.100 ;
        RECT 86.125 2.055 86.295 4.770 ;
        RECT 73.060 0.985 73.230 1.720 ;
        RECT 74.980 1.635 76.120 1.805 ;
        RECT 73.545 0.765 73.715 1.535 ;
        RECT 72.575 0.595 73.715 0.765 ;
        RECT 72.575 0.515 72.745 0.595 ;
        RECT 73.545 0.515 73.715 0.595 ;
        RECT 74.980 0.505 75.150 1.635 ;
        RECT 75.950 0.755 76.120 1.635 ;
        RECT 76.435 1.710 77.045 1.880 ;
        RECT 78.310 1.805 78.480 1.885 ;
        RECT 79.280 1.805 79.450 1.885 ;
        RECT 76.435 0.975 76.605 1.710 ;
        RECT 78.310 1.635 79.450 1.805 ;
        RECT 76.920 0.755 77.090 1.525 ;
        RECT 75.950 0.585 77.090 0.755 ;
        RECT 75.950 0.505 76.120 0.585 ;
        RECT 76.920 0.505 77.090 0.585 ;
        RECT 78.310 0.505 78.480 1.635 ;
        RECT 79.280 0.755 79.450 1.635 ;
        RECT 80.250 0.755 80.420 1.885 ;
        RECT 79.280 0.585 80.420 0.755 ;
        RECT 79.280 0.505 79.450 0.585 ;
        RECT 80.250 0.505 80.420 0.585 ;
        RECT 81.640 1.805 81.810 1.885 ;
        RECT 82.610 1.805 82.780 1.885 ;
        RECT 81.640 1.635 82.780 1.805 ;
        RECT 81.640 0.505 81.810 1.635 ;
        RECT 82.610 0.755 82.780 1.635 ;
        RECT 83.580 0.755 83.750 1.885 ;
        RECT 82.610 0.585 83.750 0.755 ;
        RECT 82.610 0.505 82.780 0.585 ;
        RECT 83.580 0.505 83.750 0.585 ;
        RECT 84.970 1.805 85.140 1.885 ;
        RECT 85.940 1.805 86.110 1.885 ;
        RECT 84.970 1.635 86.110 1.805 ;
        RECT 84.970 0.505 85.140 1.635 ;
        RECT 85.940 0.755 86.110 1.635 ;
        RECT 86.910 0.755 87.080 1.530 ;
        RECT 85.940 0.585 87.080 0.755 ;
        RECT 85.940 0.505 86.110 0.585 ;
        RECT 86.910 0.505 87.080 0.585 ;
      LAYER mcon ;
        RECT 1.025 4.355 1.195 4.525 ;
        RECT 3.245 3.615 3.415 3.785 ;
        RECT 3.985 3.985 4.155 4.155 ;
        RECT 5.835 3.985 6.005 4.155 ;
        RECT 8.795 3.615 8.965 3.785 ;
        RECT 10.645 3.615 10.815 3.785 ;
        RECT 11.385 4.355 11.555 4.525 ;
        RECT 12.125 3.615 12.295 3.785 ;
        RECT 13.975 3.615 14.145 3.785 ;
        RECT 16.935 4.355 17.105 4.525 ;
        RECT 18.785 3.985 18.955 4.155 ;
        RECT 21.005 2.875 21.175 3.045 ;
        RECT 21.745 3.985 21.915 4.155 ;
        RECT 23.595 3.985 23.765 4.155 ;
        RECT 24.335 4.355 24.505 4.525 ;
        RECT 25.075 2.875 25.245 3.045 ;
        RECT 26.925 4.355 27.095 4.525 ;
        RECT 29.145 3.615 29.315 3.785 ;
        RECT 29.885 3.985 30.055 4.155 ;
        RECT 31.735 3.985 31.905 4.155 ;
        RECT 34.695 3.615 34.865 3.785 ;
        RECT 36.545 3.615 36.715 3.785 ;
        RECT 37.285 4.355 37.455 4.525 ;
        RECT 38.025 3.615 38.195 3.785 ;
        RECT 39.875 3.615 40.045 3.785 ;
        RECT 42.835 4.355 43.005 4.525 ;
        RECT 44.685 3.985 44.855 4.155 ;
        RECT 46.905 3.245 47.075 3.415 ;
        RECT 47.645 3.985 47.815 4.155 ;
        RECT 49.495 3.985 49.665 4.155 ;
        RECT 50.235 4.355 50.405 4.525 ;
        RECT 50.975 3.245 51.145 3.415 ;
        RECT 52.825 4.355 52.995 4.525 ;
        RECT 55.045 3.615 55.215 3.785 ;
        RECT 55.785 3.985 55.955 4.155 ;
        RECT 57.635 3.985 57.805 4.155 ;
        RECT 60.595 3.615 60.765 3.785 ;
        RECT 62.445 3.615 62.615 3.785 ;
        RECT 63.185 4.355 63.355 4.525 ;
        RECT 79.725 5.355 79.895 5.525 ;
        RECT 63.925 3.615 64.095 3.785 ;
        RECT 65.775 3.615 65.945 3.785 ;
        RECT 68.735 4.355 68.905 4.525 ;
        RECT 70.585 3.985 70.755 4.155 ;
        RECT 72.805 3.615 72.975 3.785 ;
        RECT 73.545 3.985 73.715 4.155 ;
        RECT 75.395 3.985 75.565 4.155 ;
        RECT 76.135 4.355 76.305 4.525 ;
        RECT 81.725 5.355 81.895 5.525 ;
        RECT 83.045 5.355 83.215 5.525 ;
        RECT 85.065 5.355 85.235 5.525 ;
        RECT 76.875 3.615 77.045 3.785 ;
        RECT 78.355 4.725 78.525 4.895 ;
        RECT 78.355 3.245 78.525 3.415 ;
        RECT 79.465 4.355 79.635 4.525 ;
        RECT 79.465 3.615 79.635 3.785 ;
        RECT 82.055 4.725 82.225 4.895 ;
        RECT 83.535 2.875 83.705 3.045 ;
        RECT 83.535 2.135 83.705 2.305 ;
        RECT 85.015 2.135 85.185 2.305 ;
        RECT 86.125 4.355 86.295 4.525 ;
      LAYER met1 ;
        RECT 79.695 5.525 79.925 5.555 ;
        RECT 81.695 5.525 81.925 5.555 ;
        RECT 83.015 5.525 83.245 5.555 ;
        RECT 85.035 5.525 85.265 5.555 ;
        RECT 79.665 5.355 81.955 5.525 ;
        RECT 82.985 5.355 85.295 5.525 ;
        RECT 79.695 5.325 79.925 5.355 ;
        RECT 81.695 5.325 81.925 5.355 ;
        RECT 83.015 5.325 83.245 5.355 ;
        RECT 85.035 5.325 85.265 5.355 ;
        RECT 78.325 4.895 78.555 4.925 ;
        RECT 82.025 4.895 82.255 4.925 ;
        RECT 78.295 4.725 82.285 4.895 ;
        RECT 78.325 4.695 78.555 4.725 ;
        RECT 82.025 4.695 82.255 4.725 ;
        RECT 0.995 4.525 1.225 4.555 ;
        RECT 11.355 4.525 11.585 4.555 ;
        RECT 16.905 4.525 17.135 4.555 ;
        RECT 24.305 4.525 24.535 4.555 ;
        RECT 26.895 4.525 27.125 4.555 ;
        RECT 37.255 4.525 37.485 4.555 ;
        RECT 42.805 4.525 43.035 4.555 ;
        RECT 50.205 4.525 50.435 4.555 ;
        RECT 52.795 4.525 53.025 4.555 ;
        RECT 63.155 4.525 63.385 4.555 ;
        RECT 68.705 4.525 68.935 4.555 ;
        RECT 76.105 4.525 76.335 4.555 ;
        RECT 79.435 4.525 79.665 4.555 ;
        RECT 86.095 4.525 86.325 4.555 ;
        RECT 0.965 4.355 24.565 4.525 ;
        RECT 26.865 4.355 50.465 4.525 ;
        RECT 52.765 4.355 76.365 4.525 ;
        RECT 79.405 4.355 86.355 4.525 ;
        RECT 0.995 4.325 1.225 4.355 ;
        RECT 11.355 4.325 11.585 4.355 ;
        RECT 16.905 4.325 17.135 4.355 ;
        RECT 24.305 4.325 24.535 4.355 ;
        RECT 26.895 4.325 27.125 4.355 ;
        RECT 37.255 4.325 37.485 4.355 ;
        RECT 42.805 4.325 43.035 4.355 ;
        RECT 50.205 4.325 50.435 4.355 ;
        RECT 52.795 4.325 53.025 4.355 ;
        RECT 63.155 4.325 63.385 4.355 ;
        RECT 68.705 4.325 68.935 4.355 ;
        RECT 76.105 4.325 76.335 4.355 ;
        RECT 79.435 4.325 79.665 4.355 ;
        RECT 86.095 4.325 86.325 4.355 ;
        RECT 3.955 4.155 4.185 4.185 ;
        RECT 5.805 4.155 6.035 4.185 ;
        RECT 18.755 4.155 18.985 4.185 ;
        RECT 21.715 4.155 21.945 4.185 ;
        RECT 23.565 4.155 23.795 4.185 ;
        RECT 29.855 4.155 30.085 4.185 ;
        RECT 31.705 4.155 31.935 4.185 ;
        RECT 44.655 4.155 44.885 4.185 ;
        RECT 47.615 4.155 47.845 4.185 ;
        RECT 49.465 4.155 49.695 4.185 ;
        RECT 55.755 4.155 55.985 4.185 ;
        RECT 57.605 4.155 57.835 4.185 ;
        RECT 70.555 4.155 70.785 4.185 ;
        RECT 73.515 4.155 73.745 4.185 ;
        RECT 75.365 4.155 75.595 4.185 ;
        RECT 3.925 3.985 19.015 4.155 ;
        RECT 21.685 3.985 23.825 4.155 ;
        RECT 29.825 3.985 44.915 4.155 ;
        RECT 47.585 3.985 49.725 4.155 ;
        RECT 55.725 3.985 70.815 4.155 ;
        RECT 73.485 3.985 75.625 4.155 ;
        RECT 3.955 3.955 4.185 3.985 ;
        RECT 5.805 3.955 6.035 3.985 ;
        RECT 18.755 3.955 18.985 3.985 ;
        RECT 21.715 3.955 21.945 3.985 ;
        RECT 23.565 3.955 23.795 3.985 ;
        RECT 29.855 3.955 30.085 3.985 ;
        RECT 31.705 3.955 31.935 3.985 ;
        RECT 44.655 3.955 44.885 3.985 ;
        RECT 47.615 3.955 47.845 3.985 ;
        RECT 49.465 3.955 49.695 3.985 ;
        RECT 55.755 3.955 55.985 3.985 ;
        RECT 57.605 3.955 57.835 3.985 ;
        RECT 70.555 3.955 70.785 3.985 ;
        RECT 73.515 3.955 73.745 3.985 ;
        RECT 75.365 3.955 75.595 3.985 ;
        RECT 3.215 3.785 3.445 3.815 ;
        RECT 8.765 3.785 8.995 3.815 ;
        RECT 10.615 3.785 10.845 3.815 ;
        RECT 12.095 3.785 12.325 3.815 ;
        RECT 13.945 3.785 14.175 3.815 ;
        RECT 29.115 3.785 29.345 3.815 ;
        RECT 34.665 3.785 34.895 3.815 ;
        RECT 36.515 3.785 36.745 3.815 ;
        RECT 37.995 3.785 38.225 3.815 ;
        RECT 39.845 3.785 40.075 3.815 ;
        RECT 55.015 3.785 55.245 3.815 ;
        RECT 60.565 3.785 60.795 3.815 ;
        RECT 62.415 3.785 62.645 3.815 ;
        RECT 63.895 3.785 64.125 3.815 ;
        RECT 65.745 3.785 65.975 3.815 ;
        RECT 72.775 3.785 73.005 3.815 ;
        RECT 76.845 3.785 77.075 3.815 ;
        RECT 79.435 3.785 79.665 3.815 ;
        RECT 3.185 3.615 10.875 3.785 ;
        RECT 12.065 3.615 14.205 3.785 ;
        RECT 29.085 3.615 36.775 3.785 ;
        RECT 37.965 3.615 40.105 3.785 ;
        RECT 54.985 3.615 62.675 3.785 ;
        RECT 63.865 3.615 66.005 3.785 ;
        RECT 72.745 3.615 79.695 3.785 ;
        RECT 3.215 3.585 3.445 3.615 ;
        RECT 8.765 3.585 8.995 3.615 ;
        RECT 10.615 3.585 10.845 3.615 ;
        RECT 12.095 3.585 12.325 3.615 ;
        RECT 13.945 3.585 14.175 3.615 ;
        RECT 29.115 3.585 29.345 3.615 ;
        RECT 34.665 3.585 34.895 3.615 ;
        RECT 36.515 3.585 36.745 3.615 ;
        RECT 37.995 3.585 38.225 3.615 ;
        RECT 39.845 3.585 40.075 3.615 ;
        RECT 55.015 3.585 55.245 3.615 ;
        RECT 60.565 3.585 60.795 3.615 ;
        RECT 62.415 3.585 62.645 3.615 ;
        RECT 63.895 3.585 64.125 3.615 ;
        RECT 65.745 3.585 65.975 3.615 ;
        RECT 72.775 3.585 73.005 3.615 ;
        RECT 76.845 3.585 77.075 3.615 ;
        RECT 79.435 3.585 79.665 3.615 ;
        RECT 46.875 3.415 47.105 3.445 ;
        RECT 50.945 3.415 51.175 3.445 ;
        RECT 78.325 3.415 78.555 3.445 ;
        RECT 46.845 3.245 78.585 3.415 ;
        RECT 46.875 3.215 47.105 3.245 ;
        RECT 50.945 3.215 51.175 3.245 ;
        RECT 78.325 3.215 78.555 3.245 ;
        RECT 20.975 3.045 21.205 3.075 ;
        RECT 25.045 3.045 25.275 3.075 ;
        RECT 83.505 3.045 83.735 3.075 ;
        RECT 20.945 2.875 83.765 3.045 ;
        RECT 20.975 2.845 21.205 2.875 ;
        RECT 25.045 2.845 25.275 2.875 ;
        RECT 83.505 2.845 83.735 2.875 ;
        RECT 83.505 2.305 83.735 2.335 ;
        RECT 84.985 2.305 85.215 2.335 ;
        RECT 83.475 2.135 85.245 2.305 ;
        RECT 83.505 2.105 83.735 2.135 ;
        RECT 84.985 2.105 85.215 2.135 ;
  END
END TMRDFFRNQNX1






MACRO TMRDFFRNQX1
  CLASS BLOCK ;
  FOREIGN TMRDFFRNQX1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 90.750 BY 7.950 ;
  PIN Q
    ANTENNADIFFAREA 0.771900 ;
    PORT
      LAYER li1 ;
        RECT 88.715 4.895 88.885 7.250 ;
        RECT 88.715 4.725 89.255 4.895 ;
        RECT 89.085 2.305 89.255 4.725 ;
        RECT 88.715 2.135 89.255 2.305 ;
        RECT 88.715 0.975 88.885 2.135 ;
      LAYER mcon ;
        RECT 89.085 3.985 89.255 4.155 ;
      LAYER met1 ;
        RECT 89.055 4.155 89.285 4.185 ;
        RECT 89.025 3.985 89.435 4.155 ;
        RECT 89.055 3.955 89.285 3.985 ;
    END
  END Q
  PIN D
    ANTENNAGATEAREA 3.044550 ;
    PORT
      LAYER li1 ;
        RECT 6.945 2.055 7.115 5.095 ;
        RECT 32.845 2.055 33.015 5.095 ;
        RECT 58.745 2.055 58.915 5.095 ;
      LAYER mcon ;
        RECT 6.945 2.135 7.115 2.305 ;
        RECT 32.845 2.135 33.015 2.305 ;
        RECT 58.745 2.135 58.915 2.305 ;
      LAYER met1 ;
        RECT 6.915 2.305 7.145 2.335 ;
        RECT 32.815 2.305 33.045 2.335 ;
        RECT 58.715 2.305 58.945 2.335 ;
        RECT 6.885 2.135 59.095 2.305 ;
        RECT 6.915 2.105 7.145 2.135 ;
        RECT 32.815 2.105 33.045 2.135 ;
        RECT 58.715 2.105 58.945 2.135 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 6.089100 ;
    PORT
      LAYER li1 ;
        RECT 2.135 2.055 2.305 5.095 ;
        RECT 15.085 2.055 15.255 5.095 ;
        RECT 28.035 2.055 28.205 5.095 ;
        RECT 40.985 2.055 41.155 5.095 ;
        RECT 53.935 2.055 54.105 5.095 ;
        RECT 66.885 2.055 67.055 5.095 ;
      LAYER mcon ;
        RECT 2.135 4.725 2.305 4.895 ;
        RECT 15.085 4.725 15.255 4.895 ;
        RECT 28.035 4.725 28.205 4.895 ;
        RECT 40.985 4.725 41.155 4.895 ;
        RECT 53.935 4.725 54.105 4.895 ;
        RECT 66.885 4.725 67.055 4.895 ;
      LAYER met1 ;
        RECT 2.105 4.895 2.335 4.925 ;
        RECT 15.055 4.895 15.285 4.925 ;
        RECT 28.005 4.895 28.235 4.925 ;
        RECT 40.955 4.895 41.185 4.925 ;
        RECT 53.905 4.895 54.135 4.925 ;
        RECT 66.855 4.895 67.085 4.925 ;
        RECT 2.075 4.725 67.115 4.895 ;
        RECT 2.105 4.695 2.335 4.725 ;
        RECT 15.055 4.695 15.285 4.725 ;
        RECT 28.005 4.695 28.235 4.725 ;
        RECT 40.955 4.695 41.185 4.725 ;
        RECT 53.905 4.695 54.135 4.725 ;
        RECT 66.855 4.695 67.085 4.725 ;
    END
  END CLK
  PIN RN
    ANTENNAGATEAREA 9.208050 ;
    PORT
      LAYER li1 ;
        RECT 8.055 2.055 8.225 5.095 ;
        RECT 16.195 2.055 16.365 5.095 ;
        RECT 19.895 2.055 20.065 5.095 ;
        RECT 33.955 2.055 34.125 5.095 ;
        RECT 42.095 2.055 42.265 5.095 ;
        RECT 45.795 2.055 45.965 5.095 ;
        RECT 59.855 2.055 60.025 5.095 ;
        RECT 67.995 2.055 68.165 5.095 ;
        RECT 71.695 2.055 71.865 5.095 ;
      LAYER mcon ;
        RECT 8.055 2.505 8.225 2.675 ;
        RECT 16.195 2.505 16.365 2.675 ;
        RECT 19.895 2.505 20.065 2.675 ;
        RECT 33.955 2.505 34.125 2.675 ;
        RECT 42.095 2.505 42.265 2.675 ;
        RECT 45.795 2.505 45.965 2.675 ;
        RECT 59.855 2.505 60.025 2.675 ;
        RECT 67.995 2.505 68.165 2.675 ;
        RECT 71.695 2.505 71.865 2.675 ;
      LAYER met1 ;
        RECT 8.025 2.675 8.255 2.705 ;
        RECT 16.165 2.675 16.395 2.705 ;
        RECT 19.865 2.675 20.095 2.705 ;
        RECT 33.925 2.675 34.155 2.705 ;
        RECT 42.065 2.675 42.295 2.705 ;
        RECT 45.765 2.675 45.995 2.705 ;
        RECT 59.825 2.675 60.055 2.705 ;
        RECT 67.965 2.675 68.195 2.705 ;
        RECT 71.665 2.675 71.895 2.705 ;
        RECT 7.995 2.505 71.925 2.675 ;
        RECT 8.025 2.475 8.255 2.505 ;
        RECT 16.165 2.475 16.395 2.505 ;
        RECT 19.865 2.475 20.095 2.505 ;
        RECT 33.925 2.475 34.155 2.505 ;
        RECT 42.065 2.475 42.295 2.505 ;
        RECT 45.765 2.475 45.995 2.505 ;
        RECT 59.825 2.475 60.055 2.505 ;
        RECT 67.965 2.475 68.195 2.505 ;
        RECT 71.665 2.475 71.895 2.505 ;
    END
  END RN
  PIN VDD
    ANTENNADIFFAREA 103.784348 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 90.330 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 90.065 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 1.005 5.445 1.175 7.460 ;
        RECT 1.885 5.785 2.055 7.460 ;
        RECT 2.765 5.785 2.935 7.460 ;
        RECT 3.645 5.785 3.815 7.460 ;
        RECT 4.655 4.340 4.965 7.460 ;
        RECT 5.815 5.445 5.985 7.460 ;
        RECT 6.695 5.785 6.865 7.460 ;
        RECT 7.575 5.785 7.745 7.460 ;
        RECT 8.455 5.785 8.625 7.460 ;
        RECT 9.465 4.340 9.775 7.460 ;
        RECT 10.325 5.365 10.495 7.460 ;
        RECT 11.205 5.785 11.375 7.460 ;
        RECT 12.085 5.785 12.255 7.460 ;
        RECT 12.795 4.340 13.105 7.460 ;
        RECT 13.955 5.445 14.125 7.460 ;
        RECT 14.835 5.785 15.005 7.460 ;
        RECT 15.715 5.785 15.885 7.460 ;
        RECT 16.595 5.785 16.765 7.460 ;
        RECT 17.605 4.340 17.915 7.460 ;
        RECT 18.765 5.445 18.935 7.460 ;
        RECT 19.645 5.785 19.815 7.460 ;
        RECT 20.525 5.785 20.695 7.460 ;
        RECT 21.405 5.785 21.575 7.460 ;
        RECT 22.415 4.340 22.725 7.460 ;
        RECT 23.275 5.365 23.445 7.460 ;
        RECT 24.155 5.785 24.325 7.460 ;
        RECT 25.035 5.785 25.205 7.460 ;
        RECT 25.745 4.340 26.055 7.460 ;
        RECT 26.905 5.445 27.075 7.460 ;
        RECT 27.785 5.785 27.955 7.460 ;
        RECT 28.665 5.785 28.835 7.460 ;
        RECT 29.545 5.785 29.715 7.460 ;
        RECT 30.555 4.340 30.865 7.460 ;
        RECT 31.715 5.445 31.885 7.460 ;
        RECT 32.595 5.785 32.765 7.460 ;
        RECT 33.475 5.785 33.645 7.460 ;
        RECT 34.355 5.785 34.525 7.460 ;
        RECT 35.365 4.340 35.675 7.460 ;
        RECT 36.225 5.365 36.395 7.460 ;
        RECT 37.105 5.785 37.275 7.460 ;
        RECT 37.985 5.785 38.155 7.460 ;
        RECT 38.695 4.340 39.005 7.460 ;
        RECT 39.855 5.445 40.025 7.460 ;
        RECT 40.735 5.785 40.905 7.460 ;
        RECT 41.615 5.785 41.785 7.460 ;
        RECT 42.495 5.785 42.665 7.460 ;
        RECT 43.505 4.340 43.815 7.460 ;
        RECT 44.665 5.445 44.835 7.460 ;
        RECT 45.545 5.785 45.715 7.460 ;
        RECT 46.425 5.785 46.595 7.460 ;
        RECT 47.305 5.785 47.475 7.460 ;
        RECT 48.315 4.340 48.625 7.460 ;
        RECT 49.175 5.365 49.345 7.460 ;
        RECT 50.055 5.785 50.225 7.460 ;
        RECT 50.935 5.785 51.105 7.460 ;
        RECT 51.645 4.340 51.955 7.460 ;
        RECT 52.805 5.445 52.975 7.460 ;
        RECT 53.685 5.785 53.855 7.460 ;
        RECT 54.565 5.785 54.735 7.460 ;
        RECT 55.445 5.785 55.615 7.460 ;
        RECT 56.455 4.340 56.765 7.460 ;
        RECT 57.615 5.445 57.785 7.460 ;
        RECT 58.495 5.785 58.665 7.460 ;
        RECT 59.375 5.785 59.545 7.460 ;
        RECT 60.255 5.785 60.425 7.460 ;
        RECT 61.265 4.340 61.575 7.460 ;
        RECT 62.125 5.365 62.295 7.460 ;
        RECT 63.005 5.785 63.175 7.460 ;
        RECT 63.885 5.785 64.055 7.460 ;
        RECT 64.595 4.340 64.905 7.460 ;
        RECT 65.755 5.445 65.925 7.460 ;
        RECT 66.635 5.785 66.805 7.460 ;
        RECT 67.515 5.785 67.685 7.460 ;
        RECT 68.395 5.785 68.565 7.460 ;
        RECT 69.405 4.340 69.715 7.460 ;
        RECT 70.565 5.445 70.735 7.460 ;
        RECT 71.445 5.785 71.615 7.460 ;
        RECT 72.325 5.785 72.495 7.460 ;
        RECT 73.205 5.785 73.375 7.460 ;
        RECT 74.215 4.340 74.525 7.460 ;
        RECT 75.075 5.365 75.245 7.460 ;
        RECT 75.955 5.785 76.125 7.460 ;
        RECT 76.835 5.785 77.005 7.460 ;
        RECT 77.545 4.340 77.855 7.460 ;
        RECT 78.405 5.355 78.575 7.460 ;
        RECT 79.285 5.785 79.455 7.460 ;
        RECT 80.165 5.355 80.335 7.460 ;
        RECT 80.875 4.340 81.185 7.460 ;
        RECT 84.205 4.340 84.515 7.460 ;
        RECT 87.535 4.340 87.845 7.460 ;
        RECT 88.275 5.415 88.445 7.460 ;
        RECT 89.155 5.415 89.325 7.460 ;
        RECT 89.755 4.340 90.065 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 0.995 7.525 1.165 7.695 ;
        RECT 1.355 7.525 1.525 7.695 ;
        RECT 1.715 7.525 1.885 7.695 ;
        RECT 2.075 7.525 2.245 7.695 ;
        RECT 2.565 7.525 2.735 7.695 ;
        RECT 2.925 7.525 3.095 7.695 ;
        RECT 3.285 7.525 3.455 7.695 ;
        RECT 3.645 7.525 3.815 7.695 ;
        RECT 4.005 7.525 4.175 7.695 ;
        RECT 4.365 7.525 4.535 7.695 ;
        RECT 5.085 7.525 5.255 7.695 ;
        RECT 5.445 7.525 5.615 7.695 ;
        RECT 5.805 7.525 5.975 7.695 ;
        RECT 6.165 7.525 6.335 7.695 ;
        RECT 6.525 7.525 6.695 7.695 ;
        RECT 6.885 7.525 7.055 7.695 ;
        RECT 7.375 7.525 7.545 7.695 ;
        RECT 7.735 7.525 7.905 7.695 ;
        RECT 8.095 7.525 8.265 7.695 ;
        RECT 8.455 7.525 8.625 7.695 ;
        RECT 8.815 7.525 8.985 7.695 ;
        RECT 9.175 7.525 9.345 7.695 ;
        RECT 9.895 7.525 10.065 7.695 ;
        RECT 10.255 7.525 10.425 7.695 ;
        RECT 10.615 7.525 10.785 7.695 ;
        RECT 10.975 7.525 11.145 7.695 ;
        RECT 11.425 7.525 11.595 7.695 ;
        RECT 11.785 7.525 11.955 7.695 ;
        RECT 12.145 7.525 12.315 7.695 ;
        RECT 12.505 7.525 12.675 7.695 ;
        RECT 13.225 7.525 13.395 7.695 ;
        RECT 13.585 7.525 13.755 7.695 ;
        RECT 13.945 7.525 14.115 7.695 ;
        RECT 14.305 7.525 14.475 7.695 ;
        RECT 14.665 7.525 14.835 7.695 ;
        RECT 15.025 7.525 15.195 7.695 ;
        RECT 15.515 7.525 15.685 7.695 ;
        RECT 15.875 7.525 16.045 7.695 ;
        RECT 16.235 7.525 16.405 7.695 ;
        RECT 16.595 7.525 16.765 7.695 ;
        RECT 16.955 7.525 17.125 7.695 ;
        RECT 17.315 7.525 17.485 7.695 ;
        RECT 18.035 7.525 18.205 7.695 ;
        RECT 18.395 7.525 18.565 7.695 ;
        RECT 18.755 7.525 18.925 7.695 ;
        RECT 19.115 7.525 19.285 7.695 ;
        RECT 19.475 7.525 19.645 7.695 ;
        RECT 19.835 7.525 20.005 7.695 ;
        RECT 20.325 7.525 20.495 7.695 ;
        RECT 20.685 7.525 20.855 7.695 ;
        RECT 21.045 7.525 21.215 7.695 ;
        RECT 21.405 7.525 21.575 7.695 ;
        RECT 21.765 7.525 21.935 7.695 ;
        RECT 22.125 7.525 22.295 7.695 ;
        RECT 22.845 7.525 23.015 7.695 ;
        RECT 23.205 7.525 23.375 7.695 ;
        RECT 23.565 7.525 23.735 7.695 ;
        RECT 23.925 7.525 24.095 7.695 ;
        RECT 24.375 7.525 24.545 7.695 ;
        RECT 24.735 7.525 24.905 7.695 ;
        RECT 25.095 7.525 25.265 7.695 ;
        RECT 25.455 7.525 25.625 7.695 ;
        RECT 26.175 7.525 26.345 7.695 ;
        RECT 26.535 7.525 26.705 7.695 ;
        RECT 26.895 7.525 27.065 7.695 ;
        RECT 27.255 7.525 27.425 7.695 ;
        RECT 27.615 7.525 27.785 7.695 ;
        RECT 27.975 7.525 28.145 7.695 ;
        RECT 28.465 7.525 28.635 7.695 ;
        RECT 28.825 7.525 28.995 7.695 ;
        RECT 29.185 7.525 29.355 7.695 ;
        RECT 29.545 7.525 29.715 7.695 ;
        RECT 29.905 7.525 30.075 7.695 ;
        RECT 30.265 7.525 30.435 7.695 ;
        RECT 30.985 7.525 31.155 7.695 ;
        RECT 31.345 7.525 31.515 7.695 ;
        RECT 31.705 7.525 31.875 7.695 ;
        RECT 32.065 7.525 32.235 7.695 ;
        RECT 32.425 7.525 32.595 7.695 ;
        RECT 32.785 7.525 32.955 7.695 ;
        RECT 33.275 7.525 33.445 7.695 ;
        RECT 33.635 7.525 33.805 7.695 ;
        RECT 33.995 7.525 34.165 7.695 ;
        RECT 34.355 7.525 34.525 7.695 ;
        RECT 34.715 7.525 34.885 7.695 ;
        RECT 35.075 7.525 35.245 7.695 ;
        RECT 35.795 7.525 35.965 7.695 ;
        RECT 36.155 7.525 36.325 7.695 ;
        RECT 36.515 7.525 36.685 7.695 ;
        RECT 36.875 7.525 37.045 7.695 ;
        RECT 37.325 7.525 37.495 7.695 ;
        RECT 37.685 7.525 37.855 7.695 ;
        RECT 38.045 7.525 38.215 7.695 ;
        RECT 38.405 7.525 38.575 7.695 ;
        RECT 39.125 7.525 39.295 7.695 ;
        RECT 39.485 7.525 39.655 7.695 ;
        RECT 39.845 7.525 40.015 7.695 ;
        RECT 40.205 7.525 40.375 7.695 ;
        RECT 40.565 7.525 40.735 7.695 ;
        RECT 40.925 7.525 41.095 7.695 ;
        RECT 41.415 7.525 41.585 7.695 ;
        RECT 41.775 7.525 41.945 7.695 ;
        RECT 42.135 7.525 42.305 7.695 ;
        RECT 42.495 7.525 42.665 7.695 ;
        RECT 42.855 7.525 43.025 7.695 ;
        RECT 43.215 7.525 43.385 7.695 ;
        RECT 43.935 7.525 44.105 7.695 ;
        RECT 44.295 7.525 44.465 7.695 ;
        RECT 44.655 7.525 44.825 7.695 ;
        RECT 45.015 7.525 45.185 7.695 ;
        RECT 45.375 7.525 45.545 7.695 ;
        RECT 45.735 7.525 45.905 7.695 ;
        RECT 46.225 7.525 46.395 7.695 ;
        RECT 46.585 7.525 46.755 7.695 ;
        RECT 46.945 7.525 47.115 7.695 ;
        RECT 47.305 7.525 47.475 7.695 ;
        RECT 47.665 7.525 47.835 7.695 ;
        RECT 48.025 7.525 48.195 7.695 ;
        RECT 48.745 7.525 48.915 7.695 ;
        RECT 49.105 7.525 49.275 7.695 ;
        RECT 49.465 7.525 49.635 7.695 ;
        RECT 49.825 7.525 49.995 7.695 ;
        RECT 50.275 7.525 50.445 7.695 ;
        RECT 50.635 7.525 50.805 7.695 ;
        RECT 50.995 7.525 51.165 7.695 ;
        RECT 51.355 7.525 51.525 7.695 ;
        RECT 52.075 7.525 52.245 7.695 ;
        RECT 52.435 7.525 52.605 7.695 ;
        RECT 52.795 7.525 52.965 7.695 ;
        RECT 53.155 7.525 53.325 7.695 ;
        RECT 53.515 7.525 53.685 7.695 ;
        RECT 53.875 7.525 54.045 7.695 ;
        RECT 54.365 7.525 54.535 7.695 ;
        RECT 54.725 7.525 54.895 7.695 ;
        RECT 55.085 7.525 55.255 7.695 ;
        RECT 55.445 7.525 55.615 7.695 ;
        RECT 55.805 7.525 55.975 7.695 ;
        RECT 56.165 7.525 56.335 7.695 ;
        RECT 56.885 7.525 57.055 7.695 ;
        RECT 57.245 7.525 57.415 7.695 ;
        RECT 57.605 7.525 57.775 7.695 ;
        RECT 57.965 7.525 58.135 7.695 ;
        RECT 58.325 7.525 58.495 7.695 ;
        RECT 58.685 7.525 58.855 7.695 ;
        RECT 59.175 7.525 59.345 7.695 ;
        RECT 59.535 7.525 59.705 7.695 ;
        RECT 59.895 7.525 60.065 7.695 ;
        RECT 60.255 7.525 60.425 7.695 ;
        RECT 60.615 7.525 60.785 7.695 ;
        RECT 60.975 7.525 61.145 7.695 ;
        RECT 61.695 7.525 61.865 7.695 ;
        RECT 62.055 7.525 62.225 7.695 ;
        RECT 62.415 7.525 62.585 7.695 ;
        RECT 62.775 7.525 62.945 7.695 ;
        RECT 63.225 7.525 63.395 7.695 ;
        RECT 63.585 7.525 63.755 7.695 ;
        RECT 63.945 7.525 64.115 7.695 ;
        RECT 64.305 7.525 64.475 7.695 ;
        RECT 65.025 7.525 65.195 7.695 ;
        RECT 65.385 7.525 65.555 7.695 ;
        RECT 65.745 7.525 65.915 7.695 ;
        RECT 66.105 7.525 66.275 7.695 ;
        RECT 66.465 7.525 66.635 7.695 ;
        RECT 66.825 7.525 66.995 7.695 ;
        RECT 67.315 7.525 67.485 7.695 ;
        RECT 67.675 7.525 67.845 7.695 ;
        RECT 68.035 7.525 68.205 7.695 ;
        RECT 68.395 7.525 68.565 7.695 ;
        RECT 68.755 7.525 68.925 7.695 ;
        RECT 69.115 7.525 69.285 7.695 ;
        RECT 69.835 7.525 70.005 7.695 ;
        RECT 70.195 7.525 70.365 7.695 ;
        RECT 70.555 7.525 70.725 7.695 ;
        RECT 70.915 7.525 71.085 7.695 ;
        RECT 71.275 7.525 71.445 7.695 ;
        RECT 71.635 7.525 71.805 7.695 ;
        RECT 72.125 7.525 72.295 7.695 ;
        RECT 72.485 7.525 72.655 7.695 ;
        RECT 72.845 7.525 73.015 7.695 ;
        RECT 73.205 7.525 73.375 7.695 ;
        RECT 73.565 7.525 73.735 7.695 ;
        RECT 73.925 7.525 74.095 7.695 ;
        RECT 74.645 7.525 74.815 7.695 ;
        RECT 75.005 7.525 75.175 7.695 ;
        RECT 75.365 7.525 75.535 7.695 ;
        RECT 75.725 7.525 75.895 7.695 ;
        RECT 76.175 7.525 76.345 7.695 ;
        RECT 76.535 7.525 76.705 7.695 ;
        RECT 76.895 7.525 77.065 7.695 ;
        RECT 77.255 7.525 77.425 7.695 ;
        RECT 77.975 7.525 78.145 7.695 ;
        RECT 78.335 7.525 78.505 7.695 ;
        RECT 78.695 7.525 78.865 7.695 ;
        RECT 79.055 7.525 79.225 7.695 ;
        RECT 79.505 7.525 79.675 7.695 ;
        RECT 79.865 7.525 80.035 7.695 ;
        RECT 80.225 7.525 80.395 7.695 ;
        RECT 80.585 7.525 80.755 7.695 ;
        RECT 81.305 7.525 81.475 7.695 ;
        RECT 81.665 7.525 81.835 7.695 ;
        RECT 82.025 7.525 82.195 7.695 ;
        RECT 82.385 7.525 82.555 7.695 ;
        RECT 82.835 7.525 83.005 7.695 ;
        RECT 83.195 7.525 83.365 7.695 ;
        RECT 83.555 7.525 83.725 7.695 ;
        RECT 83.915 7.525 84.085 7.695 ;
        RECT 84.635 7.525 84.805 7.695 ;
        RECT 84.995 7.525 85.165 7.695 ;
        RECT 85.355 7.525 85.525 7.695 ;
        RECT 85.715 7.525 85.885 7.695 ;
        RECT 86.165 7.525 86.335 7.695 ;
        RECT 86.525 7.525 86.695 7.695 ;
        RECT 86.885 7.525 87.055 7.695 ;
        RECT 87.245 7.525 87.415 7.695 ;
        RECT 87.965 7.525 88.135 7.695 ;
        RECT 88.325 7.525 88.495 7.695 ;
        RECT 88.715 7.525 88.885 7.695 ;
        RECT 89.105 7.525 89.275 7.695 ;
        RECT 89.465 7.525 89.635 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 90.065 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 65.090500 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 90.195 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 4.525 -0.075 5.095 -0.065 ;
        RECT 9.335 -0.075 9.905 -0.065 ;
        RECT 12.665 -0.075 13.235 -0.065 ;
        RECT 17.475 -0.075 18.045 -0.065 ;
        RECT 22.285 -0.075 22.855 -0.065 ;
        RECT 25.615 -0.075 26.185 -0.065 ;
        RECT 30.425 -0.075 30.995 -0.065 ;
        RECT 35.235 -0.075 35.805 -0.065 ;
        RECT 38.565 -0.075 39.135 -0.065 ;
        RECT 43.375 -0.075 43.945 -0.065 ;
        RECT 48.185 -0.075 48.755 -0.065 ;
        RECT 51.515 -0.075 52.085 -0.065 ;
        RECT 56.325 -0.075 56.895 -0.065 ;
        RECT 61.135 -0.075 61.705 -0.065 ;
        RECT 64.465 -0.075 65.035 -0.065 ;
        RECT 69.275 -0.075 69.845 -0.065 ;
        RECT 74.085 -0.075 74.655 -0.065 ;
        RECT 77.415 -0.075 77.985 -0.065 ;
        RECT 80.745 -0.075 81.315 -0.065 ;
        RECT 84.075 -0.075 84.645 -0.065 ;
        RECT 87.405 -0.075 87.975 -0.065 ;
        RECT 89.625 -0.075 90.195 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 0.990 0.310 1.160 1.270 ;
        RECT 4.655 0.310 4.965 2.860 ;
        RECT 5.800 0.310 5.970 1.270 ;
        RECT 9.465 0.310 9.775 2.860 ;
        RECT 10.715 0.310 10.885 1.260 ;
        RECT 12.795 0.310 13.105 2.860 ;
        RECT 13.940 0.310 14.110 1.270 ;
        RECT 17.605 0.310 17.915 2.860 ;
        RECT 18.750 0.310 18.920 1.270 ;
        RECT 22.415 0.310 22.725 2.860 ;
        RECT 23.665 0.310 23.835 1.260 ;
        RECT 25.745 0.310 26.055 2.860 ;
        RECT 26.890 0.310 27.060 1.270 ;
        RECT 30.555 0.310 30.865 2.860 ;
        RECT 31.700 0.310 31.870 1.270 ;
        RECT 35.365 0.310 35.675 2.860 ;
        RECT 36.615 0.310 36.785 1.260 ;
        RECT 38.695 0.310 39.005 2.860 ;
        RECT 39.840 0.310 40.010 1.270 ;
        RECT 43.505 0.310 43.815 2.860 ;
        RECT 44.650 0.310 44.820 1.270 ;
        RECT 48.315 0.310 48.625 2.860 ;
        RECT 49.565 0.310 49.735 1.260 ;
        RECT 51.645 0.310 51.955 2.860 ;
        RECT 52.790 0.310 52.960 1.270 ;
        RECT 56.455 0.310 56.765 2.860 ;
        RECT 57.600 0.310 57.770 1.270 ;
        RECT 61.265 0.310 61.575 2.860 ;
        RECT 62.515 0.310 62.685 1.260 ;
        RECT 64.595 0.310 64.905 2.860 ;
        RECT 65.740 0.310 65.910 1.270 ;
        RECT 69.405 0.310 69.715 2.860 ;
        RECT 70.550 0.310 70.720 1.270 ;
        RECT 74.215 0.310 74.525 2.860 ;
        RECT 75.465 0.310 75.635 1.260 ;
        RECT 77.545 0.310 77.855 2.860 ;
        RECT 78.795 0.310 78.965 1.260 ;
        RECT 80.875 0.310 81.185 2.860 ;
        RECT 82.125 0.310 82.295 1.260 ;
        RECT 84.205 0.310 84.515 2.860 ;
        RECT 85.455 0.310 85.625 1.260 ;
        RECT 87.535 0.310 87.845 2.860 ;
        RECT 88.235 0.755 88.405 1.885 ;
        RECT 89.205 0.755 89.375 1.885 ;
        RECT 88.235 0.585 89.375 0.755 ;
        RECT 88.235 0.310 88.405 0.585 ;
        RECT 88.720 0.310 88.890 0.585 ;
        RECT 89.205 0.310 89.375 0.585 ;
        RECT 89.755 0.310 90.065 2.860 ;
        RECT -0.155 0.235 83.095 0.310 ;
        RECT 83.265 0.235 90.065 0.310 ;
        RECT -0.155 0.000 90.065 0.235 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 0.995 0.065 1.165 0.235 ;
        RECT 1.355 0.065 1.525 0.235 ;
        RECT 1.715 0.065 1.885 0.235 ;
        RECT 2.075 0.065 2.245 0.235 ;
        RECT 2.565 0.065 2.735 0.235 ;
        RECT 2.925 0.065 3.095 0.235 ;
        RECT 3.285 0.065 3.455 0.235 ;
        RECT 3.645 0.065 3.815 0.235 ;
        RECT 4.005 0.065 4.175 0.235 ;
        RECT 4.365 0.065 4.535 0.235 ;
        RECT 5.085 0.065 5.255 0.235 ;
        RECT 5.445 0.065 5.615 0.235 ;
        RECT 5.805 0.065 5.975 0.235 ;
        RECT 6.165 0.065 6.335 0.235 ;
        RECT 6.525 0.065 6.695 0.235 ;
        RECT 6.885 0.065 7.055 0.235 ;
        RECT 7.375 0.065 7.545 0.235 ;
        RECT 7.735 0.065 7.905 0.235 ;
        RECT 8.095 0.065 8.265 0.235 ;
        RECT 8.455 0.065 8.625 0.235 ;
        RECT 8.815 0.065 8.985 0.235 ;
        RECT 9.175 0.065 9.345 0.235 ;
        RECT 9.895 0.065 10.065 0.235 ;
        RECT 10.255 0.065 10.425 0.235 ;
        RECT 10.615 0.065 10.785 0.235 ;
        RECT 10.975 0.065 11.145 0.235 ;
        RECT 11.425 0.065 11.595 0.235 ;
        RECT 11.785 0.065 11.955 0.235 ;
        RECT 12.145 0.065 12.315 0.235 ;
        RECT 12.505 0.065 12.675 0.235 ;
        RECT 13.225 0.065 13.395 0.235 ;
        RECT 13.585 0.065 13.755 0.235 ;
        RECT 13.945 0.065 14.115 0.235 ;
        RECT 14.305 0.065 14.475 0.235 ;
        RECT 14.665 0.065 14.835 0.235 ;
        RECT 15.025 0.065 15.195 0.235 ;
        RECT 15.515 0.065 15.685 0.235 ;
        RECT 15.875 0.065 16.045 0.235 ;
        RECT 16.235 0.065 16.405 0.235 ;
        RECT 16.595 0.065 16.765 0.235 ;
        RECT 16.955 0.065 17.125 0.235 ;
        RECT 17.315 0.065 17.485 0.235 ;
        RECT 18.035 0.065 18.205 0.235 ;
        RECT 18.395 0.065 18.565 0.235 ;
        RECT 18.755 0.065 18.925 0.235 ;
        RECT 19.115 0.065 19.285 0.235 ;
        RECT 19.475 0.065 19.645 0.235 ;
        RECT 19.835 0.065 20.005 0.235 ;
        RECT 20.325 0.065 20.495 0.235 ;
        RECT 20.685 0.065 20.855 0.235 ;
        RECT 21.045 0.065 21.215 0.235 ;
        RECT 21.405 0.065 21.575 0.235 ;
        RECT 21.765 0.065 21.935 0.235 ;
        RECT 22.125 0.065 22.295 0.235 ;
        RECT 22.845 0.065 23.015 0.235 ;
        RECT 23.205 0.065 23.375 0.235 ;
        RECT 23.565 0.065 23.735 0.235 ;
        RECT 23.925 0.065 24.095 0.235 ;
        RECT 24.375 0.065 24.545 0.235 ;
        RECT 24.735 0.065 24.905 0.235 ;
        RECT 25.095 0.065 25.265 0.235 ;
        RECT 25.455 0.065 25.625 0.235 ;
        RECT 26.175 0.065 26.345 0.235 ;
        RECT 26.535 0.065 26.705 0.235 ;
        RECT 26.895 0.065 27.065 0.235 ;
        RECT 27.255 0.065 27.425 0.235 ;
        RECT 27.615 0.065 27.785 0.235 ;
        RECT 27.975 0.065 28.145 0.235 ;
        RECT 28.465 0.065 28.635 0.235 ;
        RECT 28.825 0.065 28.995 0.235 ;
        RECT 29.185 0.065 29.355 0.235 ;
        RECT 29.545 0.065 29.715 0.235 ;
        RECT 29.905 0.065 30.075 0.235 ;
        RECT 30.265 0.065 30.435 0.235 ;
        RECT 30.985 0.065 31.155 0.235 ;
        RECT 31.345 0.065 31.515 0.235 ;
        RECT 31.705 0.065 31.875 0.235 ;
        RECT 32.065 0.065 32.235 0.235 ;
        RECT 32.425 0.065 32.595 0.235 ;
        RECT 32.785 0.065 32.955 0.235 ;
        RECT 33.275 0.065 33.445 0.235 ;
        RECT 33.635 0.065 33.805 0.235 ;
        RECT 33.995 0.065 34.165 0.235 ;
        RECT 34.355 0.065 34.525 0.235 ;
        RECT 34.715 0.065 34.885 0.235 ;
        RECT 35.075 0.065 35.245 0.235 ;
        RECT 35.795 0.065 35.965 0.235 ;
        RECT 36.155 0.065 36.325 0.235 ;
        RECT 36.515 0.065 36.685 0.235 ;
        RECT 36.875 0.065 37.045 0.235 ;
        RECT 37.325 0.065 37.495 0.235 ;
        RECT 37.685 0.065 37.855 0.235 ;
        RECT 38.045 0.065 38.215 0.235 ;
        RECT 38.405 0.065 38.575 0.235 ;
        RECT 39.125 0.065 39.295 0.235 ;
        RECT 39.485 0.065 39.655 0.235 ;
        RECT 39.845 0.065 40.015 0.235 ;
        RECT 40.205 0.065 40.375 0.235 ;
        RECT 40.565 0.065 40.735 0.235 ;
        RECT 40.925 0.065 41.095 0.235 ;
        RECT 41.415 0.065 41.585 0.235 ;
        RECT 41.775 0.065 41.945 0.235 ;
        RECT 42.135 0.065 42.305 0.235 ;
        RECT 42.495 0.065 42.665 0.235 ;
        RECT 42.855 0.065 43.025 0.235 ;
        RECT 43.215 0.065 43.385 0.235 ;
        RECT 43.935 0.065 44.105 0.235 ;
        RECT 44.295 0.065 44.465 0.235 ;
        RECT 44.655 0.065 44.825 0.235 ;
        RECT 45.015 0.065 45.185 0.235 ;
        RECT 45.375 0.065 45.545 0.235 ;
        RECT 45.735 0.065 45.905 0.235 ;
        RECT 46.225 0.065 46.395 0.235 ;
        RECT 46.585 0.065 46.755 0.235 ;
        RECT 46.945 0.065 47.115 0.235 ;
        RECT 47.305 0.065 47.475 0.235 ;
        RECT 47.665 0.065 47.835 0.235 ;
        RECT 48.025 0.065 48.195 0.235 ;
        RECT 48.745 0.065 48.915 0.235 ;
        RECT 49.105 0.065 49.275 0.235 ;
        RECT 49.465 0.065 49.635 0.235 ;
        RECT 49.825 0.065 49.995 0.235 ;
        RECT 50.275 0.065 50.445 0.235 ;
        RECT 50.635 0.065 50.805 0.235 ;
        RECT 50.995 0.065 51.165 0.235 ;
        RECT 51.355 0.065 51.525 0.235 ;
        RECT 52.075 0.065 52.245 0.235 ;
        RECT 52.435 0.065 52.605 0.235 ;
        RECT 52.795 0.065 52.965 0.235 ;
        RECT 53.155 0.065 53.325 0.235 ;
        RECT 53.515 0.065 53.685 0.235 ;
        RECT 53.875 0.065 54.045 0.235 ;
        RECT 54.365 0.065 54.535 0.235 ;
        RECT 54.725 0.065 54.895 0.235 ;
        RECT 55.085 0.065 55.255 0.235 ;
        RECT 55.445 0.065 55.615 0.235 ;
        RECT 55.805 0.065 55.975 0.235 ;
        RECT 56.165 0.065 56.335 0.235 ;
        RECT 56.885 0.065 57.055 0.235 ;
        RECT 57.245 0.065 57.415 0.235 ;
        RECT 57.605 0.065 57.775 0.235 ;
        RECT 57.965 0.065 58.135 0.235 ;
        RECT 58.325 0.065 58.495 0.235 ;
        RECT 58.685 0.065 58.855 0.235 ;
        RECT 59.175 0.065 59.345 0.235 ;
        RECT 59.535 0.065 59.705 0.235 ;
        RECT 59.895 0.065 60.065 0.235 ;
        RECT 60.255 0.065 60.425 0.235 ;
        RECT 60.615 0.065 60.785 0.235 ;
        RECT 60.975 0.065 61.145 0.235 ;
        RECT 61.695 0.065 61.865 0.235 ;
        RECT 62.055 0.065 62.225 0.235 ;
        RECT 62.415 0.065 62.585 0.235 ;
        RECT 62.775 0.065 62.945 0.235 ;
        RECT 63.225 0.065 63.395 0.235 ;
        RECT 63.585 0.065 63.755 0.235 ;
        RECT 63.945 0.065 64.115 0.235 ;
        RECT 64.305 0.065 64.475 0.235 ;
        RECT 65.025 0.065 65.195 0.235 ;
        RECT 65.385 0.065 65.555 0.235 ;
        RECT 65.745 0.065 65.915 0.235 ;
        RECT 66.105 0.065 66.275 0.235 ;
        RECT 66.465 0.065 66.635 0.235 ;
        RECT 66.825 0.065 66.995 0.235 ;
        RECT 67.315 0.065 67.485 0.235 ;
        RECT 67.675 0.065 67.845 0.235 ;
        RECT 68.035 0.065 68.205 0.235 ;
        RECT 68.395 0.065 68.565 0.235 ;
        RECT 68.755 0.065 68.925 0.235 ;
        RECT 69.115 0.065 69.285 0.235 ;
        RECT 69.835 0.065 70.005 0.235 ;
        RECT 70.195 0.065 70.365 0.235 ;
        RECT 70.555 0.065 70.725 0.235 ;
        RECT 70.915 0.065 71.085 0.235 ;
        RECT 71.275 0.065 71.445 0.235 ;
        RECT 71.635 0.065 71.805 0.235 ;
        RECT 72.125 0.065 72.295 0.235 ;
        RECT 72.485 0.065 72.655 0.235 ;
        RECT 72.845 0.065 73.015 0.235 ;
        RECT 73.205 0.065 73.375 0.235 ;
        RECT 73.565 0.065 73.735 0.235 ;
        RECT 73.925 0.065 74.095 0.235 ;
        RECT 74.645 0.065 74.815 0.235 ;
        RECT 75.005 0.065 75.175 0.235 ;
        RECT 75.365 0.065 75.535 0.235 ;
        RECT 75.725 0.065 75.895 0.235 ;
        RECT 76.175 0.065 76.345 0.235 ;
        RECT 76.535 0.065 76.705 0.235 ;
        RECT 76.895 0.065 77.065 0.235 ;
        RECT 77.255 0.065 77.425 0.235 ;
        RECT 77.975 0.065 78.145 0.235 ;
        RECT 78.335 0.065 78.505 0.235 ;
        RECT 78.695 0.065 78.865 0.235 ;
        RECT 79.055 0.065 79.225 0.235 ;
        RECT 79.505 0.065 79.675 0.235 ;
        RECT 79.865 0.065 80.035 0.235 ;
        RECT 80.225 0.065 80.395 0.235 ;
        RECT 80.585 0.065 80.755 0.235 ;
        RECT 81.305 0.065 81.475 0.235 ;
        RECT 81.665 0.065 81.835 0.235 ;
        RECT 82.025 0.065 82.195 0.235 ;
        RECT 82.385 0.065 82.555 0.235 ;
        RECT 82.835 0.065 83.005 0.235 ;
        RECT 83.195 0.065 83.365 0.235 ;
        RECT 83.555 0.065 83.725 0.235 ;
        RECT 83.915 0.065 84.085 0.235 ;
        RECT 84.635 0.065 84.805 0.235 ;
        RECT 84.995 0.065 85.165 0.235 ;
        RECT 85.355 0.065 85.525 0.235 ;
        RECT 85.715 0.065 85.885 0.235 ;
        RECT 86.165 0.065 86.335 0.235 ;
        RECT 86.525 0.065 86.695 0.235 ;
        RECT 86.885 0.065 87.055 0.235 ;
        RECT 87.245 0.065 87.415 0.235 ;
        RECT 87.965 0.065 88.135 0.235 ;
        RECT 88.325 0.065 88.495 0.235 ;
        RECT 88.715 0.065 88.885 0.235 ;
        RECT 89.105 0.065 89.275 0.235 ;
        RECT 89.465 0.065 89.635 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 90.065 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 1.445 5.470 1.615 7.250 ;
        RECT 2.325 5.470 2.495 7.250 ;
        RECT 3.205 5.470 3.375 7.250 ;
        RECT 6.255 5.470 6.425 7.250 ;
        RECT 7.135 5.470 7.305 7.250 ;
        RECT 8.015 5.470 8.185 7.250 ;
        RECT 10.765 5.515 10.935 7.250 ;
        RECT 11.645 5.515 11.815 7.250 ;
        RECT 1.445 5.300 4.155 5.470 ;
        RECT 6.255 5.300 8.965 5.470 ;
        RECT 10.765 5.345 12.295 5.515 ;
        RECT 1.025 2.055 1.195 5.095 ;
        RECT 3.245 2.055 3.415 5.095 ;
        RECT 0.505 1.815 0.675 1.895 ;
        RECT 1.475 1.815 1.645 1.895 ;
        RECT 2.445 1.815 2.615 1.895 ;
        RECT 0.505 1.645 2.615 1.815 ;
        RECT 0.505 0.515 0.675 1.645 ;
        RECT 1.475 0.765 1.645 1.645 ;
        RECT 2.445 1.565 2.615 1.645 ;
        RECT 1.965 1.220 2.135 1.300 ;
        RECT 3.015 1.220 3.185 1.895 ;
        RECT 3.985 1.890 4.155 5.300 ;
        RECT 5.835 2.055 6.005 5.095 ;
        RECT 1.965 1.050 3.185 1.220 ;
        RECT 1.965 0.970 2.135 1.050 ;
        RECT 2.445 0.765 2.615 0.845 ;
        RECT 1.475 0.595 2.615 0.765 ;
        RECT 1.475 0.515 1.645 0.595 ;
        RECT 2.445 0.515 2.615 0.595 ;
        RECT 3.015 0.765 3.185 1.050 ;
        RECT 3.500 1.720 4.155 1.890 ;
        RECT 5.315 1.815 5.485 1.895 ;
        RECT 6.285 1.815 6.455 1.895 ;
        RECT 7.255 1.815 7.425 1.895 ;
        RECT 3.500 0.985 3.670 1.720 ;
        RECT 5.315 1.645 7.425 1.815 ;
        RECT 3.985 0.765 4.155 1.535 ;
        RECT 3.015 0.595 4.155 0.765 ;
        RECT 3.015 0.515 3.185 0.595 ;
        RECT 3.985 0.515 4.155 0.595 ;
        RECT 5.315 0.515 5.485 1.645 ;
        RECT 6.285 0.765 6.455 1.645 ;
        RECT 7.255 1.565 7.425 1.645 ;
        RECT 6.775 1.220 6.945 1.300 ;
        RECT 7.825 1.220 7.995 1.895 ;
        RECT 8.795 1.890 8.965 5.300 ;
        RECT 10.645 2.055 10.815 5.095 ;
        RECT 11.415 4.940 11.585 5.095 ;
        RECT 11.385 4.765 11.585 4.940 ;
        RECT 11.385 2.055 11.555 4.765 ;
        RECT 6.775 1.050 7.995 1.220 ;
        RECT 6.775 0.970 6.945 1.050 ;
        RECT 7.255 0.765 7.425 0.845 ;
        RECT 6.285 0.595 7.425 0.765 ;
        RECT 6.285 0.515 6.455 0.595 ;
        RECT 7.255 0.515 7.425 0.595 ;
        RECT 7.825 0.765 7.995 1.050 ;
        RECT 8.310 1.720 8.965 1.890 ;
        RECT 10.230 1.805 10.400 1.885 ;
        RECT 11.200 1.805 11.370 1.885 ;
        RECT 12.125 1.880 12.295 5.345 ;
        RECT 14.395 5.470 14.565 7.250 ;
        RECT 15.275 5.470 15.445 7.250 ;
        RECT 16.155 5.470 16.325 7.250 ;
        RECT 19.205 5.470 19.375 7.250 ;
        RECT 20.085 5.470 20.255 7.250 ;
        RECT 20.965 5.470 21.135 7.250 ;
        RECT 23.715 5.515 23.885 7.250 ;
        RECT 24.595 5.515 24.765 7.250 ;
        RECT 14.395 5.300 17.105 5.470 ;
        RECT 19.205 5.300 21.915 5.470 ;
        RECT 23.715 5.345 25.245 5.515 ;
        RECT 13.975 2.055 14.145 5.095 ;
        RECT 8.310 0.985 8.480 1.720 ;
        RECT 10.230 1.635 11.370 1.805 ;
        RECT 8.795 0.765 8.965 1.535 ;
        RECT 7.825 0.595 8.965 0.765 ;
        RECT 7.825 0.515 7.995 0.595 ;
        RECT 8.795 0.515 8.965 0.595 ;
        RECT 10.230 0.505 10.400 1.635 ;
        RECT 11.200 0.755 11.370 1.635 ;
        RECT 11.685 1.710 12.295 1.880 ;
        RECT 13.455 1.815 13.625 1.895 ;
        RECT 14.425 1.815 14.595 1.895 ;
        RECT 15.395 1.815 15.565 1.895 ;
        RECT 11.685 0.975 11.855 1.710 ;
        RECT 13.455 1.645 15.565 1.815 ;
        RECT 12.170 0.755 12.340 1.525 ;
        RECT 11.200 0.585 12.340 0.755 ;
        RECT 11.200 0.505 11.370 0.585 ;
        RECT 12.170 0.505 12.340 0.585 ;
        RECT 13.455 0.515 13.625 1.645 ;
        RECT 14.425 0.765 14.595 1.645 ;
        RECT 15.395 1.565 15.565 1.645 ;
        RECT 14.915 1.220 15.085 1.300 ;
        RECT 15.965 1.220 16.135 1.895 ;
        RECT 16.935 1.890 17.105 5.300 ;
        RECT 18.785 2.055 18.955 5.095 ;
        RECT 21.005 2.055 21.175 5.095 ;
        RECT 14.915 1.050 16.135 1.220 ;
        RECT 14.915 0.970 15.085 1.050 ;
        RECT 15.395 0.765 15.565 0.845 ;
        RECT 14.425 0.595 15.565 0.765 ;
        RECT 14.425 0.515 14.595 0.595 ;
        RECT 15.395 0.515 15.565 0.595 ;
        RECT 15.965 0.765 16.135 1.050 ;
        RECT 16.450 1.720 17.105 1.890 ;
        RECT 18.265 1.815 18.435 1.895 ;
        RECT 19.235 1.815 19.405 1.895 ;
        RECT 20.205 1.815 20.375 1.895 ;
        RECT 16.450 0.985 16.620 1.720 ;
        RECT 18.265 1.645 20.375 1.815 ;
        RECT 16.935 0.765 17.105 1.535 ;
        RECT 15.965 0.595 17.105 0.765 ;
        RECT 15.965 0.515 16.135 0.595 ;
        RECT 16.935 0.515 17.105 0.595 ;
        RECT 18.265 0.515 18.435 1.645 ;
        RECT 19.235 0.765 19.405 1.645 ;
        RECT 20.205 1.565 20.375 1.645 ;
        RECT 19.725 1.220 19.895 1.300 ;
        RECT 20.775 1.220 20.945 1.895 ;
        RECT 21.745 1.890 21.915 5.300 ;
        RECT 23.595 2.055 23.765 5.095 ;
        RECT 24.365 4.940 24.535 5.095 ;
        RECT 24.335 4.765 24.535 4.940 ;
        RECT 24.335 2.055 24.505 4.765 ;
        RECT 19.725 1.050 20.945 1.220 ;
        RECT 19.725 0.970 19.895 1.050 ;
        RECT 20.205 0.765 20.375 0.845 ;
        RECT 19.235 0.595 20.375 0.765 ;
        RECT 19.235 0.515 19.405 0.595 ;
        RECT 20.205 0.515 20.375 0.595 ;
        RECT 20.775 0.765 20.945 1.050 ;
        RECT 21.260 1.720 21.915 1.890 ;
        RECT 23.180 1.805 23.350 1.885 ;
        RECT 24.150 1.805 24.320 1.885 ;
        RECT 25.075 1.880 25.245 5.345 ;
        RECT 27.345 5.470 27.515 7.250 ;
        RECT 28.225 5.470 28.395 7.250 ;
        RECT 29.105 5.470 29.275 7.250 ;
        RECT 32.155 5.470 32.325 7.250 ;
        RECT 33.035 5.470 33.205 7.250 ;
        RECT 33.915 5.470 34.085 7.250 ;
        RECT 36.665 5.515 36.835 7.250 ;
        RECT 37.545 5.515 37.715 7.250 ;
        RECT 27.345 5.300 30.055 5.470 ;
        RECT 32.155 5.300 34.865 5.470 ;
        RECT 36.665 5.345 38.195 5.515 ;
        RECT 26.925 2.055 27.095 5.095 ;
        RECT 29.145 2.055 29.315 5.095 ;
        RECT 21.260 0.985 21.430 1.720 ;
        RECT 23.180 1.635 24.320 1.805 ;
        RECT 21.745 0.765 21.915 1.535 ;
        RECT 20.775 0.595 21.915 0.765 ;
        RECT 20.775 0.515 20.945 0.595 ;
        RECT 21.745 0.515 21.915 0.595 ;
        RECT 23.180 0.505 23.350 1.635 ;
        RECT 24.150 0.755 24.320 1.635 ;
        RECT 24.635 1.710 25.245 1.880 ;
        RECT 26.405 1.815 26.575 1.895 ;
        RECT 27.375 1.815 27.545 1.895 ;
        RECT 28.345 1.815 28.515 1.895 ;
        RECT 24.635 0.975 24.805 1.710 ;
        RECT 26.405 1.645 28.515 1.815 ;
        RECT 25.120 0.755 25.290 1.525 ;
        RECT 24.150 0.585 25.290 0.755 ;
        RECT 24.150 0.505 24.320 0.585 ;
        RECT 25.120 0.505 25.290 0.585 ;
        RECT 26.405 0.515 26.575 1.645 ;
        RECT 27.375 0.765 27.545 1.645 ;
        RECT 28.345 1.565 28.515 1.645 ;
        RECT 27.865 1.220 28.035 1.300 ;
        RECT 28.915 1.220 29.085 1.895 ;
        RECT 29.885 1.890 30.055 5.300 ;
        RECT 31.735 2.055 31.905 5.095 ;
        RECT 27.865 1.050 29.085 1.220 ;
        RECT 27.865 0.970 28.035 1.050 ;
        RECT 28.345 0.765 28.515 0.845 ;
        RECT 27.375 0.595 28.515 0.765 ;
        RECT 27.375 0.515 27.545 0.595 ;
        RECT 28.345 0.515 28.515 0.595 ;
        RECT 28.915 0.765 29.085 1.050 ;
        RECT 29.400 1.720 30.055 1.890 ;
        RECT 31.215 1.815 31.385 1.895 ;
        RECT 32.185 1.815 32.355 1.895 ;
        RECT 33.155 1.815 33.325 1.895 ;
        RECT 29.400 0.985 29.570 1.720 ;
        RECT 31.215 1.645 33.325 1.815 ;
        RECT 29.885 0.765 30.055 1.535 ;
        RECT 28.915 0.595 30.055 0.765 ;
        RECT 28.915 0.515 29.085 0.595 ;
        RECT 29.885 0.515 30.055 0.595 ;
        RECT 31.215 0.515 31.385 1.645 ;
        RECT 32.185 0.765 32.355 1.645 ;
        RECT 33.155 1.565 33.325 1.645 ;
        RECT 32.675 1.220 32.845 1.300 ;
        RECT 33.725 1.220 33.895 1.895 ;
        RECT 34.695 1.890 34.865 5.300 ;
        RECT 36.545 2.055 36.715 5.095 ;
        RECT 37.315 4.940 37.485 5.095 ;
        RECT 37.285 4.765 37.485 4.940 ;
        RECT 37.285 2.055 37.455 4.765 ;
        RECT 32.675 1.050 33.895 1.220 ;
        RECT 32.675 0.970 32.845 1.050 ;
        RECT 33.155 0.765 33.325 0.845 ;
        RECT 32.185 0.595 33.325 0.765 ;
        RECT 32.185 0.515 32.355 0.595 ;
        RECT 33.155 0.515 33.325 0.595 ;
        RECT 33.725 0.765 33.895 1.050 ;
        RECT 34.210 1.720 34.865 1.890 ;
        RECT 36.130 1.805 36.300 1.885 ;
        RECT 37.100 1.805 37.270 1.885 ;
        RECT 38.025 1.880 38.195 5.345 ;
        RECT 40.295 5.470 40.465 7.250 ;
        RECT 41.175 5.470 41.345 7.250 ;
        RECT 42.055 5.470 42.225 7.250 ;
        RECT 45.105 5.470 45.275 7.250 ;
        RECT 45.985 5.470 46.155 7.250 ;
        RECT 46.865 5.470 47.035 7.250 ;
        RECT 49.615 5.515 49.785 7.250 ;
        RECT 50.495 5.515 50.665 7.250 ;
        RECT 40.295 5.300 43.005 5.470 ;
        RECT 45.105 5.300 47.815 5.470 ;
        RECT 49.615 5.345 51.145 5.515 ;
        RECT 39.875 2.055 40.045 5.095 ;
        RECT 34.210 0.985 34.380 1.720 ;
        RECT 36.130 1.635 37.270 1.805 ;
        RECT 34.695 0.765 34.865 1.535 ;
        RECT 33.725 0.595 34.865 0.765 ;
        RECT 33.725 0.515 33.895 0.595 ;
        RECT 34.695 0.515 34.865 0.595 ;
        RECT 36.130 0.505 36.300 1.635 ;
        RECT 37.100 0.755 37.270 1.635 ;
        RECT 37.585 1.710 38.195 1.880 ;
        RECT 39.355 1.815 39.525 1.895 ;
        RECT 40.325 1.815 40.495 1.895 ;
        RECT 41.295 1.815 41.465 1.895 ;
        RECT 37.585 0.975 37.755 1.710 ;
        RECT 39.355 1.645 41.465 1.815 ;
        RECT 38.070 0.755 38.240 1.525 ;
        RECT 37.100 0.585 38.240 0.755 ;
        RECT 37.100 0.505 37.270 0.585 ;
        RECT 38.070 0.505 38.240 0.585 ;
        RECT 39.355 0.515 39.525 1.645 ;
        RECT 40.325 0.765 40.495 1.645 ;
        RECT 41.295 1.565 41.465 1.645 ;
        RECT 40.815 1.220 40.985 1.300 ;
        RECT 41.865 1.220 42.035 1.895 ;
        RECT 42.835 1.890 43.005 5.300 ;
        RECT 44.685 2.055 44.855 5.095 ;
        RECT 46.905 2.055 47.075 5.095 ;
        RECT 40.815 1.050 42.035 1.220 ;
        RECT 40.815 0.970 40.985 1.050 ;
        RECT 41.295 0.765 41.465 0.845 ;
        RECT 40.325 0.595 41.465 0.765 ;
        RECT 40.325 0.515 40.495 0.595 ;
        RECT 41.295 0.515 41.465 0.595 ;
        RECT 41.865 0.765 42.035 1.050 ;
        RECT 42.350 1.720 43.005 1.890 ;
        RECT 44.165 1.815 44.335 1.895 ;
        RECT 45.135 1.815 45.305 1.895 ;
        RECT 46.105 1.815 46.275 1.895 ;
        RECT 42.350 0.985 42.520 1.720 ;
        RECT 44.165 1.645 46.275 1.815 ;
        RECT 42.835 0.765 43.005 1.535 ;
        RECT 41.865 0.595 43.005 0.765 ;
        RECT 41.865 0.515 42.035 0.595 ;
        RECT 42.835 0.515 43.005 0.595 ;
        RECT 44.165 0.515 44.335 1.645 ;
        RECT 45.135 0.765 45.305 1.645 ;
        RECT 46.105 1.565 46.275 1.645 ;
        RECT 45.625 1.220 45.795 1.300 ;
        RECT 46.675 1.220 46.845 1.895 ;
        RECT 47.645 1.890 47.815 5.300 ;
        RECT 49.495 2.055 49.665 5.095 ;
        RECT 50.265 4.940 50.435 5.095 ;
        RECT 50.235 4.765 50.435 4.940 ;
        RECT 50.235 2.055 50.405 4.765 ;
        RECT 45.625 1.050 46.845 1.220 ;
        RECT 45.625 0.970 45.795 1.050 ;
        RECT 46.105 0.765 46.275 0.845 ;
        RECT 45.135 0.595 46.275 0.765 ;
        RECT 45.135 0.515 45.305 0.595 ;
        RECT 46.105 0.515 46.275 0.595 ;
        RECT 46.675 0.765 46.845 1.050 ;
        RECT 47.160 1.720 47.815 1.890 ;
        RECT 49.080 1.805 49.250 1.885 ;
        RECT 50.050 1.805 50.220 1.885 ;
        RECT 50.975 1.880 51.145 5.345 ;
        RECT 53.245 5.470 53.415 7.250 ;
        RECT 54.125 5.470 54.295 7.250 ;
        RECT 55.005 5.470 55.175 7.250 ;
        RECT 58.055 5.470 58.225 7.250 ;
        RECT 58.935 5.470 59.105 7.250 ;
        RECT 59.815 5.470 59.985 7.250 ;
        RECT 62.565 5.515 62.735 7.250 ;
        RECT 63.445 5.515 63.615 7.250 ;
        RECT 53.245 5.300 55.955 5.470 ;
        RECT 58.055 5.300 60.765 5.470 ;
        RECT 62.565 5.345 64.095 5.515 ;
        RECT 52.825 2.055 52.995 5.095 ;
        RECT 55.045 2.055 55.215 5.095 ;
        RECT 47.160 0.985 47.330 1.720 ;
        RECT 49.080 1.635 50.220 1.805 ;
        RECT 47.645 0.765 47.815 1.535 ;
        RECT 46.675 0.595 47.815 0.765 ;
        RECT 46.675 0.515 46.845 0.595 ;
        RECT 47.645 0.515 47.815 0.595 ;
        RECT 49.080 0.505 49.250 1.635 ;
        RECT 50.050 0.755 50.220 1.635 ;
        RECT 50.535 1.710 51.145 1.880 ;
        RECT 52.305 1.815 52.475 1.895 ;
        RECT 53.275 1.815 53.445 1.895 ;
        RECT 54.245 1.815 54.415 1.895 ;
        RECT 50.535 0.975 50.705 1.710 ;
        RECT 52.305 1.645 54.415 1.815 ;
        RECT 51.020 0.755 51.190 1.525 ;
        RECT 50.050 0.585 51.190 0.755 ;
        RECT 50.050 0.505 50.220 0.585 ;
        RECT 51.020 0.505 51.190 0.585 ;
        RECT 52.305 0.515 52.475 1.645 ;
        RECT 53.275 0.765 53.445 1.645 ;
        RECT 54.245 1.565 54.415 1.645 ;
        RECT 53.765 1.220 53.935 1.300 ;
        RECT 54.815 1.220 54.985 1.895 ;
        RECT 55.785 1.890 55.955 5.300 ;
        RECT 57.635 2.055 57.805 5.095 ;
        RECT 53.765 1.050 54.985 1.220 ;
        RECT 53.765 0.970 53.935 1.050 ;
        RECT 54.245 0.765 54.415 0.845 ;
        RECT 53.275 0.595 54.415 0.765 ;
        RECT 53.275 0.515 53.445 0.595 ;
        RECT 54.245 0.515 54.415 0.595 ;
        RECT 54.815 0.765 54.985 1.050 ;
        RECT 55.300 1.720 55.955 1.890 ;
        RECT 57.115 1.815 57.285 1.895 ;
        RECT 58.085 1.815 58.255 1.895 ;
        RECT 59.055 1.815 59.225 1.895 ;
        RECT 55.300 0.985 55.470 1.720 ;
        RECT 57.115 1.645 59.225 1.815 ;
        RECT 55.785 0.765 55.955 1.535 ;
        RECT 54.815 0.595 55.955 0.765 ;
        RECT 54.815 0.515 54.985 0.595 ;
        RECT 55.785 0.515 55.955 0.595 ;
        RECT 57.115 0.515 57.285 1.645 ;
        RECT 58.085 0.765 58.255 1.645 ;
        RECT 59.055 1.565 59.225 1.645 ;
        RECT 58.575 1.220 58.745 1.300 ;
        RECT 59.625 1.220 59.795 1.895 ;
        RECT 60.595 1.890 60.765 5.300 ;
        RECT 62.445 2.055 62.615 5.095 ;
        RECT 63.215 4.940 63.385 5.095 ;
        RECT 63.185 4.765 63.385 4.940 ;
        RECT 63.185 2.055 63.355 4.765 ;
        RECT 58.575 1.050 59.795 1.220 ;
        RECT 58.575 0.970 58.745 1.050 ;
        RECT 59.055 0.765 59.225 0.845 ;
        RECT 58.085 0.595 59.225 0.765 ;
        RECT 58.085 0.515 58.255 0.595 ;
        RECT 59.055 0.515 59.225 0.595 ;
        RECT 59.625 0.765 59.795 1.050 ;
        RECT 60.110 1.720 60.765 1.890 ;
        RECT 62.030 1.805 62.200 1.885 ;
        RECT 63.000 1.805 63.170 1.885 ;
        RECT 63.925 1.880 64.095 5.345 ;
        RECT 66.195 5.470 66.365 7.250 ;
        RECT 67.075 5.470 67.245 7.250 ;
        RECT 67.955 5.470 68.125 7.250 ;
        RECT 71.005 5.470 71.175 7.250 ;
        RECT 71.885 5.470 72.055 7.250 ;
        RECT 72.765 5.470 72.935 7.250 ;
        RECT 75.515 5.515 75.685 7.250 ;
        RECT 76.395 5.515 76.565 7.250 ;
        RECT 78.845 7.055 79.025 7.225 ;
        RECT 78.845 5.525 79.015 7.055 ;
        RECT 79.725 5.525 79.895 7.225 ;
        RECT 66.195 5.300 68.905 5.470 ;
        RECT 71.005 5.300 73.715 5.470 ;
        RECT 75.515 5.345 77.045 5.515 ;
        RECT 78.845 5.355 79.895 5.525 ;
        RECT 65.775 2.055 65.945 5.095 ;
        RECT 60.110 0.985 60.280 1.720 ;
        RECT 62.030 1.635 63.170 1.805 ;
        RECT 60.595 0.765 60.765 1.535 ;
        RECT 59.625 0.595 60.765 0.765 ;
        RECT 59.625 0.515 59.795 0.595 ;
        RECT 60.595 0.515 60.765 0.595 ;
        RECT 62.030 0.505 62.200 1.635 ;
        RECT 63.000 0.755 63.170 1.635 ;
        RECT 63.485 1.710 64.095 1.880 ;
        RECT 65.255 1.815 65.425 1.895 ;
        RECT 66.225 1.815 66.395 1.895 ;
        RECT 67.195 1.815 67.365 1.895 ;
        RECT 63.485 0.975 63.655 1.710 ;
        RECT 65.255 1.645 67.365 1.815 ;
        RECT 63.970 0.755 64.140 1.525 ;
        RECT 63.000 0.585 64.140 0.755 ;
        RECT 63.000 0.505 63.170 0.585 ;
        RECT 63.970 0.505 64.140 0.585 ;
        RECT 65.255 0.515 65.425 1.645 ;
        RECT 66.225 0.765 66.395 1.645 ;
        RECT 67.195 1.565 67.365 1.645 ;
        RECT 66.715 1.220 66.885 1.300 ;
        RECT 67.765 1.220 67.935 1.895 ;
        RECT 68.735 1.890 68.905 5.300 ;
        RECT 70.585 2.055 70.755 5.095 ;
        RECT 72.805 2.055 72.975 5.095 ;
        RECT 66.715 1.050 67.935 1.220 ;
        RECT 66.715 0.970 66.885 1.050 ;
        RECT 67.195 0.765 67.365 0.845 ;
        RECT 66.225 0.595 67.365 0.765 ;
        RECT 66.225 0.515 66.395 0.595 ;
        RECT 67.195 0.515 67.365 0.595 ;
        RECT 67.765 0.765 67.935 1.050 ;
        RECT 68.250 1.720 68.905 1.890 ;
        RECT 70.065 1.815 70.235 1.895 ;
        RECT 71.035 1.815 71.205 1.895 ;
        RECT 72.005 1.815 72.175 1.895 ;
        RECT 68.250 0.985 68.420 1.720 ;
        RECT 70.065 1.645 72.175 1.815 ;
        RECT 68.735 0.765 68.905 1.535 ;
        RECT 67.765 0.595 68.905 0.765 ;
        RECT 67.765 0.515 67.935 0.595 ;
        RECT 68.735 0.515 68.905 0.595 ;
        RECT 70.065 0.515 70.235 1.645 ;
        RECT 71.035 0.765 71.205 1.645 ;
        RECT 72.005 1.565 72.175 1.645 ;
        RECT 71.525 1.220 71.695 1.300 ;
        RECT 72.575 1.220 72.745 1.895 ;
        RECT 73.545 1.890 73.715 5.300 ;
        RECT 75.395 2.055 75.565 5.095 ;
        RECT 76.165 4.940 76.335 5.095 ;
        RECT 76.135 4.765 76.335 4.940 ;
        RECT 76.135 2.055 76.305 4.765 ;
        RECT 71.525 1.050 72.745 1.220 ;
        RECT 71.525 0.970 71.695 1.050 ;
        RECT 72.005 0.765 72.175 0.845 ;
        RECT 71.035 0.595 72.175 0.765 ;
        RECT 71.035 0.515 71.205 0.595 ;
        RECT 72.005 0.515 72.175 0.595 ;
        RECT 72.575 0.765 72.745 1.050 ;
        RECT 73.060 1.720 73.715 1.890 ;
        RECT 74.980 1.805 75.150 1.885 ;
        RECT 75.950 1.805 76.120 1.885 ;
        RECT 76.875 1.880 77.045 5.345 ;
        RECT 79.725 5.275 79.895 5.355 ;
        RECT 81.725 7.055 83.655 7.225 ;
        RECT 81.725 5.275 81.895 7.055 ;
        RECT 82.165 5.525 82.335 6.795 ;
        RECT 82.605 5.785 82.775 7.055 ;
        RECT 83.045 5.525 83.215 6.795 ;
        RECT 83.485 5.605 83.655 7.055 ;
        RECT 85.065 7.055 86.995 7.225 ;
        RECT 82.165 5.355 83.215 5.525 ;
        RECT 83.045 5.275 83.215 5.355 ;
        RECT 85.065 5.275 85.235 7.055 ;
        RECT 85.505 5.525 85.675 6.795 ;
        RECT 85.945 5.785 86.115 7.055 ;
        RECT 86.385 5.525 86.555 6.795 ;
        RECT 86.825 5.785 86.995 7.055 ;
        RECT 85.505 5.355 87.035 5.525 ;
        RECT 78.355 2.055 78.525 5.100 ;
        RECT 79.505 4.940 79.675 5.100 ;
        RECT 79.465 4.770 79.675 4.940 ;
        RECT 79.465 2.055 79.635 4.770 ;
        RECT 82.055 2.055 82.225 5.100 ;
        RECT 83.535 2.055 83.705 5.100 ;
        RECT 85.015 2.055 85.185 5.100 ;
        RECT 86.125 4.770 86.315 5.100 ;
        RECT 86.125 2.055 86.295 4.770 ;
        RECT 73.060 0.985 73.230 1.720 ;
        RECT 74.980 1.635 76.120 1.805 ;
        RECT 73.545 0.765 73.715 1.535 ;
        RECT 72.575 0.595 73.715 0.765 ;
        RECT 72.575 0.515 72.745 0.595 ;
        RECT 73.545 0.515 73.715 0.595 ;
        RECT 74.980 0.505 75.150 1.635 ;
        RECT 75.950 0.755 76.120 1.635 ;
        RECT 76.435 1.710 77.045 1.880 ;
        RECT 78.310 1.805 78.480 1.885 ;
        RECT 79.280 1.805 79.450 1.885 ;
        RECT 76.435 0.975 76.605 1.710 ;
        RECT 78.310 1.635 79.450 1.805 ;
        RECT 76.920 0.755 77.090 1.525 ;
        RECT 75.950 0.585 77.090 0.755 ;
        RECT 75.950 0.505 76.120 0.585 ;
        RECT 76.920 0.505 77.090 0.585 ;
        RECT 78.310 0.505 78.480 1.635 ;
        RECT 79.280 0.755 79.450 1.635 ;
        RECT 79.765 1.310 79.935 1.485 ;
        RECT 79.760 1.155 79.935 1.310 ;
        RECT 79.760 0.975 79.930 1.155 ;
        RECT 80.250 0.755 80.420 1.885 ;
        RECT 79.280 0.585 80.420 0.755 ;
        RECT 79.280 0.505 79.450 0.585 ;
        RECT 80.250 0.505 80.420 0.585 ;
        RECT 81.640 1.805 81.810 1.885 ;
        RECT 82.610 1.805 82.780 1.885 ;
        RECT 81.640 1.635 82.780 1.805 ;
        RECT 81.640 0.505 81.810 1.635 ;
        RECT 82.610 0.755 82.780 1.635 ;
        RECT 83.095 0.975 83.265 1.485 ;
        RECT 83.580 0.755 83.750 1.885 ;
        RECT 82.610 0.585 83.750 0.755 ;
        RECT 82.610 0.505 82.780 0.585 ;
        RECT 83.580 0.505 83.750 0.585 ;
        RECT 84.970 1.805 85.140 1.885 ;
        RECT 85.940 1.805 86.110 1.885 ;
        RECT 86.865 1.870 87.035 5.355 ;
        RECT 88.345 2.055 88.515 5.095 ;
        RECT 84.970 1.635 86.110 1.805 ;
        RECT 84.970 0.505 85.140 1.635 ;
        RECT 85.940 0.755 86.110 1.635 ;
        RECT 86.425 1.700 87.035 1.870 ;
        RECT 86.425 0.975 86.595 1.700 ;
        RECT 86.910 0.755 87.080 1.530 ;
        RECT 85.940 0.585 87.080 0.755 ;
        RECT 85.940 0.505 86.110 0.585 ;
        RECT 86.910 0.505 87.080 0.585 ;
      LAYER mcon ;
        RECT 1.025 4.355 1.195 4.525 ;
        RECT 3.245 3.615 3.415 3.785 ;
        RECT 3.985 3.985 4.155 4.155 ;
        RECT 5.835 3.985 6.005 4.155 ;
        RECT 8.795 3.615 8.965 3.785 ;
        RECT 10.645 3.615 10.815 3.785 ;
        RECT 11.385 4.355 11.555 4.525 ;
        RECT 12.125 3.615 12.295 3.785 ;
        RECT 13.975 3.615 14.145 3.785 ;
        RECT 16.935 4.355 17.105 4.525 ;
        RECT 18.785 3.985 18.955 4.155 ;
        RECT 21.005 2.875 21.175 3.045 ;
        RECT 21.745 3.985 21.915 4.155 ;
        RECT 23.595 3.985 23.765 4.155 ;
        RECT 24.335 4.355 24.505 4.525 ;
        RECT 25.075 2.875 25.245 3.045 ;
        RECT 26.925 4.355 27.095 4.525 ;
        RECT 29.145 3.615 29.315 3.785 ;
        RECT 29.885 3.985 30.055 4.155 ;
        RECT 31.735 3.985 31.905 4.155 ;
        RECT 34.695 3.615 34.865 3.785 ;
        RECT 36.545 3.615 36.715 3.785 ;
        RECT 37.285 4.355 37.455 4.525 ;
        RECT 38.025 3.615 38.195 3.785 ;
        RECT 39.875 3.615 40.045 3.785 ;
        RECT 42.835 4.355 43.005 4.525 ;
        RECT 44.685 3.985 44.855 4.155 ;
        RECT 46.905 3.245 47.075 3.415 ;
        RECT 47.645 3.985 47.815 4.155 ;
        RECT 49.495 3.985 49.665 4.155 ;
        RECT 50.235 4.355 50.405 4.525 ;
        RECT 50.975 3.245 51.145 3.415 ;
        RECT 52.825 4.355 52.995 4.525 ;
        RECT 55.045 3.615 55.215 3.785 ;
        RECT 55.785 3.985 55.955 4.155 ;
        RECT 57.635 3.985 57.805 4.155 ;
        RECT 60.595 3.615 60.765 3.785 ;
        RECT 62.445 3.615 62.615 3.785 ;
        RECT 63.185 4.355 63.355 4.525 ;
        RECT 79.725 5.355 79.895 5.525 ;
        RECT 63.925 3.615 64.095 3.785 ;
        RECT 65.775 3.615 65.945 3.785 ;
        RECT 68.735 4.355 68.905 4.525 ;
        RECT 70.585 3.985 70.755 4.155 ;
        RECT 72.805 3.615 72.975 3.785 ;
        RECT 73.545 3.985 73.715 4.155 ;
        RECT 75.395 3.985 75.565 4.155 ;
        RECT 76.135 4.355 76.305 4.525 ;
        RECT 81.725 5.355 81.895 5.525 ;
        RECT 83.045 5.355 83.215 5.525 ;
        RECT 85.065 5.355 85.235 5.525 ;
        RECT 76.875 3.615 77.045 3.785 ;
        RECT 78.355 4.725 78.525 4.895 ;
        RECT 78.355 3.245 78.525 3.415 ;
        RECT 79.465 4.355 79.635 4.525 ;
        RECT 79.465 3.615 79.635 3.785 ;
        RECT 82.055 4.725 82.225 4.895 ;
        RECT 83.535 2.875 83.705 3.045 ;
        RECT 83.535 2.135 83.705 2.305 ;
        RECT 85.015 2.135 85.185 2.305 ;
        RECT 86.125 4.355 86.295 4.525 ;
        RECT 86.865 3.985 87.035 4.155 ;
        RECT 79.765 1.235 79.935 1.405 ;
        RECT 83.095 1.235 83.265 1.405 ;
        RECT 88.345 3.985 88.515 4.155 ;
        RECT 86.425 1.235 86.595 1.405 ;
      LAYER met1 ;
        RECT 79.695 5.525 79.925 5.555 ;
        RECT 81.695 5.525 81.925 5.555 ;
        RECT 83.015 5.525 83.245 5.555 ;
        RECT 85.035 5.525 85.265 5.555 ;
        RECT 79.665 5.355 81.955 5.525 ;
        RECT 82.985 5.355 85.295 5.525 ;
        RECT 79.695 5.325 79.925 5.355 ;
        RECT 81.695 5.325 81.925 5.355 ;
        RECT 83.015 5.325 83.245 5.355 ;
        RECT 85.035 5.325 85.265 5.355 ;
        RECT 78.325 4.895 78.555 4.925 ;
        RECT 82.025 4.895 82.255 4.925 ;
        RECT 78.295 4.725 82.285 4.895 ;
        RECT 78.325 4.695 78.555 4.725 ;
        RECT 82.025 4.695 82.255 4.725 ;
        RECT 0.995 4.525 1.225 4.555 ;
        RECT 11.355 4.525 11.585 4.555 ;
        RECT 16.905 4.525 17.135 4.555 ;
        RECT 24.305 4.525 24.535 4.555 ;
        RECT 26.895 4.525 27.125 4.555 ;
        RECT 37.255 4.525 37.485 4.555 ;
        RECT 42.805 4.525 43.035 4.555 ;
        RECT 50.205 4.525 50.435 4.555 ;
        RECT 52.795 4.525 53.025 4.555 ;
        RECT 63.155 4.525 63.385 4.555 ;
        RECT 68.705 4.525 68.935 4.555 ;
        RECT 76.105 4.525 76.335 4.555 ;
        RECT 79.435 4.525 79.665 4.555 ;
        RECT 86.095 4.525 86.325 4.555 ;
        RECT 0.965 4.355 24.565 4.525 ;
        RECT 26.865 4.355 50.465 4.525 ;
        RECT 52.765 4.355 76.365 4.525 ;
        RECT 79.405 4.355 86.355 4.525 ;
        RECT 0.995 4.325 1.225 4.355 ;
        RECT 11.355 4.325 11.585 4.355 ;
        RECT 16.905 4.325 17.135 4.355 ;
        RECT 24.305 4.325 24.535 4.355 ;
        RECT 26.895 4.325 27.125 4.355 ;
        RECT 37.255 4.325 37.485 4.355 ;
        RECT 42.805 4.325 43.035 4.355 ;
        RECT 50.205 4.325 50.435 4.355 ;
        RECT 52.795 4.325 53.025 4.355 ;
        RECT 63.155 4.325 63.385 4.355 ;
        RECT 68.705 4.325 68.935 4.355 ;
        RECT 76.105 4.325 76.335 4.355 ;
        RECT 79.435 4.325 79.665 4.355 ;
        RECT 86.095 4.325 86.325 4.355 ;
        RECT 3.955 4.155 4.185 4.185 ;
        RECT 5.805 4.155 6.035 4.185 ;
        RECT 18.755 4.155 18.985 4.185 ;
        RECT 21.715 4.155 21.945 4.185 ;
        RECT 23.565 4.155 23.795 4.185 ;
        RECT 29.855 4.155 30.085 4.185 ;
        RECT 31.705 4.155 31.935 4.185 ;
        RECT 44.655 4.155 44.885 4.185 ;
        RECT 47.615 4.155 47.845 4.185 ;
        RECT 49.465 4.155 49.695 4.185 ;
        RECT 55.755 4.155 55.985 4.185 ;
        RECT 57.605 4.155 57.835 4.185 ;
        RECT 70.555 4.155 70.785 4.185 ;
        RECT 73.515 4.155 73.745 4.185 ;
        RECT 75.365 4.155 75.595 4.185 ;
        RECT 86.835 4.155 87.065 4.185 ;
        RECT 88.315 4.155 88.545 4.185 ;
        RECT 3.925 3.985 19.015 4.155 ;
        RECT 21.685 3.985 23.825 4.155 ;
        RECT 29.825 3.985 44.915 4.155 ;
        RECT 47.585 3.985 49.725 4.155 ;
        RECT 55.725 3.985 70.815 4.155 ;
        RECT 73.485 3.985 75.625 4.155 ;
        RECT 86.805 3.985 88.575 4.155 ;
        RECT 3.955 3.955 4.185 3.985 ;
        RECT 5.805 3.955 6.035 3.985 ;
        RECT 18.755 3.955 18.985 3.985 ;
        RECT 21.715 3.955 21.945 3.985 ;
        RECT 23.565 3.955 23.795 3.985 ;
        RECT 29.855 3.955 30.085 3.985 ;
        RECT 31.705 3.955 31.935 3.985 ;
        RECT 44.655 3.955 44.885 3.985 ;
        RECT 47.615 3.955 47.845 3.985 ;
        RECT 49.465 3.955 49.695 3.985 ;
        RECT 55.755 3.955 55.985 3.985 ;
        RECT 57.605 3.955 57.835 3.985 ;
        RECT 70.555 3.955 70.785 3.985 ;
        RECT 73.515 3.955 73.745 3.985 ;
        RECT 75.365 3.955 75.595 3.985 ;
        RECT 86.835 3.955 87.065 3.985 ;
        RECT 88.315 3.955 88.545 3.985 ;
        RECT 3.215 3.785 3.445 3.815 ;
        RECT 8.765 3.785 8.995 3.815 ;
        RECT 10.615 3.785 10.845 3.815 ;
        RECT 12.095 3.785 12.325 3.815 ;
        RECT 13.945 3.785 14.175 3.815 ;
        RECT 29.115 3.785 29.345 3.815 ;
        RECT 34.665 3.785 34.895 3.815 ;
        RECT 36.515 3.785 36.745 3.815 ;
        RECT 37.995 3.785 38.225 3.815 ;
        RECT 39.845 3.785 40.075 3.815 ;
        RECT 55.015 3.785 55.245 3.815 ;
        RECT 60.565 3.785 60.795 3.815 ;
        RECT 62.415 3.785 62.645 3.815 ;
        RECT 63.895 3.785 64.125 3.815 ;
        RECT 65.745 3.785 65.975 3.815 ;
        RECT 72.775 3.785 73.005 3.815 ;
        RECT 76.845 3.785 77.075 3.815 ;
        RECT 79.435 3.785 79.665 3.815 ;
        RECT 3.185 3.615 10.875 3.785 ;
        RECT 12.065 3.615 14.205 3.785 ;
        RECT 29.085 3.615 36.775 3.785 ;
        RECT 37.965 3.615 40.105 3.785 ;
        RECT 54.985 3.615 62.675 3.785 ;
        RECT 63.865 3.615 66.005 3.785 ;
        RECT 72.745 3.615 79.695 3.785 ;
        RECT 3.215 3.585 3.445 3.615 ;
        RECT 8.765 3.585 8.995 3.615 ;
        RECT 10.615 3.585 10.845 3.615 ;
        RECT 12.095 3.585 12.325 3.615 ;
        RECT 13.945 3.585 14.175 3.615 ;
        RECT 29.115 3.585 29.345 3.615 ;
        RECT 34.665 3.585 34.895 3.615 ;
        RECT 36.515 3.585 36.745 3.615 ;
        RECT 37.995 3.585 38.225 3.615 ;
        RECT 39.845 3.585 40.075 3.615 ;
        RECT 55.015 3.585 55.245 3.615 ;
        RECT 60.565 3.585 60.795 3.615 ;
        RECT 62.415 3.585 62.645 3.615 ;
        RECT 63.895 3.585 64.125 3.615 ;
        RECT 65.745 3.585 65.975 3.615 ;
        RECT 72.775 3.585 73.005 3.615 ;
        RECT 76.845 3.585 77.075 3.615 ;
        RECT 79.435 3.585 79.665 3.615 ;
        RECT 46.875 3.415 47.105 3.445 ;
        RECT 50.945 3.415 51.175 3.445 ;
        RECT 78.325 3.415 78.555 3.445 ;
        RECT 46.845 3.245 78.585 3.415 ;
        RECT 46.875 3.215 47.105 3.245 ;
        RECT 50.945 3.215 51.175 3.245 ;
        RECT 78.325 3.215 78.555 3.245 ;
        RECT 20.975 3.045 21.205 3.075 ;
        RECT 25.045 3.045 25.275 3.075 ;
        RECT 83.505 3.045 83.735 3.075 ;
        RECT 20.945 2.875 83.765 3.045 ;
        RECT 20.975 2.845 21.205 2.875 ;
        RECT 25.045 2.845 25.275 2.875 ;
        RECT 83.505 2.845 83.735 2.875 ;
        RECT 83.505 2.305 83.735 2.335 ;
        RECT 84.985 2.305 85.215 2.335 ;
        RECT 83.475 2.135 85.245 2.305 ;
        RECT 83.505 2.105 83.735 2.135 ;
        RECT 84.985 2.105 85.215 2.135 ;
        RECT 79.735 1.405 79.965 1.435 ;
        RECT 83.065 1.405 83.295 1.435 ;
        RECT 86.395 1.405 86.625 1.435 ;
        RECT 79.705 1.235 86.655 1.405 ;
        RECT 79.735 1.205 79.965 1.235 ;
        RECT 83.065 1.205 83.295 1.235 ;
        RECT 86.395 1.205 86.625 1.235 ;
  END
END TMRDFFRNQX1






MACRO TMRDFFSNQNX1
  CLASS BLOCK ;
  FOREIGN TMRDFFSNQNX1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 84.090 BY 7.950 ;
  PIN QN
    ANTENNADIFFAREA 1.734950 ;
    PORT
      LAYER li1 ;
        RECT 81.065 5.525 81.235 6.795 ;
        RECT 81.945 5.525 82.115 6.795 ;
        RECT 81.065 5.355 82.595 5.525 ;
        RECT 82.425 1.870 82.595 5.355 ;
        RECT 81.985 1.700 82.595 1.870 ;
        RECT 75.325 1.310 75.495 1.485 ;
        RECT 75.320 1.155 75.495 1.310 ;
        RECT 75.320 0.975 75.490 1.155 ;
        RECT 78.655 0.975 78.825 1.485 ;
        RECT 81.985 0.975 82.155 1.700 ;
      LAYER mcon ;
        RECT 82.425 3.985 82.595 4.155 ;
        RECT 75.325 1.235 75.495 1.405 ;
        RECT 78.655 1.235 78.825 1.405 ;
        RECT 81.985 1.235 82.155 1.405 ;
      LAYER met1 ;
        RECT 82.395 4.155 82.625 4.185 ;
        RECT 82.365 3.985 82.775 4.155 ;
        RECT 82.395 3.955 82.625 3.985 ;
        RECT 75.295 1.405 75.525 1.435 ;
        RECT 78.625 1.405 78.855 1.435 ;
        RECT 81.955 1.405 82.185 1.435 ;
        RECT 75.265 1.235 82.215 1.405 ;
        RECT 75.295 1.205 75.525 1.235 ;
        RECT 78.625 1.205 78.855 1.235 ;
        RECT 81.955 1.205 82.185 1.235 ;
    END
  END QN
  PIN D
    ANTENNAGATEAREA 3.099750 ;
    PORT
      LAYER li1 ;
        RECT 1.025 2.055 1.195 5.095 ;
        RECT 25.445 2.055 25.615 5.095 ;
        RECT 49.865 2.055 50.035 5.095 ;
      LAYER mcon ;
        RECT 1.025 2.135 1.195 2.305 ;
        RECT 25.445 2.135 25.615 2.305 ;
        RECT 49.865 2.135 50.035 2.305 ;
      LAYER met1 ;
        RECT 0.995 2.305 1.225 2.335 ;
        RECT 25.415 2.305 25.645 2.335 ;
        RECT 49.835 2.305 50.065 2.335 ;
        RECT 0.965 2.135 50.095 2.305 ;
        RECT 0.995 2.105 1.225 2.135 ;
        RECT 25.415 2.105 25.645 2.135 ;
        RECT 49.835 2.105 50.065 2.135 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 6.126300 ;
    PORT
      LAYER li1 ;
        RECT 5.465 2.055 5.635 5.095 ;
        RECT 14.745 4.975 14.915 5.095 ;
        RECT 14.715 4.765 14.915 4.975 ;
        RECT 14.715 2.055 14.885 4.765 ;
        RECT 29.885 2.055 30.055 5.095 ;
        RECT 39.165 4.975 39.335 5.095 ;
        RECT 39.135 4.765 39.335 4.975 ;
        RECT 39.135 2.055 39.305 4.765 ;
        RECT 54.305 2.055 54.475 5.095 ;
        RECT 63.585 4.975 63.755 5.095 ;
        RECT 63.555 4.765 63.755 4.975 ;
        RECT 63.555 2.055 63.725 4.765 ;
      LAYER mcon ;
        RECT 5.465 4.725 5.635 4.895 ;
        RECT 14.715 4.725 14.885 4.895 ;
        RECT 29.885 4.725 30.055 4.895 ;
        RECT 39.135 4.725 39.305 4.895 ;
        RECT 54.305 4.725 54.475 4.895 ;
        RECT 63.555 4.725 63.725 4.895 ;
      LAYER met1 ;
        RECT 5.435 4.895 5.665 4.925 ;
        RECT 14.685 4.895 14.915 4.925 ;
        RECT 29.855 4.895 30.085 4.925 ;
        RECT 39.105 4.895 39.335 4.925 ;
        RECT 54.275 4.895 54.505 4.925 ;
        RECT 63.525 4.895 63.755 4.925 ;
        RECT 5.405 4.725 63.785 4.895 ;
        RECT 5.435 4.695 5.665 4.725 ;
        RECT 14.685 4.695 14.915 4.725 ;
        RECT 29.855 4.695 30.085 4.725 ;
        RECT 39.105 4.695 39.335 4.725 ;
        RECT 54.275 4.695 54.505 4.725 ;
        RECT 63.525 4.695 63.755 4.725 ;
    END
  END CLK
  PIN SN
    ANTENNAGATEAREA 6.089100 ;
    PORT
      LAYER li1 ;
        RECT 10.275 2.055 10.445 5.095 ;
        RECT 21.745 2.055 21.915 5.095 ;
        RECT 34.695 2.055 34.865 5.095 ;
        RECT 46.165 2.055 46.335 5.095 ;
        RECT 59.115 2.055 59.285 5.095 ;
        RECT 70.585 2.055 70.755 5.095 ;
      LAYER mcon ;
        RECT 10.275 2.505 10.445 2.675 ;
        RECT 21.745 2.505 21.915 2.675 ;
        RECT 34.695 2.505 34.865 2.675 ;
        RECT 46.165 2.505 46.335 2.675 ;
        RECT 59.115 2.505 59.285 2.675 ;
        RECT 70.585 2.505 70.755 2.675 ;
      LAYER met1 ;
        RECT 10.245 2.675 10.475 2.705 ;
        RECT 21.715 2.675 21.945 2.705 ;
        RECT 34.665 2.675 34.895 2.705 ;
        RECT 46.135 2.675 46.365 2.705 ;
        RECT 59.085 2.675 59.315 2.705 ;
        RECT 70.555 2.675 70.785 2.705 ;
        RECT 10.215 2.505 70.815 2.675 ;
        RECT 10.245 2.475 10.475 2.505 ;
        RECT 21.715 2.475 21.945 2.505 ;
        RECT 34.665 2.475 34.895 2.505 ;
        RECT 46.135 2.475 46.365 2.505 ;
        RECT 59.085 2.475 59.315 2.505 ;
        RECT 70.555 2.475 70.785 2.505 ;
    END
  END SN
  PIN VDD
    ANTENNADIFFAREA 96.856300 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 83.670 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 83.405 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 0.705 5.365 0.875 7.460 ;
        RECT 1.585 5.785 1.755 7.460 ;
        RECT 2.465 5.785 2.635 7.460 ;
        RECT 3.175 4.340 3.485 7.460 ;
        RECT 4.335 5.445 4.505 7.460 ;
        RECT 5.215 5.785 5.385 7.460 ;
        RECT 6.095 5.785 6.265 7.460 ;
        RECT 6.975 5.785 7.145 7.460 ;
        RECT 7.985 4.340 8.295 7.460 ;
        RECT 9.145 5.445 9.315 7.460 ;
        RECT 10.025 5.785 10.195 7.460 ;
        RECT 10.905 5.785 11.075 7.460 ;
        RECT 11.785 5.785 11.955 7.460 ;
        RECT 12.795 4.340 13.105 7.460 ;
        RECT 13.655 5.365 13.825 7.460 ;
        RECT 14.535 5.785 14.705 7.460 ;
        RECT 15.415 5.785 15.585 7.460 ;
        RECT 16.125 4.340 16.435 7.460 ;
        RECT 16.985 5.365 17.155 7.460 ;
        RECT 17.865 5.785 18.035 7.460 ;
        RECT 18.745 5.785 18.915 7.460 ;
        RECT 19.455 4.340 19.765 7.460 ;
        RECT 20.615 5.445 20.785 7.460 ;
        RECT 21.495 5.785 21.665 7.460 ;
        RECT 22.375 5.785 22.545 7.460 ;
        RECT 23.255 5.785 23.425 7.460 ;
        RECT 24.265 4.340 24.575 7.460 ;
        RECT 25.125 5.365 25.295 7.460 ;
        RECT 26.005 5.785 26.175 7.460 ;
        RECT 26.885 5.785 27.055 7.460 ;
        RECT 27.595 4.340 27.905 7.460 ;
        RECT 28.755 5.445 28.925 7.460 ;
        RECT 29.635 5.785 29.805 7.460 ;
        RECT 30.515 5.785 30.685 7.460 ;
        RECT 31.395 5.785 31.565 7.460 ;
        RECT 32.405 4.340 32.715 7.460 ;
        RECT 33.565 5.445 33.735 7.460 ;
        RECT 34.445 5.785 34.615 7.460 ;
        RECT 35.325 5.785 35.495 7.460 ;
        RECT 36.205 5.785 36.375 7.460 ;
        RECT 37.215 4.340 37.525 7.460 ;
        RECT 38.075 5.365 38.245 7.460 ;
        RECT 38.955 5.785 39.125 7.460 ;
        RECT 39.835 5.785 40.005 7.460 ;
        RECT 40.545 4.340 40.855 7.460 ;
        RECT 41.405 5.365 41.575 7.460 ;
        RECT 42.285 5.785 42.455 7.460 ;
        RECT 43.165 5.785 43.335 7.460 ;
        RECT 43.875 4.340 44.185 7.460 ;
        RECT 45.035 5.445 45.205 7.460 ;
        RECT 45.915 5.785 46.085 7.460 ;
        RECT 46.795 5.785 46.965 7.460 ;
        RECT 47.675 5.785 47.845 7.460 ;
        RECT 48.685 4.340 48.995 7.460 ;
        RECT 49.545 5.365 49.715 7.460 ;
        RECT 50.425 5.785 50.595 7.460 ;
        RECT 51.305 5.785 51.475 7.460 ;
        RECT 52.015 4.340 52.325 7.460 ;
        RECT 53.175 5.445 53.345 7.460 ;
        RECT 54.055 5.785 54.225 7.460 ;
        RECT 54.935 5.785 55.105 7.460 ;
        RECT 55.815 5.785 55.985 7.460 ;
        RECT 56.825 4.340 57.135 7.460 ;
        RECT 57.985 5.445 58.155 7.460 ;
        RECT 58.865 5.785 59.035 7.460 ;
        RECT 59.745 5.785 59.915 7.460 ;
        RECT 60.625 5.785 60.795 7.460 ;
        RECT 61.635 4.340 61.945 7.460 ;
        RECT 62.495 5.365 62.665 7.460 ;
        RECT 63.375 5.785 63.545 7.460 ;
        RECT 64.255 5.785 64.425 7.460 ;
        RECT 64.965 4.340 65.275 7.460 ;
        RECT 65.825 5.365 65.995 7.460 ;
        RECT 66.705 5.785 66.875 7.460 ;
        RECT 67.585 5.785 67.755 7.460 ;
        RECT 68.295 4.340 68.605 7.460 ;
        RECT 69.455 5.445 69.625 7.460 ;
        RECT 70.335 5.785 70.505 7.460 ;
        RECT 71.215 5.785 71.385 7.460 ;
        RECT 72.095 5.785 72.265 7.460 ;
        RECT 73.105 4.340 73.415 7.460 ;
        RECT 73.965 5.355 74.135 7.460 ;
        RECT 74.845 5.785 75.015 7.460 ;
        RECT 75.725 5.355 75.895 7.460 ;
        RECT 76.435 4.340 76.745 7.460 ;
        RECT 79.765 4.340 80.075 7.460 ;
        RECT 83.095 4.340 83.405 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 0.995 7.525 1.165 7.695 ;
        RECT 1.355 7.525 1.525 7.695 ;
        RECT 1.805 7.525 1.975 7.695 ;
        RECT 2.165 7.525 2.335 7.695 ;
        RECT 2.525 7.525 2.695 7.695 ;
        RECT 2.885 7.525 3.055 7.695 ;
        RECT 3.605 7.525 3.775 7.695 ;
        RECT 3.965 7.525 4.135 7.695 ;
        RECT 4.325 7.525 4.495 7.695 ;
        RECT 4.685 7.525 4.855 7.695 ;
        RECT 5.045 7.525 5.215 7.695 ;
        RECT 5.405 7.525 5.575 7.695 ;
        RECT 5.895 7.525 6.065 7.695 ;
        RECT 6.255 7.525 6.425 7.695 ;
        RECT 6.615 7.525 6.785 7.695 ;
        RECT 6.975 7.525 7.145 7.695 ;
        RECT 7.335 7.525 7.505 7.695 ;
        RECT 7.695 7.525 7.865 7.695 ;
        RECT 8.415 7.525 8.585 7.695 ;
        RECT 8.775 7.525 8.945 7.695 ;
        RECT 9.135 7.525 9.305 7.695 ;
        RECT 9.495 7.525 9.665 7.695 ;
        RECT 9.855 7.525 10.025 7.695 ;
        RECT 10.215 7.525 10.385 7.695 ;
        RECT 10.705 7.525 10.875 7.695 ;
        RECT 11.065 7.525 11.235 7.695 ;
        RECT 11.425 7.525 11.595 7.695 ;
        RECT 11.785 7.525 11.955 7.695 ;
        RECT 12.145 7.525 12.315 7.695 ;
        RECT 12.505 7.525 12.675 7.695 ;
        RECT 13.225 7.525 13.395 7.695 ;
        RECT 13.585 7.525 13.755 7.695 ;
        RECT 13.945 7.525 14.115 7.695 ;
        RECT 14.305 7.525 14.475 7.695 ;
        RECT 14.755 7.525 14.925 7.695 ;
        RECT 15.115 7.525 15.285 7.695 ;
        RECT 15.475 7.525 15.645 7.695 ;
        RECT 15.835 7.525 16.005 7.695 ;
        RECT 16.555 7.525 16.725 7.695 ;
        RECT 16.915 7.525 17.085 7.695 ;
        RECT 17.275 7.525 17.445 7.695 ;
        RECT 17.635 7.525 17.805 7.695 ;
        RECT 18.085 7.525 18.255 7.695 ;
        RECT 18.445 7.525 18.615 7.695 ;
        RECT 18.805 7.525 18.975 7.695 ;
        RECT 19.165 7.525 19.335 7.695 ;
        RECT 19.885 7.525 20.055 7.695 ;
        RECT 20.245 7.525 20.415 7.695 ;
        RECT 20.605 7.525 20.775 7.695 ;
        RECT 20.965 7.525 21.135 7.695 ;
        RECT 21.325 7.525 21.495 7.695 ;
        RECT 21.685 7.525 21.855 7.695 ;
        RECT 22.175 7.525 22.345 7.695 ;
        RECT 22.535 7.525 22.705 7.695 ;
        RECT 22.895 7.525 23.065 7.695 ;
        RECT 23.255 7.525 23.425 7.695 ;
        RECT 23.615 7.525 23.785 7.695 ;
        RECT 23.975 7.525 24.145 7.695 ;
        RECT 24.695 7.525 24.865 7.695 ;
        RECT 25.055 7.525 25.225 7.695 ;
        RECT 25.415 7.525 25.585 7.695 ;
        RECT 25.775 7.525 25.945 7.695 ;
        RECT 26.225 7.525 26.395 7.695 ;
        RECT 26.585 7.525 26.755 7.695 ;
        RECT 26.945 7.525 27.115 7.695 ;
        RECT 27.305 7.525 27.475 7.695 ;
        RECT 28.025 7.525 28.195 7.695 ;
        RECT 28.385 7.525 28.555 7.695 ;
        RECT 28.745 7.525 28.915 7.695 ;
        RECT 29.105 7.525 29.275 7.695 ;
        RECT 29.465 7.525 29.635 7.695 ;
        RECT 29.825 7.525 29.995 7.695 ;
        RECT 30.315 7.525 30.485 7.695 ;
        RECT 30.675 7.525 30.845 7.695 ;
        RECT 31.035 7.525 31.205 7.695 ;
        RECT 31.395 7.525 31.565 7.695 ;
        RECT 31.755 7.525 31.925 7.695 ;
        RECT 32.115 7.525 32.285 7.695 ;
        RECT 32.835 7.525 33.005 7.695 ;
        RECT 33.195 7.525 33.365 7.695 ;
        RECT 33.555 7.525 33.725 7.695 ;
        RECT 33.915 7.525 34.085 7.695 ;
        RECT 34.275 7.525 34.445 7.695 ;
        RECT 34.635 7.525 34.805 7.695 ;
        RECT 35.125 7.525 35.295 7.695 ;
        RECT 35.485 7.525 35.655 7.695 ;
        RECT 35.845 7.525 36.015 7.695 ;
        RECT 36.205 7.525 36.375 7.695 ;
        RECT 36.565 7.525 36.735 7.695 ;
        RECT 36.925 7.525 37.095 7.695 ;
        RECT 37.645 7.525 37.815 7.695 ;
        RECT 38.005 7.525 38.175 7.695 ;
        RECT 38.365 7.525 38.535 7.695 ;
        RECT 38.725 7.525 38.895 7.695 ;
        RECT 39.175 7.525 39.345 7.695 ;
        RECT 39.535 7.525 39.705 7.695 ;
        RECT 39.895 7.525 40.065 7.695 ;
        RECT 40.255 7.525 40.425 7.695 ;
        RECT 40.975 7.525 41.145 7.695 ;
        RECT 41.335 7.525 41.505 7.695 ;
        RECT 41.695 7.525 41.865 7.695 ;
        RECT 42.055 7.525 42.225 7.695 ;
        RECT 42.505 7.525 42.675 7.695 ;
        RECT 42.865 7.525 43.035 7.695 ;
        RECT 43.225 7.525 43.395 7.695 ;
        RECT 43.585 7.525 43.755 7.695 ;
        RECT 44.305 7.525 44.475 7.695 ;
        RECT 44.665 7.525 44.835 7.695 ;
        RECT 45.025 7.525 45.195 7.695 ;
        RECT 45.385 7.525 45.555 7.695 ;
        RECT 45.745 7.525 45.915 7.695 ;
        RECT 46.105 7.525 46.275 7.695 ;
        RECT 46.595 7.525 46.765 7.695 ;
        RECT 46.955 7.525 47.125 7.695 ;
        RECT 47.315 7.525 47.485 7.695 ;
        RECT 47.675 7.525 47.845 7.695 ;
        RECT 48.035 7.525 48.205 7.695 ;
        RECT 48.395 7.525 48.565 7.695 ;
        RECT 49.115 7.525 49.285 7.695 ;
        RECT 49.475 7.525 49.645 7.695 ;
        RECT 49.835 7.525 50.005 7.695 ;
        RECT 50.195 7.525 50.365 7.695 ;
        RECT 50.645 7.525 50.815 7.695 ;
        RECT 51.005 7.525 51.175 7.695 ;
        RECT 51.365 7.525 51.535 7.695 ;
        RECT 51.725 7.525 51.895 7.695 ;
        RECT 52.445 7.525 52.615 7.695 ;
        RECT 52.805 7.525 52.975 7.695 ;
        RECT 53.165 7.525 53.335 7.695 ;
        RECT 53.525 7.525 53.695 7.695 ;
        RECT 53.885 7.525 54.055 7.695 ;
        RECT 54.245 7.525 54.415 7.695 ;
        RECT 54.735 7.525 54.905 7.695 ;
        RECT 55.095 7.525 55.265 7.695 ;
        RECT 55.455 7.525 55.625 7.695 ;
        RECT 55.815 7.525 55.985 7.695 ;
        RECT 56.175 7.525 56.345 7.695 ;
        RECT 56.535 7.525 56.705 7.695 ;
        RECT 57.255 7.525 57.425 7.695 ;
        RECT 57.615 7.525 57.785 7.695 ;
        RECT 57.975 7.525 58.145 7.695 ;
        RECT 58.335 7.525 58.505 7.695 ;
        RECT 58.695 7.525 58.865 7.695 ;
        RECT 59.055 7.525 59.225 7.695 ;
        RECT 59.545 7.525 59.715 7.695 ;
        RECT 59.905 7.525 60.075 7.695 ;
        RECT 60.265 7.525 60.435 7.695 ;
        RECT 60.625 7.525 60.795 7.695 ;
        RECT 60.985 7.525 61.155 7.695 ;
        RECT 61.345 7.525 61.515 7.695 ;
        RECT 62.065 7.525 62.235 7.695 ;
        RECT 62.425 7.525 62.595 7.695 ;
        RECT 62.785 7.525 62.955 7.695 ;
        RECT 63.145 7.525 63.315 7.695 ;
        RECT 63.595 7.525 63.765 7.695 ;
        RECT 63.955 7.525 64.125 7.695 ;
        RECT 64.315 7.525 64.485 7.695 ;
        RECT 64.675 7.525 64.845 7.695 ;
        RECT 65.395 7.525 65.565 7.695 ;
        RECT 65.755 7.525 65.925 7.695 ;
        RECT 66.115 7.525 66.285 7.695 ;
        RECT 66.475 7.525 66.645 7.695 ;
        RECT 66.925 7.525 67.095 7.695 ;
        RECT 67.285 7.525 67.455 7.695 ;
        RECT 67.645 7.525 67.815 7.695 ;
        RECT 68.005 7.525 68.175 7.695 ;
        RECT 68.725 7.525 68.895 7.695 ;
        RECT 69.085 7.525 69.255 7.695 ;
        RECT 69.445 7.525 69.615 7.695 ;
        RECT 69.805 7.525 69.975 7.695 ;
        RECT 70.165 7.525 70.335 7.695 ;
        RECT 70.525 7.525 70.695 7.695 ;
        RECT 71.015 7.525 71.185 7.695 ;
        RECT 71.375 7.525 71.545 7.695 ;
        RECT 71.735 7.525 71.905 7.695 ;
        RECT 72.095 7.525 72.265 7.695 ;
        RECT 72.455 7.525 72.625 7.695 ;
        RECT 72.815 7.525 72.985 7.695 ;
        RECT 73.535 7.525 73.705 7.695 ;
        RECT 73.895 7.525 74.065 7.695 ;
        RECT 74.255 7.525 74.425 7.695 ;
        RECT 74.615 7.525 74.785 7.695 ;
        RECT 75.065 7.525 75.235 7.695 ;
        RECT 75.425 7.525 75.595 7.695 ;
        RECT 75.785 7.525 75.955 7.695 ;
        RECT 76.145 7.525 76.315 7.695 ;
        RECT 76.865 7.525 77.035 7.695 ;
        RECT 77.225 7.525 77.395 7.695 ;
        RECT 77.585 7.525 77.755 7.695 ;
        RECT 77.945 7.525 78.115 7.695 ;
        RECT 78.395 7.525 78.565 7.695 ;
        RECT 78.755 7.525 78.925 7.695 ;
        RECT 79.115 7.525 79.285 7.695 ;
        RECT 79.475 7.525 79.645 7.695 ;
        RECT 80.195 7.525 80.365 7.695 ;
        RECT 80.555 7.525 80.725 7.695 ;
        RECT 80.915 7.525 81.085 7.695 ;
        RECT 81.275 7.525 81.445 7.695 ;
        RECT 81.725 7.525 81.895 7.695 ;
        RECT 82.085 7.525 82.255 7.695 ;
        RECT 82.445 7.525 82.615 7.695 ;
        RECT 82.805 7.525 82.975 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 83.405 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 59.995197 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 83.535 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 3.045 -0.075 3.615 -0.065 ;
        RECT 7.855 -0.075 8.425 -0.065 ;
        RECT 12.665 -0.075 13.235 -0.065 ;
        RECT 15.995 -0.075 16.565 -0.065 ;
        RECT 19.325 -0.075 19.895 -0.065 ;
        RECT 24.135 -0.075 24.705 -0.065 ;
        RECT 27.465 -0.075 28.035 -0.065 ;
        RECT 32.275 -0.075 32.845 -0.065 ;
        RECT 37.085 -0.075 37.655 -0.065 ;
        RECT 40.415 -0.075 40.985 -0.065 ;
        RECT 43.745 -0.075 44.315 -0.065 ;
        RECT 48.555 -0.075 49.125 -0.065 ;
        RECT 51.885 -0.075 52.455 -0.065 ;
        RECT 56.695 -0.075 57.265 -0.065 ;
        RECT 61.505 -0.075 62.075 -0.065 ;
        RECT 64.835 -0.075 65.405 -0.065 ;
        RECT 68.165 -0.075 68.735 -0.065 ;
        RECT 72.975 -0.075 73.545 -0.065 ;
        RECT 76.305 -0.075 76.875 -0.065 ;
        RECT 79.635 -0.075 80.205 -0.065 ;
        RECT 82.965 -0.075 83.535 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 1.095 0.310 1.265 1.260 ;
        RECT 3.175 0.310 3.485 2.860 ;
        RECT 4.320 0.310 4.490 1.270 ;
        RECT 7.985 0.310 8.295 2.860 ;
        RECT 9.130 0.310 9.300 1.270 ;
        RECT 12.795 0.310 13.105 2.860 ;
        RECT 14.045 0.310 14.215 1.260 ;
        RECT 16.125 0.310 16.435 2.860 ;
        RECT 17.375 0.310 17.545 1.260 ;
        RECT 19.455 0.310 19.765 2.860 ;
        RECT 20.600 0.310 20.770 1.270 ;
        RECT 24.265 0.310 24.575 2.860 ;
        RECT 25.515 0.310 25.685 1.260 ;
        RECT 27.595 0.310 27.905 2.860 ;
        RECT 28.740 0.310 28.910 1.270 ;
        RECT 32.405 0.310 32.715 2.860 ;
        RECT 33.550 0.310 33.720 1.270 ;
        RECT 37.215 0.310 37.525 2.860 ;
        RECT 38.465 0.310 38.635 1.260 ;
        RECT 40.545 0.310 40.855 2.860 ;
        RECT 41.795 0.310 41.965 1.260 ;
        RECT 43.875 0.310 44.185 2.860 ;
        RECT 45.020 0.310 45.190 1.270 ;
        RECT 48.685 0.310 48.995 2.860 ;
        RECT 49.935 0.310 50.105 1.260 ;
        RECT 52.015 0.310 52.325 2.860 ;
        RECT 53.160 0.310 53.330 1.270 ;
        RECT 56.825 0.310 57.135 2.860 ;
        RECT 57.970 0.310 58.140 1.270 ;
        RECT 61.635 0.310 61.945 2.860 ;
        RECT 62.885 0.310 63.055 1.260 ;
        RECT 64.965 0.310 65.275 2.860 ;
        RECT 66.215 0.310 66.385 1.260 ;
        RECT 68.295 0.310 68.605 2.860 ;
        RECT 69.440 0.310 69.610 1.270 ;
        RECT 73.105 0.310 73.415 2.860 ;
        RECT 74.355 0.310 74.525 1.260 ;
        RECT 76.435 0.310 76.745 2.860 ;
        RECT 77.685 0.310 77.855 1.260 ;
        RECT 79.765 0.310 80.075 2.860 ;
        RECT 81.015 0.310 81.185 1.260 ;
        RECT 83.095 0.310 83.405 2.860 ;
        RECT -0.155 0.235 78.655 0.310 ;
        RECT 78.825 0.235 83.405 0.310 ;
        RECT -0.155 0.000 83.405 0.235 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 0.995 0.065 1.165 0.235 ;
        RECT 1.355 0.065 1.525 0.235 ;
        RECT 1.805 0.065 1.975 0.235 ;
        RECT 2.165 0.065 2.335 0.235 ;
        RECT 2.525 0.065 2.695 0.235 ;
        RECT 2.885 0.065 3.055 0.235 ;
        RECT 3.605 0.065 3.775 0.235 ;
        RECT 3.965 0.065 4.135 0.235 ;
        RECT 4.325 0.065 4.495 0.235 ;
        RECT 4.685 0.065 4.855 0.235 ;
        RECT 5.045 0.065 5.215 0.235 ;
        RECT 5.405 0.065 5.575 0.235 ;
        RECT 5.895 0.065 6.065 0.235 ;
        RECT 6.255 0.065 6.425 0.235 ;
        RECT 6.615 0.065 6.785 0.235 ;
        RECT 6.975 0.065 7.145 0.235 ;
        RECT 7.335 0.065 7.505 0.235 ;
        RECT 7.695 0.065 7.865 0.235 ;
        RECT 8.415 0.065 8.585 0.235 ;
        RECT 8.775 0.065 8.945 0.235 ;
        RECT 9.135 0.065 9.305 0.235 ;
        RECT 9.495 0.065 9.665 0.235 ;
        RECT 9.855 0.065 10.025 0.235 ;
        RECT 10.215 0.065 10.385 0.235 ;
        RECT 10.705 0.065 10.875 0.235 ;
        RECT 11.065 0.065 11.235 0.235 ;
        RECT 11.425 0.065 11.595 0.235 ;
        RECT 11.785 0.065 11.955 0.235 ;
        RECT 12.145 0.065 12.315 0.235 ;
        RECT 12.505 0.065 12.675 0.235 ;
        RECT 13.225 0.065 13.395 0.235 ;
        RECT 13.585 0.065 13.755 0.235 ;
        RECT 13.945 0.065 14.115 0.235 ;
        RECT 14.305 0.065 14.475 0.235 ;
        RECT 14.755 0.065 14.925 0.235 ;
        RECT 15.115 0.065 15.285 0.235 ;
        RECT 15.475 0.065 15.645 0.235 ;
        RECT 15.835 0.065 16.005 0.235 ;
        RECT 16.555 0.065 16.725 0.235 ;
        RECT 16.915 0.065 17.085 0.235 ;
        RECT 17.275 0.065 17.445 0.235 ;
        RECT 17.635 0.065 17.805 0.235 ;
        RECT 18.085 0.065 18.255 0.235 ;
        RECT 18.445 0.065 18.615 0.235 ;
        RECT 18.805 0.065 18.975 0.235 ;
        RECT 19.165 0.065 19.335 0.235 ;
        RECT 19.885 0.065 20.055 0.235 ;
        RECT 20.245 0.065 20.415 0.235 ;
        RECT 20.605 0.065 20.775 0.235 ;
        RECT 20.965 0.065 21.135 0.235 ;
        RECT 21.325 0.065 21.495 0.235 ;
        RECT 21.685 0.065 21.855 0.235 ;
        RECT 22.175 0.065 22.345 0.235 ;
        RECT 22.535 0.065 22.705 0.235 ;
        RECT 22.895 0.065 23.065 0.235 ;
        RECT 23.255 0.065 23.425 0.235 ;
        RECT 23.615 0.065 23.785 0.235 ;
        RECT 23.975 0.065 24.145 0.235 ;
        RECT 24.695 0.065 24.865 0.235 ;
        RECT 25.055 0.065 25.225 0.235 ;
        RECT 25.415 0.065 25.585 0.235 ;
        RECT 25.775 0.065 25.945 0.235 ;
        RECT 26.225 0.065 26.395 0.235 ;
        RECT 26.585 0.065 26.755 0.235 ;
        RECT 26.945 0.065 27.115 0.235 ;
        RECT 27.305 0.065 27.475 0.235 ;
        RECT 28.025 0.065 28.195 0.235 ;
        RECT 28.385 0.065 28.555 0.235 ;
        RECT 28.745 0.065 28.915 0.235 ;
        RECT 29.105 0.065 29.275 0.235 ;
        RECT 29.465 0.065 29.635 0.235 ;
        RECT 29.825 0.065 29.995 0.235 ;
        RECT 30.315 0.065 30.485 0.235 ;
        RECT 30.675 0.065 30.845 0.235 ;
        RECT 31.035 0.065 31.205 0.235 ;
        RECT 31.395 0.065 31.565 0.235 ;
        RECT 31.755 0.065 31.925 0.235 ;
        RECT 32.115 0.065 32.285 0.235 ;
        RECT 32.835 0.065 33.005 0.235 ;
        RECT 33.195 0.065 33.365 0.235 ;
        RECT 33.555 0.065 33.725 0.235 ;
        RECT 33.915 0.065 34.085 0.235 ;
        RECT 34.275 0.065 34.445 0.235 ;
        RECT 34.635 0.065 34.805 0.235 ;
        RECT 35.125 0.065 35.295 0.235 ;
        RECT 35.485 0.065 35.655 0.235 ;
        RECT 35.845 0.065 36.015 0.235 ;
        RECT 36.205 0.065 36.375 0.235 ;
        RECT 36.565 0.065 36.735 0.235 ;
        RECT 36.925 0.065 37.095 0.235 ;
        RECT 37.645 0.065 37.815 0.235 ;
        RECT 38.005 0.065 38.175 0.235 ;
        RECT 38.365 0.065 38.535 0.235 ;
        RECT 38.725 0.065 38.895 0.235 ;
        RECT 39.175 0.065 39.345 0.235 ;
        RECT 39.535 0.065 39.705 0.235 ;
        RECT 39.895 0.065 40.065 0.235 ;
        RECT 40.255 0.065 40.425 0.235 ;
        RECT 40.975 0.065 41.145 0.235 ;
        RECT 41.335 0.065 41.505 0.235 ;
        RECT 41.695 0.065 41.865 0.235 ;
        RECT 42.055 0.065 42.225 0.235 ;
        RECT 42.505 0.065 42.675 0.235 ;
        RECT 42.865 0.065 43.035 0.235 ;
        RECT 43.225 0.065 43.395 0.235 ;
        RECT 43.585 0.065 43.755 0.235 ;
        RECT 44.305 0.065 44.475 0.235 ;
        RECT 44.665 0.065 44.835 0.235 ;
        RECT 45.025 0.065 45.195 0.235 ;
        RECT 45.385 0.065 45.555 0.235 ;
        RECT 45.745 0.065 45.915 0.235 ;
        RECT 46.105 0.065 46.275 0.235 ;
        RECT 46.595 0.065 46.765 0.235 ;
        RECT 46.955 0.065 47.125 0.235 ;
        RECT 47.315 0.065 47.485 0.235 ;
        RECT 47.675 0.065 47.845 0.235 ;
        RECT 48.035 0.065 48.205 0.235 ;
        RECT 48.395 0.065 48.565 0.235 ;
        RECT 49.115 0.065 49.285 0.235 ;
        RECT 49.475 0.065 49.645 0.235 ;
        RECT 49.835 0.065 50.005 0.235 ;
        RECT 50.195 0.065 50.365 0.235 ;
        RECT 50.645 0.065 50.815 0.235 ;
        RECT 51.005 0.065 51.175 0.235 ;
        RECT 51.365 0.065 51.535 0.235 ;
        RECT 51.725 0.065 51.895 0.235 ;
        RECT 52.445 0.065 52.615 0.235 ;
        RECT 52.805 0.065 52.975 0.235 ;
        RECT 53.165 0.065 53.335 0.235 ;
        RECT 53.525 0.065 53.695 0.235 ;
        RECT 53.885 0.065 54.055 0.235 ;
        RECT 54.245 0.065 54.415 0.235 ;
        RECT 54.735 0.065 54.905 0.235 ;
        RECT 55.095 0.065 55.265 0.235 ;
        RECT 55.455 0.065 55.625 0.235 ;
        RECT 55.815 0.065 55.985 0.235 ;
        RECT 56.175 0.065 56.345 0.235 ;
        RECT 56.535 0.065 56.705 0.235 ;
        RECT 57.255 0.065 57.425 0.235 ;
        RECT 57.615 0.065 57.785 0.235 ;
        RECT 57.975 0.065 58.145 0.235 ;
        RECT 58.335 0.065 58.505 0.235 ;
        RECT 58.695 0.065 58.865 0.235 ;
        RECT 59.055 0.065 59.225 0.235 ;
        RECT 59.545 0.065 59.715 0.235 ;
        RECT 59.905 0.065 60.075 0.235 ;
        RECT 60.265 0.065 60.435 0.235 ;
        RECT 60.625 0.065 60.795 0.235 ;
        RECT 60.985 0.065 61.155 0.235 ;
        RECT 61.345 0.065 61.515 0.235 ;
        RECT 62.065 0.065 62.235 0.235 ;
        RECT 62.425 0.065 62.595 0.235 ;
        RECT 62.785 0.065 62.955 0.235 ;
        RECT 63.145 0.065 63.315 0.235 ;
        RECT 63.595 0.065 63.765 0.235 ;
        RECT 63.955 0.065 64.125 0.235 ;
        RECT 64.315 0.065 64.485 0.235 ;
        RECT 64.675 0.065 64.845 0.235 ;
        RECT 65.395 0.065 65.565 0.235 ;
        RECT 65.755 0.065 65.925 0.235 ;
        RECT 66.115 0.065 66.285 0.235 ;
        RECT 66.475 0.065 66.645 0.235 ;
        RECT 66.925 0.065 67.095 0.235 ;
        RECT 67.285 0.065 67.455 0.235 ;
        RECT 67.645 0.065 67.815 0.235 ;
        RECT 68.005 0.065 68.175 0.235 ;
        RECT 68.725 0.065 68.895 0.235 ;
        RECT 69.085 0.065 69.255 0.235 ;
        RECT 69.445 0.065 69.615 0.235 ;
        RECT 69.805 0.065 69.975 0.235 ;
        RECT 70.165 0.065 70.335 0.235 ;
        RECT 70.525 0.065 70.695 0.235 ;
        RECT 71.015 0.065 71.185 0.235 ;
        RECT 71.375 0.065 71.545 0.235 ;
        RECT 71.735 0.065 71.905 0.235 ;
        RECT 72.095 0.065 72.265 0.235 ;
        RECT 72.455 0.065 72.625 0.235 ;
        RECT 72.815 0.065 72.985 0.235 ;
        RECT 73.535 0.065 73.705 0.235 ;
        RECT 73.895 0.065 74.065 0.235 ;
        RECT 74.255 0.065 74.425 0.235 ;
        RECT 74.615 0.065 74.785 0.235 ;
        RECT 75.065 0.065 75.235 0.235 ;
        RECT 75.425 0.065 75.595 0.235 ;
        RECT 75.785 0.065 75.955 0.235 ;
        RECT 76.145 0.065 76.315 0.235 ;
        RECT 76.865 0.065 77.035 0.235 ;
        RECT 77.225 0.065 77.395 0.235 ;
        RECT 77.585 0.065 77.755 0.235 ;
        RECT 77.945 0.065 78.115 0.235 ;
        RECT 78.395 0.065 78.565 0.235 ;
        RECT 78.755 0.065 78.925 0.235 ;
        RECT 79.115 0.065 79.285 0.235 ;
        RECT 79.475 0.065 79.645 0.235 ;
        RECT 80.195 0.065 80.365 0.235 ;
        RECT 80.555 0.065 80.725 0.235 ;
        RECT 80.915 0.065 81.085 0.235 ;
        RECT 81.275 0.065 81.445 0.235 ;
        RECT 81.725 0.065 81.895 0.235 ;
        RECT 82.085 0.065 82.255 0.235 ;
        RECT 82.445 0.065 82.615 0.235 ;
        RECT 82.805 0.065 82.975 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 83.405 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 1.145 5.515 1.315 7.250 ;
        RECT 2.025 5.515 2.195 7.250 ;
        RECT 1.145 5.345 2.675 5.515 ;
        RECT 1.795 4.940 1.965 5.095 ;
        RECT 1.765 4.765 1.965 4.940 ;
        RECT 1.765 2.055 1.935 4.765 ;
        RECT 0.610 1.805 0.780 1.885 ;
        RECT 1.580 1.805 1.750 1.885 ;
        RECT 2.505 1.880 2.675 5.345 ;
        RECT 4.775 5.470 4.945 7.250 ;
        RECT 5.655 5.470 5.825 7.250 ;
        RECT 6.535 5.470 6.705 7.250 ;
        RECT 9.585 5.470 9.755 7.250 ;
        RECT 10.465 5.470 10.635 7.250 ;
        RECT 11.345 5.470 11.515 7.250 ;
        RECT 14.095 5.515 14.265 7.250 ;
        RECT 14.975 5.515 15.145 7.250 ;
        RECT 17.425 5.515 17.595 7.250 ;
        RECT 18.305 5.515 18.475 7.250 ;
        RECT 4.775 5.300 7.485 5.470 ;
        RECT 9.585 5.300 12.295 5.470 ;
        RECT 14.095 5.345 15.625 5.515 ;
        RECT 17.425 5.345 18.955 5.515 ;
        RECT 4.355 2.055 4.525 5.095 ;
        RECT 6.575 2.055 6.745 5.095 ;
        RECT 7.315 4.605 7.485 5.300 ;
        RECT 7.310 4.275 7.485 4.605 ;
        RECT 0.610 1.635 1.750 1.805 ;
        RECT 0.610 0.505 0.780 1.635 ;
        RECT 1.580 0.755 1.750 1.635 ;
        RECT 2.065 1.710 2.675 1.880 ;
        RECT 3.835 1.815 4.005 1.895 ;
        RECT 4.805 1.815 4.975 1.895 ;
        RECT 5.775 1.815 5.945 1.895 ;
        RECT 2.065 0.975 2.235 1.710 ;
        RECT 3.835 1.645 5.945 1.815 ;
        RECT 2.550 0.755 2.720 1.525 ;
        RECT 1.580 0.585 2.720 0.755 ;
        RECT 1.580 0.505 1.750 0.585 ;
        RECT 2.550 0.505 2.720 0.585 ;
        RECT 3.835 0.515 4.005 1.645 ;
        RECT 4.805 0.765 4.975 1.645 ;
        RECT 5.775 1.565 5.945 1.645 ;
        RECT 5.295 1.220 5.465 1.300 ;
        RECT 6.345 1.220 6.515 1.895 ;
        RECT 7.315 1.890 7.485 4.275 ;
        RECT 9.165 2.055 9.335 5.095 ;
        RECT 11.385 2.055 11.555 5.095 ;
        RECT 5.295 1.050 6.515 1.220 ;
        RECT 5.295 0.970 5.465 1.050 ;
        RECT 5.775 0.765 5.945 0.845 ;
        RECT 4.805 0.595 5.945 0.765 ;
        RECT 4.805 0.515 4.975 0.595 ;
        RECT 5.775 0.515 5.945 0.595 ;
        RECT 6.345 0.765 6.515 1.050 ;
        RECT 6.830 1.720 7.485 1.890 ;
        RECT 8.645 1.815 8.815 1.895 ;
        RECT 9.615 1.815 9.785 1.895 ;
        RECT 10.585 1.815 10.755 1.895 ;
        RECT 6.830 0.985 7.000 1.720 ;
        RECT 8.645 1.645 10.755 1.815 ;
        RECT 7.315 0.765 7.485 1.535 ;
        RECT 6.345 0.595 7.485 0.765 ;
        RECT 6.345 0.515 6.515 0.595 ;
        RECT 7.315 0.515 7.485 0.595 ;
        RECT 8.645 0.515 8.815 1.645 ;
        RECT 9.615 0.765 9.785 1.645 ;
        RECT 10.585 1.565 10.755 1.645 ;
        RECT 10.105 1.220 10.275 1.300 ;
        RECT 11.155 1.220 11.325 1.895 ;
        RECT 12.125 1.890 12.295 5.300 ;
        RECT 13.975 2.055 14.145 5.095 ;
        RECT 10.105 1.050 11.325 1.220 ;
        RECT 10.105 0.970 10.275 1.050 ;
        RECT 10.585 0.765 10.755 0.845 ;
        RECT 9.615 0.595 10.755 0.765 ;
        RECT 9.615 0.515 9.785 0.595 ;
        RECT 10.585 0.515 10.755 0.595 ;
        RECT 11.155 0.765 11.325 1.050 ;
        RECT 11.640 1.720 12.295 1.890 ;
        RECT 13.560 1.805 13.730 1.885 ;
        RECT 14.530 1.805 14.700 1.885 ;
        RECT 15.455 1.880 15.625 5.345 ;
        RECT 17.305 2.055 17.475 5.095 ;
        RECT 18.075 4.940 18.245 5.095 ;
        RECT 18.045 4.765 18.245 4.940 ;
        RECT 18.045 2.055 18.215 4.765 ;
        RECT 11.640 0.985 11.810 1.720 ;
        RECT 13.560 1.635 14.700 1.805 ;
        RECT 12.125 0.765 12.295 1.535 ;
        RECT 11.155 0.595 12.295 0.765 ;
        RECT 11.155 0.515 11.325 0.595 ;
        RECT 12.125 0.515 12.295 0.595 ;
        RECT 13.560 0.505 13.730 1.635 ;
        RECT 14.530 0.755 14.700 1.635 ;
        RECT 15.015 1.710 15.625 1.880 ;
        RECT 16.890 1.805 17.060 1.885 ;
        RECT 17.860 1.805 18.030 1.885 ;
        RECT 18.785 1.880 18.955 5.345 ;
        RECT 21.055 5.470 21.225 7.250 ;
        RECT 21.935 5.470 22.105 7.250 ;
        RECT 22.815 5.470 22.985 7.250 ;
        RECT 25.565 5.515 25.735 7.250 ;
        RECT 26.445 5.515 26.615 7.250 ;
        RECT 21.055 5.300 23.765 5.470 ;
        RECT 25.565 5.345 27.095 5.515 ;
        RECT 20.635 2.055 20.805 5.095 ;
        RECT 22.855 2.055 23.025 5.095 ;
        RECT 15.015 0.975 15.185 1.710 ;
        RECT 16.890 1.635 18.030 1.805 ;
        RECT 15.500 0.755 15.670 1.525 ;
        RECT 14.530 0.585 15.670 0.755 ;
        RECT 14.530 0.505 14.700 0.585 ;
        RECT 15.500 0.505 15.670 0.585 ;
        RECT 16.890 0.505 17.060 1.635 ;
        RECT 17.860 0.755 18.030 1.635 ;
        RECT 18.345 1.710 18.955 1.880 ;
        RECT 20.115 1.815 20.285 1.895 ;
        RECT 21.085 1.815 21.255 1.895 ;
        RECT 22.055 1.815 22.225 1.895 ;
        RECT 18.345 0.975 18.515 1.710 ;
        RECT 20.115 1.645 22.225 1.815 ;
        RECT 18.830 0.755 19.000 1.525 ;
        RECT 17.860 0.585 19.000 0.755 ;
        RECT 17.860 0.505 18.030 0.585 ;
        RECT 18.830 0.505 19.000 0.585 ;
        RECT 20.115 0.515 20.285 1.645 ;
        RECT 21.085 0.765 21.255 1.645 ;
        RECT 22.055 1.565 22.225 1.645 ;
        RECT 21.575 1.220 21.745 1.300 ;
        RECT 22.625 1.220 22.795 1.895 ;
        RECT 23.595 1.890 23.765 5.300 ;
        RECT 26.215 4.940 26.385 5.095 ;
        RECT 26.185 4.765 26.385 4.940 ;
        RECT 26.185 2.055 26.355 4.765 ;
        RECT 21.575 1.050 22.795 1.220 ;
        RECT 21.575 0.970 21.745 1.050 ;
        RECT 22.055 0.765 22.225 0.845 ;
        RECT 21.085 0.595 22.225 0.765 ;
        RECT 21.085 0.515 21.255 0.595 ;
        RECT 22.055 0.515 22.225 0.595 ;
        RECT 22.625 0.765 22.795 1.050 ;
        RECT 23.110 1.720 23.765 1.890 ;
        RECT 25.030 1.805 25.200 1.885 ;
        RECT 26.000 1.805 26.170 1.885 ;
        RECT 26.925 1.880 27.095 5.345 ;
        RECT 29.195 5.470 29.365 7.250 ;
        RECT 30.075 5.470 30.245 7.250 ;
        RECT 30.955 5.470 31.125 7.250 ;
        RECT 34.005 5.470 34.175 7.250 ;
        RECT 34.885 5.470 35.055 7.250 ;
        RECT 35.765 5.470 35.935 7.250 ;
        RECT 38.515 5.515 38.685 7.250 ;
        RECT 39.395 5.515 39.565 7.250 ;
        RECT 41.845 5.515 42.015 7.250 ;
        RECT 42.725 5.515 42.895 7.250 ;
        RECT 29.195 5.300 31.905 5.470 ;
        RECT 34.005 5.300 36.715 5.470 ;
        RECT 38.515 5.345 40.045 5.515 ;
        RECT 41.845 5.345 43.375 5.515 ;
        RECT 28.775 2.055 28.945 5.095 ;
        RECT 30.995 2.055 31.165 5.095 ;
        RECT 31.735 4.605 31.905 5.300 ;
        RECT 31.730 4.275 31.905 4.605 ;
        RECT 23.110 0.985 23.280 1.720 ;
        RECT 25.030 1.635 26.170 1.805 ;
        RECT 23.595 0.765 23.765 1.535 ;
        RECT 22.625 0.595 23.765 0.765 ;
        RECT 22.625 0.515 22.795 0.595 ;
        RECT 23.595 0.515 23.765 0.595 ;
        RECT 25.030 0.505 25.200 1.635 ;
        RECT 26.000 0.755 26.170 1.635 ;
        RECT 26.485 1.710 27.095 1.880 ;
        RECT 28.255 1.815 28.425 1.895 ;
        RECT 29.225 1.815 29.395 1.895 ;
        RECT 30.195 1.815 30.365 1.895 ;
        RECT 26.485 0.975 26.655 1.710 ;
        RECT 28.255 1.645 30.365 1.815 ;
        RECT 26.970 0.755 27.140 1.525 ;
        RECT 26.000 0.585 27.140 0.755 ;
        RECT 26.000 0.505 26.170 0.585 ;
        RECT 26.970 0.505 27.140 0.585 ;
        RECT 28.255 0.515 28.425 1.645 ;
        RECT 29.225 0.765 29.395 1.645 ;
        RECT 30.195 1.565 30.365 1.645 ;
        RECT 29.715 1.220 29.885 1.300 ;
        RECT 30.765 1.220 30.935 1.895 ;
        RECT 31.735 1.890 31.905 4.275 ;
        RECT 33.585 2.055 33.755 5.095 ;
        RECT 35.805 2.055 35.975 5.095 ;
        RECT 29.715 1.050 30.935 1.220 ;
        RECT 29.715 0.970 29.885 1.050 ;
        RECT 30.195 0.765 30.365 0.845 ;
        RECT 29.225 0.595 30.365 0.765 ;
        RECT 29.225 0.515 29.395 0.595 ;
        RECT 30.195 0.515 30.365 0.595 ;
        RECT 30.765 0.765 30.935 1.050 ;
        RECT 31.250 1.720 31.905 1.890 ;
        RECT 33.065 1.815 33.235 1.895 ;
        RECT 34.035 1.815 34.205 1.895 ;
        RECT 35.005 1.815 35.175 1.895 ;
        RECT 31.250 0.985 31.420 1.720 ;
        RECT 33.065 1.645 35.175 1.815 ;
        RECT 31.735 0.765 31.905 1.535 ;
        RECT 30.765 0.595 31.905 0.765 ;
        RECT 30.765 0.515 30.935 0.595 ;
        RECT 31.735 0.515 31.905 0.595 ;
        RECT 33.065 0.515 33.235 1.645 ;
        RECT 34.035 0.765 34.205 1.645 ;
        RECT 35.005 1.565 35.175 1.645 ;
        RECT 34.525 1.220 34.695 1.300 ;
        RECT 35.575 1.220 35.745 1.895 ;
        RECT 36.545 1.890 36.715 5.300 ;
        RECT 38.395 2.055 38.565 5.095 ;
        RECT 34.525 1.050 35.745 1.220 ;
        RECT 34.525 0.970 34.695 1.050 ;
        RECT 35.005 0.765 35.175 0.845 ;
        RECT 34.035 0.595 35.175 0.765 ;
        RECT 34.035 0.515 34.205 0.595 ;
        RECT 35.005 0.515 35.175 0.595 ;
        RECT 35.575 0.765 35.745 1.050 ;
        RECT 36.060 1.720 36.715 1.890 ;
        RECT 37.980 1.805 38.150 1.885 ;
        RECT 38.950 1.805 39.120 1.885 ;
        RECT 39.875 1.880 40.045 5.345 ;
        RECT 41.725 2.055 41.895 5.095 ;
        RECT 42.495 4.940 42.665 5.095 ;
        RECT 42.465 4.765 42.665 4.940 ;
        RECT 42.465 2.055 42.635 4.765 ;
        RECT 36.060 0.985 36.230 1.720 ;
        RECT 37.980 1.635 39.120 1.805 ;
        RECT 36.545 0.765 36.715 1.535 ;
        RECT 35.575 0.595 36.715 0.765 ;
        RECT 35.575 0.515 35.745 0.595 ;
        RECT 36.545 0.515 36.715 0.595 ;
        RECT 37.980 0.505 38.150 1.635 ;
        RECT 38.950 0.755 39.120 1.635 ;
        RECT 39.435 1.710 40.045 1.880 ;
        RECT 41.310 1.805 41.480 1.885 ;
        RECT 42.280 1.805 42.450 1.885 ;
        RECT 43.205 1.880 43.375 5.345 ;
        RECT 45.475 5.470 45.645 7.250 ;
        RECT 46.355 5.470 46.525 7.250 ;
        RECT 47.235 5.470 47.405 7.250 ;
        RECT 49.985 5.515 50.155 7.250 ;
        RECT 50.865 5.515 51.035 7.250 ;
        RECT 45.475 5.300 48.185 5.470 ;
        RECT 49.985 5.345 51.515 5.515 ;
        RECT 45.055 2.055 45.225 5.095 ;
        RECT 47.275 2.055 47.445 5.095 ;
        RECT 39.435 0.975 39.605 1.710 ;
        RECT 41.310 1.635 42.450 1.805 ;
        RECT 39.920 0.755 40.090 1.525 ;
        RECT 38.950 0.585 40.090 0.755 ;
        RECT 38.950 0.505 39.120 0.585 ;
        RECT 39.920 0.505 40.090 0.585 ;
        RECT 41.310 0.505 41.480 1.635 ;
        RECT 42.280 0.755 42.450 1.635 ;
        RECT 42.765 1.710 43.375 1.880 ;
        RECT 44.535 1.815 44.705 1.895 ;
        RECT 45.505 1.815 45.675 1.895 ;
        RECT 46.475 1.815 46.645 1.895 ;
        RECT 42.765 0.975 42.935 1.710 ;
        RECT 44.535 1.645 46.645 1.815 ;
        RECT 43.250 0.755 43.420 1.525 ;
        RECT 42.280 0.585 43.420 0.755 ;
        RECT 42.280 0.505 42.450 0.585 ;
        RECT 43.250 0.505 43.420 0.585 ;
        RECT 44.535 0.515 44.705 1.645 ;
        RECT 45.505 0.765 45.675 1.645 ;
        RECT 46.475 1.565 46.645 1.645 ;
        RECT 45.995 1.220 46.165 1.300 ;
        RECT 47.045 1.220 47.215 1.895 ;
        RECT 48.015 1.890 48.185 5.300 ;
        RECT 50.635 4.940 50.805 5.095 ;
        RECT 50.605 4.765 50.805 4.940 ;
        RECT 50.605 2.055 50.775 4.765 ;
        RECT 45.995 1.050 47.215 1.220 ;
        RECT 45.995 0.970 46.165 1.050 ;
        RECT 46.475 0.765 46.645 0.845 ;
        RECT 45.505 0.595 46.645 0.765 ;
        RECT 45.505 0.515 45.675 0.595 ;
        RECT 46.475 0.515 46.645 0.595 ;
        RECT 47.045 0.765 47.215 1.050 ;
        RECT 47.530 1.720 48.185 1.890 ;
        RECT 49.450 1.805 49.620 1.885 ;
        RECT 50.420 1.805 50.590 1.885 ;
        RECT 51.345 1.880 51.515 5.345 ;
        RECT 53.615 5.470 53.785 7.250 ;
        RECT 54.495 5.470 54.665 7.250 ;
        RECT 55.375 5.470 55.545 7.250 ;
        RECT 58.425 5.470 58.595 7.250 ;
        RECT 59.305 5.470 59.475 7.250 ;
        RECT 60.185 5.470 60.355 7.250 ;
        RECT 62.935 5.515 63.105 7.250 ;
        RECT 63.815 5.515 63.985 7.250 ;
        RECT 66.265 5.515 66.435 7.250 ;
        RECT 67.145 5.515 67.315 7.250 ;
        RECT 53.615 5.300 56.325 5.470 ;
        RECT 58.425 5.300 61.135 5.470 ;
        RECT 62.935 5.345 64.465 5.515 ;
        RECT 66.265 5.345 67.795 5.515 ;
        RECT 53.195 2.055 53.365 5.095 ;
        RECT 55.415 2.055 55.585 5.095 ;
        RECT 56.155 4.605 56.325 5.300 ;
        RECT 56.150 4.275 56.325 4.605 ;
        RECT 47.530 0.985 47.700 1.720 ;
        RECT 49.450 1.635 50.590 1.805 ;
        RECT 48.015 0.765 48.185 1.535 ;
        RECT 47.045 0.595 48.185 0.765 ;
        RECT 47.045 0.515 47.215 0.595 ;
        RECT 48.015 0.515 48.185 0.595 ;
        RECT 49.450 0.505 49.620 1.635 ;
        RECT 50.420 0.755 50.590 1.635 ;
        RECT 50.905 1.710 51.515 1.880 ;
        RECT 52.675 1.815 52.845 1.895 ;
        RECT 53.645 1.815 53.815 1.895 ;
        RECT 54.615 1.815 54.785 1.895 ;
        RECT 50.905 0.975 51.075 1.710 ;
        RECT 52.675 1.645 54.785 1.815 ;
        RECT 51.390 0.755 51.560 1.525 ;
        RECT 50.420 0.585 51.560 0.755 ;
        RECT 50.420 0.505 50.590 0.585 ;
        RECT 51.390 0.505 51.560 0.585 ;
        RECT 52.675 0.515 52.845 1.645 ;
        RECT 53.645 0.765 53.815 1.645 ;
        RECT 54.615 1.565 54.785 1.645 ;
        RECT 54.135 1.220 54.305 1.300 ;
        RECT 55.185 1.220 55.355 1.895 ;
        RECT 56.155 1.890 56.325 4.275 ;
        RECT 58.005 2.055 58.175 5.095 ;
        RECT 60.225 2.055 60.395 5.095 ;
        RECT 54.135 1.050 55.355 1.220 ;
        RECT 54.135 0.970 54.305 1.050 ;
        RECT 54.615 0.765 54.785 0.845 ;
        RECT 53.645 0.595 54.785 0.765 ;
        RECT 53.645 0.515 53.815 0.595 ;
        RECT 54.615 0.515 54.785 0.595 ;
        RECT 55.185 0.765 55.355 1.050 ;
        RECT 55.670 1.720 56.325 1.890 ;
        RECT 57.485 1.815 57.655 1.895 ;
        RECT 58.455 1.815 58.625 1.895 ;
        RECT 59.425 1.815 59.595 1.895 ;
        RECT 55.670 0.985 55.840 1.720 ;
        RECT 57.485 1.645 59.595 1.815 ;
        RECT 56.155 0.765 56.325 1.535 ;
        RECT 55.185 0.595 56.325 0.765 ;
        RECT 55.185 0.515 55.355 0.595 ;
        RECT 56.155 0.515 56.325 0.595 ;
        RECT 57.485 0.515 57.655 1.645 ;
        RECT 58.455 0.765 58.625 1.645 ;
        RECT 59.425 1.565 59.595 1.645 ;
        RECT 58.945 1.220 59.115 1.300 ;
        RECT 59.995 1.220 60.165 1.895 ;
        RECT 60.965 1.890 61.135 5.300 ;
        RECT 62.815 2.055 62.985 5.095 ;
        RECT 58.945 1.050 60.165 1.220 ;
        RECT 58.945 0.970 59.115 1.050 ;
        RECT 59.425 0.765 59.595 0.845 ;
        RECT 58.455 0.595 59.595 0.765 ;
        RECT 58.455 0.515 58.625 0.595 ;
        RECT 59.425 0.515 59.595 0.595 ;
        RECT 59.995 0.765 60.165 1.050 ;
        RECT 60.480 1.720 61.135 1.890 ;
        RECT 62.400 1.805 62.570 1.885 ;
        RECT 63.370 1.805 63.540 1.885 ;
        RECT 64.295 1.880 64.465 5.345 ;
        RECT 66.145 2.055 66.315 5.095 ;
        RECT 66.915 4.940 67.085 5.095 ;
        RECT 66.885 4.765 67.085 4.940 ;
        RECT 66.885 2.055 67.055 4.765 ;
        RECT 60.480 0.985 60.650 1.720 ;
        RECT 62.400 1.635 63.540 1.805 ;
        RECT 60.965 0.765 61.135 1.535 ;
        RECT 59.995 0.595 61.135 0.765 ;
        RECT 59.995 0.515 60.165 0.595 ;
        RECT 60.965 0.515 61.135 0.595 ;
        RECT 62.400 0.505 62.570 1.635 ;
        RECT 63.370 0.755 63.540 1.635 ;
        RECT 63.855 1.710 64.465 1.880 ;
        RECT 65.730 1.805 65.900 1.885 ;
        RECT 66.700 1.805 66.870 1.885 ;
        RECT 67.625 1.880 67.795 5.345 ;
        RECT 69.895 5.470 70.065 7.250 ;
        RECT 70.775 5.470 70.945 7.250 ;
        RECT 71.655 5.470 71.825 7.250 ;
        RECT 74.405 7.055 74.585 7.225 ;
        RECT 74.405 5.525 74.575 7.055 ;
        RECT 75.285 5.525 75.455 7.225 ;
        RECT 69.895 5.300 72.605 5.470 ;
        RECT 74.405 5.355 75.455 5.525 ;
        RECT 69.475 2.055 69.645 5.095 ;
        RECT 71.695 2.055 71.865 5.095 ;
        RECT 63.855 0.975 64.025 1.710 ;
        RECT 65.730 1.635 66.870 1.805 ;
        RECT 64.340 0.755 64.510 1.525 ;
        RECT 63.370 0.585 64.510 0.755 ;
        RECT 63.370 0.505 63.540 0.585 ;
        RECT 64.340 0.505 64.510 0.585 ;
        RECT 65.730 0.505 65.900 1.635 ;
        RECT 66.700 0.755 66.870 1.635 ;
        RECT 67.185 1.710 67.795 1.880 ;
        RECT 68.955 1.815 69.125 1.895 ;
        RECT 69.925 1.815 70.095 1.895 ;
        RECT 70.895 1.815 71.065 1.895 ;
        RECT 67.185 0.975 67.355 1.710 ;
        RECT 68.955 1.645 71.065 1.815 ;
        RECT 67.670 0.755 67.840 1.525 ;
        RECT 66.700 0.585 67.840 0.755 ;
        RECT 66.700 0.505 66.870 0.585 ;
        RECT 67.670 0.505 67.840 0.585 ;
        RECT 68.955 0.515 69.125 1.645 ;
        RECT 69.925 0.765 70.095 1.645 ;
        RECT 70.895 1.565 71.065 1.645 ;
        RECT 70.415 1.220 70.585 1.300 ;
        RECT 71.465 1.220 71.635 1.895 ;
        RECT 72.435 1.890 72.605 5.300 ;
        RECT 75.285 5.275 75.455 5.355 ;
        RECT 77.285 7.055 79.215 7.225 ;
        RECT 77.285 5.275 77.455 7.055 ;
        RECT 77.725 5.525 77.895 6.795 ;
        RECT 78.165 5.785 78.335 7.055 ;
        RECT 78.605 5.525 78.775 6.795 ;
        RECT 79.045 5.605 79.215 7.055 ;
        RECT 80.625 7.055 82.555 7.225 ;
        RECT 77.725 5.355 78.775 5.525 ;
        RECT 78.605 5.275 78.775 5.355 ;
        RECT 80.625 5.275 80.795 7.055 ;
        RECT 81.505 5.785 81.675 7.055 ;
        RECT 82.385 5.785 82.555 7.055 ;
        RECT 73.915 2.055 74.085 5.100 ;
        RECT 75.065 4.940 75.235 5.100 ;
        RECT 75.025 4.770 75.235 4.940 ;
        RECT 75.025 2.055 75.195 4.770 ;
        RECT 77.615 2.055 77.785 5.100 ;
        RECT 79.095 2.055 79.265 5.100 ;
        RECT 80.575 2.055 80.745 5.100 ;
        RECT 81.685 4.770 81.875 5.100 ;
        RECT 81.685 2.055 81.855 4.770 ;
        RECT 70.415 1.050 71.635 1.220 ;
        RECT 70.415 0.970 70.585 1.050 ;
        RECT 70.895 0.765 71.065 0.845 ;
        RECT 69.925 0.595 71.065 0.765 ;
        RECT 69.925 0.515 70.095 0.595 ;
        RECT 70.895 0.515 71.065 0.595 ;
        RECT 71.465 0.765 71.635 1.050 ;
        RECT 71.950 1.720 72.605 1.890 ;
        RECT 73.870 1.805 74.040 1.885 ;
        RECT 74.840 1.805 75.010 1.885 ;
        RECT 71.950 0.985 72.120 1.720 ;
        RECT 73.870 1.635 75.010 1.805 ;
        RECT 72.435 0.765 72.605 1.535 ;
        RECT 71.465 0.595 72.605 0.765 ;
        RECT 71.465 0.515 71.635 0.595 ;
        RECT 72.435 0.515 72.605 0.595 ;
        RECT 73.870 0.505 74.040 1.635 ;
        RECT 74.840 0.755 75.010 1.635 ;
        RECT 75.810 0.755 75.980 1.885 ;
        RECT 74.840 0.585 75.980 0.755 ;
        RECT 74.840 0.505 75.010 0.585 ;
        RECT 75.810 0.505 75.980 0.585 ;
        RECT 77.200 1.805 77.370 1.885 ;
        RECT 78.170 1.805 78.340 1.885 ;
        RECT 77.200 1.635 78.340 1.805 ;
        RECT 77.200 0.505 77.370 1.635 ;
        RECT 78.170 0.755 78.340 1.635 ;
        RECT 79.140 0.755 79.310 1.885 ;
        RECT 78.170 0.585 79.310 0.755 ;
        RECT 78.170 0.505 78.340 0.585 ;
        RECT 79.140 0.505 79.310 0.585 ;
        RECT 80.530 1.805 80.700 1.885 ;
        RECT 81.500 1.805 81.670 1.885 ;
        RECT 80.530 1.635 81.670 1.805 ;
        RECT 80.530 0.505 80.700 1.635 ;
        RECT 81.500 0.755 81.670 1.635 ;
        RECT 82.470 0.755 82.640 1.530 ;
        RECT 81.500 0.585 82.640 0.755 ;
        RECT 81.500 0.505 81.670 0.585 ;
        RECT 82.470 0.505 82.640 0.585 ;
      LAYER mcon ;
        RECT 1.765 4.355 1.935 4.525 ;
        RECT 2.505 2.875 2.675 3.045 ;
        RECT 4.355 2.870 4.525 3.040 ;
        RECT 7.310 4.355 7.480 4.525 ;
        RECT 6.575 3.985 6.745 4.155 ;
        RECT 9.165 2.875 9.335 3.045 ;
        RECT 11.385 3.985 11.555 4.155 ;
        RECT 12.125 2.875 12.295 3.045 ;
        RECT 13.975 2.875 14.145 3.045 ;
        RECT 15.455 3.985 15.625 4.155 ;
        RECT 17.305 4.355 17.475 4.525 ;
        RECT 18.045 3.245 18.215 3.415 ;
        RECT 18.785 4.355 18.955 4.525 ;
        RECT 20.635 4.355 20.805 4.525 ;
        RECT 22.855 3.985 23.025 4.155 ;
        RECT 23.595 3.245 23.765 3.415 ;
        RECT 26.185 4.355 26.355 4.525 ;
        RECT 26.925 2.875 27.095 3.045 ;
        RECT 28.775 2.870 28.945 3.040 ;
        RECT 31.730 4.355 31.900 4.525 ;
        RECT 30.995 3.985 31.165 4.155 ;
        RECT 33.585 2.875 33.755 3.045 ;
        RECT 35.805 3.985 35.975 4.155 ;
        RECT 36.545 2.875 36.715 3.045 ;
        RECT 38.395 2.875 38.565 3.045 ;
        RECT 39.875 3.985 40.045 4.155 ;
        RECT 41.725 4.355 41.895 4.525 ;
        RECT 42.465 3.615 42.635 3.785 ;
        RECT 43.205 4.355 43.375 4.525 ;
        RECT 45.055 4.355 45.225 4.525 ;
        RECT 47.275 3.985 47.445 4.155 ;
        RECT 48.015 3.615 48.185 3.785 ;
        RECT 50.605 4.355 50.775 4.525 ;
        RECT 51.345 2.875 51.515 3.045 ;
        RECT 53.195 2.870 53.365 3.040 ;
        RECT 56.150 4.355 56.320 4.525 ;
        RECT 55.415 3.985 55.585 4.155 ;
        RECT 58.005 2.875 58.175 3.045 ;
        RECT 60.225 3.985 60.395 4.155 ;
        RECT 60.965 2.875 61.135 3.045 ;
        RECT 62.815 2.875 62.985 3.045 ;
        RECT 64.295 3.985 64.465 4.155 ;
        RECT 66.145 4.355 66.315 4.525 ;
        RECT 75.285 5.355 75.455 5.525 ;
        RECT 66.885 4.355 67.055 4.525 ;
        RECT 67.625 4.725 67.795 4.895 ;
        RECT 69.475 4.725 69.645 4.895 ;
        RECT 71.695 3.985 71.865 4.155 ;
        RECT 77.285 5.355 77.455 5.525 ;
        RECT 78.605 5.355 78.775 5.525 ;
        RECT 80.625 5.355 80.795 5.525 ;
        RECT 72.435 4.355 72.605 4.525 ;
        RECT 73.915 4.725 74.085 4.895 ;
        RECT 73.915 3.615 74.085 3.785 ;
        RECT 75.025 4.355 75.195 4.525 ;
        RECT 77.615 4.725 77.785 4.895 ;
        RECT 79.095 3.245 79.265 3.415 ;
        RECT 79.095 2.135 79.265 2.305 ;
        RECT 80.575 2.135 80.745 2.305 ;
        RECT 81.685 4.355 81.855 4.525 ;
      LAYER met1 ;
        RECT 75.255 5.525 75.485 5.555 ;
        RECT 77.255 5.525 77.485 5.555 ;
        RECT 78.575 5.525 78.805 5.555 ;
        RECT 80.595 5.525 80.825 5.555 ;
        RECT 75.225 5.355 77.515 5.525 ;
        RECT 78.545 5.355 80.855 5.525 ;
        RECT 75.255 5.325 75.485 5.355 ;
        RECT 77.255 5.325 77.485 5.355 ;
        RECT 78.575 5.325 78.805 5.355 ;
        RECT 80.595 5.325 80.825 5.355 ;
        RECT 67.595 4.895 67.825 4.925 ;
        RECT 69.445 4.895 69.675 4.925 ;
        RECT 73.885 4.895 74.115 4.925 ;
        RECT 77.585 4.895 77.815 4.925 ;
        RECT 67.565 4.725 69.705 4.895 ;
        RECT 73.855 4.725 77.845 4.895 ;
        RECT 67.595 4.695 67.825 4.725 ;
        RECT 69.445 4.695 69.675 4.725 ;
        RECT 73.885 4.695 74.115 4.725 ;
        RECT 77.585 4.695 77.815 4.725 ;
        RECT 1.735 4.525 1.965 4.555 ;
        RECT 7.280 4.525 7.510 4.555 ;
        RECT 17.275 4.525 17.505 4.555 ;
        RECT 18.755 4.525 18.985 4.555 ;
        RECT 20.605 4.525 20.835 4.555 ;
        RECT 26.155 4.525 26.385 4.555 ;
        RECT 31.700 4.525 31.930 4.555 ;
        RECT 41.695 4.525 41.925 4.555 ;
        RECT 43.175 4.525 43.405 4.555 ;
        RECT 45.025 4.525 45.255 4.555 ;
        RECT 50.575 4.525 50.805 4.555 ;
        RECT 56.120 4.525 56.350 4.555 ;
        RECT 66.115 4.525 66.345 4.555 ;
        RECT 66.855 4.525 67.085 4.555 ;
        RECT 72.405 4.525 72.635 4.555 ;
        RECT 74.995 4.525 75.225 4.555 ;
        RECT 81.655 4.525 81.885 4.555 ;
        RECT 1.705 4.355 17.535 4.525 ;
        RECT 18.725 4.355 20.865 4.525 ;
        RECT 26.125 4.355 41.955 4.525 ;
        RECT 43.145 4.355 45.285 4.525 ;
        RECT 50.545 4.355 66.375 4.525 ;
        RECT 66.825 4.355 81.915 4.525 ;
        RECT 1.735 4.325 1.965 4.355 ;
        RECT 7.280 4.325 7.510 4.355 ;
        RECT 17.275 4.325 17.505 4.355 ;
        RECT 18.755 4.325 18.985 4.355 ;
        RECT 20.605 4.325 20.835 4.355 ;
        RECT 26.155 4.325 26.385 4.355 ;
        RECT 31.700 4.325 31.930 4.355 ;
        RECT 41.695 4.325 41.925 4.355 ;
        RECT 43.175 4.325 43.405 4.355 ;
        RECT 45.025 4.325 45.255 4.355 ;
        RECT 50.575 4.325 50.805 4.355 ;
        RECT 56.120 4.325 56.350 4.355 ;
        RECT 66.115 4.325 66.345 4.355 ;
        RECT 66.855 4.325 67.085 4.355 ;
        RECT 72.405 4.325 72.635 4.355 ;
        RECT 74.995 4.325 75.225 4.355 ;
        RECT 81.655 4.325 81.885 4.355 ;
        RECT 6.545 4.155 6.775 4.185 ;
        RECT 11.355 4.155 11.585 4.185 ;
        RECT 15.425 4.155 15.655 4.185 ;
        RECT 22.825 4.155 23.055 4.185 ;
        RECT 30.965 4.155 31.195 4.185 ;
        RECT 35.775 4.155 36.005 4.185 ;
        RECT 39.845 4.155 40.075 4.185 ;
        RECT 47.245 4.155 47.475 4.185 ;
        RECT 55.385 4.155 55.615 4.185 ;
        RECT 60.195 4.155 60.425 4.185 ;
        RECT 64.265 4.155 64.495 4.185 ;
        RECT 71.665 4.155 71.895 4.185 ;
        RECT 6.515 3.985 23.085 4.155 ;
        RECT 30.935 3.985 47.505 4.155 ;
        RECT 55.355 3.985 71.925 4.155 ;
        RECT 6.545 3.955 6.775 3.985 ;
        RECT 11.355 3.955 11.585 3.985 ;
        RECT 15.425 3.955 15.655 3.985 ;
        RECT 22.825 3.955 23.055 3.985 ;
        RECT 30.965 3.955 31.195 3.985 ;
        RECT 35.775 3.955 36.005 3.985 ;
        RECT 39.845 3.955 40.075 3.985 ;
        RECT 47.245 3.955 47.475 3.985 ;
        RECT 55.385 3.955 55.615 3.985 ;
        RECT 60.195 3.955 60.425 3.985 ;
        RECT 64.265 3.955 64.495 3.985 ;
        RECT 71.665 3.955 71.895 3.985 ;
        RECT 42.435 3.785 42.665 3.815 ;
        RECT 47.985 3.785 48.215 3.815 ;
        RECT 73.885 3.785 74.115 3.815 ;
        RECT 42.405 3.615 74.145 3.785 ;
        RECT 42.435 3.585 42.665 3.615 ;
        RECT 47.985 3.585 48.215 3.615 ;
        RECT 73.885 3.585 74.115 3.615 ;
        RECT 18.015 3.415 18.245 3.445 ;
        RECT 23.565 3.415 23.795 3.445 ;
        RECT 79.065 3.415 79.295 3.445 ;
        RECT 17.985 3.245 79.325 3.415 ;
        RECT 18.015 3.215 18.245 3.245 ;
        RECT 23.565 3.215 23.795 3.245 ;
        RECT 79.065 3.215 79.295 3.245 ;
        RECT 2.475 3.045 2.705 3.075 ;
        RECT 4.325 3.045 4.555 3.070 ;
        RECT 9.135 3.045 9.365 3.075 ;
        RECT 12.095 3.045 12.325 3.075 ;
        RECT 13.945 3.045 14.175 3.075 ;
        RECT 26.895 3.045 27.125 3.075 ;
        RECT 28.745 3.045 28.975 3.070 ;
        RECT 33.555 3.045 33.785 3.075 ;
        RECT 36.515 3.045 36.745 3.075 ;
        RECT 38.365 3.045 38.595 3.075 ;
        RECT 51.315 3.045 51.545 3.075 ;
        RECT 53.165 3.045 53.395 3.070 ;
        RECT 57.975 3.045 58.205 3.075 ;
        RECT 60.935 3.045 61.165 3.075 ;
        RECT 62.785 3.045 63.015 3.075 ;
        RECT 2.445 2.875 9.395 3.045 ;
        RECT 12.065 2.875 14.205 3.045 ;
        RECT 26.865 2.875 33.815 3.045 ;
        RECT 36.485 2.875 38.625 3.045 ;
        RECT 51.285 2.875 58.235 3.045 ;
        RECT 60.905 2.875 63.045 3.045 ;
        RECT 2.475 2.845 2.705 2.875 ;
        RECT 4.295 2.870 4.705 2.875 ;
        RECT 4.325 2.840 4.555 2.870 ;
        RECT 9.135 2.845 9.365 2.875 ;
        RECT 12.095 2.845 12.325 2.875 ;
        RECT 13.945 2.845 14.175 2.875 ;
        RECT 26.895 2.845 27.125 2.875 ;
        RECT 28.715 2.870 29.125 2.875 ;
        RECT 28.745 2.840 28.975 2.870 ;
        RECT 33.555 2.845 33.785 2.875 ;
        RECT 36.515 2.845 36.745 2.875 ;
        RECT 38.365 2.845 38.595 2.875 ;
        RECT 51.315 2.845 51.545 2.875 ;
        RECT 53.135 2.870 53.545 2.875 ;
        RECT 53.165 2.840 53.395 2.870 ;
        RECT 57.975 2.845 58.205 2.875 ;
        RECT 60.935 2.845 61.165 2.875 ;
        RECT 62.785 2.845 63.015 2.875 ;
        RECT 79.065 2.305 79.295 2.335 ;
        RECT 80.545 2.305 80.775 2.335 ;
        RECT 79.035 2.135 80.805 2.305 ;
        RECT 79.065 2.105 79.295 2.135 ;
        RECT 80.545 2.105 80.775 2.135 ;
  END
END TMRDFFSNQNX1






MACRO TMRDFFSNQX1
  CLASS BLOCK ;
  FOREIGN TMRDFFSNQX1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 86.310 BY 7.950 ;
  PIN Q
    ANTENNADIFFAREA 0.771900 ;
    PORT
      LAYER li1 ;
        RECT 84.275 4.895 84.445 7.250 ;
        RECT 84.275 4.725 84.815 4.895 ;
        RECT 84.645 2.305 84.815 4.725 ;
        RECT 84.275 2.135 84.815 2.305 ;
        RECT 84.275 0.975 84.445 2.135 ;
      LAYER mcon ;
        RECT 84.645 3.985 84.815 4.155 ;
      LAYER met1 ;
        RECT 84.615 4.155 84.845 4.185 ;
        RECT 84.585 3.985 84.995 4.155 ;
        RECT 84.615 3.955 84.845 3.985 ;
    END
  END Q
  PIN D
    ANTENNAGATEAREA 3.099750 ;
    PORT
      LAYER li1 ;
        RECT 1.025 2.055 1.195 5.095 ;
        RECT 25.445 2.055 25.615 5.095 ;
        RECT 49.865 2.055 50.035 5.095 ;
      LAYER mcon ;
        RECT 1.025 2.135 1.195 2.305 ;
        RECT 25.445 2.135 25.615 2.305 ;
        RECT 49.865 2.135 50.035 2.305 ;
      LAYER met1 ;
        RECT 0.995 2.305 1.225 2.335 ;
        RECT 25.415 2.305 25.645 2.335 ;
        RECT 49.835 2.305 50.065 2.335 ;
        RECT 0.965 2.135 50.095 2.305 ;
        RECT 0.995 2.105 1.225 2.135 ;
        RECT 25.415 2.105 25.645 2.135 ;
        RECT 49.835 2.105 50.065 2.135 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 6.126300 ;
    PORT
      LAYER li1 ;
        RECT 5.465 2.055 5.635 5.095 ;
        RECT 14.745 4.975 14.915 5.095 ;
        RECT 14.715 4.765 14.915 4.975 ;
        RECT 14.715 2.055 14.885 4.765 ;
        RECT 29.885 2.055 30.055 5.095 ;
        RECT 39.165 4.975 39.335 5.095 ;
        RECT 39.135 4.765 39.335 4.975 ;
        RECT 39.135 2.055 39.305 4.765 ;
        RECT 54.305 2.055 54.475 5.095 ;
        RECT 63.585 4.975 63.755 5.095 ;
        RECT 63.555 4.765 63.755 4.975 ;
        RECT 63.555 2.055 63.725 4.765 ;
      LAYER mcon ;
        RECT 5.465 4.725 5.635 4.895 ;
        RECT 14.715 4.725 14.885 4.895 ;
        RECT 29.885 4.725 30.055 4.895 ;
        RECT 39.135 4.725 39.305 4.895 ;
        RECT 54.305 4.725 54.475 4.895 ;
        RECT 63.555 4.725 63.725 4.895 ;
      LAYER met1 ;
        RECT 5.435 4.895 5.665 4.925 ;
        RECT 14.685 4.895 14.915 4.925 ;
        RECT 29.855 4.895 30.085 4.925 ;
        RECT 39.105 4.895 39.335 4.925 ;
        RECT 54.275 4.895 54.505 4.925 ;
        RECT 63.525 4.895 63.755 4.925 ;
        RECT 5.405 4.725 63.785 4.895 ;
        RECT 5.435 4.695 5.665 4.725 ;
        RECT 14.685 4.695 14.915 4.725 ;
        RECT 29.855 4.695 30.085 4.725 ;
        RECT 39.105 4.695 39.335 4.725 ;
        RECT 54.275 4.695 54.505 4.725 ;
        RECT 63.525 4.695 63.755 4.725 ;
    END
  END CLK
  PIN SN
    ANTENNAGATEAREA 6.089100 ;
    PORT
      LAYER li1 ;
        RECT 10.275 2.055 10.445 5.095 ;
        RECT 21.745 2.055 21.915 5.095 ;
        RECT 34.695 2.055 34.865 5.095 ;
        RECT 46.165 2.055 46.335 5.095 ;
        RECT 59.115 2.055 59.285 5.095 ;
        RECT 70.585 2.055 70.755 5.095 ;
      LAYER mcon ;
        RECT 10.275 2.505 10.445 2.675 ;
        RECT 21.745 2.505 21.915 2.675 ;
        RECT 34.695 2.505 34.865 2.675 ;
        RECT 46.165 2.505 46.335 2.675 ;
        RECT 59.115 2.505 59.285 2.675 ;
        RECT 70.585 2.505 70.755 2.675 ;
      LAYER met1 ;
        RECT 10.245 2.675 10.475 2.705 ;
        RECT 21.715 2.675 21.945 2.705 ;
        RECT 34.665 2.675 34.895 2.705 ;
        RECT 46.135 2.675 46.365 2.705 ;
        RECT 59.085 2.675 59.315 2.705 ;
        RECT 70.555 2.675 70.785 2.705 ;
        RECT 10.215 2.505 70.815 2.675 ;
        RECT 10.245 2.475 10.475 2.505 ;
        RECT 21.715 2.475 21.945 2.505 ;
        RECT 34.665 2.475 34.895 2.505 ;
        RECT 46.135 2.475 46.365 2.505 ;
        RECT 59.085 2.475 59.315 2.505 ;
        RECT 70.555 2.475 70.785 2.505 ;
    END
  END SN
  PIN VDD
    ANTENNADIFFAREA 99.913147 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 85.890 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 85.625 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 0.705 5.365 0.875 7.460 ;
        RECT 1.585 5.785 1.755 7.460 ;
        RECT 2.465 5.785 2.635 7.460 ;
        RECT 3.175 4.340 3.485 7.460 ;
        RECT 4.335 5.445 4.505 7.460 ;
        RECT 5.215 5.785 5.385 7.460 ;
        RECT 6.095 5.785 6.265 7.460 ;
        RECT 6.975 5.785 7.145 7.460 ;
        RECT 7.985 4.340 8.295 7.460 ;
        RECT 9.145 5.445 9.315 7.460 ;
        RECT 10.025 5.785 10.195 7.460 ;
        RECT 10.905 5.785 11.075 7.460 ;
        RECT 11.785 5.785 11.955 7.460 ;
        RECT 12.795 4.340 13.105 7.460 ;
        RECT 13.655 5.365 13.825 7.460 ;
        RECT 14.535 5.785 14.705 7.460 ;
        RECT 15.415 5.785 15.585 7.460 ;
        RECT 16.125 4.340 16.435 7.460 ;
        RECT 16.985 5.365 17.155 7.460 ;
        RECT 17.865 5.785 18.035 7.460 ;
        RECT 18.745 5.785 18.915 7.460 ;
        RECT 19.455 4.340 19.765 7.460 ;
        RECT 20.615 5.445 20.785 7.460 ;
        RECT 21.495 5.785 21.665 7.460 ;
        RECT 22.375 5.785 22.545 7.460 ;
        RECT 23.255 5.785 23.425 7.460 ;
        RECT 24.265 4.340 24.575 7.460 ;
        RECT 25.125 5.365 25.295 7.460 ;
        RECT 26.005 5.785 26.175 7.460 ;
        RECT 26.885 5.785 27.055 7.460 ;
        RECT 27.595 4.340 27.905 7.460 ;
        RECT 28.755 5.445 28.925 7.460 ;
        RECT 29.635 5.785 29.805 7.460 ;
        RECT 30.515 5.785 30.685 7.460 ;
        RECT 31.395 5.785 31.565 7.460 ;
        RECT 32.405 4.340 32.715 7.460 ;
        RECT 33.565 5.445 33.735 7.460 ;
        RECT 34.445 5.785 34.615 7.460 ;
        RECT 35.325 5.785 35.495 7.460 ;
        RECT 36.205 5.785 36.375 7.460 ;
        RECT 37.215 4.340 37.525 7.460 ;
        RECT 38.075 5.365 38.245 7.460 ;
        RECT 38.955 5.785 39.125 7.460 ;
        RECT 39.835 5.785 40.005 7.460 ;
        RECT 40.545 4.340 40.855 7.460 ;
        RECT 41.405 5.365 41.575 7.460 ;
        RECT 42.285 5.785 42.455 7.460 ;
        RECT 43.165 5.785 43.335 7.460 ;
        RECT 43.875 4.340 44.185 7.460 ;
        RECT 45.035 5.445 45.205 7.460 ;
        RECT 45.915 5.785 46.085 7.460 ;
        RECT 46.795 5.785 46.965 7.460 ;
        RECT 47.675 5.785 47.845 7.460 ;
        RECT 48.685 4.340 48.995 7.460 ;
        RECT 49.545 5.365 49.715 7.460 ;
        RECT 50.425 5.785 50.595 7.460 ;
        RECT 51.305 5.785 51.475 7.460 ;
        RECT 52.015 4.340 52.325 7.460 ;
        RECT 53.175 5.445 53.345 7.460 ;
        RECT 54.055 5.785 54.225 7.460 ;
        RECT 54.935 5.785 55.105 7.460 ;
        RECT 55.815 5.785 55.985 7.460 ;
        RECT 56.825 4.340 57.135 7.460 ;
        RECT 57.985 5.445 58.155 7.460 ;
        RECT 58.865 5.785 59.035 7.460 ;
        RECT 59.745 5.785 59.915 7.460 ;
        RECT 60.625 5.785 60.795 7.460 ;
        RECT 61.635 4.340 61.945 7.460 ;
        RECT 62.495 5.365 62.665 7.460 ;
        RECT 63.375 5.785 63.545 7.460 ;
        RECT 64.255 5.785 64.425 7.460 ;
        RECT 64.965 4.340 65.275 7.460 ;
        RECT 65.825 5.365 65.995 7.460 ;
        RECT 66.705 5.785 66.875 7.460 ;
        RECT 67.585 5.785 67.755 7.460 ;
        RECT 68.295 4.340 68.605 7.460 ;
        RECT 69.455 5.445 69.625 7.460 ;
        RECT 70.335 5.785 70.505 7.460 ;
        RECT 71.215 5.785 71.385 7.460 ;
        RECT 72.095 5.785 72.265 7.460 ;
        RECT 73.105 4.340 73.415 7.460 ;
        RECT 73.965 5.355 74.135 7.460 ;
        RECT 74.845 5.785 75.015 7.460 ;
        RECT 75.725 5.355 75.895 7.460 ;
        RECT 76.435 4.340 76.745 7.460 ;
        RECT 79.765 4.340 80.075 7.460 ;
        RECT 83.095 4.340 83.405 7.460 ;
        RECT 83.835 5.415 84.005 7.460 ;
        RECT 84.715 5.415 84.885 7.460 ;
        RECT 85.315 4.340 85.625 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 0.995 7.525 1.165 7.695 ;
        RECT 1.355 7.525 1.525 7.695 ;
        RECT 1.805 7.525 1.975 7.695 ;
        RECT 2.165 7.525 2.335 7.695 ;
        RECT 2.525 7.525 2.695 7.695 ;
        RECT 2.885 7.525 3.055 7.695 ;
        RECT 3.605 7.525 3.775 7.695 ;
        RECT 3.965 7.525 4.135 7.695 ;
        RECT 4.325 7.525 4.495 7.695 ;
        RECT 4.685 7.525 4.855 7.695 ;
        RECT 5.045 7.525 5.215 7.695 ;
        RECT 5.405 7.525 5.575 7.695 ;
        RECT 5.895 7.525 6.065 7.695 ;
        RECT 6.255 7.525 6.425 7.695 ;
        RECT 6.615 7.525 6.785 7.695 ;
        RECT 6.975 7.525 7.145 7.695 ;
        RECT 7.335 7.525 7.505 7.695 ;
        RECT 7.695 7.525 7.865 7.695 ;
        RECT 8.415 7.525 8.585 7.695 ;
        RECT 8.775 7.525 8.945 7.695 ;
        RECT 9.135 7.525 9.305 7.695 ;
        RECT 9.495 7.525 9.665 7.695 ;
        RECT 9.855 7.525 10.025 7.695 ;
        RECT 10.215 7.525 10.385 7.695 ;
        RECT 10.705 7.525 10.875 7.695 ;
        RECT 11.065 7.525 11.235 7.695 ;
        RECT 11.425 7.525 11.595 7.695 ;
        RECT 11.785 7.525 11.955 7.695 ;
        RECT 12.145 7.525 12.315 7.695 ;
        RECT 12.505 7.525 12.675 7.695 ;
        RECT 13.225 7.525 13.395 7.695 ;
        RECT 13.585 7.525 13.755 7.695 ;
        RECT 13.945 7.525 14.115 7.695 ;
        RECT 14.305 7.525 14.475 7.695 ;
        RECT 14.755 7.525 14.925 7.695 ;
        RECT 15.115 7.525 15.285 7.695 ;
        RECT 15.475 7.525 15.645 7.695 ;
        RECT 15.835 7.525 16.005 7.695 ;
        RECT 16.555 7.525 16.725 7.695 ;
        RECT 16.915 7.525 17.085 7.695 ;
        RECT 17.275 7.525 17.445 7.695 ;
        RECT 17.635 7.525 17.805 7.695 ;
        RECT 18.085 7.525 18.255 7.695 ;
        RECT 18.445 7.525 18.615 7.695 ;
        RECT 18.805 7.525 18.975 7.695 ;
        RECT 19.165 7.525 19.335 7.695 ;
        RECT 19.885 7.525 20.055 7.695 ;
        RECT 20.245 7.525 20.415 7.695 ;
        RECT 20.605 7.525 20.775 7.695 ;
        RECT 20.965 7.525 21.135 7.695 ;
        RECT 21.325 7.525 21.495 7.695 ;
        RECT 21.685 7.525 21.855 7.695 ;
        RECT 22.175 7.525 22.345 7.695 ;
        RECT 22.535 7.525 22.705 7.695 ;
        RECT 22.895 7.525 23.065 7.695 ;
        RECT 23.255 7.525 23.425 7.695 ;
        RECT 23.615 7.525 23.785 7.695 ;
        RECT 23.975 7.525 24.145 7.695 ;
        RECT 24.695 7.525 24.865 7.695 ;
        RECT 25.055 7.525 25.225 7.695 ;
        RECT 25.415 7.525 25.585 7.695 ;
        RECT 25.775 7.525 25.945 7.695 ;
        RECT 26.225 7.525 26.395 7.695 ;
        RECT 26.585 7.525 26.755 7.695 ;
        RECT 26.945 7.525 27.115 7.695 ;
        RECT 27.305 7.525 27.475 7.695 ;
        RECT 28.025 7.525 28.195 7.695 ;
        RECT 28.385 7.525 28.555 7.695 ;
        RECT 28.745 7.525 28.915 7.695 ;
        RECT 29.105 7.525 29.275 7.695 ;
        RECT 29.465 7.525 29.635 7.695 ;
        RECT 29.825 7.525 29.995 7.695 ;
        RECT 30.315 7.525 30.485 7.695 ;
        RECT 30.675 7.525 30.845 7.695 ;
        RECT 31.035 7.525 31.205 7.695 ;
        RECT 31.395 7.525 31.565 7.695 ;
        RECT 31.755 7.525 31.925 7.695 ;
        RECT 32.115 7.525 32.285 7.695 ;
        RECT 32.835 7.525 33.005 7.695 ;
        RECT 33.195 7.525 33.365 7.695 ;
        RECT 33.555 7.525 33.725 7.695 ;
        RECT 33.915 7.525 34.085 7.695 ;
        RECT 34.275 7.525 34.445 7.695 ;
        RECT 34.635 7.525 34.805 7.695 ;
        RECT 35.125 7.525 35.295 7.695 ;
        RECT 35.485 7.525 35.655 7.695 ;
        RECT 35.845 7.525 36.015 7.695 ;
        RECT 36.205 7.525 36.375 7.695 ;
        RECT 36.565 7.525 36.735 7.695 ;
        RECT 36.925 7.525 37.095 7.695 ;
        RECT 37.645 7.525 37.815 7.695 ;
        RECT 38.005 7.525 38.175 7.695 ;
        RECT 38.365 7.525 38.535 7.695 ;
        RECT 38.725 7.525 38.895 7.695 ;
        RECT 39.175 7.525 39.345 7.695 ;
        RECT 39.535 7.525 39.705 7.695 ;
        RECT 39.895 7.525 40.065 7.695 ;
        RECT 40.255 7.525 40.425 7.695 ;
        RECT 40.975 7.525 41.145 7.695 ;
        RECT 41.335 7.525 41.505 7.695 ;
        RECT 41.695 7.525 41.865 7.695 ;
        RECT 42.055 7.525 42.225 7.695 ;
        RECT 42.505 7.525 42.675 7.695 ;
        RECT 42.865 7.525 43.035 7.695 ;
        RECT 43.225 7.525 43.395 7.695 ;
        RECT 43.585 7.525 43.755 7.695 ;
        RECT 44.305 7.525 44.475 7.695 ;
        RECT 44.665 7.525 44.835 7.695 ;
        RECT 45.025 7.525 45.195 7.695 ;
        RECT 45.385 7.525 45.555 7.695 ;
        RECT 45.745 7.525 45.915 7.695 ;
        RECT 46.105 7.525 46.275 7.695 ;
        RECT 46.595 7.525 46.765 7.695 ;
        RECT 46.955 7.525 47.125 7.695 ;
        RECT 47.315 7.525 47.485 7.695 ;
        RECT 47.675 7.525 47.845 7.695 ;
        RECT 48.035 7.525 48.205 7.695 ;
        RECT 48.395 7.525 48.565 7.695 ;
        RECT 49.115 7.525 49.285 7.695 ;
        RECT 49.475 7.525 49.645 7.695 ;
        RECT 49.835 7.525 50.005 7.695 ;
        RECT 50.195 7.525 50.365 7.695 ;
        RECT 50.645 7.525 50.815 7.695 ;
        RECT 51.005 7.525 51.175 7.695 ;
        RECT 51.365 7.525 51.535 7.695 ;
        RECT 51.725 7.525 51.895 7.695 ;
        RECT 52.445 7.525 52.615 7.695 ;
        RECT 52.805 7.525 52.975 7.695 ;
        RECT 53.165 7.525 53.335 7.695 ;
        RECT 53.525 7.525 53.695 7.695 ;
        RECT 53.885 7.525 54.055 7.695 ;
        RECT 54.245 7.525 54.415 7.695 ;
        RECT 54.735 7.525 54.905 7.695 ;
        RECT 55.095 7.525 55.265 7.695 ;
        RECT 55.455 7.525 55.625 7.695 ;
        RECT 55.815 7.525 55.985 7.695 ;
        RECT 56.175 7.525 56.345 7.695 ;
        RECT 56.535 7.525 56.705 7.695 ;
        RECT 57.255 7.525 57.425 7.695 ;
        RECT 57.615 7.525 57.785 7.695 ;
        RECT 57.975 7.525 58.145 7.695 ;
        RECT 58.335 7.525 58.505 7.695 ;
        RECT 58.695 7.525 58.865 7.695 ;
        RECT 59.055 7.525 59.225 7.695 ;
        RECT 59.545 7.525 59.715 7.695 ;
        RECT 59.905 7.525 60.075 7.695 ;
        RECT 60.265 7.525 60.435 7.695 ;
        RECT 60.625 7.525 60.795 7.695 ;
        RECT 60.985 7.525 61.155 7.695 ;
        RECT 61.345 7.525 61.515 7.695 ;
        RECT 62.065 7.525 62.235 7.695 ;
        RECT 62.425 7.525 62.595 7.695 ;
        RECT 62.785 7.525 62.955 7.695 ;
        RECT 63.145 7.525 63.315 7.695 ;
        RECT 63.595 7.525 63.765 7.695 ;
        RECT 63.955 7.525 64.125 7.695 ;
        RECT 64.315 7.525 64.485 7.695 ;
        RECT 64.675 7.525 64.845 7.695 ;
        RECT 65.395 7.525 65.565 7.695 ;
        RECT 65.755 7.525 65.925 7.695 ;
        RECT 66.115 7.525 66.285 7.695 ;
        RECT 66.475 7.525 66.645 7.695 ;
        RECT 66.925 7.525 67.095 7.695 ;
        RECT 67.285 7.525 67.455 7.695 ;
        RECT 67.645 7.525 67.815 7.695 ;
        RECT 68.005 7.525 68.175 7.695 ;
        RECT 68.725 7.525 68.895 7.695 ;
        RECT 69.085 7.525 69.255 7.695 ;
        RECT 69.445 7.525 69.615 7.695 ;
        RECT 69.805 7.525 69.975 7.695 ;
        RECT 70.165 7.525 70.335 7.695 ;
        RECT 70.525 7.525 70.695 7.695 ;
        RECT 71.015 7.525 71.185 7.695 ;
        RECT 71.375 7.525 71.545 7.695 ;
        RECT 71.735 7.525 71.905 7.695 ;
        RECT 72.095 7.525 72.265 7.695 ;
        RECT 72.455 7.525 72.625 7.695 ;
        RECT 72.815 7.525 72.985 7.695 ;
        RECT 73.535 7.525 73.705 7.695 ;
        RECT 73.895 7.525 74.065 7.695 ;
        RECT 74.255 7.525 74.425 7.695 ;
        RECT 74.615 7.525 74.785 7.695 ;
        RECT 75.065 7.525 75.235 7.695 ;
        RECT 75.425 7.525 75.595 7.695 ;
        RECT 75.785 7.525 75.955 7.695 ;
        RECT 76.145 7.525 76.315 7.695 ;
        RECT 76.865 7.525 77.035 7.695 ;
        RECT 77.225 7.525 77.395 7.695 ;
        RECT 77.585 7.525 77.755 7.695 ;
        RECT 77.945 7.525 78.115 7.695 ;
        RECT 78.395 7.525 78.565 7.695 ;
        RECT 78.755 7.525 78.925 7.695 ;
        RECT 79.115 7.525 79.285 7.695 ;
        RECT 79.475 7.525 79.645 7.695 ;
        RECT 80.195 7.525 80.365 7.695 ;
        RECT 80.555 7.525 80.725 7.695 ;
        RECT 80.915 7.525 81.085 7.695 ;
        RECT 81.275 7.525 81.445 7.695 ;
        RECT 81.725 7.525 81.895 7.695 ;
        RECT 82.085 7.525 82.255 7.695 ;
        RECT 82.445 7.525 82.615 7.695 ;
        RECT 82.805 7.525 82.975 7.695 ;
        RECT 83.525 7.525 83.695 7.695 ;
        RECT 83.885 7.525 84.055 7.695 ;
        RECT 84.275 7.525 84.445 7.695 ;
        RECT 84.665 7.525 84.835 7.695 ;
        RECT 85.025 7.525 85.195 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 85.625 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 62.959297 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 85.755 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 3.045 -0.075 3.615 -0.065 ;
        RECT 7.855 -0.075 8.425 -0.065 ;
        RECT 12.665 -0.075 13.235 -0.065 ;
        RECT 15.995 -0.075 16.565 -0.065 ;
        RECT 19.325 -0.075 19.895 -0.065 ;
        RECT 24.135 -0.075 24.705 -0.065 ;
        RECT 27.465 -0.075 28.035 -0.065 ;
        RECT 32.275 -0.075 32.845 -0.065 ;
        RECT 37.085 -0.075 37.655 -0.065 ;
        RECT 40.415 -0.075 40.985 -0.065 ;
        RECT 43.745 -0.075 44.315 -0.065 ;
        RECT 48.555 -0.075 49.125 -0.065 ;
        RECT 51.885 -0.075 52.455 -0.065 ;
        RECT 56.695 -0.075 57.265 -0.065 ;
        RECT 61.505 -0.075 62.075 -0.065 ;
        RECT 64.835 -0.075 65.405 -0.065 ;
        RECT 68.165 -0.075 68.735 -0.065 ;
        RECT 72.975 -0.075 73.545 -0.065 ;
        RECT 76.305 -0.075 76.875 -0.065 ;
        RECT 79.635 -0.075 80.205 -0.065 ;
        RECT 82.965 -0.075 83.535 -0.065 ;
        RECT 85.185 -0.075 85.755 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 1.095 0.310 1.265 1.260 ;
        RECT 3.175 0.310 3.485 2.860 ;
        RECT 4.320 0.310 4.490 1.270 ;
        RECT 7.985 0.310 8.295 2.860 ;
        RECT 9.130 0.310 9.300 1.270 ;
        RECT 12.795 0.310 13.105 2.860 ;
        RECT 14.045 0.310 14.215 1.260 ;
        RECT 16.125 0.310 16.435 2.860 ;
        RECT 17.375 0.310 17.545 1.260 ;
        RECT 19.455 0.310 19.765 2.860 ;
        RECT 20.600 0.310 20.770 1.270 ;
        RECT 24.265 0.310 24.575 2.860 ;
        RECT 25.515 0.310 25.685 1.260 ;
        RECT 27.595 0.310 27.905 2.860 ;
        RECT 28.740 0.310 28.910 1.270 ;
        RECT 32.405 0.310 32.715 2.860 ;
        RECT 33.550 0.310 33.720 1.270 ;
        RECT 37.215 0.310 37.525 2.860 ;
        RECT 38.465 0.310 38.635 1.260 ;
        RECT 40.545 0.310 40.855 2.860 ;
        RECT 41.795 0.310 41.965 1.260 ;
        RECT 43.875 0.310 44.185 2.860 ;
        RECT 45.020 0.310 45.190 1.270 ;
        RECT 48.685 0.310 48.995 2.860 ;
        RECT 49.935 0.310 50.105 1.260 ;
        RECT 52.015 0.310 52.325 2.860 ;
        RECT 53.160 0.310 53.330 1.270 ;
        RECT 56.825 0.310 57.135 2.860 ;
        RECT 57.970 0.310 58.140 1.270 ;
        RECT 61.635 0.310 61.945 2.860 ;
        RECT 62.885 0.310 63.055 1.260 ;
        RECT 64.965 0.310 65.275 2.860 ;
        RECT 66.215 0.310 66.385 1.260 ;
        RECT 68.295 0.310 68.605 2.860 ;
        RECT 69.440 0.310 69.610 1.270 ;
        RECT 73.105 0.310 73.415 2.860 ;
        RECT 74.355 0.310 74.525 1.260 ;
        RECT 76.435 0.310 76.745 2.860 ;
        RECT 77.685 0.310 77.855 1.260 ;
        RECT 79.765 0.310 80.075 2.860 ;
        RECT 81.015 0.310 81.185 1.260 ;
        RECT 83.095 0.310 83.405 2.860 ;
        RECT 83.795 0.755 83.965 1.885 ;
        RECT 84.765 0.755 84.935 1.885 ;
        RECT 83.795 0.585 84.935 0.755 ;
        RECT 83.795 0.310 83.965 0.585 ;
        RECT 84.280 0.310 84.450 0.585 ;
        RECT 84.765 0.310 84.935 0.585 ;
        RECT 85.315 0.310 85.625 2.860 ;
        RECT -0.155 0.235 78.655 0.310 ;
        RECT 78.825 0.235 85.625 0.310 ;
        RECT -0.155 0.000 85.625 0.235 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 0.995 0.065 1.165 0.235 ;
        RECT 1.355 0.065 1.525 0.235 ;
        RECT 1.805 0.065 1.975 0.235 ;
        RECT 2.165 0.065 2.335 0.235 ;
        RECT 2.525 0.065 2.695 0.235 ;
        RECT 2.885 0.065 3.055 0.235 ;
        RECT 3.605 0.065 3.775 0.235 ;
        RECT 3.965 0.065 4.135 0.235 ;
        RECT 4.325 0.065 4.495 0.235 ;
        RECT 4.685 0.065 4.855 0.235 ;
        RECT 5.045 0.065 5.215 0.235 ;
        RECT 5.405 0.065 5.575 0.235 ;
        RECT 5.895 0.065 6.065 0.235 ;
        RECT 6.255 0.065 6.425 0.235 ;
        RECT 6.615 0.065 6.785 0.235 ;
        RECT 6.975 0.065 7.145 0.235 ;
        RECT 7.335 0.065 7.505 0.235 ;
        RECT 7.695 0.065 7.865 0.235 ;
        RECT 8.415 0.065 8.585 0.235 ;
        RECT 8.775 0.065 8.945 0.235 ;
        RECT 9.135 0.065 9.305 0.235 ;
        RECT 9.495 0.065 9.665 0.235 ;
        RECT 9.855 0.065 10.025 0.235 ;
        RECT 10.215 0.065 10.385 0.235 ;
        RECT 10.705 0.065 10.875 0.235 ;
        RECT 11.065 0.065 11.235 0.235 ;
        RECT 11.425 0.065 11.595 0.235 ;
        RECT 11.785 0.065 11.955 0.235 ;
        RECT 12.145 0.065 12.315 0.235 ;
        RECT 12.505 0.065 12.675 0.235 ;
        RECT 13.225 0.065 13.395 0.235 ;
        RECT 13.585 0.065 13.755 0.235 ;
        RECT 13.945 0.065 14.115 0.235 ;
        RECT 14.305 0.065 14.475 0.235 ;
        RECT 14.755 0.065 14.925 0.235 ;
        RECT 15.115 0.065 15.285 0.235 ;
        RECT 15.475 0.065 15.645 0.235 ;
        RECT 15.835 0.065 16.005 0.235 ;
        RECT 16.555 0.065 16.725 0.235 ;
        RECT 16.915 0.065 17.085 0.235 ;
        RECT 17.275 0.065 17.445 0.235 ;
        RECT 17.635 0.065 17.805 0.235 ;
        RECT 18.085 0.065 18.255 0.235 ;
        RECT 18.445 0.065 18.615 0.235 ;
        RECT 18.805 0.065 18.975 0.235 ;
        RECT 19.165 0.065 19.335 0.235 ;
        RECT 19.885 0.065 20.055 0.235 ;
        RECT 20.245 0.065 20.415 0.235 ;
        RECT 20.605 0.065 20.775 0.235 ;
        RECT 20.965 0.065 21.135 0.235 ;
        RECT 21.325 0.065 21.495 0.235 ;
        RECT 21.685 0.065 21.855 0.235 ;
        RECT 22.175 0.065 22.345 0.235 ;
        RECT 22.535 0.065 22.705 0.235 ;
        RECT 22.895 0.065 23.065 0.235 ;
        RECT 23.255 0.065 23.425 0.235 ;
        RECT 23.615 0.065 23.785 0.235 ;
        RECT 23.975 0.065 24.145 0.235 ;
        RECT 24.695 0.065 24.865 0.235 ;
        RECT 25.055 0.065 25.225 0.235 ;
        RECT 25.415 0.065 25.585 0.235 ;
        RECT 25.775 0.065 25.945 0.235 ;
        RECT 26.225 0.065 26.395 0.235 ;
        RECT 26.585 0.065 26.755 0.235 ;
        RECT 26.945 0.065 27.115 0.235 ;
        RECT 27.305 0.065 27.475 0.235 ;
        RECT 28.025 0.065 28.195 0.235 ;
        RECT 28.385 0.065 28.555 0.235 ;
        RECT 28.745 0.065 28.915 0.235 ;
        RECT 29.105 0.065 29.275 0.235 ;
        RECT 29.465 0.065 29.635 0.235 ;
        RECT 29.825 0.065 29.995 0.235 ;
        RECT 30.315 0.065 30.485 0.235 ;
        RECT 30.675 0.065 30.845 0.235 ;
        RECT 31.035 0.065 31.205 0.235 ;
        RECT 31.395 0.065 31.565 0.235 ;
        RECT 31.755 0.065 31.925 0.235 ;
        RECT 32.115 0.065 32.285 0.235 ;
        RECT 32.835 0.065 33.005 0.235 ;
        RECT 33.195 0.065 33.365 0.235 ;
        RECT 33.555 0.065 33.725 0.235 ;
        RECT 33.915 0.065 34.085 0.235 ;
        RECT 34.275 0.065 34.445 0.235 ;
        RECT 34.635 0.065 34.805 0.235 ;
        RECT 35.125 0.065 35.295 0.235 ;
        RECT 35.485 0.065 35.655 0.235 ;
        RECT 35.845 0.065 36.015 0.235 ;
        RECT 36.205 0.065 36.375 0.235 ;
        RECT 36.565 0.065 36.735 0.235 ;
        RECT 36.925 0.065 37.095 0.235 ;
        RECT 37.645 0.065 37.815 0.235 ;
        RECT 38.005 0.065 38.175 0.235 ;
        RECT 38.365 0.065 38.535 0.235 ;
        RECT 38.725 0.065 38.895 0.235 ;
        RECT 39.175 0.065 39.345 0.235 ;
        RECT 39.535 0.065 39.705 0.235 ;
        RECT 39.895 0.065 40.065 0.235 ;
        RECT 40.255 0.065 40.425 0.235 ;
        RECT 40.975 0.065 41.145 0.235 ;
        RECT 41.335 0.065 41.505 0.235 ;
        RECT 41.695 0.065 41.865 0.235 ;
        RECT 42.055 0.065 42.225 0.235 ;
        RECT 42.505 0.065 42.675 0.235 ;
        RECT 42.865 0.065 43.035 0.235 ;
        RECT 43.225 0.065 43.395 0.235 ;
        RECT 43.585 0.065 43.755 0.235 ;
        RECT 44.305 0.065 44.475 0.235 ;
        RECT 44.665 0.065 44.835 0.235 ;
        RECT 45.025 0.065 45.195 0.235 ;
        RECT 45.385 0.065 45.555 0.235 ;
        RECT 45.745 0.065 45.915 0.235 ;
        RECT 46.105 0.065 46.275 0.235 ;
        RECT 46.595 0.065 46.765 0.235 ;
        RECT 46.955 0.065 47.125 0.235 ;
        RECT 47.315 0.065 47.485 0.235 ;
        RECT 47.675 0.065 47.845 0.235 ;
        RECT 48.035 0.065 48.205 0.235 ;
        RECT 48.395 0.065 48.565 0.235 ;
        RECT 49.115 0.065 49.285 0.235 ;
        RECT 49.475 0.065 49.645 0.235 ;
        RECT 49.835 0.065 50.005 0.235 ;
        RECT 50.195 0.065 50.365 0.235 ;
        RECT 50.645 0.065 50.815 0.235 ;
        RECT 51.005 0.065 51.175 0.235 ;
        RECT 51.365 0.065 51.535 0.235 ;
        RECT 51.725 0.065 51.895 0.235 ;
        RECT 52.445 0.065 52.615 0.235 ;
        RECT 52.805 0.065 52.975 0.235 ;
        RECT 53.165 0.065 53.335 0.235 ;
        RECT 53.525 0.065 53.695 0.235 ;
        RECT 53.885 0.065 54.055 0.235 ;
        RECT 54.245 0.065 54.415 0.235 ;
        RECT 54.735 0.065 54.905 0.235 ;
        RECT 55.095 0.065 55.265 0.235 ;
        RECT 55.455 0.065 55.625 0.235 ;
        RECT 55.815 0.065 55.985 0.235 ;
        RECT 56.175 0.065 56.345 0.235 ;
        RECT 56.535 0.065 56.705 0.235 ;
        RECT 57.255 0.065 57.425 0.235 ;
        RECT 57.615 0.065 57.785 0.235 ;
        RECT 57.975 0.065 58.145 0.235 ;
        RECT 58.335 0.065 58.505 0.235 ;
        RECT 58.695 0.065 58.865 0.235 ;
        RECT 59.055 0.065 59.225 0.235 ;
        RECT 59.545 0.065 59.715 0.235 ;
        RECT 59.905 0.065 60.075 0.235 ;
        RECT 60.265 0.065 60.435 0.235 ;
        RECT 60.625 0.065 60.795 0.235 ;
        RECT 60.985 0.065 61.155 0.235 ;
        RECT 61.345 0.065 61.515 0.235 ;
        RECT 62.065 0.065 62.235 0.235 ;
        RECT 62.425 0.065 62.595 0.235 ;
        RECT 62.785 0.065 62.955 0.235 ;
        RECT 63.145 0.065 63.315 0.235 ;
        RECT 63.595 0.065 63.765 0.235 ;
        RECT 63.955 0.065 64.125 0.235 ;
        RECT 64.315 0.065 64.485 0.235 ;
        RECT 64.675 0.065 64.845 0.235 ;
        RECT 65.395 0.065 65.565 0.235 ;
        RECT 65.755 0.065 65.925 0.235 ;
        RECT 66.115 0.065 66.285 0.235 ;
        RECT 66.475 0.065 66.645 0.235 ;
        RECT 66.925 0.065 67.095 0.235 ;
        RECT 67.285 0.065 67.455 0.235 ;
        RECT 67.645 0.065 67.815 0.235 ;
        RECT 68.005 0.065 68.175 0.235 ;
        RECT 68.725 0.065 68.895 0.235 ;
        RECT 69.085 0.065 69.255 0.235 ;
        RECT 69.445 0.065 69.615 0.235 ;
        RECT 69.805 0.065 69.975 0.235 ;
        RECT 70.165 0.065 70.335 0.235 ;
        RECT 70.525 0.065 70.695 0.235 ;
        RECT 71.015 0.065 71.185 0.235 ;
        RECT 71.375 0.065 71.545 0.235 ;
        RECT 71.735 0.065 71.905 0.235 ;
        RECT 72.095 0.065 72.265 0.235 ;
        RECT 72.455 0.065 72.625 0.235 ;
        RECT 72.815 0.065 72.985 0.235 ;
        RECT 73.535 0.065 73.705 0.235 ;
        RECT 73.895 0.065 74.065 0.235 ;
        RECT 74.255 0.065 74.425 0.235 ;
        RECT 74.615 0.065 74.785 0.235 ;
        RECT 75.065 0.065 75.235 0.235 ;
        RECT 75.425 0.065 75.595 0.235 ;
        RECT 75.785 0.065 75.955 0.235 ;
        RECT 76.145 0.065 76.315 0.235 ;
        RECT 76.865 0.065 77.035 0.235 ;
        RECT 77.225 0.065 77.395 0.235 ;
        RECT 77.585 0.065 77.755 0.235 ;
        RECT 77.945 0.065 78.115 0.235 ;
        RECT 78.395 0.065 78.565 0.235 ;
        RECT 78.755 0.065 78.925 0.235 ;
        RECT 79.115 0.065 79.285 0.235 ;
        RECT 79.475 0.065 79.645 0.235 ;
        RECT 80.195 0.065 80.365 0.235 ;
        RECT 80.555 0.065 80.725 0.235 ;
        RECT 80.915 0.065 81.085 0.235 ;
        RECT 81.275 0.065 81.445 0.235 ;
        RECT 81.725 0.065 81.895 0.235 ;
        RECT 82.085 0.065 82.255 0.235 ;
        RECT 82.445 0.065 82.615 0.235 ;
        RECT 82.805 0.065 82.975 0.235 ;
        RECT 83.525 0.065 83.695 0.235 ;
        RECT 83.885 0.065 84.055 0.235 ;
        RECT 84.275 0.065 84.445 0.235 ;
        RECT 84.665 0.065 84.835 0.235 ;
        RECT 85.025 0.065 85.195 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 85.625 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 1.145 5.515 1.315 7.250 ;
        RECT 2.025 5.515 2.195 7.250 ;
        RECT 1.145 5.345 2.675 5.515 ;
        RECT 1.795 4.940 1.965 5.095 ;
        RECT 1.765 4.765 1.965 4.940 ;
        RECT 1.765 2.055 1.935 4.765 ;
        RECT 0.610 1.805 0.780 1.885 ;
        RECT 1.580 1.805 1.750 1.885 ;
        RECT 2.505 1.880 2.675 5.345 ;
        RECT 4.775 5.470 4.945 7.250 ;
        RECT 5.655 5.470 5.825 7.250 ;
        RECT 6.535 5.470 6.705 7.250 ;
        RECT 9.585 5.470 9.755 7.250 ;
        RECT 10.465 5.470 10.635 7.250 ;
        RECT 11.345 5.470 11.515 7.250 ;
        RECT 14.095 5.515 14.265 7.250 ;
        RECT 14.975 5.515 15.145 7.250 ;
        RECT 17.425 5.515 17.595 7.250 ;
        RECT 18.305 5.515 18.475 7.250 ;
        RECT 4.775 5.300 7.485 5.470 ;
        RECT 9.585 5.300 12.295 5.470 ;
        RECT 14.095 5.345 15.625 5.515 ;
        RECT 17.425 5.345 18.955 5.515 ;
        RECT 4.355 2.055 4.525 5.095 ;
        RECT 6.575 2.055 6.745 5.095 ;
        RECT 7.315 4.605 7.485 5.300 ;
        RECT 7.310 4.275 7.485 4.605 ;
        RECT 0.610 1.635 1.750 1.805 ;
        RECT 0.610 0.505 0.780 1.635 ;
        RECT 1.580 0.755 1.750 1.635 ;
        RECT 2.065 1.710 2.675 1.880 ;
        RECT 3.835 1.815 4.005 1.895 ;
        RECT 4.805 1.815 4.975 1.895 ;
        RECT 5.775 1.815 5.945 1.895 ;
        RECT 2.065 0.975 2.235 1.710 ;
        RECT 3.835 1.645 5.945 1.815 ;
        RECT 2.550 0.755 2.720 1.525 ;
        RECT 1.580 0.585 2.720 0.755 ;
        RECT 1.580 0.505 1.750 0.585 ;
        RECT 2.550 0.505 2.720 0.585 ;
        RECT 3.835 0.515 4.005 1.645 ;
        RECT 4.805 0.765 4.975 1.645 ;
        RECT 5.775 1.565 5.945 1.645 ;
        RECT 5.295 1.220 5.465 1.300 ;
        RECT 6.345 1.220 6.515 1.895 ;
        RECT 7.315 1.890 7.485 4.275 ;
        RECT 9.165 2.055 9.335 5.095 ;
        RECT 11.385 2.055 11.555 5.095 ;
        RECT 5.295 1.050 6.515 1.220 ;
        RECT 5.295 0.970 5.465 1.050 ;
        RECT 5.775 0.765 5.945 0.845 ;
        RECT 4.805 0.595 5.945 0.765 ;
        RECT 4.805 0.515 4.975 0.595 ;
        RECT 5.775 0.515 5.945 0.595 ;
        RECT 6.345 0.765 6.515 1.050 ;
        RECT 6.830 1.720 7.485 1.890 ;
        RECT 8.645 1.815 8.815 1.895 ;
        RECT 9.615 1.815 9.785 1.895 ;
        RECT 10.585 1.815 10.755 1.895 ;
        RECT 6.830 0.985 7.000 1.720 ;
        RECT 8.645 1.645 10.755 1.815 ;
        RECT 7.315 0.765 7.485 1.535 ;
        RECT 6.345 0.595 7.485 0.765 ;
        RECT 6.345 0.515 6.515 0.595 ;
        RECT 7.315 0.515 7.485 0.595 ;
        RECT 8.645 0.515 8.815 1.645 ;
        RECT 9.615 0.765 9.785 1.645 ;
        RECT 10.585 1.565 10.755 1.645 ;
        RECT 10.105 1.220 10.275 1.300 ;
        RECT 11.155 1.220 11.325 1.895 ;
        RECT 12.125 1.890 12.295 5.300 ;
        RECT 13.975 2.055 14.145 5.095 ;
        RECT 10.105 1.050 11.325 1.220 ;
        RECT 10.105 0.970 10.275 1.050 ;
        RECT 10.585 0.765 10.755 0.845 ;
        RECT 9.615 0.595 10.755 0.765 ;
        RECT 9.615 0.515 9.785 0.595 ;
        RECT 10.585 0.515 10.755 0.595 ;
        RECT 11.155 0.765 11.325 1.050 ;
        RECT 11.640 1.720 12.295 1.890 ;
        RECT 13.560 1.805 13.730 1.885 ;
        RECT 14.530 1.805 14.700 1.885 ;
        RECT 15.455 1.880 15.625 5.345 ;
        RECT 17.305 2.055 17.475 5.095 ;
        RECT 18.075 4.940 18.245 5.095 ;
        RECT 18.045 4.765 18.245 4.940 ;
        RECT 18.045 2.055 18.215 4.765 ;
        RECT 11.640 0.985 11.810 1.720 ;
        RECT 13.560 1.635 14.700 1.805 ;
        RECT 12.125 0.765 12.295 1.535 ;
        RECT 11.155 0.595 12.295 0.765 ;
        RECT 11.155 0.515 11.325 0.595 ;
        RECT 12.125 0.515 12.295 0.595 ;
        RECT 13.560 0.505 13.730 1.635 ;
        RECT 14.530 0.755 14.700 1.635 ;
        RECT 15.015 1.710 15.625 1.880 ;
        RECT 16.890 1.805 17.060 1.885 ;
        RECT 17.860 1.805 18.030 1.885 ;
        RECT 18.785 1.880 18.955 5.345 ;
        RECT 21.055 5.470 21.225 7.250 ;
        RECT 21.935 5.470 22.105 7.250 ;
        RECT 22.815 5.470 22.985 7.250 ;
        RECT 25.565 5.515 25.735 7.250 ;
        RECT 26.445 5.515 26.615 7.250 ;
        RECT 21.055 5.300 23.765 5.470 ;
        RECT 25.565 5.345 27.095 5.515 ;
        RECT 20.635 2.055 20.805 5.095 ;
        RECT 22.855 2.055 23.025 5.095 ;
        RECT 15.015 0.975 15.185 1.710 ;
        RECT 16.890 1.635 18.030 1.805 ;
        RECT 15.500 0.755 15.670 1.525 ;
        RECT 14.530 0.585 15.670 0.755 ;
        RECT 14.530 0.505 14.700 0.585 ;
        RECT 15.500 0.505 15.670 0.585 ;
        RECT 16.890 0.505 17.060 1.635 ;
        RECT 17.860 0.755 18.030 1.635 ;
        RECT 18.345 1.710 18.955 1.880 ;
        RECT 20.115 1.815 20.285 1.895 ;
        RECT 21.085 1.815 21.255 1.895 ;
        RECT 22.055 1.815 22.225 1.895 ;
        RECT 18.345 0.975 18.515 1.710 ;
        RECT 20.115 1.645 22.225 1.815 ;
        RECT 18.830 0.755 19.000 1.525 ;
        RECT 17.860 0.585 19.000 0.755 ;
        RECT 17.860 0.505 18.030 0.585 ;
        RECT 18.830 0.505 19.000 0.585 ;
        RECT 20.115 0.515 20.285 1.645 ;
        RECT 21.085 0.765 21.255 1.645 ;
        RECT 22.055 1.565 22.225 1.645 ;
        RECT 21.575 1.220 21.745 1.300 ;
        RECT 22.625 1.220 22.795 1.895 ;
        RECT 23.595 1.890 23.765 5.300 ;
        RECT 26.215 4.940 26.385 5.095 ;
        RECT 26.185 4.765 26.385 4.940 ;
        RECT 26.185 2.055 26.355 4.765 ;
        RECT 21.575 1.050 22.795 1.220 ;
        RECT 21.575 0.970 21.745 1.050 ;
        RECT 22.055 0.765 22.225 0.845 ;
        RECT 21.085 0.595 22.225 0.765 ;
        RECT 21.085 0.515 21.255 0.595 ;
        RECT 22.055 0.515 22.225 0.595 ;
        RECT 22.625 0.765 22.795 1.050 ;
        RECT 23.110 1.720 23.765 1.890 ;
        RECT 25.030 1.805 25.200 1.885 ;
        RECT 26.000 1.805 26.170 1.885 ;
        RECT 26.925 1.880 27.095 5.345 ;
        RECT 29.195 5.470 29.365 7.250 ;
        RECT 30.075 5.470 30.245 7.250 ;
        RECT 30.955 5.470 31.125 7.250 ;
        RECT 34.005 5.470 34.175 7.250 ;
        RECT 34.885 5.470 35.055 7.250 ;
        RECT 35.765 5.470 35.935 7.250 ;
        RECT 38.515 5.515 38.685 7.250 ;
        RECT 39.395 5.515 39.565 7.250 ;
        RECT 41.845 5.515 42.015 7.250 ;
        RECT 42.725 5.515 42.895 7.250 ;
        RECT 29.195 5.300 31.905 5.470 ;
        RECT 34.005 5.300 36.715 5.470 ;
        RECT 38.515 5.345 40.045 5.515 ;
        RECT 41.845 5.345 43.375 5.515 ;
        RECT 28.775 2.055 28.945 5.095 ;
        RECT 30.995 2.055 31.165 5.095 ;
        RECT 31.735 4.605 31.905 5.300 ;
        RECT 31.730 4.275 31.905 4.605 ;
        RECT 23.110 0.985 23.280 1.720 ;
        RECT 25.030 1.635 26.170 1.805 ;
        RECT 23.595 0.765 23.765 1.535 ;
        RECT 22.625 0.595 23.765 0.765 ;
        RECT 22.625 0.515 22.795 0.595 ;
        RECT 23.595 0.515 23.765 0.595 ;
        RECT 25.030 0.505 25.200 1.635 ;
        RECT 26.000 0.755 26.170 1.635 ;
        RECT 26.485 1.710 27.095 1.880 ;
        RECT 28.255 1.815 28.425 1.895 ;
        RECT 29.225 1.815 29.395 1.895 ;
        RECT 30.195 1.815 30.365 1.895 ;
        RECT 26.485 0.975 26.655 1.710 ;
        RECT 28.255 1.645 30.365 1.815 ;
        RECT 26.970 0.755 27.140 1.525 ;
        RECT 26.000 0.585 27.140 0.755 ;
        RECT 26.000 0.505 26.170 0.585 ;
        RECT 26.970 0.505 27.140 0.585 ;
        RECT 28.255 0.515 28.425 1.645 ;
        RECT 29.225 0.765 29.395 1.645 ;
        RECT 30.195 1.565 30.365 1.645 ;
        RECT 29.715 1.220 29.885 1.300 ;
        RECT 30.765 1.220 30.935 1.895 ;
        RECT 31.735 1.890 31.905 4.275 ;
        RECT 33.585 2.055 33.755 5.095 ;
        RECT 35.805 2.055 35.975 5.095 ;
        RECT 29.715 1.050 30.935 1.220 ;
        RECT 29.715 0.970 29.885 1.050 ;
        RECT 30.195 0.765 30.365 0.845 ;
        RECT 29.225 0.595 30.365 0.765 ;
        RECT 29.225 0.515 29.395 0.595 ;
        RECT 30.195 0.515 30.365 0.595 ;
        RECT 30.765 0.765 30.935 1.050 ;
        RECT 31.250 1.720 31.905 1.890 ;
        RECT 33.065 1.815 33.235 1.895 ;
        RECT 34.035 1.815 34.205 1.895 ;
        RECT 35.005 1.815 35.175 1.895 ;
        RECT 31.250 0.985 31.420 1.720 ;
        RECT 33.065 1.645 35.175 1.815 ;
        RECT 31.735 0.765 31.905 1.535 ;
        RECT 30.765 0.595 31.905 0.765 ;
        RECT 30.765 0.515 30.935 0.595 ;
        RECT 31.735 0.515 31.905 0.595 ;
        RECT 33.065 0.515 33.235 1.645 ;
        RECT 34.035 0.765 34.205 1.645 ;
        RECT 35.005 1.565 35.175 1.645 ;
        RECT 34.525 1.220 34.695 1.300 ;
        RECT 35.575 1.220 35.745 1.895 ;
        RECT 36.545 1.890 36.715 5.300 ;
        RECT 38.395 2.055 38.565 5.095 ;
        RECT 34.525 1.050 35.745 1.220 ;
        RECT 34.525 0.970 34.695 1.050 ;
        RECT 35.005 0.765 35.175 0.845 ;
        RECT 34.035 0.595 35.175 0.765 ;
        RECT 34.035 0.515 34.205 0.595 ;
        RECT 35.005 0.515 35.175 0.595 ;
        RECT 35.575 0.765 35.745 1.050 ;
        RECT 36.060 1.720 36.715 1.890 ;
        RECT 37.980 1.805 38.150 1.885 ;
        RECT 38.950 1.805 39.120 1.885 ;
        RECT 39.875 1.880 40.045 5.345 ;
        RECT 41.725 2.055 41.895 5.095 ;
        RECT 42.495 4.940 42.665 5.095 ;
        RECT 42.465 4.765 42.665 4.940 ;
        RECT 42.465 2.055 42.635 4.765 ;
        RECT 36.060 0.985 36.230 1.720 ;
        RECT 37.980 1.635 39.120 1.805 ;
        RECT 36.545 0.765 36.715 1.535 ;
        RECT 35.575 0.595 36.715 0.765 ;
        RECT 35.575 0.515 35.745 0.595 ;
        RECT 36.545 0.515 36.715 0.595 ;
        RECT 37.980 0.505 38.150 1.635 ;
        RECT 38.950 0.755 39.120 1.635 ;
        RECT 39.435 1.710 40.045 1.880 ;
        RECT 41.310 1.805 41.480 1.885 ;
        RECT 42.280 1.805 42.450 1.885 ;
        RECT 43.205 1.880 43.375 5.345 ;
        RECT 45.475 5.470 45.645 7.250 ;
        RECT 46.355 5.470 46.525 7.250 ;
        RECT 47.235 5.470 47.405 7.250 ;
        RECT 49.985 5.515 50.155 7.250 ;
        RECT 50.865 5.515 51.035 7.250 ;
        RECT 45.475 5.300 48.185 5.470 ;
        RECT 49.985 5.345 51.515 5.515 ;
        RECT 45.055 2.055 45.225 5.095 ;
        RECT 47.275 2.055 47.445 5.095 ;
        RECT 39.435 0.975 39.605 1.710 ;
        RECT 41.310 1.635 42.450 1.805 ;
        RECT 39.920 0.755 40.090 1.525 ;
        RECT 38.950 0.585 40.090 0.755 ;
        RECT 38.950 0.505 39.120 0.585 ;
        RECT 39.920 0.505 40.090 0.585 ;
        RECT 41.310 0.505 41.480 1.635 ;
        RECT 42.280 0.755 42.450 1.635 ;
        RECT 42.765 1.710 43.375 1.880 ;
        RECT 44.535 1.815 44.705 1.895 ;
        RECT 45.505 1.815 45.675 1.895 ;
        RECT 46.475 1.815 46.645 1.895 ;
        RECT 42.765 0.975 42.935 1.710 ;
        RECT 44.535 1.645 46.645 1.815 ;
        RECT 43.250 0.755 43.420 1.525 ;
        RECT 42.280 0.585 43.420 0.755 ;
        RECT 42.280 0.505 42.450 0.585 ;
        RECT 43.250 0.505 43.420 0.585 ;
        RECT 44.535 0.515 44.705 1.645 ;
        RECT 45.505 0.765 45.675 1.645 ;
        RECT 46.475 1.565 46.645 1.645 ;
        RECT 45.995 1.220 46.165 1.300 ;
        RECT 47.045 1.220 47.215 1.895 ;
        RECT 48.015 1.890 48.185 5.300 ;
        RECT 50.635 4.940 50.805 5.095 ;
        RECT 50.605 4.765 50.805 4.940 ;
        RECT 50.605 2.055 50.775 4.765 ;
        RECT 45.995 1.050 47.215 1.220 ;
        RECT 45.995 0.970 46.165 1.050 ;
        RECT 46.475 0.765 46.645 0.845 ;
        RECT 45.505 0.595 46.645 0.765 ;
        RECT 45.505 0.515 45.675 0.595 ;
        RECT 46.475 0.515 46.645 0.595 ;
        RECT 47.045 0.765 47.215 1.050 ;
        RECT 47.530 1.720 48.185 1.890 ;
        RECT 49.450 1.805 49.620 1.885 ;
        RECT 50.420 1.805 50.590 1.885 ;
        RECT 51.345 1.880 51.515 5.345 ;
        RECT 53.615 5.470 53.785 7.250 ;
        RECT 54.495 5.470 54.665 7.250 ;
        RECT 55.375 5.470 55.545 7.250 ;
        RECT 58.425 5.470 58.595 7.250 ;
        RECT 59.305 5.470 59.475 7.250 ;
        RECT 60.185 5.470 60.355 7.250 ;
        RECT 62.935 5.515 63.105 7.250 ;
        RECT 63.815 5.515 63.985 7.250 ;
        RECT 66.265 5.515 66.435 7.250 ;
        RECT 67.145 5.515 67.315 7.250 ;
        RECT 53.615 5.300 56.325 5.470 ;
        RECT 58.425 5.300 61.135 5.470 ;
        RECT 62.935 5.345 64.465 5.515 ;
        RECT 66.265 5.345 67.795 5.515 ;
        RECT 53.195 2.055 53.365 5.095 ;
        RECT 55.415 2.055 55.585 5.095 ;
        RECT 56.155 4.605 56.325 5.300 ;
        RECT 56.150 4.275 56.325 4.605 ;
        RECT 47.530 0.985 47.700 1.720 ;
        RECT 49.450 1.635 50.590 1.805 ;
        RECT 48.015 0.765 48.185 1.535 ;
        RECT 47.045 0.595 48.185 0.765 ;
        RECT 47.045 0.515 47.215 0.595 ;
        RECT 48.015 0.515 48.185 0.595 ;
        RECT 49.450 0.505 49.620 1.635 ;
        RECT 50.420 0.755 50.590 1.635 ;
        RECT 50.905 1.710 51.515 1.880 ;
        RECT 52.675 1.815 52.845 1.895 ;
        RECT 53.645 1.815 53.815 1.895 ;
        RECT 54.615 1.815 54.785 1.895 ;
        RECT 50.905 0.975 51.075 1.710 ;
        RECT 52.675 1.645 54.785 1.815 ;
        RECT 51.390 0.755 51.560 1.525 ;
        RECT 50.420 0.585 51.560 0.755 ;
        RECT 50.420 0.505 50.590 0.585 ;
        RECT 51.390 0.505 51.560 0.585 ;
        RECT 52.675 0.515 52.845 1.645 ;
        RECT 53.645 0.765 53.815 1.645 ;
        RECT 54.615 1.565 54.785 1.645 ;
        RECT 54.135 1.220 54.305 1.300 ;
        RECT 55.185 1.220 55.355 1.895 ;
        RECT 56.155 1.890 56.325 4.275 ;
        RECT 58.005 2.055 58.175 5.095 ;
        RECT 60.225 2.055 60.395 5.095 ;
        RECT 54.135 1.050 55.355 1.220 ;
        RECT 54.135 0.970 54.305 1.050 ;
        RECT 54.615 0.765 54.785 0.845 ;
        RECT 53.645 0.595 54.785 0.765 ;
        RECT 53.645 0.515 53.815 0.595 ;
        RECT 54.615 0.515 54.785 0.595 ;
        RECT 55.185 0.765 55.355 1.050 ;
        RECT 55.670 1.720 56.325 1.890 ;
        RECT 57.485 1.815 57.655 1.895 ;
        RECT 58.455 1.815 58.625 1.895 ;
        RECT 59.425 1.815 59.595 1.895 ;
        RECT 55.670 0.985 55.840 1.720 ;
        RECT 57.485 1.645 59.595 1.815 ;
        RECT 56.155 0.765 56.325 1.535 ;
        RECT 55.185 0.595 56.325 0.765 ;
        RECT 55.185 0.515 55.355 0.595 ;
        RECT 56.155 0.515 56.325 0.595 ;
        RECT 57.485 0.515 57.655 1.645 ;
        RECT 58.455 0.765 58.625 1.645 ;
        RECT 59.425 1.565 59.595 1.645 ;
        RECT 58.945 1.220 59.115 1.300 ;
        RECT 59.995 1.220 60.165 1.895 ;
        RECT 60.965 1.890 61.135 5.300 ;
        RECT 62.815 2.055 62.985 5.095 ;
        RECT 58.945 1.050 60.165 1.220 ;
        RECT 58.945 0.970 59.115 1.050 ;
        RECT 59.425 0.765 59.595 0.845 ;
        RECT 58.455 0.595 59.595 0.765 ;
        RECT 58.455 0.515 58.625 0.595 ;
        RECT 59.425 0.515 59.595 0.595 ;
        RECT 59.995 0.765 60.165 1.050 ;
        RECT 60.480 1.720 61.135 1.890 ;
        RECT 62.400 1.805 62.570 1.885 ;
        RECT 63.370 1.805 63.540 1.885 ;
        RECT 64.295 1.880 64.465 5.345 ;
        RECT 66.145 2.055 66.315 5.095 ;
        RECT 66.915 4.940 67.085 5.095 ;
        RECT 66.885 4.765 67.085 4.940 ;
        RECT 66.885 2.055 67.055 4.765 ;
        RECT 60.480 0.985 60.650 1.720 ;
        RECT 62.400 1.635 63.540 1.805 ;
        RECT 60.965 0.765 61.135 1.535 ;
        RECT 59.995 0.595 61.135 0.765 ;
        RECT 59.995 0.515 60.165 0.595 ;
        RECT 60.965 0.515 61.135 0.595 ;
        RECT 62.400 0.505 62.570 1.635 ;
        RECT 63.370 0.755 63.540 1.635 ;
        RECT 63.855 1.710 64.465 1.880 ;
        RECT 65.730 1.805 65.900 1.885 ;
        RECT 66.700 1.805 66.870 1.885 ;
        RECT 67.625 1.880 67.795 5.345 ;
        RECT 69.895 5.470 70.065 7.250 ;
        RECT 70.775 5.470 70.945 7.250 ;
        RECT 71.655 5.470 71.825 7.250 ;
        RECT 74.405 7.055 74.585 7.225 ;
        RECT 74.405 5.525 74.575 7.055 ;
        RECT 75.285 5.525 75.455 7.225 ;
        RECT 69.895 5.300 72.605 5.470 ;
        RECT 74.405 5.355 75.455 5.525 ;
        RECT 69.475 2.055 69.645 5.095 ;
        RECT 71.695 2.055 71.865 5.095 ;
        RECT 63.855 0.975 64.025 1.710 ;
        RECT 65.730 1.635 66.870 1.805 ;
        RECT 64.340 0.755 64.510 1.525 ;
        RECT 63.370 0.585 64.510 0.755 ;
        RECT 63.370 0.505 63.540 0.585 ;
        RECT 64.340 0.505 64.510 0.585 ;
        RECT 65.730 0.505 65.900 1.635 ;
        RECT 66.700 0.755 66.870 1.635 ;
        RECT 67.185 1.710 67.795 1.880 ;
        RECT 68.955 1.815 69.125 1.895 ;
        RECT 69.925 1.815 70.095 1.895 ;
        RECT 70.895 1.815 71.065 1.895 ;
        RECT 67.185 0.975 67.355 1.710 ;
        RECT 68.955 1.645 71.065 1.815 ;
        RECT 67.670 0.755 67.840 1.525 ;
        RECT 66.700 0.585 67.840 0.755 ;
        RECT 66.700 0.505 66.870 0.585 ;
        RECT 67.670 0.505 67.840 0.585 ;
        RECT 68.955 0.515 69.125 1.645 ;
        RECT 69.925 0.765 70.095 1.645 ;
        RECT 70.895 1.565 71.065 1.645 ;
        RECT 70.415 1.220 70.585 1.300 ;
        RECT 71.465 1.220 71.635 1.895 ;
        RECT 72.435 1.890 72.605 5.300 ;
        RECT 75.285 5.275 75.455 5.355 ;
        RECT 77.285 7.055 79.215 7.225 ;
        RECT 77.285 5.275 77.455 7.055 ;
        RECT 77.725 5.525 77.895 6.795 ;
        RECT 78.165 5.785 78.335 7.055 ;
        RECT 78.605 5.525 78.775 6.795 ;
        RECT 79.045 5.605 79.215 7.055 ;
        RECT 80.625 7.055 82.555 7.225 ;
        RECT 77.725 5.355 78.775 5.525 ;
        RECT 78.605 5.275 78.775 5.355 ;
        RECT 80.625 5.275 80.795 7.055 ;
        RECT 81.065 5.525 81.235 6.795 ;
        RECT 81.505 5.785 81.675 7.055 ;
        RECT 81.945 5.525 82.115 6.795 ;
        RECT 82.385 5.785 82.555 7.055 ;
        RECT 81.065 5.355 82.595 5.525 ;
        RECT 73.915 2.055 74.085 5.100 ;
        RECT 75.065 4.940 75.235 5.100 ;
        RECT 75.025 4.770 75.235 4.940 ;
        RECT 75.025 2.055 75.195 4.770 ;
        RECT 77.615 2.055 77.785 5.100 ;
        RECT 79.095 2.055 79.265 5.100 ;
        RECT 80.575 2.055 80.745 5.100 ;
        RECT 81.685 4.770 81.875 5.100 ;
        RECT 81.685 2.055 81.855 4.770 ;
        RECT 70.415 1.050 71.635 1.220 ;
        RECT 70.415 0.970 70.585 1.050 ;
        RECT 70.895 0.765 71.065 0.845 ;
        RECT 69.925 0.595 71.065 0.765 ;
        RECT 69.925 0.515 70.095 0.595 ;
        RECT 70.895 0.515 71.065 0.595 ;
        RECT 71.465 0.765 71.635 1.050 ;
        RECT 71.950 1.720 72.605 1.890 ;
        RECT 73.870 1.805 74.040 1.885 ;
        RECT 74.840 1.805 75.010 1.885 ;
        RECT 71.950 0.985 72.120 1.720 ;
        RECT 73.870 1.635 75.010 1.805 ;
        RECT 72.435 0.765 72.605 1.535 ;
        RECT 71.465 0.595 72.605 0.765 ;
        RECT 71.465 0.515 71.635 0.595 ;
        RECT 72.435 0.515 72.605 0.595 ;
        RECT 73.870 0.505 74.040 1.635 ;
        RECT 74.840 0.755 75.010 1.635 ;
        RECT 75.325 1.310 75.495 1.485 ;
        RECT 75.320 1.155 75.495 1.310 ;
        RECT 75.320 0.975 75.490 1.155 ;
        RECT 75.810 0.755 75.980 1.885 ;
        RECT 74.840 0.585 75.980 0.755 ;
        RECT 74.840 0.505 75.010 0.585 ;
        RECT 75.810 0.505 75.980 0.585 ;
        RECT 77.200 1.805 77.370 1.885 ;
        RECT 78.170 1.805 78.340 1.885 ;
        RECT 77.200 1.635 78.340 1.805 ;
        RECT 77.200 0.505 77.370 1.635 ;
        RECT 78.170 0.755 78.340 1.635 ;
        RECT 78.655 0.975 78.825 1.485 ;
        RECT 79.140 0.755 79.310 1.885 ;
        RECT 78.170 0.585 79.310 0.755 ;
        RECT 78.170 0.505 78.340 0.585 ;
        RECT 79.140 0.505 79.310 0.585 ;
        RECT 80.530 1.805 80.700 1.885 ;
        RECT 81.500 1.805 81.670 1.885 ;
        RECT 82.425 1.870 82.595 5.355 ;
        RECT 83.905 2.055 84.075 5.095 ;
        RECT 80.530 1.635 81.670 1.805 ;
        RECT 80.530 0.505 80.700 1.635 ;
        RECT 81.500 0.755 81.670 1.635 ;
        RECT 81.985 1.700 82.595 1.870 ;
        RECT 81.985 0.975 82.155 1.700 ;
        RECT 82.470 0.755 82.640 1.530 ;
        RECT 81.500 0.585 82.640 0.755 ;
        RECT 81.500 0.505 81.670 0.585 ;
        RECT 82.470 0.505 82.640 0.585 ;
      LAYER mcon ;
        RECT 1.765 4.355 1.935 4.525 ;
        RECT 2.505 2.875 2.675 3.045 ;
        RECT 4.355 2.870 4.525 3.040 ;
        RECT 7.310 4.355 7.480 4.525 ;
        RECT 6.575 3.985 6.745 4.155 ;
        RECT 9.165 2.875 9.335 3.045 ;
        RECT 11.385 3.985 11.555 4.155 ;
        RECT 12.125 2.875 12.295 3.045 ;
        RECT 13.975 2.875 14.145 3.045 ;
        RECT 15.455 3.985 15.625 4.155 ;
        RECT 17.305 4.355 17.475 4.525 ;
        RECT 18.045 3.245 18.215 3.415 ;
        RECT 18.785 4.355 18.955 4.525 ;
        RECT 20.635 4.355 20.805 4.525 ;
        RECT 22.855 3.985 23.025 4.155 ;
        RECT 23.595 3.245 23.765 3.415 ;
        RECT 26.185 4.355 26.355 4.525 ;
        RECT 26.925 2.875 27.095 3.045 ;
        RECT 28.775 2.870 28.945 3.040 ;
        RECT 31.730 4.355 31.900 4.525 ;
        RECT 30.995 3.985 31.165 4.155 ;
        RECT 33.585 2.875 33.755 3.045 ;
        RECT 35.805 3.985 35.975 4.155 ;
        RECT 36.545 2.875 36.715 3.045 ;
        RECT 38.395 2.875 38.565 3.045 ;
        RECT 39.875 3.985 40.045 4.155 ;
        RECT 41.725 4.355 41.895 4.525 ;
        RECT 42.465 3.615 42.635 3.785 ;
        RECT 43.205 4.355 43.375 4.525 ;
        RECT 45.055 4.355 45.225 4.525 ;
        RECT 47.275 3.985 47.445 4.155 ;
        RECT 48.015 3.615 48.185 3.785 ;
        RECT 50.605 4.355 50.775 4.525 ;
        RECT 51.345 2.875 51.515 3.045 ;
        RECT 53.195 2.870 53.365 3.040 ;
        RECT 56.150 4.355 56.320 4.525 ;
        RECT 55.415 3.985 55.585 4.155 ;
        RECT 58.005 2.875 58.175 3.045 ;
        RECT 60.225 3.985 60.395 4.155 ;
        RECT 60.965 2.875 61.135 3.045 ;
        RECT 62.815 2.875 62.985 3.045 ;
        RECT 64.295 3.985 64.465 4.155 ;
        RECT 66.145 4.355 66.315 4.525 ;
        RECT 75.285 5.355 75.455 5.525 ;
        RECT 66.885 4.355 67.055 4.525 ;
        RECT 67.625 4.725 67.795 4.895 ;
        RECT 69.475 4.725 69.645 4.895 ;
        RECT 71.695 3.985 71.865 4.155 ;
        RECT 77.285 5.355 77.455 5.525 ;
        RECT 78.605 5.355 78.775 5.525 ;
        RECT 80.625 5.355 80.795 5.525 ;
        RECT 72.435 4.355 72.605 4.525 ;
        RECT 73.915 4.725 74.085 4.895 ;
        RECT 73.915 3.615 74.085 3.785 ;
        RECT 75.025 4.355 75.195 4.525 ;
        RECT 77.615 4.725 77.785 4.895 ;
        RECT 79.095 3.245 79.265 3.415 ;
        RECT 79.095 2.135 79.265 2.305 ;
        RECT 80.575 2.135 80.745 2.305 ;
        RECT 81.685 4.355 81.855 4.525 ;
        RECT 82.425 3.985 82.595 4.155 ;
        RECT 75.325 1.235 75.495 1.405 ;
        RECT 78.655 1.235 78.825 1.405 ;
        RECT 83.905 3.985 84.075 4.155 ;
        RECT 81.985 1.235 82.155 1.405 ;
      LAYER met1 ;
        RECT 75.255 5.525 75.485 5.555 ;
        RECT 77.255 5.525 77.485 5.555 ;
        RECT 78.575 5.525 78.805 5.555 ;
        RECT 80.595 5.525 80.825 5.555 ;
        RECT 75.225 5.355 77.515 5.525 ;
        RECT 78.545 5.355 80.855 5.525 ;
        RECT 75.255 5.325 75.485 5.355 ;
        RECT 77.255 5.325 77.485 5.355 ;
        RECT 78.575 5.325 78.805 5.355 ;
        RECT 80.595 5.325 80.825 5.355 ;
        RECT 67.595 4.895 67.825 4.925 ;
        RECT 69.445 4.895 69.675 4.925 ;
        RECT 73.885 4.895 74.115 4.925 ;
        RECT 77.585 4.895 77.815 4.925 ;
        RECT 67.565 4.725 69.705 4.895 ;
        RECT 73.855 4.725 77.845 4.895 ;
        RECT 67.595 4.695 67.825 4.725 ;
        RECT 69.445 4.695 69.675 4.725 ;
        RECT 73.885 4.695 74.115 4.725 ;
        RECT 77.585 4.695 77.815 4.725 ;
        RECT 1.735 4.525 1.965 4.555 ;
        RECT 7.280 4.525 7.510 4.555 ;
        RECT 17.275 4.525 17.505 4.555 ;
        RECT 18.755 4.525 18.985 4.555 ;
        RECT 20.605 4.525 20.835 4.555 ;
        RECT 26.155 4.525 26.385 4.555 ;
        RECT 31.700 4.525 31.930 4.555 ;
        RECT 41.695 4.525 41.925 4.555 ;
        RECT 43.175 4.525 43.405 4.555 ;
        RECT 45.025 4.525 45.255 4.555 ;
        RECT 50.575 4.525 50.805 4.555 ;
        RECT 56.120 4.525 56.350 4.555 ;
        RECT 66.115 4.525 66.345 4.555 ;
        RECT 66.855 4.525 67.085 4.555 ;
        RECT 72.405 4.525 72.635 4.555 ;
        RECT 74.995 4.525 75.225 4.555 ;
        RECT 81.655 4.525 81.885 4.555 ;
        RECT 1.705 4.355 17.535 4.525 ;
        RECT 18.725 4.355 20.865 4.525 ;
        RECT 26.125 4.355 41.955 4.525 ;
        RECT 43.145 4.355 45.285 4.525 ;
        RECT 50.545 4.355 66.375 4.525 ;
        RECT 66.825 4.355 81.915 4.525 ;
        RECT 1.735 4.325 1.965 4.355 ;
        RECT 7.280 4.325 7.510 4.355 ;
        RECT 17.275 4.325 17.505 4.355 ;
        RECT 18.755 4.325 18.985 4.355 ;
        RECT 20.605 4.325 20.835 4.355 ;
        RECT 26.155 4.325 26.385 4.355 ;
        RECT 31.700 4.325 31.930 4.355 ;
        RECT 41.695 4.325 41.925 4.355 ;
        RECT 43.175 4.325 43.405 4.355 ;
        RECT 45.025 4.325 45.255 4.355 ;
        RECT 50.575 4.325 50.805 4.355 ;
        RECT 56.120 4.325 56.350 4.355 ;
        RECT 66.115 4.325 66.345 4.355 ;
        RECT 66.855 4.325 67.085 4.355 ;
        RECT 72.405 4.325 72.635 4.355 ;
        RECT 74.995 4.325 75.225 4.355 ;
        RECT 81.655 4.325 81.885 4.355 ;
        RECT 6.545 4.155 6.775 4.185 ;
        RECT 11.355 4.155 11.585 4.185 ;
        RECT 15.425 4.155 15.655 4.185 ;
        RECT 22.825 4.155 23.055 4.185 ;
        RECT 30.965 4.155 31.195 4.185 ;
        RECT 35.775 4.155 36.005 4.185 ;
        RECT 39.845 4.155 40.075 4.185 ;
        RECT 47.245 4.155 47.475 4.185 ;
        RECT 55.385 4.155 55.615 4.185 ;
        RECT 60.195 4.155 60.425 4.185 ;
        RECT 64.265 4.155 64.495 4.185 ;
        RECT 71.665 4.155 71.895 4.185 ;
        RECT 82.395 4.155 82.625 4.185 ;
        RECT 83.875 4.155 84.105 4.185 ;
        RECT 6.515 3.985 23.085 4.155 ;
        RECT 30.935 3.985 47.505 4.155 ;
        RECT 55.355 3.985 71.925 4.155 ;
        RECT 82.365 3.985 84.135 4.155 ;
        RECT 6.545 3.955 6.775 3.985 ;
        RECT 11.355 3.955 11.585 3.985 ;
        RECT 15.425 3.955 15.655 3.985 ;
        RECT 22.825 3.955 23.055 3.985 ;
        RECT 30.965 3.955 31.195 3.985 ;
        RECT 35.775 3.955 36.005 3.985 ;
        RECT 39.845 3.955 40.075 3.985 ;
        RECT 47.245 3.955 47.475 3.985 ;
        RECT 55.385 3.955 55.615 3.985 ;
        RECT 60.195 3.955 60.425 3.985 ;
        RECT 64.265 3.955 64.495 3.985 ;
        RECT 71.665 3.955 71.895 3.985 ;
        RECT 82.395 3.955 82.625 3.985 ;
        RECT 83.875 3.955 84.105 3.985 ;
        RECT 42.435 3.785 42.665 3.815 ;
        RECT 47.985 3.785 48.215 3.815 ;
        RECT 73.885 3.785 74.115 3.815 ;
        RECT 42.405 3.615 74.145 3.785 ;
        RECT 42.435 3.585 42.665 3.615 ;
        RECT 47.985 3.585 48.215 3.615 ;
        RECT 73.885 3.585 74.115 3.615 ;
        RECT 18.015 3.415 18.245 3.445 ;
        RECT 23.565 3.415 23.795 3.445 ;
        RECT 79.065 3.415 79.295 3.445 ;
        RECT 17.985 3.245 79.325 3.415 ;
        RECT 18.015 3.215 18.245 3.245 ;
        RECT 23.565 3.215 23.795 3.245 ;
        RECT 79.065 3.215 79.295 3.245 ;
        RECT 2.475 3.045 2.705 3.075 ;
        RECT 4.325 3.045 4.555 3.070 ;
        RECT 9.135 3.045 9.365 3.075 ;
        RECT 12.095 3.045 12.325 3.075 ;
        RECT 13.945 3.045 14.175 3.075 ;
        RECT 26.895 3.045 27.125 3.075 ;
        RECT 28.745 3.045 28.975 3.070 ;
        RECT 33.555 3.045 33.785 3.075 ;
        RECT 36.515 3.045 36.745 3.075 ;
        RECT 38.365 3.045 38.595 3.075 ;
        RECT 51.315 3.045 51.545 3.075 ;
        RECT 53.165 3.045 53.395 3.070 ;
        RECT 57.975 3.045 58.205 3.075 ;
        RECT 60.935 3.045 61.165 3.075 ;
        RECT 62.785 3.045 63.015 3.075 ;
        RECT 2.445 2.875 9.395 3.045 ;
        RECT 12.065 2.875 14.205 3.045 ;
        RECT 26.865 2.875 33.815 3.045 ;
        RECT 36.485 2.875 38.625 3.045 ;
        RECT 51.285 2.875 58.235 3.045 ;
        RECT 60.905 2.875 63.045 3.045 ;
        RECT 2.475 2.845 2.705 2.875 ;
        RECT 4.295 2.870 4.705 2.875 ;
        RECT 4.325 2.840 4.555 2.870 ;
        RECT 9.135 2.845 9.365 2.875 ;
        RECT 12.095 2.845 12.325 2.875 ;
        RECT 13.945 2.845 14.175 2.875 ;
        RECT 26.895 2.845 27.125 2.875 ;
        RECT 28.715 2.870 29.125 2.875 ;
        RECT 28.745 2.840 28.975 2.870 ;
        RECT 33.555 2.845 33.785 2.875 ;
        RECT 36.515 2.845 36.745 2.875 ;
        RECT 38.365 2.845 38.595 2.875 ;
        RECT 51.315 2.845 51.545 2.875 ;
        RECT 53.135 2.870 53.545 2.875 ;
        RECT 53.165 2.840 53.395 2.870 ;
        RECT 57.975 2.845 58.205 2.875 ;
        RECT 60.935 2.845 61.165 2.875 ;
        RECT 62.785 2.845 63.015 2.875 ;
        RECT 79.065 2.305 79.295 2.335 ;
        RECT 80.545 2.305 80.775 2.335 ;
        RECT 79.035 2.135 80.805 2.305 ;
        RECT 79.065 2.105 79.295 2.135 ;
        RECT 80.545 2.105 80.775 2.135 ;
        RECT 75.295 1.405 75.525 1.435 ;
        RECT 78.625 1.405 78.855 1.435 ;
        RECT 81.955 1.405 82.185 1.435 ;
        RECT 75.265 1.235 82.215 1.405 ;
        RECT 75.295 1.205 75.525 1.235 ;
        RECT 78.625 1.205 78.855 1.235 ;
        RECT 81.955 1.205 82.185 1.235 ;
  END
END TMRDFFSNQX1






MACRO TMRDFFSNRNQNX1
  CLASS BLOCK ;
  FOREIGN TMRDFFSNRNQNX1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 97.410 BY 7.950 ;
  PIN QN
    ANTENNADIFFAREA 1.734950 ;
    PORT
      LAYER li1 ;
        RECT 94.385 5.525 94.555 6.795 ;
        RECT 95.265 5.525 95.435 6.795 ;
        RECT 94.385 5.355 95.915 5.525 ;
        RECT 95.745 1.870 95.915 5.355 ;
        RECT 95.305 1.700 95.915 1.870 ;
        RECT 88.645 1.310 88.815 1.485 ;
        RECT 88.640 1.155 88.815 1.310 ;
        RECT 88.640 0.975 88.810 1.155 ;
        RECT 91.975 0.975 92.145 1.485 ;
        RECT 95.305 0.975 95.475 1.700 ;
      LAYER mcon ;
        RECT 95.745 3.985 95.915 4.155 ;
        RECT 88.645 1.235 88.815 1.405 ;
        RECT 91.975 1.235 92.145 1.405 ;
        RECT 95.305 1.235 95.475 1.405 ;
      LAYER met1 ;
        RECT 95.715 4.155 95.945 4.185 ;
        RECT 95.685 3.985 96.095 4.155 ;
        RECT 95.715 3.955 95.945 3.985 ;
        RECT 88.615 1.405 88.845 1.435 ;
        RECT 91.945 1.405 92.175 1.435 ;
        RECT 95.275 1.405 95.505 1.435 ;
        RECT 88.585 1.235 95.535 1.405 ;
        RECT 88.615 1.205 88.845 1.235 ;
        RECT 91.945 1.205 92.175 1.235 ;
        RECT 95.275 1.205 95.505 1.235 ;
    END
  END QN
  PIN D
    ANTENNAGATEAREA 3.099750 ;
    PORT
      LAYER li1 ;
        RECT 1.025 2.055 1.195 5.095 ;
        RECT 29.885 2.055 30.055 5.095 ;
        RECT 58.745 2.055 58.915 5.095 ;
      LAYER mcon ;
        RECT 1.025 4.355 1.195 4.525 ;
        RECT 29.885 4.355 30.055 4.525 ;
        RECT 58.745 4.355 58.915 4.525 ;
      LAYER met1 ;
        RECT 0.995 4.525 1.225 4.555 ;
        RECT 29.855 4.525 30.085 4.555 ;
        RECT 58.715 4.525 58.945 4.555 ;
        RECT 0.845 4.355 59.095 4.525 ;
        RECT 0.995 4.325 1.225 4.355 ;
        RECT 29.855 4.325 30.085 4.355 ;
        RECT 58.715 4.325 58.945 4.355 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 6.089100 ;
    PORT
      LAYER li1 ;
        RECT 6.945 4.975 7.115 5.095 ;
        RECT 6.940 4.645 7.115 4.975 ;
        RECT 6.945 2.055 7.115 4.645 ;
        RECT 16.565 2.055 16.735 5.095 ;
        RECT 35.805 4.975 35.975 5.095 ;
        RECT 35.800 4.645 35.975 4.975 ;
        RECT 35.805 2.055 35.975 4.645 ;
        RECT 45.425 2.055 45.595 5.095 ;
        RECT 64.665 4.975 64.835 5.095 ;
        RECT 64.660 4.645 64.835 4.975 ;
        RECT 64.665 2.055 64.835 4.645 ;
        RECT 74.285 2.055 74.455 5.095 ;
      LAYER mcon ;
        RECT 6.940 4.725 7.110 4.895 ;
        RECT 16.565 4.725 16.735 4.895 ;
        RECT 35.800 4.725 35.970 4.895 ;
        RECT 45.425 4.725 45.595 4.895 ;
        RECT 64.660 4.725 64.830 4.895 ;
        RECT 74.285 4.725 74.455 4.895 ;
      LAYER met1 ;
        RECT 6.910 4.895 7.140 4.925 ;
        RECT 16.535 4.895 16.765 4.925 ;
        RECT 35.770 4.895 36.000 4.925 ;
        RECT 45.395 4.895 45.625 4.925 ;
        RECT 64.630 4.895 64.860 4.925 ;
        RECT 74.255 4.895 74.485 4.925 ;
        RECT 6.880 4.725 74.515 4.895 ;
        RECT 6.910 4.695 7.140 4.725 ;
        RECT 16.535 4.695 16.765 4.725 ;
        RECT 35.770 4.695 36.000 4.725 ;
        RECT 45.395 4.695 45.625 4.725 ;
        RECT 64.630 4.695 64.860 4.725 ;
        RECT 74.255 4.695 74.485 4.725 ;
    END
  END CLK
  PIN SN
    ANTENNAGATEAREA 6.089100 ;
    PORT
      LAYER li1 ;
        RECT 11.755 2.055 11.925 5.095 ;
        RECT 26.185 2.055 26.355 5.095 ;
        RECT 40.615 2.055 40.785 5.095 ;
        RECT 55.045 2.055 55.215 5.095 ;
        RECT 69.475 2.055 69.645 5.095 ;
        RECT 83.905 2.055 84.075 5.095 ;
      LAYER mcon ;
        RECT 11.755 2.140 11.925 2.310 ;
        RECT 26.185 2.135 26.355 2.305 ;
        RECT 40.615 2.140 40.785 2.310 ;
        RECT 55.045 2.135 55.215 2.305 ;
        RECT 69.475 2.140 69.645 2.310 ;
        RECT 83.905 2.135 84.075 2.305 ;
      LAYER met1 ;
        RECT 11.725 2.310 11.955 2.340 ;
        RECT 11.695 2.305 12.105 2.310 ;
        RECT 26.155 2.305 26.385 2.335 ;
        RECT 40.585 2.310 40.815 2.340 ;
        RECT 40.555 2.305 40.965 2.310 ;
        RECT 55.015 2.305 55.245 2.335 ;
        RECT 69.445 2.310 69.675 2.340 ;
        RECT 69.415 2.305 69.825 2.310 ;
        RECT 83.875 2.305 84.105 2.335 ;
        RECT 11.695 2.140 84.135 2.305 ;
        RECT 11.720 2.135 84.135 2.140 ;
        RECT 11.725 2.110 11.955 2.135 ;
        RECT 26.155 2.105 26.385 2.135 ;
        RECT 40.585 2.110 40.815 2.135 ;
        RECT 55.015 2.105 55.245 2.135 ;
        RECT 69.445 2.110 69.675 2.135 ;
        RECT 83.875 2.105 84.105 2.135 ;
    END
  END SN
  PIN RN
    ANTENNAGATEAREA 9.170850 ;
    PORT
      LAYER li1 ;
        RECT 2.135 2.055 2.305 5.095 ;
        RECT 17.675 2.055 17.845 5.095 ;
        RECT 21.375 2.055 21.545 5.095 ;
        RECT 30.995 2.055 31.165 5.095 ;
        RECT 46.535 2.055 46.705 5.095 ;
        RECT 50.235 2.055 50.405 5.095 ;
        RECT 59.855 2.055 60.025 5.095 ;
        RECT 75.395 2.055 75.565 5.095 ;
        RECT 79.095 2.055 79.265 5.095 ;
      LAYER mcon ;
        RECT 2.135 2.505 2.305 2.675 ;
        RECT 17.675 2.505 17.845 2.675 ;
        RECT 21.375 2.505 21.545 2.675 ;
        RECT 30.995 2.505 31.165 2.675 ;
        RECT 46.535 2.505 46.705 2.675 ;
        RECT 50.235 2.505 50.405 2.675 ;
        RECT 59.855 2.505 60.025 2.675 ;
        RECT 75.395 2.505 75.565 2.675 ;
        RECT 79.095 2.505 79.265 2.675 ;
      LAYER met1 ;
        RECT 2.105 2.675 2.335 2.705 ;
        RECT 17.645 2.675 17.875 2.705 ;
        RECT 21.345 2.675 21.575 2.705 ;
        RECT 30.965 2.675 31.195 2.705 ;
        RECT 46.505 2.675 46.735 2.705 ;
        RECT 50.205 2.675 50.435 2.705 ;
        RECT 59.825 2.675 60.055 2.705 ;
        RECT 75.365 2.675 75.595 2.705 ;
        RECT 79.065 2.675 79.295 2.705 ;
        RECT 2.075 2.505 79.325 2.675 ;
        RECT 2.105 2.475 2.335 2.505 ;
        RECT 17.645 2.475 17.875 2.505 ;
        RECT 21.345 2.475 21.575 2.505 ;
        RECT 30.965 2.475 31.195 2.505 ;
        RECT 46.505 2.475 46.735 2.505 ;
        RECT 50.205 2.475 50.435 2.505 ;
        RECT 59.825 2.475 60.055 2.505 ;
        RECT 75.365 2.475 75.595 2.505 ;
        RECT 79.065 2.475 79.295 2.505 ;
    END
  END RN
  PIN VDD
    ANTENNADIFFAREA 108.469894 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 96.990 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 96.725 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 1.005 5.445 1.175 7.460 ;
        RECT 1.885 5.785 2.055 7.460 ;
        RECT 2.765 5.785 2.935 7.460 ;
        RECT 3.645 5.785 3.815 7.460 ;
        RECT 4.655 4.340 4.965 7.460 ;
        RECT 5.815 5.445 5.985 7.460 ;
        RECT 6.695 5.785 6.865 7.460 ;
        RECT 7.575 5.785 7.745 7.460 ;
        RECT 8.455 5.785 8.625 7.460 ;
        RECT 9.465 4.340 9.775 7.460 ;
        RECT 10.625 5.445 10.795 7.460 ;
        RECT 11.505 5.785 11.675 7.460 ;
        RECT 12.385 5.785 12.555 7.460 ;
        RECT 13.265 5.785 13.435 7.460 ;
        RECT 14.275 4.340 14.585 7.460 ;
        RECT 15.435 5.445 15.605 7.460 ;
        RECT 16.315 5.785 16.485 7.460 ;
        RECT 17.195 5.785 17.365 7.460 ;
        RECT 18.075 5.785 18.245 7.460 ;
        RECT 19.085 4.340 19.395 7.460 ;
        RECT 20.245 5.445 20.415 7.460 ;
        RECT 21.125 5.785 21.295 7.460 ;
        RECT 22.005 5.785 22.175 7.460 ;
        RECT 22.885 5.785 23.055 7.460 ;
        RECT 23.895 4.340 24.205 7.460 ;
        RECT 25.055 5.445 25.225 7.460 ;
        RECT 25.935 5.785 26.105 7.460 ;
        RECT 26.815 5.785 26.985 7.460 ;
        RECT 27.695 5.785 27.865 7.460 ;
        RECT 28.705 4.340 29.015 7.460 ;
        RECT 29.865 5.445 30.035 7.460 ;
        RECT 30.745 5.785 30.915 7.460 ;
        RECT 31.625 5.785 31.795 7.460 ;
        RECT 32.505 5.785 32.675 7.460 ;
        RECT 33.515 4.340 33.825 7.460 ;
        RECT 34.675 5.445 34.845 7.460 ;
        RECT 35.555 5.785 35.725 7.460 ;
        RECT 36.435 5.785 36.605 7.460 ;
        RECT 37.315 5.785 37.485 7.460 ;
        RECT 38.325 4.340 38.635 7.460 ;
        RECT 39.485 5.445 39.655 7.460 ;
        RECT 40.365 5.785 40.535 7.460 ;
        RECT 41.245 5.785 41.415 7.460 ;
        RECT 42.125 5.785 42.295 7.460 ;
        RECT 43.135 4.340 43.445 7.460 ;
        RECT 44.295 5.445 44.465 7.460 ;
        RECT 45.175 5.785 45.345 7.460 ;
        RECT 46.055 5.785 46.225 7.460 ;
        RECT 46.935 5.785 47.105 7.460 ;
        RECT 47.945 4.340 48.255 7.460 ;
        RECT 49.105 5.445 49.275 7.460 ;
        RECT 49.985 5.785 50.155 7.460 ;
        RECT 50.865 5.785 51.035 7.460 ;
        RECT 51.745 5.785 51.915 7.460 ;
        RECT 52.755 4.340 53.065 7.460 ;
        RECT 53.915 5.445 54.085 7.460 ;
        RECT 54.795 5.785 54.965 7.460 ;
        RECT 55.675 5.785 55.845 7.460 ;
        RECT 56.555 5.785 56.725 7.460 ;
        RECT 57.565 4.340 57.875 7.460 ;
        RECT 58.725 5.445 58.895 7.460 ;
        RECT 59.605 5.785 59.775 7.460 ;
        RECT 60.485 5.785 60.655 7.460 ;
        RECT 61.365 5.785 61.535 7.460 ;
        RECT 62.375 4.340 62.685 7.460 ;
        RECT 63.535 5.445 63.705 7.460 ;
        RECT 64.415 5.785 64.585 7.460 ;
        RECT 65.295 5.785 65.465 7.460 ;
        RECT 66.175 5.785 66.345 7.460 ;
        RECT 67.185 4.340 67.495 7.460 ;
        RECT 68.345 5.445 68.515 7.460 ;
        RECT 69.225 5.785 69.395 7.460 ;
        RECT 70.105 5.785 70.275 7.460 ;
        RECT 70.985 5.785 71.155 7.460 ;
        RECT 71.995 4.340 72.305 7.460 ;
        RECT 73.155 5.445 73.325 7.460 ;
        RECT 74.035 5.785 74.205 7.460 ;
        RECT 74.915 5.785 75.085 7.460 ;
        RECT 75.795 5.785 75.965 7.460 ;
        RECT 76.805 4.340 77.115 7.460 ;
        RECT 77.965 5.445 78.135 7.460 ;
        RECT 78.845 5.785 79.015 7.460 ;
        RECT 79.725 5.785 79.895 7.460 ;
        RECT 80.605 5.785 80.775 7.460 ;
        RECT 81.615 4.340 81.925 7.460 ;
        RECT 82.775 5.445 82.945 7.460 ;
        RECT 83.655 5.785 83.825 7.460 ;
        RECT 84.535 5.785 84.705 7.460 ;
        RECT 85.415 5.785 85.585 7.460 ;
        RECT 86.425 4.340 86.735 7.460 ;
        RECT 87.285 5.355 87.455 7.460 ;
        RECT 88.165 5.785 88.335 7.460 ;
        RECT 89.045 5.355 89.215 7.460 ;
        RECT 89.755 4.340 90.065 7.460 ;
        RECT 93.085 4.340 93.395 7.460 ;
        RECT 96.415 4.340 96.725 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 0.995 7.525 1.165 7.695 ;
        RECT 1.355 7.525 1.525 7.695 ;
        RECT 1.715 7.525 1.885 7.695 ;
        RECT 2.075 7.525 2.245 7.695 ;
        RECT 2.565 7.525 2.735 7.695 ;
        RECT 2.925 7.525 3.095 7.695 ;
        RECT 3.285 7.525 3.455 7.695 ;
        RECT 3.645 7.525 3.815 7.695 ;
        RECT 4.005 7.525 4.175 7.695 ;
        RECT 4.365 7.525 4.535 7.695 ;
        RECT 5.085 7.525 5.255 7.695 ;
        RECT 5.445 7.525 5.615 7.695 ;
        RECT 5.805 7.525 5.975 7.695 ;
        RECT 6.165 7.525 6.335 7.695 ;
        RECT 6.525 7.525 6.695 7.695 ;
        RECT 6.885 7.525 7.055 7.695 ;
        RECT 7.375 7.525 7.545 7.695 ;
        RECT 7.735 7.525 7.905 7.695 ;
        RECT 8.095 7.525 8.265 7.695 ;
        RECT 8.455 7.525 8.625 7.695 ;
        RECT 8.815 7.525 8.985 7.695 ;
        RECT 9.175 7.525 9.345 7.695 ;
        RECT 9.895 7.525 10.065 7.695 ;
        RECT 10.255 7.525 10.425 7.695 ;
        RECT 10.615 7.525 10.785 7.695 ;
        RECT 10.975 7.525 11.145 7.695 ;
        RECT 11.335 7.525 11.505 7.695 ;
        RECT 11.695 7.525 11.865 7.695 ;
        RECT 12.185 7.525 12.355 7.695 ;
        RECT 12.545 7.525 12.715 7.695 ;
        RECT 12.905 7.525 13.075 7.695 ;
        RECT 13.265 7.525 13.435 7.695 ;
        RECT 13.625 7.525 13.795 7.695 ;
        RECT 13.985 7.525 14.155 7.695 ;
        RECT 14.705 7.525 14.875 7.695 ;
        RECT 15.065 7.525 15.235 7.695 ;
        RECT 15.425 7.525 15.595 7.695 ;
        RECT 15.785 7.525 15.955 7.695 ;
        RECT 16.145 7.525 16.315 7.695 ;
        RECT 16.505 7.525 16.675 7.695 ;
        RECT 16.995 7.525 17.165 7.695 ;
        RECT 17.355 7.525 17.525 7.695 ;
        RECT 17.715 7.525 17.885 7.695 ;
        RECT 18.075 7.525 18.245 7.695 ;
        RECT 18.435 7.525 18.605 7.695 ;
        RECT 18.795 7.525 18.965 7.695 ;
        RECT 19.515 7.525 19.685 7.695 ;
        RECT 19.875 7.525 20.045 7.695 ;
        RECT 20.235 7.525 20.405 7.695 ;
        RECT 20.595 7.525 20.765 7.695 ;
        RECT 20.955 7.525 21.125 7.695 ;
        RECT 21.315 7.525 21.485 7.695 ;
        RECT 21.805 7.525 21.975 7.695 ;
        RECT 22.165 7.525 22.335 7.695 ;
        RECT 22.525 7.525 22.695 7.695 ;
        RECT 22.885 7.525 23.055 7.695 ;
        RECT 23.245 7.525 23.415 7.695 ;
        RECT 23.605 7.525 23.775 7.695 ;
        RECT 24.325 7.525 24.495 7.695 ;
        RECT 24.685 7.525 24.855 7.695 ;
        RECT 25.045 7.525 25.215 7.695 ;
        RECT 25.405 7.525 25.575 7.695 ;
        RECT 25.765 7.525 25.935 7.695 ;
        RECT 26.125 7.525 26.295 7.695 ;
        RECT 26.615 7.525 26.785 7.695 ;
        RECT 26.975 7.525 27.145 7.695 ;
        RECT 27.335 7.525 27.505 7.695 ;
        RECT 27.695 7.525 27.865 7.695 ;
        RECT 28.055 7.525 28.225 7.695 ;
        RECT 28.415 7.525 28.585 7.695 ;
        RECT 29.135 7.525 29.305 7.695 ;
        RECT 29.495 7.525 29.665 7.695 ;
        RECT 29.855 7.525 30.025 7.695 ;
        RECT 30.215 7.525 30.385 7.695 ;
        RECT 30.575 7.525 30.745 7.695 ;
        RECT 30.935 7.525 31.105 7.695 ;
        RECT 31.425 7.525 31.595 7.695 ;
        RECT 31.785 7.525 31.955 7.695 ;
        RECT 32.145 7.525 32.315 7.695 ;
        RECT 32.505 7.525 32.675 7.695 ;
        RECT 32.865 7.525 33.035 7.695 ;
        RECT 33.225 7.525 33.395 7.695 ;
        RECT 33.945 7.525 34.115 7.695 ;
        RECT 34.305 7.525 34.475 7.695 ;
        RECT 34.665 7.525 34.835 7.695 ;
        RECT 35.025 7.525 35.195 7.695 ;
        RECT 35.385 7.525 35.555 7.695 ;
        RECT 35.745 7.525 35.915 7.695 ;
        RECT 36.235 7.525 36.405 7.695 ;
        RECT 36.595 7.525 36.765 7.695 ;
        RECT 36.955 7.525 37.125 7.695 ;
        RECT 37.315 7.525 37.485 7.695 ;
        RECT 37.675 7.525 37.845 7.695 ;
        RECT 38.035 7.525 38.205 7.695 ;
        RECT 38.755 7.525 38.925 7.695 ;
        RECT 39.115 7.525 39.285 7.695 ;
        RECT 39.475 7.525 39.645 7.695 ;
        RECT 39.835 7.525 40.005 7.695 ;
        RECT 40.195 7.525 40.365 7.695 ;
        RECT 40.555 7.525 40.725 7.695 ;
        RECT 41.045 7.525 41.215 7.695 ;
        RECT 41.405 7.525 41.575 7.695 ;
        RECT 41.765 7.525 41.935 7.695 ;
        RECT 42.125 7.525 42.295 7.695 ;
        RECT 42.485 7.525 42.655 7.695 ;
        RECT 42.845 7.525 43.015 7.695 ;
        RECT 43.565 7.525 43.735 7.695 ;
        RECT 43.925 7.525 44.095 7.695 ;
        RECT 44.285 7.525 44.455 7.695 ;
        RECT 44.645 7.525 44.815 7.695 ;
        RECT 45.005 7.525 45.175 7.695 ;
        RECT 45.365 7.525 45.535 7.695 ;
        RECT 45.855 7.525 46.025 7.695 ;
        RECT 46.215 7.525 46.385 7.695 ;
        RECT 46.575 7.525 46.745 7.695 ;
        RECT 46.935 7.525 47.105 7.695 ;
        RECT 47.295 7.525 47.465 7.695 ;
        RECT 47.655 7.525 47.825 7.695 ;
        RECT 48.375 7.525 48.545 7.695 ;
        RECT 48.735 7.525 48.905 7.695 ;
        RECT 49.095 7.525 49.265 7.695 ;
        RECT 49.455 7.525 49.625 7.695 ;
        RECT 49.815 7.525 49.985 7.695 ;
        RECT 50.175 7.525 50.345 7.695 ;
        RECT 50.665 7.525 50.835 7.695 ;
        RECT 51.025 7.525 51.195 7.695 ;
        RECT 51.385 7.525 51.555 7.695 ;
        RECT 51.745 7.525 51.915 7.695 ;
        RECT 52.105 7.525 52.275 7.695 ;
        RECT 52.465 7.525 52.635 7.695 ;
        RECT 53.185 7.525 53.355 7.695 ;
        RECT 53.545 7.525 53.715 7.695 ;
        RECT 53.905 7.525 54.075 7.695 ;
        RECT 54.265 7.525 54.435 7.695 ;
        RECT 54.625 7.525 54.795 7.695 ;
        RECT 54.985 7.525 55.155 7.695 ;
        RECT 55.475 7.525 55.645 7.695 ;
        RECT 55.835 7.525 56.005 7.695 ;
        RECT 56.195 7.525 56.365 7.695 ;
        RECT 56.555 7.525 56.725 7.695 ;
        RECT 56.915 7.525 57.085 7.695 ;
        RECT 57.275 7.525 57.445 7.695 ;
        RECT 57.995 7.525 58.165 7.695 ;
        RECT 58.355 7.525 58.525 7.695 ;
        RECT 58.715 7.525 58.885 7.695 ;
        RECT 59.075 7.525 59.245 7.695 ;
        RECT 59.435 7.525 59.605 7.695 ;
        RECT 59.795 7.525 59.965 7.695 ;
        RECT 60.285 7.525 60.455 7.695 ;
        RECT 60.645 7.525 60.815 7.695 ;
        RECT 61.005 7.525 61.175 7.695 ;
        RECT 61.365 7.525 61.535 7.695 ;
        RECT 61.725 7.525 61.895 7.695 ;
        RECT 62.085 7.525 62.255 7.695 ;
        RECT 62.805 7.525 62.975 7.695 ;
        RECT 63.165 7.525 63.335 7.695 ;
        RECT 63.525 7.525 63.695 7.695 ;
        RECT 63.885 7.525 64.055 7.695 ;
        RECT 64.245 7.525 64.415 7.695 ;
        RECT 64.605 7.525 64.775 7.695 ;
        RECT 65.095 7.525 65.265 7.695 ;
        RECT 65.455 7.525 65.625 7.695 ;
        RECT 65.815 7.525 65.985 7.695 ;
        RECT 66.175 7.525 66.345 7.695 ;
        RECT 66.535 7.525 66.705 7.695 ;
        RECT 66.895 7.525 67.065 7.695 ;
        RECT 67.615 7.525 67.785 7.695 ;
        RECT 67.975 7.525 68.145 7.695 ;
        RECT 68.335 7.525 68.505 7.695 ;
        RECT 68.695 7.525 68.865 7.695 ;
        RECT 69.055 7.525 69.225 7.695 ;
        RECT 69.415 7.525 69.585 7.695 ;
        RECT 69.905 7.525 70.075 7.695 ;
        RECT 70.265 7.525 70.435 7.695 ;
        RECT 70.625 7.525 70.795 7.695 ;
        RECT 70.985 7.525 71.155 7.695 ;
        RECT 71.345 7.525 71.515 7.695 ;
        RECT 71.705 7.525 71.875 7.695 ;
        RECT 72.425 7.525 72.595 7.695 ;
        RECT 72.785 7.525 72.955 7.695 ;
        RECT 73.145 7.525 73.315 7.695 ;
        RECT 73.505 7.525 73.675 7.695 ;
        RECT 73.865 7.525 74.035 7.695 ;
        RECT 74.225 7.525 74.395 7.695 ;
        RECT 74.715 7.525 74.885 7.695 ;
        RECT 75.075 7.525 75.245 7.695 ;
        RECT 75.435 7.525 75.605 7.695 ;
        RECT 75.795 7.525 75.965 7.695 ;
        RECT 76.155 7.525 76.325 7.695 ;
        RECT 76.515 7.525 76.685 7.695 ;
        RECT 77.235 7.525 77.405 7.695 ;
        RECT 77.595 7.525 77.765 7.695 ;
        RECT 77.955 7.525 78.125 7.695 ;
        RECT 78.315 7.525 78.485 7.695 ;
        RECT 78.675 7.525 78.845 7.695 ;
        RECT 79.035 7.525 79.205 7.695 ;
        RECT 79.525 7.525 79.695 7.695 ;
        RECT 79.885 7.525 80.055 7.695 ;
        RECT 80.245 7.525 80.415 7.695 ;
        RECT 80.605 7.525 80.775 7.695 ;
        RECT 80.965 7.525 81.135 7.695 ;
        RECT 81.325 7.525 81.495 7.695 ;
        RECT 82.045 7.525 82.215 7.695 ;
        RECT 82.405 7.525 82.575 7.695 ;
        RECT 82.765 7.525 82.935 7.695 ;
        RECT 83.125 7.525 83.295 7.695 ;
        RECT 83.485 7.525 83.655 7.695 ;
        RECT 83.845 7.525 84.015 7.695 ;
        RECT 84.335 7.525 84.505 7.695 ;
        RECT 84.695 7.525 84.865 7.695 ;
        RECT 85.055 7.525 85.225 7.695 ;
        RECT 85.415 7.525 85.585 7.695 ;
        RECT 85.775 7.525 85.945 7.695 ;
        RECT 86.135 7.525 86.305 7.695 ;
        RECT 86.855 7.525 87.025 7.695 ;
        RECT 87.215 7.525 87.385 7.695 ;
        RECT 87.575 7.525 87.745 7.695 ;
        RECT 87.935 7.525 88.105 7.695 ;
        RECT 88.385 7.525 88.555 7.695 ;
        RECT 88.745 7.525 88.915 7.695 ;
        RECT 89.105 7.525 89.275 7.695 ;
        RECT 89.465 7.525 89.635 7.695 ;
        RECT 90.185 7.525 90.355 7.695 ;
        RECT 90.545 7.525 90.715 7.695 ;
        RECT 90.905 7.525 91.075 7.695 ;
        RECT 91.265 7.525 91.435 7.695 ;
        RECT 91.715 7.525 91.885 7.695 ;
        RECT 92.075 7.525 92.245 7.695 ;
        RECT 92.435 7.525 92.605 7.695 ;
        RECT 92.795 7.525 92.965 7.695 ;
        RECT 93.515 7.525 93.685 7.695 ;
        RECT 93.875 7.525 94.045 7.695 ;
        RECT 94.235 7.525 94.405 7.695 ;
        RECT 94.595 7.525 94.765 7.695 ;
        RECT 95.045 7.525 95.215 7.695 ;
        RECT 95.405 7.525 95.575 7.695 ;
        RECT 95.765 7.525 95.935 7.695 ;
        RECT 96.125 7.525 96.295 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 96.725 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 66.388802 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 96.855 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 4.525 -0.075 5.095 -0.065 ;
        RECT 9.335 -0.075 9.905 -0.065 ;
        RECT 14.145 -0.075 14.715 -0.065 ;
        RECT 18.955 -0.075 19.525 -0.065 ;
        RECT 23.765 -0.075 24.335 -0.065 ;
        RECT 28.575 -0.075 29.145 -0.065 ;
        RECT 33.385 -0.075 33.955 -0.065 ;
        RECT 38.195 -0.075 38.765 -0.065 ;
        RECT 43.005 -0.075 43.575 -0.065 ;
        RECT 47.815 -0.075 48.385 -0.065 ;
        RECT 52.625 -0.075 53.195 -0.065 ;
        RECT 57.435 -0.075 58.005 -0.065 ;
        RECT 62.245 -0.075 62.815 -0.065 ;
        RECT 67.055 -0.075 67.625 -0.065 ;
        RECT 71.865 -0.075 72.435 -0.065 ;
        RECT 76.675 -0.075 77.245 -0.065 ;
        RECT 81.485 -0.075 82.055 -0.065 ;
        RECT 86.295 -0.075 86.865 -0.065 ;
        RECT 89.625 -0.075 90.195 -0.065 ;
        RECT 92.955 -0.075 93.525 -0.065 ;
        RECT 96.285 -0.075 96.855 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 0.990 0.310 1.160 1.270 ;
        RECT 4.655 0.310 4.965 2.860 ;
        RECT 5.800 0.310 5.970 1.270 ;
        RECT 9.465 0.310 9.775 2.860 ;
        RECT 10.610 0.310 10.780 1.270 ;
        RECT 14.275 0.310 14.585 2.860 ;
        RECT 15.420 0.310 15.590 1.270 ;
        RECT 19.085 0.310 19.395 2.860 ;
        RECT 20.230 0.310 20.400 1.270 ;
        RECT 23.895 0.310 24.205 2.860 ;
        RECT 25.040 0.310 25.210 1.270 ;
        RECT 28.705 0.310 29.015 2.860 ;
        RECT 29.850 0.310 30.020 1.270 ;
        RECT 33.515 0.310 33.825 2.860 ;
        RECT 34.660 0.310 34.830 1.270 ;
        RECT 38.325 0.310 38.635 2.860 ;
        RECT 39.470 0.310 39.640 1.270 ;
        RECT 43.135 0.310 43.445 2.860 ;
        RECT 44.280 0.310 44.450 1.270 ;
        RECT 47.945 0.310 48.255 2.860 ;
        RECT 49.090 0.310 49.260 1.270 ;
        RECT 52.755 0.310 53.065 2.860 ;
        RECT 53.900 0.310 54.070 1.270 ;
        RECT 57.565 0.310 57.875 2.860 ;
        RECT 58.710 0.310 58.880 1.270 ;
        RECT 62.375 0.310 62.685 2.860 ;
        RECT 63.520 0.310 63.690 1.270 ;
        RECT 67.185 0.310 67.495 2.860 ;
        RECT 68.330 0.310 68.500 1.270 ;
        RECT 71.995 0.310 72.305 2.860 ;
        RECT 73.140 0.310 73.310 1.270 ;
        RECT 76.805 0.310 77.115 2.860 ;
        RECT 77.950 0.310 78.120 1.270 ;
        RECT 81.615 0.310 81.925 2.860 ;
        RECT 82.760 0.310 82.930 1.270 ;
        RECT 86.425 0.310 86.735 2.860 ;
        RECT 87.675 0.310 87.845 1.260 ;
        RECT 89.755 0.310 90.065 2.860 ;
        RECT 91.005 0.310 91.175 1.260 ;
        RECT 93.085 0.310 93.395 2.860 ;
        RECT 94.335 0.310 94.505 1.260 ;
        RECT 96.415 0.310 96.725 2.860 ;
        RECT -0.155 0.235 91.975 0.310 ;
        RECT 92.145 0.235 96.725 0.310 ;
        RECT -0.155 0.000 96.725 0.235 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 0.995 0.065 1.165 0.235 ;
        RECT 1.355 0.065 1.525 0.235 ;
        RECT 1.715 0.065 1.885 0.235 ;
        RECT 2.075 0.065 2.245 0.235 ;
        RECT 2.565 0.065 2.735 0.235 ;
        RECT 2.925 0.065 3.095 0.235 ;
        RECT 3.285 0.065 3.455 0.235 ;
        RECT 3.645 0.065 3.815 0.235 ;
        RECT 4.005 0.065 4.175 0.235 ;
        RECT 4.365 0.065 4.535 0.235 ;
        RECT 5.085 0.065 5.255 0.235 ;
        RECT 5.445 0.065 5.615 0.235 ;
        RECT 5.805 0.065 5.975 0.235 ;
        RECT 6.165 0.065 6.335 0.235 ;
        RECT 6.525 0.065 6.695 0.235 ;
        RECT 6.885 0.065 7.055 0.235 ;
        RECT 7.375 0.065 7.545 0.235 ;
        RECT 7.735 0.065 7.905 0.235 ;
        RECT 8.095 0.065 8.265 0.235 ;
        RECT 8.455 0.065 8.625 0.235 ;
        RECT 8.815 0.065 8.985 0.235 ;
        RECT 9.175 0.065 9.345 0.235 ;
        RECT 9.895 0.065 10.065 0.235 ;
        RECT 10.255 0.065 10.425 0.235 ;
        RECT 10.615 0.065 10.785 0.235 ;
        RECT 10.975 0.065 11.145 0.235 ;
        RECT 11.335 0.065 11.505 0.235 ;
        RECT 11.695 0.065 11.865 0.235 ;
        RECT 12.185 0.065 12.355 0.235 ;
        RECT 12.545 0.065 12.715 0.235 ;
        RECT 12.905 0.065 13.075 0.235 ;
        RECT 13.265 0.065 13.435 0.235 ;
        RECT 13.625 0.065 13.795 0.235 ;
        RECT 13.985 0.065 14.155 0.235 ;
        RECT 14.705 0.065 14.875 0.235 ;
        RECT 15.065 0.065 15.235 0.235 ;
        RECT 15.425 0.065 15.595 0.235 ;
        RECT 15.785 0.065 15.955 0.235 ;
        RECT 16.145 0.065 16.315 0.235 ;
        RECT 16.505 0.065 16.675 0.235 ;
        RECT 16.995 0.065 17.165 0.235 ;
        RECT 17.355 0.065 17.525 0.235 ;
        RECT 17.715 0.065 17.885 0.235 ;
        RECT 18.075 0.065 18.245 0.235 ;
        RECT 18.435 0.065 18.605 0.235 ;
        RECT 18.795 0.065 18.965 0.235 ;
        RECT 19.515 0.065 19.685 0.235 ;
        RECT 19.875 0.065 20.045 0.235 ;
        RECT 20.235 0.065 20.405 0.235 ;
        RECT 20.595 0.065 20.765 0.235 ;
        RECT 20.955 0.065 21.125 0.235 ;
        RECT 21.315 0.065 21.485 0.235 ;
        RECT 21.805 0.065 21.975 0.235 ;
        RECT 22.165 0.065 22.335 0.235 ;
        RECT 22.525 0.065 22.695 0.235 ;
        RECT 22.885 0.065 23.055 0.235 ;
        RECT 23.245 0.065 23.415 0.235 ;
        RECT 23.605 0.065 23.775 0.235 ;
        RECT 24.325 0.065 24.495 0.235 ;
        RECT 24.685 0.065 24.855 0.235 ;
        RECT 25.045 0.065 25.215 0.235 ;
        RECT 25.405 0.065 25.575 0.235 ;
        RECT 25.765 0.065 25.935 0.235 ;
        RECT 26.125 0.065 26.295 0.235 ;
        RECT 26.615 0.065 26.785 0.235 ;
        RECT 26.975 0.065 27.145 0.235 ;
        RECT 27.335 0.065 27.505 0.235 ;
        RECT 27.695 0.065 27.865 0.235 ;
        RECT 28.055 0.065 28.225 0.235 ;
        RECT 28.415 0.065 28.585 0.235 ;
        RECT 29.135 0.065 29.305 0.235 ;
        RECT 29.495 0.065 29.665 0.235 ;
        RECT 29.855 0.065 30.025 0.235 ;
        RECT 30.215 0.065 30.385 0.235 ;
        RECT 30.575 0.065 30.745 0.235 ;
        RECT 30.935 0.065 31.105 0.235 ;
        RECT 31.425 0.065 31.595 0.235 ;
        RECT 31.785 0.065 31.955 0.235 ;
        RECT 32.145 0.065 32.315 0.235 ;
        RECT 32.505 0.065 32.675 0.235 ;
        RECT 32.865 0.065 33.035 0.235 ;
        RECT 33.225 0.065 33.395 0.235 ;
        RECT 33.945 0.065 34.115 0.235 ;
        RECT 34.305 0.065 34.475 0.235 ;
        RECT 34.665 0.065 34.835 0.235 ;
        RECT 35.025 0.065 35.195 0.235 ;
        RECT 35.385 0.065 35.555 0.235 ;
        RECT 35.745 0.065 35.915 0.235 ;
        RECT 36.235 0.065 36.405 0.235 ;
        RECT 36.595 0.065 36.765 0.235 ;
        RECT 36.955 0.065 37.125 0.235 ;
        RECT 37.315 0.065 37.485 0.235 ;
        RECT 37.675 0.065 37.845 0.235 ;
        RECT 38.035 0.065 38.205 0.235 ;
        RECT 38.755 0.065 38.925 0.235 ;
        RECT 39.115 0.065 39.285 0.235 ;
        RECT 39.475 0.065 39.645 0.235 ;
        RECT 39.835 0.065 40.005 0.235 ;
        RECT 40.195 0.065 40.365 0.235 ;
        RECT 40.555 0.065 40.725 0.235 ;
        RECT 41.045 0.065 41.215 0.235 ;
        RECT 41.405 0.065 41.575 0.235 ;
        RECT 41.765 0.065 41.935 0.235 ;
        RECT 42.125 0.065 42.295 0.235 ;
        RECT 42.485 0.065 42.655 0.235 ;
        RECT 42.845 0.065 43.015 0.235 ;
        RECT 43.565 0.065 43.735 0.235 ;
        RECT 43.925 0.065 44.095 0.235 ;
        RECT 44.285 0.065 44.455 0.235 ;
        RECT 44.645 0.065 44.815 0.235 ;
        RECT 45.005 0.065 45.175 0.235 ;
        RECT 45.365 0.065 45.535 0.235 ;
        RECT 45.855 0.065 46.025 0.235 ;
        RECT 46.215 0.065 46.385 0.235 ;
        RECT 46.575 0.065 46.745 0.235 ;
        RECT 46.935 0.065 47.105 0.235 ;
        RECT 47.295 0.065 47.465 0.235 ;
        RECT 47.655 0.065 47.825 0.235 ;
        RECT 48.375 0.065 48.545 0.235 ;
        RECT 48.735 0.065 48.905 0.235 ;
        RECT 49.095 0.065 49.265 0.235 ;
        RECT 49.455 0.065 49.625 0.235 ;
        RECT 49.815 0.065 49.985 0.235 ;
        RECT 50.175 0.065 50.345 0.235 ;
        RECT 50.665 0.065 50.835 0.235 ;
        RECT 51.025 0.065 51.195 0.235 ;
        RECT 51.385 0.065 51.555 0.235 ;
        RECT 51.745 0.065 51.915 0.235 ;
        RECT 52.105 0.065 52.275 0.235 ;
        RECT 52.465 0.065 52.635 0.235 ;
        RECT 53.185 0.065 53.355 0.235 ;
        RECT 53.545 0.065 53.715 0.235 ;
        RECT 53.905 0.065 54.075 0.235 ;
        RECT 54.265 0.065 54.435 0.235 ;
        RECT 54.625 0.065 54.795 0.235 ;
        RECT 54.985 0.065 55.155 0.235 ;
        RECT 55.475 0.065 55.645 0.235 ;
        RECT 55.835 0.065 56.005 0.235 ;
        RECT 56.195 0.065 56.365 0.235 ;
        RECT 56.555 0.065 56.725 0.235 ;
        RECT 56.915 0.065 57.085 0.235 ;
        RECT 57.275 0.065 57.445 0.235 ;
        RECT 57.995 0.065 58.165 0.235 ;
        RECT 58.355 0.065 58.525 0.235 ;
        RECT 58.715 0.065 58.885 0.235 ;
        RECT 59.075 0.065 59.245 0.235 ;
        RECT 59.435 0.065 59.605 0.235 ;
        RECT 59.795 0.065 59.965 0.235 ;
        RECT 60.285 0.065 60.455 0.235 ;
        RECT 60.645 0.065 60.815 0.235 ;
        RECT 61.005 0.065 61.175 0.235 ;
        RECT 61.365 0.065 61.535 0.235 ;
        RECT 61.725 0.065 61.895 0.235 ;
        RECT 62.085 0.065 62.255 0.235 ;
        RECT 62.805 0.065 62.975 0.235 ;
        RECT 63.165 0.065 63.335 0.235 ;
        RECT 63.525 0.065 63.695 0.235 ;
        RECT 63.885 0.065 64.055 0.235 ;
        RECT 64.245 0.065 64.415 0.235 ;
        RECT 64.605 0.065 64.775 0.235 ;
        RECT 65.095 0.065 65.265 0.235 ;
        RECT 65.455 0.065 65.625 0.235 ;
        RECT 65.815 0.065 65.985 0.235 ;
        RECT 66.175 0.065 66.345 0.235 ;
        RECT 66.535 0.065 66.705 0.235 ;
        RECT 66.895 0.065 67.065 0.235 ;
        RECT 67.615 0.065 67.785 0.235 ;
        RECT 67.975 0.065 68.145 0.235 ;
        RECT 68.335 0.065 68.505 0.235 ;
        RECT 68.695 0.065 68.865 0.235 ;
        RECT 69.055 0.065 69.225 0.235 ;
        RECT 69.415 0.065 69.585 0.235 ;
        RECT 69.905 0.065 70.075 0.235 ;
        RECT 70.265 0.065 70.435 0.235 ;
        RECT 70.625 0.065 70.795 0.235 ;
        RECT 70.985 0.065 71.155 0.235 ;
        RECT 71.345 0.065 71.515 0.235 ;
        RECT 71.705 0.065 71.875 0.235 ;
        RECT 72.425 0.065 72.595 0.235 ;
        RECT 72.785 0.065 72.955 0.235 ;
        RECT 73.145 0.065 73.315 0.235 ;
        RECT 73.505 0.065 73.675 0.235 ;
        RECT 73.865 0.065 74.035 0.235 ;
        RECT 74.225 0.065 74.395 0.235 ;
        RECT 74.715 0.065 74.885 0.235 ;
        RECT 75.075 0.065 75.245 0.235 ;
        RECT 75.435 0.065 75.605 0.235 ;
        RECT 75.795 0.065 75.965 0.235 ;
        RECT 76.155 0.065 76.325 0.235 ;
        RECT 76.515 0.065 76.685 0.235 ;
        RECT 77.235 0.065 77.405 0.235 ;
        RECT 77.595 0.065 77.765 0.235 ;
        RECT 77.955 0.065 78.125 0.235 ;
        RECT 78.315 0.065 78.485 0.235 ;
        RECT 78.675 0.065 78.845 0.235 ;
        RECT 79.035 0.065 79.205 0.235 ;
        RECT 79.525 0.065 79.695 0.235 ;
        RECT 79.885 0.065 80.055 0.235 ;
        RECT 80.245 0.065 80.415 0.235 ;
        RECT 80.605 0.065 80.775 0.235 ;
        RECT 80.965 0.065 81.135 0.235 ;
        RECT 81.325 0.065 81.495 0.235 ;
        RECT 82.045 0.065 82.215 0.235 ;
        RECT 82.405 0.065 82.575 0.235 ;
        RECT 82.765 0.065 82.935 0.235 ;
        RECT 83.125 0.065 83.295 0.235 ;
        RECT 83.485 0.065 83.655 0.235 ;
        RECT 83.845 0.065 84.015 0.235 ;
        RECT 84.335 0.065 84.505 0.235 ;
        RECT 84.695 0.065 84.865 0.235 ;
        RECT 85.055 0.065 85.225 0.235 ;
        RECT 85.415 0.065 85.585 0.235 ;
        RECT 85.775 0.065 85.945 0.235 ;
        RECT 86.135 0.065 86.305 0.235 ;
        RECT 86.855 0.065 87.025 0.235 ;
        RECT 87.215 0.065 87.385 0.235 ;
        RECT 87.575 0.065 87.745 0.235 ;
        RECT 87.935 0.065 88.105 0.235 ;
        RECT 88.385 0.065 88.555 0.235 ;
        RECT 88.745 0.065 88.915 0.235 ;
        RECT 89.105 0.065 89.275 0.235 ;
        RECT 89.465 0.065 89.635 0.235 ;
        RECT 90.185 0.065 90.355 0.235 ;
        RECT 90.545 0.065 90.715 0.235 ;
        RECT 90.905 0.065 91.075 0.235 ;
        RECT 91.265 0.065 91.435 0.235 ;
        RECT 91.715 0.065 91.885 0.235 ;
        RECT 92.075 0.065 92.245 0.235 ;
        RECT 92.435 0.065 92.605 0.235 ;
        RECT 92.795 0.065 92.965 0.235 ;
        RECT 93.515 0.065 93.685 0.235 ;
        RECT 93.875 0.065 94.045 0.235 ;
        RECT 94.235 0.065 94.405 0.235 ;
        RECT 94.595 0.065 94.765 0.235 ;
        RECT 95.045 0.065 95.215 0.235 ;
        RECT 95.405 0.065 95.575 0.235 ;
        RECT 95.765 0.065 95.935 0.235 ;
        RECT 96.125 0.065 96.295 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 96.725 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 1.445 5.470 1.615 7.250 ;
        RECT 2.325 5.470 2.495 7.250 ;
        RECT 3.205 5.470 3.375 7.250 ;
        RECT 6.255 5.470 6.425 7.250 ;
        RECT 7.135 5.470 7.305 7.250 ;
        RECT 8.015 5.470 8.185 7.250 ;
        RECT 11.065 5.470 11.235 7.250 ;
        RECT 11.945 5.470 12.115 7.250 ;
        RECT 12.825 5.470 12.995 7.250 ;
        RECT 15.875 5.470 16.045 7.250 ;
        RECT 16.755 5.470 16.925 7.250 ;
        RECT 17.635 5.470 17.805 7.250 ;
        RECT 20.685 5.470 20.855 7.250 ;
        RECT 21.565 5.470 21.735 7.250 ;
        RECT 22.445 5.470 22.615 7.250 ;
        RECT 25.495 5.470 25.665 7.250 ;
        RECT 26.375 5.470 26.545 7.250 ;
        RECT 27.255 5.470 27.425 7.250 ;
        RECT 30.305 5.470 30.475 7.250 ;
        RECT 31.185 5.470 31.355 7.250 ;
        RECT 32.065 5.470 32.235 7.250 ;
        RECT 35.115 5.470 35.285 7.250 ;
        RECT 35.995 5.470 36.165 7.250 ;
        RECT 36.875 5.470 37.045 7.250 ;
        RECT 39.925 5.470 40.095 7.250 ;
        RECT 40.805 5.470 40.975 7.250 ;
        RECT 41.685 5.470 41.855 7.250 ;
        RECT 44.735 5.470 44.905 7.250 ;
        RECT 45.615 5.470 45.785 7.250 ;
        RECT 46.495 5.470 46.665 7.250 ;
        RECT 49.545 5.470 49.715 7.250 ;
        RECT 50.425 5.470 50.595 7.250 ;
        RECT 51.305 5.470 51.475 7.250 ;
        RECT 54.355 5.470 54.525 7.250 ;
        RECT 55.235 5.470 55.405 7.250 ;
        RECT 56.115 5.470 56.285 7.250 ;
        RECT 59.165 5.470 59.335 7.250 ;
        RECT 60.045 5.470 60.215 7.250 ;
        RECT 60.925 5.470 61.095 7.250 ;
        RECT 63.975 5.470 64.145 7.250 ;
        RECT 64.855 5.470 65.025 7.250 ;
        RECT 65.735 5.470 65.905 7.250 ;
        RECT 68.785 5.470 68.955 7.250 ;
        RECT 69.665 5.470 69.835 7.250 ;
        RECT 70.545 5.470 70.715 7.250 ;
        RECT 73.595 5.470 73.765 7.250 ;
        RECT 74.475 5.470 74.645 7.250 ;
        RECT 75.355 5.470 75.525 7.250 ;
        RECT 78.405 5.470 78.575 7.250 ;
        RECT 79.285 5.470 79.455 7.250 ;
        RECT 80.165 5.470 80.335 7.250 ;
        RECT 83.215 5.470 83.385 7.250 ;
        RECT 84.095 5.470 84.265 7.250 ;
        RECT 84.975 5.470 85.145 7.250 ;
        RECT 87.725 7.055 87.905 7.225 ;
        RECT 87.725 5.525 87.895 7.055 ;
        RECT 88.605 5.525 88.775 7.225 ;
        RECT 1.445 5.300 4.155 5.470 ;
        RECT 6.255 5.300 8.965 5.470 ;
        RECT 11.065 5.300 13.775 5.470 ;
        RECT 15.875 5.300 18.585 5.470 ;
        RECT 20.685 5.300 23.395 5.470 ;
        RECT 25.495 5.300 28.205 5.470 ;
        RECT 30.305 5.300 33.015 5.470 ;
        RECT 35.115 5.300 37.825 5.470 ;
        RECT 39.925 5.300 42.635 5.470 ;
        RECT 44.735 5.300 47.445 5.470 ;
        RECT 49.545 5.300 52.255 5.470 ;
        RECT 54.355 5.300 57.065 5.470 ;
        RECT 59.165 5.300 61.875 5.470 ;
        RECT 63.975 5.300 66.685 5.470 ;
        RECT 68.785 5.300 71.495 5.470 ;
        RECT 73.595 5.300 76.305 5.470 ;
        RECT 78.405 5.300 81.115 5.470 ;
        RECT 83.215 5.300 85.925 5.470 ;
        RECT 87.725 5.355 88.775 5.525 ;
        RECT 3.245 2.055 3.415 5.095 ;
        RECT 0.505 1.815 0.675 1.895 ;
        RECT 1.475 1.815 1.645 1.895 ;
        RECT 2.445 1.815 2.615 1.895 ;
        RECT 0.505 1.645 2.615 1.815 ;
        RECT 0.505 0.515 0.675 1.645 ;
        RECT 1.475 0.765 1.645 1.645 ;
        RECT 2.445 1.565 2.615 1.645 ;
        RECT 1.965 1.220 2.135 1.300 ;
        RECT 3.015 1.220 3.185 1.895 ;
        RECT 3.985 1.890 4.155 5.300 ;
        RECT 5.835 2.055 6.005 5.095 ;
        RECT 8.055 4.235 8.225 5.095 ;
        RECT 8.050 3.905 8.225 4.235 ;
        RECT 8.055 2.055 8.225 3.905 ;
        RECT 1.965 1.050 3.185 1.220 ;
        RECT 1.965 0.970 2.135 1.050 ;
        RECT 2.445 0.765 2.615 0.845 ;
        RECT 1.475 0.595 2.615 0.765 ;
        RECT 1.475 0.515 1.645 0.595 ;
        RECT 2.445 0.515 2.615 0.595 ;
        RECT 3.015 0.765 3.185 1.050 ;
        RECT 3.500 1.720 4.155 1.890 ;
        RECT 5.315 1.815 5.485 1.895 ;
        RECT 6.285 1.815 6.455 1.895 ;
        RECT 7.255 1.815 7.425 1.895 ;
        RECT 3.500 0.985 3.670 1.720 ;
        RECT 5.315 1.645 7.425 1.815 ;
        RECT 3.985 0.765 4.155 1.535 ;
        RECT 3.015 0.595 4.155 0.765 ;
        RECT 3.015 0.515 3.185 0.595 ;
        RECT 3.985 0.515 4.155 0.595 ;
        RECT 5.315 0.515 5.485 1.645 ;
        RECT 6.285 0.765 6.455 1.645 ;
        RECT 7.255 1.565 7.425 1.645 ;
        RECT 6.775 1.220 6.945 1.300 ;
        RECT 7.825 1.220 7.995 1.895 ;
        RECT 8.795 1.890 8.965 5.300 ;
        RECT 10.645 2.055 10.815 5.095 ;
        RECT 12.865 2.055 13.035 5.095 ;
        RECT 6.775 1.050 7.995 1.220 ;
        RECT 6.775 0.970 6.945 1.050 ;
        RECT 7.255 0.765 7.425 0.845 ;
        RECT 6.285 0.595 7.425 0.765 ;
        RECT 6.285 0.515 6.455 0.595 ;
        RECT 7.255 0.515 7.425 0.595 ;
        RECT 7.825 0.765 7.995 1.050 ;
        RECT 8.310 1.720 8.965 1.890 ;
        RECT 10.125 1.815 10.295 1.895 ;
        RECT 11.095 1.815 11.265 1.895 ;
        RECT 12.065 1.815 12.235 1.895 ;
        RECT 8.310 0.985 8.480 1.720 ;
        RECT 10.125 1.645 12.235 1.815 ;
        RECT 8.795 0.765 8.965 1.535 ;
        RECT 7.825 0.595 8.965 0.765 ;
        RECT 7.825 0.515 7.995 0.595 ;
        RECT 8.795 0.515 8.965 0.595 ;
        RECT 10.125 0.515 10.295 1.645 ;
        RECT 11.095 0.765 11.265 1.645 ;
        RECT 12.065 1.565 12.235 1.645 ;
        RECT 11.585 1.220 11.755 1.300 ;
        RECT 12.635 1.220 12.805 1.895 ;
        RECT 13.605 1.890 13.775 5.300 ;
        RECT 15.455 2.055 15.625 5.095 ;
        RECT 11.585 1.050 12.805 1.220 ;
        RECT 11.585 0.970 11.755 1.050 ;
        RECT 12.065 0.765 12.235 0.845 ;
        RECT 11.095 0.595 12.235 0.765 ;
        RECT 11.095 0.515 11.265 0.595 ;
        RECT 12.065 0.515 12.235 0.595 ;
        RECT 12.635 0.765 12.805 1.050 ;
        RECT 13.120 1.720 13.775 1.890 ;
        RECT 14.935 1.815 15.105 1.895 ;
        RECT 15.905 1.815 16.075 1.895 ;
        RECT 16.875 1.815 17.045 1.895 ;
        RECT 13.120 0.985 13.290 1.720 ;
        RECT 14.935 1.645 17.045 1.815 ;
        RECT 13.605 0.765 13.775 1.535 ;
        RECT 12.635 0.595 13.775 0.765 ;
        RECT 12.635 0.515 12.805 0.595 ;
        RECT 13.605 0.515 13.775 0.595 ;
        RECT 14.935 0.515 15.105 1.645 ;
        RECT 15.905 0.765 16.075 1.645 ;
        RECT 16.875 1.565 17.045 1.645 ;
        RECT 16.395 1.220 16.565 1.300 ;
        RECT 17.445 1.220 17.615 1.895 ;
        RECT 18.415 1.890 18.585 5.300 ;
        RECT 20.265 2.055 20.435 5.095 ;
        RECT 22.485 2.055 22.655 5.095 ;
        RECT 16.395 1.050 17.615 1.220 ;
        RECT 16.395 0.970 16.565 1.050 ;
        RECT 16.875 0.765 17.045 0.845 ;
        RECT 15.905 0.595 17.045 0.765 ;
        RECT 15.905 0.515 16.075 0.595 ;
        RECT 16.875 0.515 17.045 0.595 ;
        RECT 17.445 0.765 17.615 1.050 ;
        RECT 17.930 1.720 18.585 1.890 ;
        RECT 19.745 1.815 19.915 1.895 ;
        RECT 20.715 1.815 20.885 1.895 ;
        RECT 21.685 1.815 21.855 1.895 ;
        RECT 17.930 0.985 18.100 1.720 ;
        RECT 19.745 1.645 21.855 1.815 ;
        RECT 18.415 0.765 18.585 1.535 ;
        RECT 17.445 0.595 18.585 0.765 ;
        RECT 17.445 0.515 17.615 0.595 ;
        RECT 18.415 0.515 18.585 0.595 ;
        RECT 19.745 0.515 19.915 1.645 ;
        RECT 20.715 0.765 20.885 1.645 ;
        RECT 21.685 1.565 21.855 1.645 ;
        RECT 21.205 1.220 21.375 1.300 ;
        RECT 22.255 1.220 22.425 1.895 ;
        RECT 23.225 1.890 23.395 5.300 ;
        RECT 25.075 2.055 25.245 5.095 ;
        RECT 27.295 2.055 27.465 5.095 ;
        RECT 21.205 1.050 22.425 1.220 ;
        RECT 21.205 0.970 21.375 1.050 ;
        RECT 21.685 0.765 21.855 0.845 ;
        RECT 20.715 0.595 21.855 0.765 ;
        RECT 20.715 0.515 20.885 0.595 ;
        RECT 21.685 0.515 21.855 0.595 ;
        RECT 22.255 0.765 22.425 1.050 ;
        RECT 22.740 1.720 23.395 1.890 ;
        RECT 24.555 1.815 24.725 1.895 ;
        RECT 25.525 1.815 25.695 1.895 ;
        RECT 26.495 1.815 26.665 1.895 ;
        RECT 22.740 0.985 22.910 1.720 ;
        RECT 24.555 1.645 26.665 1.815 ;
        RECT 23.225 0.765 23.395 1.535 ;
        RECT 22.255 0.595 23.395 0.765 ;
        RECT 22.255 0.515 22.425 0.595 ;
        RECT 23.225 0.515 23.395 0.595 ;
        RECT 24.555 0.515 24.725 1.645 ;
        RECT 25.525 0.765 25.695 1.645 ;
        RECT 26.495 1.565 26.665 1.645 ;
        RECT 26.015 1.220 26.185 1.300 ;
        RECT 27.065 1.220 27.235 1.895 ;
        RECT 28.035 1.890 28.205 5.300 ;
        RECT 32.105 2.055 32.275 5.095 ;
        RECT 26.015 1.050 27.235 1.220 ;
        RECT 26.015 0.970 26.185 1.050 ;
        RECT 26.495 0.765 26.665 0.845 ;
        RECT 25.525 0.595 26.665 0.765 ;
        RECT 25.525 0.515 25.695 0.595 ;
        RECT 26.495 0.515 26.665 0.595 ;
        RECT 27.065 0.765 27.235 1.050 ;
        RECT 27.550 1.720 28.205 1.890 ;
        RECT 29.365 1.815 29.535 1.895 ;
        RECT 30.335 1.815 30.505 1.895 ;
        RECT 31.305 1.815 31.475 1.895 ;
        RECT 27.550 0.985 27.720 1.720 ;
        RECT 29.365 1.645 31.475 1.815 ;
        RECT 28.035 0.765 28.205 1.535 ;
        RECT 27.065 0.595 28.205 0.765 ;
        RECT 27.065 0.515 27.235 0.595 ;
        RECT 28.035 0.515 28.205 0.595 ;
        RECT 29.365 0.515 29.535 1.645 ;
        RECT 30.335 0.765 30.505 1.645 ;
        RECT 31.305 1.565 31.475 1.645 ;
        RECT 30.825 1.220 30.995 1.300 ;
        RECT 31.875 1.220 32.045 1.895 ;
        RECT 32.845 1.890 33.015 5.300 ;
        RECT 34.695 2.055 34.865 5.095 ;
        RECT 36.915 4.235 37.085 5.095 ;
        RECT 36.910 3.905 37.085 4.235 ;
        RECT 36.915 2.055 37.085 3.905 ;
        RECT 30.825 1.050 32.045 1.220 ;
        RECT 30.825 0.970 30.995 1.050 ;
        RECT 31.305 0.765 31.475 0.845 ;
        RECT 30.335 0.595 31.475 0.765 ;
        RECT 30.335 0.515 30.505 0.595 ;
        RECT 31.305 0.515 31.475 0.595 ;
        RECT 31.875 0.765 32.045 1.050 ;
        RECT 32.360 1.720 33.015 1.890 ;
        RECT 34.175 1.815 34.345 1.895 ;
        RECT 35.145 1.815 35.315 1.895 ;
        RECT 36.115 1.815 36.285 1.895 ;
        RECT 32.360 0.985 32.530 1.720 ;
        RECT 34.175 1.645 36.285 1.815 ;
        RECT 32.845 0.765 33.015 1.535 ;
        RECT 31.875 0.595 33.015 0.765 ;
        RECT 31.875 0.515 32.045 0.595 ;
        RECT 32.845 0.515 33.015 0.595 ;
        RECT 34.175 0.515 34.345 1.645 ;
        RECT 35.145 0.765 35.315 1.645 ;
        RECT 36.115 1.565 36.285 1.645 ;
        RECT 35.635 1.220 35.805 1.300 ;
        RECT 36.685 1.220 36.855 1.895 ;
        RECT 37.655 1.890 37.825 5.300 ;
        RECT 39.505 2.055 39.675 5.095 ;
        RECT 41.725 2.055 41.895 5.095 ;
        RECT 35.635 1.050 36.855 1.220 ;
        RECT 35.635 0.970 35.805 1.050 ;
        RECT 36.115 0.765 36.285 0.845 ;
        RECT 35.145 0.595 36.285 0.765 ;
        RECT 35.145 0.515 35.315 0.595 ;
        RECT 36.115 0.515 36.285 0.595 ;
        RECT 36.685 0.765 36.855 1.050 ;
        RECT 37.170 1.720 37.825 1.890 ;
        RECT 38.985 1.815 39.155 1.895 ;
        RECT 39.955 1.815 40.125 1.895 ;
        RECT 40.925 1.815 41.095 1.895 ;
        RECT 37.170 0.985 37.340 1.720 ;
        RECT 38.985 1.645 41.095 1.815 ;
        RECT 37.655 0.765 37.825 1.535 ;
        RECT 36.685 0.595 37.825 0.765 ;
        RECT 36.685 0.515 36.855 0.595 ;
        RECT 37.655 0.515 37.825 0.595 ;
        RECT 38.985 0.515 39.155 1.645 ;
        RECT 39.955 0.765 40.125 1.645 ;
        RECT 40.925 1.565 41.095 1.645 ;
        RECT 40.445 1.220 40.615 1.300 ;
        RECT 41.495 1.220 41.665 1.895 ;
        RECT 42.465 1.890 42.635 5.300 ;
        RECT 44.315 2.055 44.485 5.095 ;
        RECT 40.445 1.050 41.665 1.220 ;
        RECT 40.445 0.970 40.615 1.050 ;
        RECT 40.925 0.765 41.095 0.845 ;
        RECT 39.955 0.595 41.095 0.765 ;
        RECT 39.955 0.515 40.125 0.595 ;
        RECT 40.925 0.515 41.095 0.595 ;
        RECT 41.495 0.765 41.665 1.050 ;
        RECT 41.980 1.720 42.635 1.890 ;
        RECT 43.795 1.815 43.965 1.895 ;
        RECT 44.765 1.815 44.935 1.895 ;
        RECT 45.735 1.815 45.905 1.895 ;
        RECT 41.980 0.985 42.150 1.720 ;
        RECT 43.795 1.645 45.905 1.815 ;
        RECT 42.465 0.765 42.635 1.535 ;
        RECT 41.495 0.595 42.635 0.765 ;
        RECT 41.495 0.515 41.665 0.595 ;
        RECT 42.465 0.515 42.635 0.595 ;
        RECT 43.795 0.515 43.965 1.645 ;
        RECT 44.765 0.765 44.935 1.645 ;
        RECT 45.735 1.565 45.905 1.645 ;
        RECT 45.255 1.220 45.425 1.300 ;
        RECT 46.305 1.220 46.475 1.895 ;
        RECT 47.275 1.890 47.445 5.300 ;
        RECT 49.125 2.055 49.295 5.095 ;
        RECT 51.345 2.055 51.515 5.095 ;
        RECT 45.255 1.050 46.475 1.220 ;
        RECT 45.255 0.970 45.425 1.050 ;
        RECT 45.735 0.765 45.905 0.845 ;
        RECT 44.765 0.595 45.905 0.765 ;
        RECT 44.765 0.515 44.935 0.595 ;
        RECT 45.735 0.515 45.905 0.595 ;
        RECT 46.305 0.765 46.475 1.050 ;
        RECT 46.790 1.720 47.445 1.890 ;
        RECT 48.605 1.815 48.775 1.895 ;
        RECT 49.575 1.815 49.745 1.895 ;
        RECT 50.545 1.815 50.715 1.895 ;
        RECT 46.790 0.985 46.960 1.720 ;
        RECT 48.605 1.645 50.715 1.815 ;
        RECT 47.275 0.765 47.445 1.535 ;
        RECT 46.305 0.595 47.445 0.765 ;
        RECT 46.305 0.515 46.475 0.595 ;
        RECT 47.275 0.515 47.445 0.595 ;
        RECT 48.605 0.515 48.775 1.645 ;
        RECT 49.575 0.765 49.745 1.645 ;
        RECT 50.545 1.565 50.715 1.645 ;
        RECT 50.065 1.220 50.235 1.300 ;
        RECT 51.115 1.220 51.285 1.895 ;
        RECT 52.085 1.890 52.255 5.300 ;
        RECT 53.935 2.055 54.105 5.095 ;
        RECT 56.155 2.055 56.325 5.095 ;
        RECT 50.065 1.050 51.285 1.220 ;
        RECT 50.065 0.970 50.235 1.050 ;
        RECT 50.545 0.765 50.715 0.845 ;
        RECT 49.575 0.595 50.715 0.765 ;
        RECT 49.575 0.515 49.745 0.595 ;
        RECT 50.545 0.515 50.715 0.595 ;
        RECT 51.115 0.765 51.285 1.050 ;
        RECT 51.600 1.720 52.255 1.890 ;
        RECT 53.415 1.815 53.585 1.895 ;
        RECT 54.385 1.815 54.555 1.895 ;
        RECT 55.355 1.815 55.525 1.895 ;
        RECT 51.600 0.985 51.770 1.720 ;
        RECT 53.415 1.645 55.525 1.815 ;
        RECT 52.085 0.765 52.255 1.535 ;
        RECT 51.115 0.595 52.255 0.765 ;
        RECT 51.115 0.515 51.285 0.595 ;
        RECT 52.085 0.515 52.255 0.595 ;
        RECT 53.415 0.515 53.585 1.645 ;
        RECT 54.385 0.765 54.555 1.645 ;
        RECT 55.355 1.565 55.525 1.645 ;
        RECT 54.875 1.220 55.045 1.300 ;
        RECT 55.925 1.220 56.095 1.895 ;
        RECT 56.895 1.890 57.065 5.300 ;
        RECT 60.965 2.055 61.135 5.095 ;
        RECT 54.875 1.050 56.095 1.220 ;
        RECT 54.875 0.970 55.045 1.050 ;
        RECT 55.355 0.765 55.525 0.845 ;
        RECT 54.385 0.595 55.525 0.765 ;
        RECT 54.385 0.515 54.555 0.595 ;
        RECT 55.355 0.515 55.525 0.595 ;
        RECT 55.925 0.765 56.095 1.050 ;
        RECT 56.410 1.720 57.065 1.890 ;
        RECT 58.225 1.815 58.395 1.895 ;
        RECT 59.195 1.815 59.365 1.895 ;
        RECT 60.165 1.815 60.335 1.895 ;
        RECT 56.410 0.985 56.580 1.720 ;
        RECT 58.225 1.645 60.335 1.815 ;
        RECT 56.895 0.765 57.065 1.535 ;
        RECT 55.925 0.595 57.065 0.765 ;
        RECT 55.925 0.515 56.095 0.595 ;
        RECT 56.895 0.515 57.065 0.595 ;
        RECT 58.225 0.515 58.395 1.645 ;
        RECT 59.195 0.765 59.365 1.645 ;
        RECT 60.165 1.565 60.335 1.645 ;
        RECT 59.685 1.220 59.855 1.300 ;
        RECT 60.735 1.220 60.905 1.895 ;
        RECT 61.705 1.890 61.875 5.300 ;
        RECT 63.555 2.055 63.725 5.095 ;
        RECT 65.775 4.235 65.945 5.095 ;
        RECT 65.770 3.905 65.945 4.235 ;
        RECT 65.775 2.055 65.945 3.905 ;
        RECT 59.685 1.050 60.905 1.220 ;
        RECT 59.685 0.970 59.855 1.050 ;
        RECT 60.165 0.765 60.335 0.845 ;
        RECT 59.195 0.595 60.335 0.765 ;
        RECT 59.195 0.515 59.365 0.595 ;
        RECT 60.165 0.515 60.335 0.595 ;
        RECT 60.735 0.765 60.905 1.050 ;
        RECT 61.220 1.720 61.875 1.890 ;
        RECT 63.035 1.815 63.205 1.895 ;
        RECT 64.005 1.815 64.175 1.895 ;
        RECT 64.975 1.815 65.145 1.895 ;
        RECT 61.220 0.985 61.390 1.720 ;
        RECT 63.035 1.645 65.145 1.815 ;
        RECT 61.705 0.765 61.875 1.535 ;
        RECT 60.735 0.595 61.875 0.765 ;
        RECT 60.735 0.515 60.905 0.595 ;
        RECT 61.705 0.515 61.875 0.595 ;
        RECT 63.035 0.515 63.205 1.645 ;
        RECT 64.005 0.765 64.175 1.645 ;
        RECT 64.975 1.565 65.145 1.645 ;
        RECT 64.495 1.220 64.665 1.300 ;
        RECT 65.545 1.220 65.715 1.895 ;
        RECT 66.515 1.890 66.685 5.300 ;
        RECT 68.365 2.055 68.535 5.095 ;
        RECT 70.585 2.055 70.755 5.095 ;
        RECT 64.495 1.050 65.715 1.220 ;
        RECT 64.495 0.970 64.665 1.050 ;
        RECT 64.975 0.765 65.145 0.845 ;
        RECT 64.005 0.595 65.145 0.765 ;
        RECT 64.005 0.515 64.175 0.595 ;
        RECT 64.975 0.515 65.145 0.595 ;
        RECT 65.545 0.765 65.715 1.050 ;
        RECT 66.030 1.720 66.685 1.890 ;
        RECT 67.845 1.815 68.015 1.895 ;
        RECT 68.815 1.815 68.985 1.895 ;
        RECT 69.785 1.815 69.955 1.895 ;
        RECT 66.030 0.985 66.200 1.720 ;
        RECT 67.845 1.645 69.955 1.815 ;
        RECT 66.515 0.765 66.685 1.535 ;
        RECT 65.545 0.595 66.685 0.765 ;
        RECT 65.545 0.515 65.715 0.595 ;
        RECT 66.515 0.515 66.685 0.595 ;
        RECT 67.845 0.515 68.015 1.645 ;
        RECT 68.815 0.765 68.985 1.645 ;
        RECT 69.785 1.565 69.955 1.645 ;
        RECT 69.305 1.220 69.475 1.300 ;
        RECT 70.355 1.220 70.525 1.895 ;
        RECT 71.325 1.890 71.495 5.300 ;
        RECT 73.175 2.055 73.345 5.095 ;
        RECT 69.305 1.050 70.525 1.220 ;
        RECT 69.305 0.970 69.475 1.050 ;
        RECT 69.785 0.765 69.955 0.845 ;
        RECT 68.815 0.595 69.955 0.765 ;
        RECT 68.815 0.515 68.985 0.595 ;
        RECT 69.785 0.515 69.955 0.595 ;
        RECT 70.355 0.765 70.525 1.050 ;
        RECT 70.840 1.720 71.495 1.890 ;
        RECT 72.655 1.815 72.825 1.895 ;
        RECT 73.625 1.815 73.795 1.895 ;
        RECT 74.595 1.815 74.765 1.895 ;
        RECT 70.840 0.985 71.010 1.720 ;
        RECT 72.655 1.645 74.765 1.815 ;
        RECT 71.325 0.765 71.495 1.535 ;
        RECT 70.355 0.595 71.495 0.765 ;
        RECT 70.355 0.515 70.525 0.595 ;
        RECT 71.325 0.515 71.495 0.595 ;
        RECT 72.655 0.515 72.825 1.645 ;
        RECT 73.625 0.765 73.795 1.645 ;
        RECT 74.595 1.565 74.765 1.645 ;
        RECT 74.115 1.220 74.285 1.300 ;
        RECT 75.165 1.220 75.335 1.895 ;
        RECT 76.135 1.890 76.305 5.300 ;
        RECT 77.985 2.055 78.155 5.095 ;
        RECT 80.205 2.055 80.375 5.095 ;
        RECT 74.115 1.050 75.335 1.220 ;
        RECT 74.115 0.970 74.285 1.050 ;
        RECT 74.595 0.765 74.765 0.845 ;
        RECT 73.625 0.595 74.765 0.765 ;
        RECT 73.625 0.515 73.795 0.595 ;
        RECT 74.595 0.515 74.765 0.595 ;
        RECT 75.165 0.765 75.335 1.050 ;
        RECT 75.650 1.720 76.305 1.890 ;
        RECT 77.465 1.815 77.635 1.895 ;
        RECT 78.435 1.815 78.605 1.895 ;
        RECT 79.405 1.815 79.575 1.895 ;
        RECT 75.650 0.985 75.820 1.720 ;
        RECT 77.465 1.645 79.575 1.815 ;
        RECT 76.135 0.765 76.305 1.535 ;
        RECT 75.165 0.595 76.305 0.765 ;
        RECT 75.165 0.515 75.335 0.595 ;
        RECT 76.135 0.515 76.305 0.595 ;
        RECT 77.465 0.515 77.635 1.645 ;
        RECT 78.435 0.765 78.605 1.645 ;
        RECT 79.405 1.565 79.575 1.645 ;
        RECT 78.925 1.220 79.095 1.300 ;
        RECT 79.975 1.220 80.145 1.895 ;
        RECT 80.945 1.890 81.115 5.300 ;
        RECT 82.795 2.055 82.965 5.095 ;
        RECT 85.015 2.055 85.185 5.095 ;
        RECT 78.925 1.050 80.145 1.220 ;
        RECT 78.925 0.970 79.095 1.050 ;
        RECT 79.405 0.765 79.575 0.845 ;
        RECT 78.435 0.595 79.575 0.765 ;
        RECT 78.435 0.515 78.605 0.595 ;
        RECT 79.405 0.515 79.575 0.595 ;
        RECT 79.975 0.765 80.145 1.050 ;
        RECT 80.460 1.720 81.115 1.890 ;
        RECT 82.275 1.815 82.445 1.895 ;
        RECT 83.245 1.815 83.415 1.895 ;
        RECT 84.215 1.815 84.385 1.895 ;
        RECT 80.460 0.985 80.630 1.720 ;
        RECT 82.275 1.645 84.385 1.815 ;
        RECT 80.945 0.765 81.115 1.535 ;
        RECT 79.975 0.595 81.115 0.765 ;
        RECT 79.975 0.515 80.145 0.595 ;
        RECT 80.945 0.515 81.115 0.595 ;
        RECT 82.275 0.515 82.445 1.645 ;
        RECT 83.245 0.765 83.415 1.645 ;
        RECT 84.215 1.565 84.385 1.645 ;
        RECT 83.735 1.220 83.905 1.300 ;
        RECT 84.785 1.220 84.955 1.895 ;
        RECT 85.755 1.890 85.925 5.300 ;
        RECT 88.605 5.275 88.775 5.355 ;
        RECT 90.605 7.055 92.535 7.225 ;
        RECT 90.605 5.275 90.775 7.055 ;
        RECT 91.045 5.525 91.215 6.795 ;
        RECT 91.485 5.785 91.655 7.055 ;
        RECT 91.925 5.525 92.095 6.795 ;
        RECT 92.365 5.605 92.535 7.055 ;
        RECT 93.945 7.055 95.875 7.225 ;
        RECT 91.045 5.355 92.095 5.525 ;
        RECT 91.925 5.275 92.095 5.355 ;
        RECT 93.945 5.275 94.115 7.055 ;
        RECT 94.825 5.785 94.995 7.055 ;
        RECT 95.705 5.785 95.875 7.055 ;
        RECT 87.235 2.055 87.405 5.100 ;
        RECT 88.385 4.940 88.555 5.100 ;
        RECT 88.345 4.770 88.555 4.940 ;
        RECT 88.345 2.055 88.515 4.770 ;
        RECT 90.935 2.055 91.105 5.100 ;
        RECT 92.415 2.055 92.585 5.100 ;
        RECT 93.895 2.055 94.065 5.100 ;
        RECT 95.005 4.770 95.195 5.100 ;
        RECT 95.005 2.055 95.175 4.770 ;
        RECT 83.735 1.050 84.955 1.220 ;
        RECT 83.735 0.970 83.905 1.050 ;
        RECT 84.215 0.765 84.385 0.845 ;
        RECT 83.245 0.595 84.385 0.765 ;
        RECT 83.245 0.515 83.415 0.595 ;
        RECT 84.215 0.515 84.385 0.595 ;
        RECT 84.785 0.765 84.955 1.050 ;
        RECT 85.270 1.720 85.925 1.890 ;
        RECT 87.190 1.805 87.360 1.885 ;
        RECT 88.160 1.805 88.330 1.885 ;
        RECT 85.270 0.985 85.440 1.720 ;
        RECT 87.190 1.635 88.330 1.805 ;
        RECT 85.755 0.765 85.925 1.535 ;
        RECT 84.785 0.595 85.925 0.765 ;
        RECT 84.785 0.515 84.955 0.595 ;
        RECT 85.755 0.515 85.925 0.595 ;
        RECT 87.190 0.505 87.360 1.635 ;
        RECT 88.160 0.755 88.330 1.635 ;
        RECT 89.130 0.755 89.300 1.885 ;
        RECT 88.160 0.585 89.300 0.755 ;
        RECT 88.160 0.505 88.330 0.585 ;
        RECT 89.130 0.505 89.300 0.585 ;
        RECT 90.520 1.805 90.690 1.885 ;
        RECT 91.490 1.805 91.660 1.885 ;
        RECT 90.520 1.635 91.660 1.805 ;
        RECT 90.520 0.505 90.690 1.635 ;
        RECT 91.490 0.755 91.660 1.635 ;
        RECT 92.460 0.755 92.630 1.885 ;
        RECT 91.490 0.585 92.630 0.755 ;
        RECT 91.490 0.505 91.660 0.585 ;
        RECT 92.460 0.505 92.630 0.585 ;
        RECT 93.850 1.805 94.020 1.885 ;
        RECT 94.820 1.805 94.990 1.885 ;
        RECT 93.850 1.635 94.990 1.805 ;
        RECT 93.850 0.505 94.020 1.635 ;
        RECT 94.820 0.755 94.990 1.635 ;
        RECT 95.790 0.755 95.960 1.530 ;
        RECT 94.820 0.585 95.960 0.755 ;
        RECT 94.820 0.505 94.990 0.585 ;
        RECT 95.790 0.505 95.960 0.585 ;
      LAYER mcon ;
        RECT 88.605 5.355 88.775 5.525 ;
        RECT 3.245 3.615 3.415 3.785 ;
        RECT 3.985 2.880 4.155 3.050 ;
        RECT 8.050 3.985 8.220 4.155 ;
        RECT 5.835 2.880 6.005 3.050 ;
        RECT 8.795 3.615 8.965 3.785 ;
        RECT 10.645 2.880 10.815 3.050 ;
        RECT 12.865 3.985 13.035 4.155 ;
        RECT 13.605 2.875 13.775 3.045 ;
        RECT 15.455 2.875 15.625 3.045 ;
        RECT 18.415 3.985 18.585 4.155 ;
        RECT 20.265 3.615 20.435 3.785 ;
        RECT 22.485 3.245 22.655 3.415 ;
        RECT 23.225 3.615 23.395 3.785 ;
        RECT 25.075 3.615 25.245 3.785 ;
        RECT 27.295 3.985 27.465 4.155 ;
        RECT 28.035 3.245 28.205 3.415 ;
        RECT 32.105 3.615 32.275 3.785 ;
        RECT 32.845 2.880 33.015 3.050 ;
        RECT 36.910 3.985 37.080 4.155 ;
        RECT 34.695 2.880 34.865 3.050 ;
        RECT 37.655 3.615 37.825 3.785 ;
        RECT 39.505 2.880 39.675 3.050 ;
        RECT 41.725 3.985 41.895 4.155 ;
        RECT 42.465 2.875 42.635 3.045 ;
        RECT 44.315 2.875 44.485 3.045 ;
        RECT 47.275 3.985 47.445 4.155 ;
        RECT 49.125 3.615 49.295 3.785 ;
        RECT 51.345 2.875 51.515 3.045 ;
        RECT 52.085 3.615 52.255 3.785 ;
        RECT 53.935 3.615 54.105 3.785 ;
        RECT 56.155 3.985 56.325 4.155 ;
        RECT 56.895 3.985 57.065 4.155 ;
        RECT 56.895 2.875 57.065 3.045 ;
        RECT 60.965 3.615 61.135 3.785 ;
        RECT 61.705 2.880 61.875 3.050 ;
        RECT 65.770 3.985 65.940 4.155 ;
        RECT 63.555 2.880 63.725 3.050 ;
        RECT 66.515 3.615 66.685 3.785 ;
        RECT 68.365 2.880 68.535 3.050 ;
        RECT 70.585 3.985 70.755 4.155 ;
        RECT 71.325 2.875 71.495 3.045 ;
        RECT 73.175 2.875 73.345 3.045 ;
        RECT 76.135 3.985 76.305 4.155 ;
        RECT 77.985 3.615 78.155 3.785 ;
        RECT 80.205 2.875 80.375 3.045 ;
        RECT 80.945 3.615 81.115 3.785 ;
        RECT 82.795 3.615 82.965 3.785 ;
        RECT 85.015 3.985 85.185 4.155 ;
        RECT 90.605 5.355 90.775 5.525 ;
        RECT 91.925 5.355 92.095 5.525 ;
        RECT 93.945 5.355 94.115 5.525 ;
        RECT 85.755 3.985 85.925 4.155 ;
        RECT 85.755 2.875 85.925 3.045 ;
        RECT 87.235 4.725 87.405 4.895 ;
        RECT 87.235 3.985 87.405 4.155 ;
        RECT 88.345 4.355 88.515 4.525 ;
        RECT 90.935 4.725 91.105 4.895 ;
        RECT 92.415 3.245 92.585 3.415 ;
        RECT 92.415 2.135 92.585 2.305 ;
        RECT 93.895 2.135 94.065 2.305 ;
        RECT 95.005 4.355 95.175 4.525 ;
      LAYER met1 ;
        RECT 88.575 5.525 88.805 5.555 ;
        RECT 90.575 5.525 90.805 5.555 ;
        RECT 91.895 5.525 92.125 5.555 ;
        RECT 93.915 5.525 94.145 5.555 ;
        RECT 88.545 5.355 90.835 5.525 ;
        RECT 91.865 5.355 94.175 5.525 ;
        RECT 88.575 5.325 88.805 5.355 ;
        RECT 90.575 5.325 90.805 5.355 ;
        RECT 91.895 5.325 92.125 5.355 ;
        RECT 93.915 5.325 94.145 5.355 ;
        RECT 87.205 4.895 87.435 4.925 ;
        RECT 90.905 4.895 91.135 4.925 ;
        RECT 87.175 4.725 91.165 4.895 ;
        RECT 87.205 4.695 87.435 4.725 ;
        RECT 90.905 4.695 91.135 4.725 ;
        RECT 88.315 4.525 88.545 4.555 ;
        RECT 94.975 4.525 95.205 4.555 ;
        RECT 59.855 4.355 95.235 4.525 ;
        RECT 8.020 4.155 8.250 4.185 ;
        RECT 12.835 4.155 13.065 4.185 ;
        RECT 18.385 4.155 18.615 4.185 ;
        RECT 27.265 4.155 27.495 4.185 ;
        RECT 36.880 4.155 37.110 4.185 ;
        RECT 41.695 4.155 41.925 4.185 ;
        RECT 47.245 4.155 47.475 4.185 ;
        RECT 56.125 4.155 56.355 4.185 ;
        RECT 56.865 4.155 57.095 4.185 ;
        RECT 59.855 4.155 60.025 4.355 ;
        RECT 88.315 4.325 88.545 4.355 ;
        RECT 94.975 4.325 95.205 4.355 ;
        RECT 65.740 4.155 65.970 4.185 ;
        RECT 70.555 4.155 70.785 4.185 ;
        RECT 76.105 4.155 76.335 4.185 ;
        RECT 84.985 4.155 85.215 4.185 ;
        RECT 85.725 4.155 85.955 4.185 ;
        RECT 87.205 4.155 87.435 4.185 ;
        RECT 7.990 3.985 27.525 4.155 ;
        RECT 36.850 3.985 56.385 4.155 ;
        RECT 56.835 3.985 60.025 4.155 ;
        RECT 65.710 3.985 85.245 4.155 ;
        RECT 85.695 3.985 87.465 4.155 ;
        RECT 8.020 3.955 8.250 3.985 ;
        RECT 12.835 3.955 13.065 3.985 ;
        RECT 18.385 3.955 18.615 3.985 ;
        RECT 27.265 3.955 27.495 3.985 ;
        RECT 36.880 3.955 37.110 3.985 ;
        RECT 41.695 3.955 41.925 3.985 ;
        RECT 47.245 3.955 47.475 3.985 ;
        RECT 56.125 3.955 56.355 3.985 ;
        RECT 56.865 3.955 57.095 3.985 ;
        RECT 65.740 3.955 65.970 3.985 ;
        RECT 70.555 3.955 70.785 3.985 ;
        RECT 76.105 3.955 76.335 3.985 ;
        RECT 84.985 3.955 85.215 3.985 ;
        RECT 85.725 3.955 85.955 3.985 ;
        RECT 87.205 3.955 87.435 3.985 ;
        RECT 3.215 3.785 3.445 3.815 ;
        RECT 8.765 3.785 8.995 3.815 ;
        RECT 20.235 3.785 20.465 3.815 ;
        RECT 23.195 3.785 23.425 3.815 ;
        RECT 25.045 3.785 25.275 3.815 ;
        RECT 32.075 3.785 32.305 3.815 ;
        RECT 37.625 3.785 37.855 3.815 ;
        RECT 49.095 3.785 49.325 3.815 ;
        RECT 52.055 3.785 52.285 3.815 ;
        RECT 53.905 3.785 54.135 3.815 ;
        RECT 60.935 3.785 61.165 3.815 ;
        RECT 66.485 3.785 66.715 3.815 ;
        RECT 77.955 3.785 78.185 3.815 ;
        RECT 80.915 3.785 81.145 3.815 ;
        RECT 82.765 3.785 82.995 3.815 ;
        RECT 3.185 3.615 20.495 3.785 ;
        RECT 23.165 3.615 25.305 3.785 ;
        RECT 32.045 3.615 49.355 3.785 ;
        RECT 52.025 3.615 54.165 3.785 ;
        RECT 60.905 3.615 78.215 3.785 ;
        RECT 80.885 3.615 83.025 3.785 ;
        RECT 3.215 3.585 3.445 3.615 ;
        RECT 8.765 3.585 8.995 3.615 ;
        RECT 20.235 3.585 20.465 3.615 ;
        RECT 23.195 3.585 23.425 3.615 ;
        RECT 25.045 3.585 25.275 3.615 ;
        RECT 32.075 3.585 32.305 3.615 ;
        RECT 37.625 3.585 37.855 3.615 ;
        RECT 49.095 3.585 49.325 3.615 ;
        RECT 52.055 3.585 52.285 3.615 ;
        RECT 53.905 3.585 54.135 3.615 ;
        RECT 60.935 3.585 61.165 3.615 ;
        RECT 66.485 3.585 66.715 3.615 ;
        RECT 77.955 3.585 78.185 3.615 ;
        RECT 80.915 3.585 81.145 3.615 ;
        RECT 82.765 3.585 82.995 3.615 ;
        RECT 22.455 3.415 22.685 3.445 ;
        RECT 28.005 3.415 28.235 3.445 ;
        RECT 92.385 3.415 92.615 3.445 ;
        RECT 22.425 3.245 92.645 3.415 ;
        RECT 22.455 3.215 22.685 3.245 ;
        RECT 28.005 3.215 28.235 3.245 ;
        RECT 92.385 3.215 92.615 3.245 ;
        RECT 3.955 3.050 4.185 3.080 ;
        RECT 5.805 3.050 6.035 3.080 ;
        RECT 10.615 3.050 10.845 3.080 ;
        RECT 3.925 2.880 10.875 3.050 ;
        RECT 13.575 3.045 13.805 3.075 ;
        RECT 15.425 3.045 15.655 3.075 ;
        RECT 32.815 3.050 33.045 3.080 ;
        RECT 34.665 3.050 34.895 3.080 ;
        RECT 39.475 3.050 39.705 3.080 ;
        RECT 3.955 2.850 4.185 2.880 ;
        RECT 5.805 2.850 6.035 2.880 ;
        RECT 10.615 2.850 10.845 2.880 ;
        RECT 13.545 2.875 15.685 3.045 ;
        RECT 32.785 2.880 39.735 3.050 ;
        RECT 42.435 3.045 42.665 3.075 ;
        RECT 44.285 3.045 44.515 3.075 ;
        RECT 51.315 3.045 51.545 3.075 ;
        RECT 56.865 3.045 57.095 3.075 ;
        RECT 61.675 3.050 61.905 3.080 ;
        RECT 63.525 3.050 63.755 3.080 ;
        RECT 68.335 3.050 68.565 3.080 ;
        RECT 13.575 2.845 13.805 2.875 ;
        RECT 15.425 2.845 15.655 2.875 ;
        RECT 32.815 2.850 33.045 2.880 ;
        RECT 34.665 2.850 34.895 2.880 ;
        RECT 39.475 2.850 39.705 2.880 ;
        RECT 42.405 2.875 44.545 3.045 ;
        RECT 51.285 2.875 57.125 3.045 ;
        RECT 61.645 2.880 68.595 3.050 ;
        RECT 71.295 3.045 71.525 3.075 ;
        RECT 73.145 3.045 73.375 3.075 ;
        RECT 80.175 3.045 80.405 3.075 ;
        RECT 85.725 3.045 85.955 3.075 ;
        RECT 42.435 2.845 42.665 2.875 ;
        RECT 44.285 2.845 44.515 2.875 ;
        RECT 51.315 2.845 51.545 2.875 ;
        RECT 56.865 2.845 57.095 2.875 ;
        RECT 61.675 2.850 61.905 2.880 ;
        RECT 63.525 2.850 63.755 2.880 ;
        RECT 68.335 2.850 68.565 2.880 ;
        RECT 71.265 2.875 73.405 3.045 ;
        RECT 80.145 2.875 85.985 3.045 ;
        RECT 71.295 2.845 71.525 2.875 ;
        RECT 73.145 2.845 73.375 2.875 ;
        RECT 80.175 2.845 80.405 2.875 ;
        RECT 85.725 2.845 85.955 2.875 ;
        RECT 92.385 2.305 92.615 2.335 ;
        RECT 93.865 2.305 94.095 2.335 ;
        RECT 92.355 2.135 94.125 2.305 ;
        RECT 92.385 2.105 92.615 2.135 ;
        RECT 93.865 2.105 94.095 2.135 ;
  END
END TMRDFFSNRNQNX1






MACRO TMRDFFSNRNQX1
  CLASS BLOCK ;
  FOREIGN TMRDFFSNRNQX1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 99.630 BY 7.950 ;
  PIN Q
    ANTENNADIFFAREA 0.771900 ;
    PORT
      LAYER li1 ;
        RECT 97.595 4.895 97.765 7.250 ;
        RECT 97.595 4.725 98.135 4.895 ;
        RECT 97.965 2.305 98.135 4.725 ;
        RECT 97.595 2.135 98.135 2.305 ;
        RECT 97.595 0.975 97.765 2.135 ;
      LAYER mcon ;
        RECT 97.965 3.985 98.135 4.155 ;
      LAYER met1 ;
        RECT 97.935 4.155 98.165 4.185 ;
        RECT 97.905 3.985 98.315 4.155 ;
        RECT 97.935 3.955 98.165 3.985 ;
    END
  END Q
  PIN D
    ANTENNAGATEAREA 3.099750 ;
    PORT
      LAYER li1 ;
        RECT 1.025 2.055 1.195 5.095 ;
        RECT 29.885 2.055 30.055 5.095 ;
        RECT 58.745 2.055 58.915 5.095 ;
      LAYER mcon ;
        RECT 1.025 4.355 1.195 4.525 ;
        RECT 29.885 4.355 30.055 4.525 ;
        RECT 58.745 4.355 58.915 4.525 ;
      LAYER met1 ;
        RECT 0.995 4.525 1.225 4.555 ;
        RECT 29.855 4.525 30.085 4.555 ;
        RECT 58.715 4.525 58.945 4.555 ;
        RECT 0.845 4.355 59.095 4.525 ;
        RECT 0.995 4.325 1.225 4.355 ;
        RECT 29.855 4.325 30.085 4.355 ;
        RECT 58.715 4.325 58.945 4.355 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 6.089100 ;
    PORT
      LAYER li1 ;
        RECT 6.945 4.975 7.115 5.095 ;
        RECT 6.940 4.645 7.115 4.975 ;
        RECT 6.945 2.055 7.115 4.645 ;
        RECT 16.565 2.055 16.735 5.095 ;
        RECT 35.805 4.975 35.975 5.095 ;
        RECT 35.800 4.645 35.975 4.975 ;
        RECT 35.805 2.055 35.975 4.645 ;
        RECT 45.425 2.055 45.595 5.095 ;
        RECT 64.665 4.975 64.835 5.095 ;
        RECT 64.660 4.645 64.835 4.975 ;
        RECT 64.665 2.055 64.835 4.645 ;
        RECT 74.285 2.055 74.455 5.095 ;
      LAYER mcon ;
        RECT 6.940 4.725 7.110 4.895 ;
        RECT 16.565 4.725 16.735 4.895 ;
        RECT 35.800 4.725 35.970 4.895 ;
        RECT 45.425 4.725 45.595 4.895 ;
        RECT 64.660 4.725 64.830 4.895 ;
        RECT 74.285 4.725 74.455 4.895 ;
      LAYER met1 ;
        RECT 6.910 4.895 7.140 4.925 ;
        RECT 16.535 4.895 16.765 4.925 ;
        RECT 35.770 4.895 36.000 4.925 ;
        RECT 45.395 4.895 45.625 4.925 ;
        RECT 64.630 4.895 64.860 4.925 ;
        RECT 74.255 4.895 74.485 4.925 ;
        RECT 6.880 4.725 74.515 4.895 ;
        RECT 6.910 4.695 7.140 4.725 ;
        RECT 16.535 4.695 16.765 4.725 ;
        RECT 35.770 4.695 36.000 4.725 ;
        RECT 45.395 4.695 45.625 4.725 ;
        RECT 64.630 4.695 64.860 4.725 ;
        RECT 74.255 4.695 74.485 4.725 ;
    END
  END CLK
  PIN SN
    ANTENNAGATEAREA 6.089100 ;
    PORT
      LAYER li1 ;
        RECT 11.755 2.055 11.925 5.095 ;
        RECT 26.185 2.055 26.355 5.095 ;
        RECT 40.615 2.055 40.785 5.095 ;
        RECT 55.045 2.055 55.215 5.095 ;
        RECT 69.475 2.055 69.645 5.095 ;
        RECT 83.905 2.055 84.075 5.095 ;
      LAYER mcon ;
        RECT 11.755 2.140 11.925 2.310 ;
        RECT 26.185 2.135 26.355 2.305 ;
        RECT 40.615 2.140 40.785 2.310 ;
        RECT 55.045 2.135 55.215 2.305 ;
        RECT 69.475 2.140 69.645 2.310 ;
        RECT 83.905 2.135 84.075 2.305 ;
      LAYER met1 ;
        RECT 11.725 2.310 11.955 2.340 ;
        RECT 11.695 2.305 12.105 2.310 ;
        RECT 26.155 2.305 26.385 2.335 ;
        RECT 40.585 2.310 40.815 2.340 ;
        RECT 40.555 2.305 40.965 2.310 ;
        RECT 55.015 2.305 55.245 2.335 ;
        RECT 69.445 2.310 69.675 2.340 ;
        RECT 69.415 2.305 69.825 2.310 ;
        RECT 83.875 2.305 84.105 2.335 ;
        RECT 11.695 2.140 84.135 2.305 ;
        RECT 11.720 2.135 84.135 2.140 ;
        RECT 11.725 2.110 11.955 2.135 ;
        RECT 26.155 2.105 26.385 2.135 ;
        RECT 40.585 2.110 40.815 2.135 ;
        RECT 55.015 2.105 55.245 2.135 ;
        RECT 69.445 2.110 69.675 2.135 ;
        RECT 83.875 2.105 84.105 2.135 ;
    END
  END SN
  PIN RN
    ANTENNAGATEAREA 9.170850 ;
    PORT
      LAYER li1 ;
        RECT 2.135 2.055 2.305 5.095 ;
        RECT 17.675 2.055 17.845 5.095 ;
        RECT 21.375 2.055 21.545 5.095 ;
        RECT 30.995 2.055 31.165 5.095 ;
        RECT 46.535 2.055 46.705 5.095 ;
        RECT 50.235 2.055 50.405 5.095 ;
        RECT 59.855 2.055 60.025 5.095 ;
        RECT 75.395 2.055 75.565 5.095 ;
        RECT 79.095 2.055 79.265 5.095 ;
      LAYER mcon ;
        RECT 2.135 2.505 2.305 2.675 ;
        RECT 17.675 2.505 17.845 2.675 ;
        RECT 21.375 2.505 21.545 2.675 ;
        RECT 30.995 2.505 31.165 2.675 ;
        RECT 46.535 2.505 46.705 2.675 ;
        RECT 50.235 2.505 50.405 2.675 ;
        RECT 59.855 2.505 60.025 2.675 ;
        RECT 75.395 2.505 75.565 2.675 ;
        RECT 79.095 2.505 79.265 2.675 ;
      LAYER met1 ;
        RECT 2.105 2.675 2.335 2.705 ;
        RECT 17.645 2.675 17.875 2.705 ;
        RECT 21.345 2.675 21.575 2.705 ;
        RECT 30.965 2.675 31.195 2.705 ;
        RECT 46.505 2.675 46.735 2.705 ;
        RECT 50.205 2.675 50.435 2.705 ;
        RECT 59.825 2.675 60.055 2.705 ;
        RECT 75.365 2.675 75.595 2.705 ;
        RECT 79.065 2.675 79.295 2.705 ;
        RECT 2.075 2.505 79.325 2.675 ;
        RECT 2.105 2.475 2.335 2.505 ;
        RECT 17.645 2.475 17.875 2.505 ;
        RECT 21.345 2.475 21.575 2.505 ;
        RECT 30.965 2.475 31.195 2.505 ;
        RECT 46.505 2.475 46.735 2.505 ;
        RECT 50.205 2.475 50.435 2.505 ;
        RECT 59.825 2.475 60.055 2.505 ;
        RECT 75.365 2.475 75.595 2.505 ;
        RECT 79.065 2.475 79.295 2.505 ;
    END
  END RN
  PIN VDD
    ANTENNADIFFAREA 111.526749 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 99.210 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 98.945 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 1.005 5.445 1.175 7.460 ;
        RECT 1.885 5.785 2.055 7.460 ;
        RECT 2.765 5.785 2.935 7.460 ;
        RECT 3.645 5.785 3.815 7.460 ;
        RECT 4.655 4.340 4.965 7.460 ;
        RECT 5.815 5.445 5.985 7.460 ;
        RECT 6.695 5.785 6.865 7.460 ;
        RECT 7.575 5.785 7.745 7.460 ;
        RECT 8.455 5.785 8.625 7.460 ;
        RECT 9.465 4.340 9.775 7.460 ;
        RECT 10.625 5.445 10.795 7.460 ;
        RECT 11.505 5.785 11.675 7.460 ;
        RECT 12.385 5.785 12.555 7.460 ;
        RECT 13.265 5.785 13.435 7.460 ;
        RECT 14.275 4.340 14.585 7.460 ;
        RECT 15.435 5.445 15.605 7.460 ;
        RECT 16.315 5.785 16.485 7.460 ;
        RECT 17.195 5.785 17.365 7.460 ;
        RECT 18.075 5.785 18.245 7.460 ;
        RECT 19.085 4.340 19.395 7.460 ;
        RECT 20.245 5.445 20.415 7.460 ;
        RECT 21.125 5.785 21.295 7.460 ;
        RECT 22.005 5.785 22.175 7.460 ;
        RECT 22.885 5.785 23.055 7.460 ;
        RECT 23.895 4.340 24.205 7.460 ;
        RECT 25.055 5.445 25.225 7.460 ;
        RECT 25.935 5.785 26.105 7.460 ;
        RECT 26.815 5.785 26.985 7.460 ;
        RECT 27.695 5.785 27.865 7.460 ;
        RECT 28.705 4.340 29.015 7.460 ;
        RECT 29.865 5.445 30.035 7.460 ;
        RECT 30.745 5.785 30.915 7.460 ;
        RECT 31.625 5.785 31.795 7.460 ;
        RECT 32.505 5.785 32.675 7.460 ;
        RECT 33.515 4.340 33.825 7.460 ;
        RECT 34.675 5.445 34.845 7.460 ;
        RECT 35.555 5.785 35.725 7.460 ;
        RECT 36.435 5.785 36.605 7.460 ;
        RECT 37.315 5.785 37.485 7.460 ;
        RECT 38.325 4.340 38.635 7.460 ;
        RECT 39.485 5.445 39.655 7.460 ;
        RECT 40.365 5.785 40.535 7.460 ;
        RECT 41.245 5.785 41.415 7.460 ;
        RECT 42.125 5.785 42.295 7.460 ;
        RECT 43.135 4.340 43.445 7.460 ;
        RECT 44.295 5.445 44.465 7.460 ;
        RECT 45.175 5.785 45.345 7.460 ;
        RECT 46.055 5.785 46.225 7.460 ;
        RECT 46.935 5.785 47.105 7.460 ;
        RECT 47.945 4.340 48.255 7.460 ;
        RECT 49.105 5.445 49.275 7.460 ;
        RECT 49.985 5.785 50.155 7.460 ;
        RECT 50.865 5.785 51.035 7.460 ;
        RECT 51.745 5.785 51.915 7.460 ;
        RECT 52.755 4.340 53.065 7.460 ;
        RECT 53.915 5.445 54.085 7.460 ;
        RECT 54.795 5.785 54.965 7.460 ;
        RECT 55.675 5.785 55.845 7.460 ;
        RECT 56.555 5.785 56.725 7.460 ;
        RECT 57.565 4.340 57.875 7.460 ;
        RECT 58.725 5.445 58.895 7.460 ;
        RECT 59.605 5.785 59.775 7.460 ;
        RECT 60.485 5.785 60.655 7.460 ;
        RECT 61.365 5.785 61.535 7.460 ;
        RECT 62.375 4.340 62.685 7.460 ;
        RECT 63.535 5.445 63.705 7.460 ;
        RECT 64.415 5.785 64.585 7.460 ;
        RECT 65.295 5.785 65.465 7.460 ;
        RECT 66.175 5.785 66.345 7.460 ;
        RECT 67.185 4.340 67.495 7.460 ;
        RECT 68.345 5.445 68.515 7.460 ;
        RECT 69.225 5.785 69.395 7.460 ;
        RECT 70.105 5.785 70.275 7.460 ;
        RECT 70.985 5.785 71.155 7.460 ;
        RECT 71.995 4.340 72.305 7.460 ;
        RECT 73.155 5.445 73.325 7.460 ;
        RECT 74.035 5.785 74.205 7.460 ;
        RECT 74.915 5.785 75.085 7.460 ;
        RECT 75.795 5.785 75.965 7.460 ;
        RECT 76.805 4.340 77.115 7.460 ;
        RECT 77.965 5.445 78.135 7.460 ;
        RECT 78.845 5.785 79.015 7.460 ;
        RECT 79.725 5.785 79.895 7.460 ;
        RECT 80.605 5.785 80.775 7.460 ;
        RECT 81.615 4.340 81.925 7.460 ;
        RECT 82.775 5.445 82.945 7.460 ;
        RECT 83.655 5.785 83.825 7.460 ;
        RECT 84.535 5.785 84.705 7.460 ;
        RECT 85.415 5.785 85.585 7.460 ;
        RECT 86.425 4.340 86.735 7.460 ;
        RECT 87.285 5.355 87.455 7.460 ;
        RECT 88.165 5.785 88.335 7.460 ;
        RECT 89.045 5.355 89.215 7.460 ;
        RECT 89.755 4.340 90.065 7.460 ;
        RECT 93.085 4.340 93.395 7.460 ;
        RECT 96.415 4.340 96.725 7.460 ;
        RECT 97.155 5.415 97.325 7.460 ;
        RECT 98.035 5.415 98.205 7.460 ;
        RECT 98.635 4.340 98.945 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 0.995 7.525 1.165 7.695 ;
        RECT 1.355 7.525 1.525 7.695 ;
        RECT 1.715 7.525 1.885 7.695 ;
        RECT 2.075 7.525 2.245 7.695 ;
        RECT 2.565 7.525 2.735 7.695 ;
        RECT 2.925 7.525 3.095 7.695 ;
        RECT 3.285 7.525 3.455 7.695 ;
        RECT 3.645 7.525 3.815 7.695 ;
        RECT 4.005 7.525 4.175 7.695 ;
        RECT 4.365 7.525 4.535 7.695 ;
        RECT 5.085 7.525 5.255 7.695 ;
        RECT 5.445 7.525 5.615 7.695 ;
        RECT 5.805 7.525 5.975 7.695 ;
        RECT 6.165 7.525 6.335 7.695 ;
        RECT 6.525 7.525 6.695 7.695 ;
        RECT 6.885 7.525 7.055 7.695 ;
        RECT 7.375 7.525 7.545 7.695 ;
        RECT 7.735 7.525 7.905 7.695 ;
        RECT 8.095 7.525 8.265 7.695 ;
        RECT 8.455 7.525 8.625 7.695 ;
        RECT 8.815 7.525 8.985 7.695 ;
        RECT 9.175 7.525 9.345 7.695 ;
        RECT 9.895 7.525 10.065 7.695 ;
        RECT 10.255 7.525 10.425 7.695 ;
        RECT 10.615 7.525 10.785 7.695 ;
        RECT 10.975 7.525 11.145 7.695 ;
        RECT 11.335 7.525 11.505 7.695 ;
        RECT 11.695 7.525 11.865 7.695 ;
        RECT 12.185 7.525 12.355 7.695 ;
        RECT 12.545 7.525 12.715 7.695 ;
        RECT 12.905 7.525 13.075 7.695 ;
        RECT 13.265 7.525 13.435 7.695 ;
        RECT 13.625 7.525 13.795 7.695 ;
        RECT 13.985 7.525 14.155 7.695 ;
        RECT 14.705 7.525 14.875 7.695 ;
        RECT 15.065 7.525 15.235 7.695 ;
        RECT 15.425 7.525 15.595 7.695 ;
        RECT 15.785 7.525 15.955 7.695 ;
        RECT 16.145 7.525 16.315 7.695 ;
        RECT 16.505 7.525 16.675 7.695 ;
        RECT 16.995 7.525 17.165 7.695 ;
        RECT 17.355 7.525 17.525 7.695 ;
        RECT 17.715 7.525 17.885 7.695 ;
        RECT 18.075 7.525 18.245 7.695 ;
        RECT 18.435 7.525 18.605 7.695 ;
        RECT 18.795 7.525 18.965 7.695 ;
        RECT 19.515 7.525 19.685 7.695 ;
        RECT 19.875 7.525 20.045 7.695 ;
        RECT 20.235 7.525 20.405 7.695 ;
        RECT 20.595 7.525 20.765 7.695 ;
        RECT 20.955 7.525 21.125 7.695 ;
        RECT 21.315 7.525 21.485 7.695 ;
        RECT 21.805 7.525 21.975 7.695 ;
        RECT 22.165 7.525 22.335 7.695 ;
        RECT 22.525 7.525 22.695 7.695 ;
        RECT 22.885 7.525 23.055 7.695 ;
        RECT 23.245 7.525 23.415 7.695 ;
        RECT 23.605 7.525 23.775 7.695 ;
        RECT 24.325 7.525 24.495 7.695 ;
        RECT 24.685 7.525 24.855 7.695 ;
        RECT 25.045 7.525 25.215 7.695 ;
        RECT 25.405 7.525 25.575 7.695 ;
        RECT 25.765 7.525 25.935 7.695 ;
        RECT 26.125 7.525 26.295 7.695 ;
        RECT 26.615 7.525 26.785 7.695 ;
        RECT 26.975 7.525 27.145 7.695 ;
        RECT 27.335 7.525 27.505 7.695 ;
        RECT 27.695 7.525 27.865 7.695 ;
        RECT 28.055 7.525 28.225 7.695 ;
        RECT 28.415 7.525 28.585 7.695 ;
        RECT 29.135 7.525 29.305 7.695 ;
        RECT 29.495 7.525 29.665 7.695 ;
        RECT 29.855 7.525 30.025 7.695 ;
        RECT 30.215 7.525 30.385 7.695 ;
        RECT 30.575 7.525 30.745 7.695 ;
        RECT 30.935 7.525 31.105 7.695 ;
        RECT 31.425 7.525 31.595 7.695 ;
        RECT 31.785 7.525 31.955 7.695 ;
        RECT 32.145 7.525 32.315 7.695 ;
        RECT 32.505 7.525 32.675 7.695 ;
        RECT 32.865 7.525 33.035 7.695 ;
        RECT 33.225 7.525 33.395 7.695 ;
        RECT 33.945 7.525 34.115 7.695 ;
        RECT 34.305 7.525 34.475 7.695 ;
        RECT 34.665 7.525 34.835 7.695 ;
        RECT 35.025 7.525 35.195 7.695 ;
        RECT 35.385 7.525 35.555 7.695 ;
        RECT 35.745 7.525 35.915 7.695 ;
        RECT 36.235 7.525 36.405 7.695 ;
        RECT 36.595 7.525 36.765 7.695 ;
        RECT 36.955 7.525 37.125 7.695 ;
        RECT 37.315 7.525 37.485 7.695 ;
        RECT 37.675 7.525 37.845 7.695 ;
        RECT 38.035 7.525 38.205 7.695 ;
        RECT 38.755 7.525 38.925 7.695 ;
        RECT 39.115 7.525 39.285 7.695 ;
        RECT 39.475 7.525 39.645 7.695 ;
        RECT 39.835 7.525 40.005 7.695 ;
        RECT 40.195 7.525 40.365 7.695 ;
        RECT 40.555 7.525 40.725 7.695 ;
        RECT 41.045 7.525 41.215 7.695 ;
        RECT 41.405 7.525 41.575 7.695 ;
        RECT 41.765 7.525 41.935 7.695 ;
        RECT 42.125 7.525 42.295 7.695 ;
        RECT 42.485 7.525 42.655 7.695 ;
        RECT 42.845 7.525 43.015 7.695 ;
        RECT 43.565 7.525 43.735 7.695 ;
        RECT 43.925 7.525 44.095 7.695 ;
        RECT 44.285 7.525 44.455 7.695 ;
        RECT 44.645 7.525 44.815 7.695 ;
        RECT 45.005 7.525 45.175 7.695 ;
        RECT 45.365 7.525 45.535 7.695 ;
        RECT 45.855 7.525 46.025 7.695 ;
        RECT 46.215 7.525 46.385 7.695 ;
        RECT 46.575 7.525 46.745 7.695 ;
        RECT 46.935 7.525 47.105 7.695 ;
        RECT 47.295 7.525 47.465 7.695 ;
        RECT 47.655 7.525 47.825 7.695 ;
        RECT 48.375 7.525 48.545 7.695 ;
        RECT 48.735 7.525 48.905 7.695 ;
        RECT 49.095 7.525 49.265 7.695 ;
        RECT 49.455 7.525 49.625 7.695 ;
        RECT 49.815 7.525 49.985 7.695 ;
        RECT 50.175 7.525 50.345 7.695 ;
        RECT 50.665 7.525 50.835 7.695 ;
        RECT 51.025 7.525 51.195 7.695 ;
        RECT 51.385 7.525 51.555 7.695 ;
        RECT 51.745 7.525 51.915 7.695 ;
        RECT 52.105 7.525 52.275 7.695 ;
        RECT 52.465 7.525 52.635 7.695 ;
        RECT 53.185 7.525 53.355 7.695 ;
        RECT 53.545 7.525 53.715 7.695 ;
        RECT 53.905 7.525 54.075 7.695 ;
        RECT 54.265 7.525 54.435 7.695 ;
        RECT 54.625 7.525 54.795 7.695 ;
        RECT 54.985 7.525 55.155 7.695 ;
        RECT 55.475 7.525 55.645 7.695 ;
        RECT 55.835 7.525 56.005 7.695 ;
        RECT 56.195 7.525 56.365 7.695 ;
        RECT 56.555 7.525 56.725 7.695 ;
        RECT 56.915 7.525 57.085 7.695 ;
        RECT 57.275 7.525 57.445 7.695 ;
        RECT 57.995 7.525 58.165 7.695 ;
        RECT 58.355 7.525 58.525 7.695 ;
        RECT 58.715 7.525 58.885 7.695 ;
        RECT 59.075 7.525 59.245 7.695 ;
        RECT 59.435 7.525 59.605 7.695 ;
        RECT 59.795 7.525 59.965 7.695 ;
        RECT 60.285 7.525 60.455 7.695 ;
        RECT 60.645 7.525 60.815 7.695 ;
        RECT 61.005 7.525 61.175 7.695 ;
        RECT 61.365 7.525 61.535 7.695 ;
        RECT 61.725 7.525 61.895 7.695 ;
        RECT 62.085 7.525 62.255 7.695 ;
        RECT 62.805 7.525 62.975 7.695 ;
        RECT 63.165 7.525 63.335 7.695 ;
        RECT 63.525 7.525 63.695 7.695 ;
        RECT 63.885 7.525 64.055 7.695 ;
        RECT 64.245 7.525 64.415 7.695 ;
        RECT 64.605 7.525 64.775 7.695 ;
        RECT 65.095 7.525 65.265 7.695 ;
        RECT 65.455 7.525 65.625 7.695 ;
        RECT 65.815 7.525 65.985 7.695 ;
        RECT 66.175 7.525 66.345 7.695 ;
        RECT 66.535 7.525 66.705 7.695 ;
        RECT 66.895 7.525 67.065 7.695 ;
        RECT 67.615 7.525 67.785 7.695 ;
        RECT 67.975 7.525 68.145 7.695 ;
        RECT 68.335 7.525 68.505 7.695 ;
        RECT 68.695 7.525 68.865 7.695 ;
        RECT 69.055 7.525 69.225 7.695 ;
        RECT 69.415 7.525 69.585 7.695 ;
        RECT 69.905 7.525 70.075 7.695 ;
        RECT 70.265 7.525 70.435 7.695 ;
        RECT 70.625 7.525 70.795 7.695 ;
        RECT 70.985 7.525 71.155 7.695 ;
        RECT 71.345 7.525 71.515 7.695 ;
        RECT 71.705 7.525 71.875 7.695 ;
        RECT 72.425 7.525 72.595 7.695 ;
        RECT 72.785 7.525 72.955 7.695 ;
        RECT 73.145 7.525 73.315 7.695 ;
        RECT 73.505 7.525 73.675 7.695 ;
        RECT 73.865 7.525 74.035 7.695 ;
        RECT 74.225 7.525 74.395 7.695 ;
        RECT 74.715 7.525 74.885 7.695 ;
        RECT 75.075 7.525 75.245 7.695 ;
        RECT 75.435 7.525 75.605 7.695 ;
        RECT 75.795 7.525 75.965 7.695 ;
        RECT 76.155 7.525 76.325 7.695 ;
        RECT 76.515 7.525 76.685 7.695 ;
        RECT 77.235 7.525 77.405 7.695 ;
        RECT 77.595 7.525 77.765 7.695 ;
        RECT 77.955 7.525 78.125 7.695 ;
        RECT 78.315 7.525 78.485 7.695 ;
        RECT 78.675 7.525 78.845 7.695 ;
        RECT 79.035 7.525 79.205 7.695 ;
        RECT 79.525 7.525 79.695 7.695 ;
        RECT 79.885 7.525 80.055 7.695 ;
        RECT 80.245 7.525 80.415 7.695 ;
        RECT 80.605 7.525 80.775 7.695 ;
        RECT 80.965 7.525 81.135 7.695 ;
        RECT 81.325 7.525 81.495 7.695 ;
        RECT 82.045 7.525 82.215 7.695 ;
        RECT 82.405 7.525 82.575 7.695 ;
        RECT 82.765 7.525 82.935 7.695 ;
        RECT 83.125 7.525 83.295 7.695 ;
        RECT 83.485 7.525 83.655 7.695 ;
        RECT 83.845 7.525 84.015 7.695 ;
        RECT 84.335 7.525 84.505 7.695 ;
        RECT 84.695 7.525 84.865 7.695 ;
        RECT 85.055 7.525 85.225 7.695 ;
        RECT 85.415 7.525 85.585 7.695 ;
        RECT 85.775 7.525 85.945 7.695 ;
        RECT 86.135 7.525 86.305 7.695 ;
        RECT 86.855 7.525 87.025 7.695 ;
        RECT 87.215 7.525 87.385 7.695 ;
        RECT 87.575 7.525 87.745 7.695 ;
        RECT 87.935 7.525 88.105 7.695 ;
        RECT 88.385 7.525 88.555 7.695 ;
        RECT 88.745 7.525 88.915 7.695 ;
        RECT 89.105 7.525 89.275 7.695 ;
        RECT 89.465 7.525 89.635 7.695 ;
        RECT 90.185 7.525 90.355 7.695 ;
        RECT 90.545 7.525 90.715 7.695 ;
        RECT 90.905 7.525 91.075 7.695 ;
        RECT 91.265 7.525 91.435 7.695 ;
        RECT 91.715 7.525 91.885 7.695 ;
        RECT 92.075 7.525 92.245 7.695 ;
        RECT 92.435 7.525 92.605 7.695 ;
        RECT 92.795 7.525 92.965 7.695 ;
        RECT 93.515 7.525 93.685 7.695 ;
        RECT 93.875 7.525 94.045 7.695 ;
        RECT 94.235 7.525 94.405 7.695 ;
        RECT 94.595 7.525 94.765 7.695 ;
        RECT 95.045 7.525 95.215 7.695 ;
        RECT 95.405 7.525 95.575 7.695 ;
        RECT 95.765 7.525 95.935 7.695 ;
        RECT 96.125 7.525 96.295 7.695 ;
        RECT 96.845 7.525 97.015 7.695 ;
        RECT 97.205 7.525 97.375 7.695 ;
        RECT 97.595 7.525 97.765 7.695 ;
        RECT 97.985 7.525 98.155 7.695 ;
        RECT 98.345 7.525 98.515 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 98.945 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 69.352898 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 99.075 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 4.525 -0.075 5.095 -0.065 ;
        RECT 9.335 -0.075 9.905 -0.065 ;
        RECT 14.145 -0.075 14.715 -0.065 ;
        RECT 18.955 -0.075 19.525 -0.065 ;
        RECT 23.765 -0.075 24.335 -0.065 ;
        RECT 28.575 -0.075 29.145 -0.065 ;
        RECT 33.385 -0.075 33.955 -0.065 ;
        RECT 38.195 -0.075 38.765 -0.065 ;
        RECT 43.005 -0.075 43.575 -0.065 ;
        RECT 47.815 -0.075 48.385 -0.065 ;
        RECT 52.625 -0.075 53.195 -0.065 ;
        RECT 57.435 -0.075 58.005 -0.065 ;
        RECT 62.245 -0.075 62.815 -0.065 ;
        RECT 67.055 -0.075 67.625 -0.065 ;
        RECT 71.865 -0.075 72.435 -0.065 ;
        RECT 76.675 -0.075 77.245 -0.065 ;
        RECT 81.485 -0.075 82.055 -0.065 ;
        RECT 86.295 -0.075 86.865 -0.065 ;
        RECT 89.625 -0.075 90.195 -0.065 ;
        RECT 92.955 -0.075 93.525 -0.065 ;
        RECT 96.285 -0.075 96.855 -0.065 ;
        RECT 98.505 -0.075 99.075 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 0.990 0.310 1.160 1.270 ;
        RECT 4.655 0.310 4.965 2.860 ;
        RECT 5.800 0.310 5.970 1.270 ;
        RECT 9.465 0.310 9.775 2.860 ;
        RECT 10.610 0.310 10.780 1.270 ;
        RECT 14.275 0.310 14.585 2.860 ;
        RECT 15.420 0.310 15.590 1.270 ;
        RECT 19.085 0.310 19.395 2.860 ;
        RECT 20.230 0.310 20.400 1.270 ;
        RECT 23.895 0.310 24.205 2.860 ;
        RECT 25.040 0.310 25.210 1.270 ;
        RECT 28.705 0.310 29.015 2.860 ;
        RECT 29.850 0.310 30.020 1.270 ;
        RECT 33.515 0.310 33.825 2.860 ;
        RECT 34.660 0.310 34.830 1.270 ;
        RECT 38.325 0.310 38.635 2.860 ;
        RECT 39.470 0.310 39.640 1.270 ;
        RECT 43.135 0.310 43.445 2.860 ;
        RECT 44.280 0.310 44.450 1.270 ;
        RECT 47.945 0.310 48.255 2.860 ;
        RECT 49.090 0.310 49.260 1.270 ;
        RECT 52.755 0.310 53.065 2.860 ;
        RECT 53.900 0.310 54.070 1.270 ;
        RECT 57.565 0.310 57.875 2.860 ;
        RECT 58.710 0.310 58.880 1.270 ;
        RECT 62.375 0.310 62.685 2.860 ;
        RECT 63.520 0.310 63.690 1.270 ;
        RECT 67.185 0.310 67.495 2.860 ;
        RECT 68.330 0.310 68.500 1.270 ;
        RECT 71.995 0.310 72.305 2.860 ;
        RECT 73.140 0.310 73.310 1.270 ;
        RECT 76.805 0.310 77.115 2.860 ;
        RECT 77.950 0.310 78.120 1.270 ;
        RECT 81.615 0.310 81.925 2.860 ;
        RECT 82.760 0.310 82.930 1.270 ;
        RECT 86.425 0.310 86.735 2.860 ;
        RECT 87.675 0.310 87.845 1.260 ;
        RECT 89.755 0.310 90.065 2.860 ;
        RECT 91.005 0.310 91.175 1.260 ;
        RECT 93.085 0.310 93.395 2.860 ;
        RECT 94.335 0.310 94.505 1.260 ;
        RECT 96.415 0.310 96.725 2.860 ;
        RECT 97.115 0.755 97.285 1.885 ;
        RECT 98.085 0.755 98.255 1.885 ;
        RECT 97.115 0.585 98.255 0.755 ;
        RECT 97.115 0.310 97.285 0.585 ;
        RECT 97.600 0.310 97.770 0.585 ;
        RECT 98.085 0.310 98.255 0.585 ;
        RECT 98.635 0.310 98.945 2.860 ;
        RECT -0.155 0.235 91.975 0.310 ;
        RECT 92.145 0.235 98.945 0.310 ;
        RECT -0.155 0.000 98.945 0.235 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 0.995 0.065 1.165 0.235 ;
        RECT 1.355 0.065 1.525 0.235 ;
        RECT 1.715 0.065 1.885 0.235 ;
        RECT 2.075 0.065 2.245 0.235 ;
        RECT 2.565 0.065 2.735 0.235 ;
        RECT 2.925 0.065 3.095 0.235 ;
        RECT 3.285 0.065 3.455 0.235 ;
        RECT 3.645 0.065 3.815 0.235 ;
        RECT 4.005 0.065 4.175 0.235 ;
        RECT 4.365 0.065 4.535 0.235 ;
        RECT 5.085 0.065 5.255 0.235 ;
        RECT 5.445 0.065 5.615 0.235 ;
        RECT 5.805 0.065 5.975 0.235 ;
        RECT 6.165 0.065 6.335 0.235 ;
        RECT 6.525 0.065 6.695 0.235 ;
        RECT 6.885 0.065 7.055 0.235 ;
        RECT 7.375 0.065 7.545 0.235 ;
        RECT 7.735 0.065 7.905 0.235 ;
        RECT 8.095 0.065 8.265 0.235 ;
        RECT 8.455 0.065 8.625 0.235 ;
        RECT 8.815 0.065 8.985 0.235 ;
        RECT 9.175 0.065 9.345 0.235 ;
        RECT 9.895 0.065 10.065 0.235 ;
        RECT 10.255 0.065 10.425 0.235 ;
        RECT 10.615 0.065 10.785 0.235 ;
        RECT 10.975 0.065 11.145 0.235 ;
        RECT 11.335 0.065 11.505 0.235 ;
        RECT 11.695 0.065 11.865 0.235 ;
        RECT 12.185 0.065 12.355 0.235 ;
        RECT 12.545 0.065 12.715 0.235 ;
        RECT 12.905 0.065 13.075 0.235 ;
        RECT 13.265 0.065 13.435 0.235 ;
        RECT 13.625 0.065 13.795 0.235 ;
        RECT 13.985 0.065 14.155 0.235 ;
        RECT 14.705 0.065 14.875 0.235 ;
        RECT 15.065 0.065 15.235 0.235 ;
        RECT 15.425 0.065 15.595 0.235 ;
        RECT 15.785 0.065 15.955 0.235 ;
        RECT 16.145 0.065 16.315 0.235 ;
        RECT 16.505 0.065 16.675 0.235 ;
        RECT 16.995 0.065 17.165 0.235 ;
        RECT 17.355 0.065 17.525 0.235 ;
        RECT 17.715 0.065 17.885 0.235 ;
        RECT 18.075 0.065 18.245 0.235 ;
        RECT 18.435 0.065 18.605 0.235 ;
        RECT 18.795 0.065 18.965 0.235 ;
        RECT 19.515 0.065 19.685 0.235 ;
        RECT 19.875 0.065 20.045 0.235 ;
        RECT 20.235 0.065 20.405 0.235 ;
        RECT 20.595 0.065 20.765 0.235 ;
        RECT 20.955 0.065 21.125 0.235 ;
        RECT 21.315 0.065 21.485 0.235 ;
        RECT 21.805 0.065 21.975 0.235 ;
        RECT 22.165 0.065 22.335 0.235 ;
        RECT 22.525 0.065 22.695 0.235 ;
        RECT 22.885 0.065 23.055 0.235 ;
        RECT 23.245 0.065 23.415 0.235 ;
        RECT 23.605 0.065 23.775 0.235 ;
        RECT 24.325 0.065 24.495 0.235 ;
        RECT 24.685 0.065 24.855 0.235 ;
        RECT 25.045 0.065 25.215 0.235 ;
        RECT 25.405 0.065 25.575 0.235 ;
        RECT 25.765 0.065 25.935 0.235 ;
        RECT 26.125 0.065 26.295 0.235 ;
        RECT 26.615 0.065 26.785 0.235 ;
        RECT 26.975 0.065 27.145 0.235 ;
        RECT 27.335 0.065 27.505 0.235 ;
        RECT 27.695 0.065 27.865 0.235 ;
        RECT 28.055 0.065 28.225 0.235 ;
        RECT 28.415 0.065 28.585 0.235 ;
        RECT 29.135 0.065 29.305 0.235 ;
        RECT 29.495 0.065 29.665 0.235 ;
        RECT 29.855 0.065 30.025 0.235 ;
        RECT 30.215 0.065 30.385 0.235 ;
        RECT 30.575 0.065 30.745 0.235 ;
        RECT 30.935 0.065 31.105 0.235 ;
        RECT 31.425 0.065 31.595 0.235 ;
        RECT 31.785 0.065 31.955 0.235 ;
        RECT 32.145 0.065 32.315 0.235 ;
        RECT 32.505 0.065 32.675 0.235 ;
        RECT 32.865 0.065 33.035 0.235 ;
        RECT 33.225 0.065 33.395 0.235 ;
        RECT 33.945 0.065 34.115 0.235 ;
        RECT 34.305 0.065 34.475 0.235 ;
        RECT 34.665 0.065 34.835 0.235 ;
        RECT 35.025 0.065 35.195 0.235 ;
        RECT 35.385 0.065 35.555 0.235 ;
        RECT 35.745 0.065 35.915 0.235 ;
        RECT 36.235 0.065 36.405 0.235 ;
        RECT 36.595 0.065 36.765 0.235 ;
        RECT 36.955 0.065 37.125 0.235 ;
        RECT 37.315 0.065 37.485 0.235 ;
        RECT 37.675 0.065 37.845 0.235 ;
        RECT 38.035 0.065 38.205 0.235 ;
        RECT 38.755 0.065 38.925 0.235 ;
        RECT 39.115 0.065 39.285 0.235 ;
        RECT 39.475 0.065 39.645 0.235 ;
        RECT 39.835 0.065 40.005 0.235 ;
        RECT 40.195 0.065 40.365 0.235 ;
        RECT 40.555 0.065 40.725 0.235 ;
        RECT 41.045 0.065 41.215 0.235 ;
        RECT 41.405 0.065 41.575 0.235 ;
        RECT 41.765 0.065 41.935 0.235 ;
        RECT 42.125 0.065 42.295 0.235 ;
        RECT 42.485 0.065 42.655 0.235 ;
        RECT 42.845 0.065 43.015 0.235 ;
        RECT 43.565 0.065 43.735 0.235 ;
        RECT 43.925 0.065 44.095 0.235 ;
        RECT 44.285 0.065 44.455 0.235 ;
        RECT 44.645 0.065 44.815 0.235 ;
        RECT 45.005 0.065 45.175 0.235 ;
        RECT 45.365 0.065 45.535 0.235 ;
        RECT 45.855 0.065 46.025 0.235 ;
        RECT 46.215 0.065 46.385 0.235 ;
        RECT 46.575 0.065 46.745 0.235 ;
        RECT 46.935 0.065 47.105 0.235 ;
        RECT 47.295 0.065 47.465 0.235 ;
        RECT 47.655 0.065 47.825 0.235 ;
        RECT 48.375 0.065 48.545 0.235 ;
        RECT 48.735 0.065 48.905 0.235 ;
        RECT 49.095 0.065 49.265 0.235 ;
        RECT 49.455 0.065 49.625 0.235 ;
        RECT 49.815 0.065 49.985 0.235 ;
        RECT 50.175 0.065 50.345 0.235 ;
        RECT 50.665 0.065 50.835 0.235 ;
        RECT 51.025 0.065 51.195 0.235 ;
        RECT 51.385 0.065 51.555 0.235 ;
        RECT 51.745 0.065 51.915 0.235 ;
        RECT 52.105 0.065 52.275 0.235 ;
        RECT 52.465 0.065 52.635 0.235 ;
        RECT 53.185 0.065 53.355 0.235 ;
        RECT 53.545 0.065 53.715 0.235 ;
        RECT 53.905 0.065 54.075 0.235 ;
        RECT 54.265 0.065 54.435 0.235 ;
        RECT 54.625 0.065 54.795 0.235 ;
        RECT 54.985 0.065 55.155 0.235 ;
        RECT 55.475 0.065 55.645 0.235 ;
        RECT 55.835 0.065 56.005 0.235 ;
        RECT 56.195 0.065 56.365 0.235 ;
        RECT 56.555 0.065 56.725 0.235 ;
        RECT 56.915 0.065 57.085 0.235 ;
        RECT 57.275 0.065 57.445 0.235 ;
        RECT 57.995 0.065 58.165 0.235 ;
        RECT 58.355 0.065 58.525 0.235 ;
        RECT 58.715 0.065 58.885 0.235 ;
        RECT 59.075 0.065 59.245 0.235 ;
        RECT 59.435 0.065 59.605 0.235 ;
        RECT 59.795 0.065 59.965 0.235 ;
        RECT 60.285 0.065 60.455 0.235 ;
        RECT 60.645 0.065 60.815 0.235 ;
        RECT 61.005 0.065 61.175 0.235 ;
        RECT 61.365 0.065 61.535 0.235 ;
        RECT 61.725 0.065 61.895 0.235 ;
        RECT 62.085 0.065 62.255 0.235 ;
        RECT 62.805 0.065 62.975 0.235 ;
        RECT 63.165 0.065 63.335 0.235 ;
        RECT 63.525 0.065 63.695 0.235 ;
        RECT 63.885 0.065 64.055 0.235 ;
        RECT 64.245 0.065 64.415 0.235 ;
        RECT 64.605 0.065 64.775 0.235 ;
        RECT 65.095 0.065 65.265 0.235 ;
        RECT 65.455 0.065 65.625 0.235 ;
        RECT 65.815 0.065 65.985 0.235 ;
        RECT 66.175 0.065 66.345 0.235 ;
        RECT 66.535 0.065 66.705 0.235 ;
        RECT 66.895 0.065 67.065 0.235 ;
        RECT 67.615 0.065 67.785 0.235 ;
        RECT 67.975 0.065 68.145 0.235 ;
        RECT 68.335 0.065 68.505 0.235 ;
        RECT 68.695 0.065 68.865 0.235 ;
        RECT 69.055 0.065 69.225 0.235 ;
        RECT 69.415 0.065 69.585 0.235 ;
        RECT 69.905 0.065 70.075 0.235 ;
        RECT 70.265 0.065 70.435 0.235 ;
        RECT 70.625 0.065 70.795 0.235 ;
        RECT 70.985 0.065 71.155 0.235 ;
        RECT 71.345 0.065 71.515 0.235 ;
        RECT 71.705 0.065 71.875 0.235 ;
        RECT 72.425 0.065 72.595 0.235 ;
        RECT 72.785 0.065 72.955 0.235 ;
        RECT 73.145 0.065 73.315 0.235 ;
        RECT 73.505 0.065 73.675 0.235 ;
        RECT 73.865 0.065 74.035 0.235 ;
        RECT 74.225 0.065 74.395 0.235 ;
        RECT 74.715 0.065 74.885 0.235 ;
        RECT 75.075 0.065 75.245 0.235 ;
        RECT 75.435 0.065 75.605 0.235 ;
        RECT 75.795 0.065 75.965 0.235 ;
        RECT 76.155 0.065 76.325 0.235 ;
        RECT 76.515 0.065 76.685 0.235 ;
        RECT 77.235 0.065 77.405 0.235 ;
        RECT 77.595 0.065 77.765 0.235 ;
        RECT 77.955 0.065 78.125 0.235 ;
        RECT 78.315 0.065 78.485 0.235 ;
        RECT 78.675 0.065 78.845 0.235 ;
        RECT 79.035 0.065 79.205 0.235 ;
        RECT 79.525 0.065 79.695 0.235 ;
        RECT 79.885 0.065 80.055 0.235 ;
        RECT 80.245 0.065 80.415 0.235 ;
        RECT 80.605 0.065 80.775 0.235 ;
        RECT 80.965 0.065 81.135 0.235 ;
        RECT 81.325 0.065 81.495 0.235 ;
        RECT 82.045 0.065 82.215 0.235 ;
        RECT 82.405 0.065 82.575 0.235 ;
        RECT 82.765 0.065 82.935 0.235 ;
        RECT 83.125 0.065 83.295 0.235 ;
        RECT 83.485 0.065 83.655 0.235 ;
        RECT 83.845 0.065 84.015 0.235 ;
        RECT 84.335 0.065 84.505 0.235 ;
        RECT 84.695 0.065 84.865 0.235 ;
        RECT 85.055 0.065 85.225 0.235 ;
        RECT 85.415 0.065 85.585 0.235 ;
        RECT 85.775 0.065 85.945 0.235 ;
        RECT 86.135 0.065 86.305 0.235 ;
        RECT 86.855 0.065 87.025 0.235 ;
        RECT 87.215 0.065 87.385 0.235 ;
        RECT 87.575 0.065 87.745 0.235 ;
        RECT 87.935 0.065 88.105 0.235 ;
        RECT 88.385 0.065 88.555 0.235 ;
        RECT 88.745 0.065 88.915 0.235 ;
        RECT 89.105 0.065 89.275 0.235 ;
        RECT 89.465 0.065 89.635 0.235 ;
        RECT 90.185 0.065 90.355 0.235 ;
        RECT 90.545 0.065 90.715 0.235 ;
        RECT 90.905 0.065 91.075 0.235 ;
        RECT 91.265 0.065 91.435 0.235 ;
        RECT 91.715 0.065 91.885 0.235 ;
        RECT 92.075 0.065 92.245 0.235 ;
        RECT 92.435 0.065 92.605 0.235 ;
        RECT 92.795 0.065 92.965 0.235 ;
        RECT 93.515 0.065 93.685 0.235 ;
        RECT 93.875 0.065 94.045 0.235 ;
        RECT 94.235 0.065 94.405 0.235 ;
        RECT 94.595 0.065 94.765 0.235 ;
        RECT 95.045 0.065 95.215 0.235 ;
        RECT 95.405 0.065 95.575 0.235 ;
        RECT 95.765 0.065 95.935 0.235 ;
        RECT 96.125 0.065 96.295 0.235 ;
        RECT 96.845 0.065 97.015 0.235 ;
        RECT 97.205 0.065 97.375 0.235 ;
        RECT 97.595 0.065 97.765 0.235 ;
        RECT 97.985 0.065 98.155 0.235 ;
        RECT 98.345 0.065 98.515 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 98.945 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 1.445 5.470 1.615 7.250 ;
        RECT 2.325 5.470 2.495 7.250 ;
        RECT 3.205 5.470 3.375 7.250 ;
        RECT 6.255 5.470 6.425 7.250 ;
        RECT 7.135 5.470 7.305 7.250 ;
        RECT 8.015 5.470 8.185 7.250 ;
        RECT 11.065 5.470 11.235 7.250 ;
        RECT 11.945 5.470 12.115 7.250 ;
        RECT 12.825 5.470 12.995 7.250 ;
        RECT 15.875 5.470 16.045 7.250 ;
        RECT 16.755 5.470 16.925 7.250 ;
        RECT 17.635 5.470 17.805 7.250 ;
        RECT 20.685 5.470 20.855 7.250 ;
        RECT 21.565 5.470 21.735 7.250 ;
        RECT 22.445 5.470 22.615 7.250 ;
        RECT 25.495 5.470 25.665 7.250 ;
        RECT 26.375 5.470 26.545 7.250 ;
        RECT 27.255 5.470 27.425 7.250 ;
        RECT 30.305 5.470 30.475 7.250 ;
        RECT 31.185 5.470 31.355 7.250 ;
        RECT 32.065 5.470 32.235 7.250 ;
        RECT 35.115 5.470 35.285 7.250 ;
        RECT 35.995 5.470 36.165 7.250 ;
        RECT 36.875 5.470 37.045 7.250 ;
        RECT 39.925 5.470 40.095 7.250 ;
        RECT 40.805 5.470 40.975 7.250 ;
        RECT 41.685 5.470 41.855 7.250 ;
        RECT 44.735 5.470 44.905 7.250 ;
        RECT 45.615 5.470 45.785 7.250 ;
        RECT 46.495 5.470 46.665 7.250 ;
        RECT 49.545 5.470 49.715 7.250 ;
        RECT 50.425 5.470 50.595 7.250 ;
        RECT 51.305 5.470 51.475 7.250 ;
        RECT 54.355 5.470 54.525 7.250 ;
        RECT 55.235 5.470 55.405 7.250 ;
        RECT 56.115 5.470 56.285 7.250 ;
        RECT 59.165 5.470 59.335 7.250 ;
        RECT 60.045 5.470 60.215 7.250 ;
        RECT 60.925 5.470 61.095 7.250 ;
        RECT 63.975 5.470 64.145 7.250 ;
        RECT 64.855 5.470 65.025 7.250 ;
        RECT 65.735 5.470 65.905 7.250 ;
        RECT 68.785 5.470 68.955 7.250 ;
        RECT 69.665 5.470 69.835 7.250 ;
        RECT 70.545 5.470 70.715 7.250 ;
        RECT 73.595 5.470 73.765 7.250 ;
        RECT 74.475 5.470 74.645 7.250 ;
        RECT 75.355 5.470 75.525 7.250 ;
        RECT 78.405 5.470 78.575 7.250 ;
        RECT 79.285 5.470 79.455 7.250 ;
        RECT 80.165 5.470 80.335 7.250 ;
        RECT 83.215 5.470 83.385 7.250 ;
        RECT 84.095 5.470 84.265 7.250 ;
        RECT 84.975 5.470 85.145 7.250 ;
        RECT 87.725 7.055 87.905 7.225 ;
        RECT 87.725 5.525 87.895 7.055 ;
        RECT 88.605 5.525 88.775 7.225 ;
        RECT 1.445 5.300 4.155 5.470 ;
        RECT 6.255 5.300 8.965 5.470 ;
        RECT 11.065 5.300 13.775 5.470 ;
        RECT 15.875 5.300 18.585 5.470 ;
        RECT 20.685 5.300 23.395 5.470 ;
        RECT 25.495 5.300 28.205 5.470 ;
        RECT 30.305 5.300 33.015 5.470 ;
        RECT 35.115 5.300 37.825 5.470 ;
        RECT 39.925 5.300 42.635 5.470 ;
        RECT 44.735 5.300 47.445 5.470 ;
        RECT 49.545 5.300 52.255 5.470 ;
        RECT 54.355 5.300 57.065 5.470 ;
        RECT 59.165 5.300 61.875 5.470 ;
        RECT 63.975 5.300 66.685 5.470 ;
        RECT 68.785 5.300 71.495 5.470 ;
        RECT 73.595 5.300 76.305 5.470 ;
        RECT 78.405 5.300 81.115 5.470 ;
        RECT 83.215 5.300 85.925 5.470 ;
        RECT 87.725 5.355 88.775 5.525 ;
        RECT 3.245 2.055 3.415 5.095 ;
        RECT 0.505 1.815 0.675 1.895 ;
        RECT 1.475 1.815 1.645 1.895 ;
        RECT 2.445 1.815 2.615 1.895 ;
        RECT 0.505 1.645 2.615 1.815 ;
        RECT 0.505 0.515 0.675 1.645 ;
        RECT 1.475 0.765 1.645 1.645 ;
        RECT 2.445 1.565 2.615 1.645 ;
        RECT 1.965 1.220 2.135 1.300 ;
        RECT 3.015 1.220 3.185 1.895 ;
        RECT 3.985 1.890 4.155 5.300 ;
        RECT 5.835 2.055 6.005 5.095 ;
        RECT 8.055 4.235 8.225 5.095 ;
        RECT 8.050 3.905 8.225 4.235 ;
        RECT 8.055 2.055 8.225 3.905 ;
        RECT 1.965 1.050 3.185 1.220 ;
        RECT 1.965 0.970 2.135 1.050 ;
        RECT 2.445 0.765 2.615 0.845 ;
        RECT 1.475 0.595 2.615 0.765 ;
        RECT 1.475 0.515 1.645 0.595 ;
        RECT 2.445 0.515 2.615 0.595 ;
        RECT 3.015 0.765 3.185 1.050 ;
        RECT 3.500 1.720 4.155 1.890 ;
        RECT 5.315 1.815 5.485 1.895 ;
        RECT 6.285 1.815 6.455 1.895 ;
        RECT 7.255 1.815 7.425 1.895 ;
        RECT 3.500 0.985 3.670 1.720 ;
        RECT 5.315 1.645 7.425 1.815 ;
        RECT 3.985 0.765 4.155 1.535 ;
        RECT 3.015 0.595 4.155 0.765 ;
        RECT 3.015 0.515 3.185 0.595 ;
        RECT 3.985 0.515 4.155 0.595 ;
        RECT 5.315 0.515 5.485 1.645 ;
        RECT 6.285 0.765 6.455 1.645 ;
        RECT 7.255 1.565 7.425 1.645 ;
        RECT 6.775 1.220 6.945 1.300 ;
        RECT 7.825 1.220 7.995 1.895 ;
        RECT 8.795 1.890 8.965 5.300 ;
        RECT 10.645 2.055 10.815 5.095 ;
        RECT 12.865 2.055 13.035 5.095 ;
        RECT 6.775 1.050 7.995 1.220 ;
        RECT 6.775 0.970 6.945 1.050 ;
        RECT 7.255 0.765 7.425 0.845 ;
        RECT 6.285 0.595 7.425 0.765 ;
        RECT 6.285 0.515 6.455 0.595 ;
        RECT 7.255 0.515 7.425 0.595 ;
        RECT 7.825 0.765 7.995 1.050 ;
        RECT 8.310 1.720 8.965 1.890 ;
        RECT 10.125 1.815 10.295 1.895 ;
        RECT 11.095 1.815 11.265 1.895 ;
        RECT 12.065 1.815 12.235 1.895 ;
        RECT 8.310 0.985 8.480 1.720 ;
        RECT 10.125 1.645 12.235 1.815 ;
        RECT 8.795 0.765 8.965 1.535 ;
        RECT 7.825 0.595 8.965 0.765 ;
        RECT 7.825 0.515 7.995 0.595 ;
        RECT 8.795 0.515 8.965 0.595 ;
        RECT 10.125 0.515 10.295 1.645 ;
        RECT 11.095 0.765 11.265 1.645 ;
        RECT 12.065 1.565 12.235 1.645 ;
        RECT 11.585 1.220 11.755 1.300 ;
        RECT 12.635 1.220 12.805 1.895 ;
        RECT 13.605 1.890 13.775 5.300 ;
        RECT 15.455 2.055 15.625 5.095 ;
        RECT 11.585 1.050 12.805 1.220 ;
        RECT 11.585 0.970 11.755 1.050 ;
        RECT 12.065 0.765 12.235 0.845 ;
        RECT 11.095 0.595 12.235 0.765 ;
        RECT 11.095 0.515 11.265 0.595 ;
        RECT 12.065 0.515 12.235 0.595 ;
        RECT 12.635 0.765 12.805 1.050 ;
        RECT 13.120 1.720 13.775 1.890 ;
        RECT 14.935 1.815 15.105 1.895 ;
        RECT 15.905 1.815 16.075 1.895 ;
        RECT 16.875 1.815 17.045 1.895 ;
        RECT 13.120 0.985 13.290 1.720 ;
        RECT 14.935 1.645 17.045 1.815 ;
        RECT 13.605 0.765 13.775 1.535 ;
        RECT 12.635 0.595 13.775 0.765 ;
        RECT 12.635 0.515 12.805 0.595 ;
        RECT 13.605 0.515 13.775 0.595 ;
        RECT 14.935 0.515 15.105 1.645 ;
        RECT 15.905 0.765 16.075 1.645 ;
        RECT 16.875 1.565 17.045 1.645 ;
        RECT 16.395 1.220 16.565 1.300 ;
        RECT 17.445 1.220 17.615 1.895 ;
        RECT 18.415 1.890 18.585 5.300 ;
        RECT 20.265 2.055 20.435 5.095 ;
        RECT 22.485 2.055 22.655 5.095 ;
        RECT 16.395 1.050 17.615 1.220 ;
        RECT 16.395 0.970 16.565 1.050 ;
        RECT 16.875 0.765 17.045 0.845 ;
        RECT 15.905 0.595 17.045 0.765 ;
        RECT 15.905 0.515 16.075 0.595 ;
        RECT 16.875 0.515 17.045 0.595 ;
        RECT 17.445 0.765 17.615 1.050 ;
        RECT 17.930 1.720 18.585 1.890 ;
        RECT 19.745 1.815 19.915 1.895 ;
        RECT 20.715 1.815 20.885 1.895 ;
        RECT 21.685 1.815 21.855 1.895 ;
        RECT 17.930 0.985 18.100 1.720 ;
        RECT 19.745 1.645 21.855 1.815 ;
        RECT 18.415 0.765 18.585 1.535 ;
        RECT 17.445 0.595 18.585 0.765 ;
        RECT 17.445 0.515 17.615 0.595 ;
        RECT 18.415 0.515 18.585 0.595 ;
        RECT 19.745 0.515 19.915 1.645 ;
        RECT 20.715 0.765 20.885 1.645 ;
        RECT 21.685 1.565 21.855 1.645 ;
        RECT 21.205 1.220 21.375 1.300 ;
        RECT 22.255 1.220 22.425 1.895 ;
        RECT 23.225 1.890 23.395 5.300 ;
        RECT 25.075 2.055 25.245 5.095 ;
        RECT 27.295 2.055 27.465 5.095 ;
        RECT 21.205 1.050 22.425 1.220 ;
        RECT 21.205 0.970 21.375 1.050 ;
        RECT 21.685 0.765 21.855 0.845 ;
        RECT 20.715 0.595 21.855 0.765 ;
        RECT 20.715 0.515 20.885 0.595 ;
        RECT 21.685 0.515 21.855 0.595 ;
        RECT 22.255 0.765 22.425 1.050 ;
        RECT 22.740 1.720 23.395 1.890 ;
        RECT 24.555 1.815 24.725 1.895 ;
        RECT 25.525 1.815 25.695 1.895 ;
        RECT 26.495 1.815 26.665 1.895 ;
        RECT 22.740 0.985 22.910 1.720 ;
        RECT 24.555 1.645 26.665 1.815 ;
        RECT 23.225 0.765 23.395 1.535 ;
        RECT 22.255 0.595 23.395 0.765 ;
        RECT 22.255 0.515 22.425 0.595 ;
        RECT 23.225 0.515 23.395 0.595 ;
        RECT 24.555 0.515 24.725 1.645 ;
        RECT 25.525 0.765 25.695 1.645 ;
        RECT 26.495 1.565 26.665 1.645 ;
        RECT 26.015 1.220 26.185 1.300 ;
        RECT 27.065 1.220 27.235 1.895 ;
        RECT 28.035 1.890 28.205 5.300 ;
        RECT 32.105 2.055 32.275 5.095 ;
        RECT 26.015 1.050 27.235 1.220 ;
        RECT 26.015 0.970 26.185 1.050 ;
        RECT 26.495 0.765 26.665 0.845 ;
        RECT 25.525 0.595 26.665 0.765 ;
        RECT 25.525 0.515 25.695 0.595 ;
        RECT 26.495 0.515 26.665 0.595 ;
        RECT 27.065 0.765 27.235 1.050 ;
        RECT 27.550 1.720 28.205 1.890 ;
        RECT 29.365 1.815 29.535 1.895 ;
        RECT 30.335 1.815 30.505 1.895 ;
        RECT 31.305 1.815 31.475 1.895 ;
        RECT 27.550 0.985 27.720 1.720 ;
        RECT 29.365 1.645 31.475 1.815 ;
        RECT 28.035 0.765 28.205 1.535 ;
        RECT 27.065 0.595 28.205 0.765 ;
        RECT 27.065 0.515 27.235 0.595 ;
        RECT 28.035 0.515 28.205 0.595 ;
        RECT 29.365 0.515 29.535 1.645 ;
        RECT 30.335 0.765 30.505 1.645 ;
        RECT 31.305 1.565 31.475 1.645 ;
        RECT 30.825 1.220 30.995 1.300 ;
        RECT 31.875 1.220 32.045 1.895 ;
        RECT 32.845 1.890 33.015 5.300 ;
        RECT 34.695 2.055 34.865 5.095 ;
        RECT 36.915 4.235 37.085 5.095 ;
        RECT 36.910 3.905 37.085 4.235 ;
        RECT 36.915 2.055 37.085 3.905 ;
        RECT 30.825 1.050 32.045 1.220 ;
        RECT 30.825 0.970 30.995 1.050 ;
        RECT 31.305 0.765 31.475 0.845 ;
        RECT 30.335 0.595 31.475 0.765 ;
        RECT 30.335 0.515 30.505 0.595 ;
        RECT 31.305 0.515 31.475 0.595 ;
        RECT 31.875 0.765 32.045 1.050 ;
        RECT 32.360 1.720 33.015 1.890 ;
        RECT 34.175 1.815 34.345 1.895 ;
        RECT 35.145 1.815 35.315 1.895 ;
        RECT 36.115 1.815 36.285 1.895 ;
        RECT 32.360 0.985 32.530 1.720 ;
        RECT 34.175 1.645 36.285 1.815 ;
        RECT 32.845 0.765 33.015 1.535 ;
        RECT 31.875 0.595 33.015 0.765 ;
        RECT 31.875 0.515 32.045 0.595 ;
        RECT 32.845 0.515 33.015 0.595 ;
        RECT 34.175 0.515 34.345 1.645 ;
        RECT 35.145 0.765 35.315 1.645 ;
        RECT 36.115 1.565 36.285 1.645 ;
        RECT 35.635 1.220 35.805 1.300 ;
        RECT 36.685 1.220 36.855 1.895 ;
        RECT 37.655 1.890 37.825 5.300 ;
        RECT 39.505 2.055 39.675 5.095 ;
        RECT 41.725 2.055 41.895 5.095 ;
        RECT 35.635 1.050 36.855 1.220 ;
        RECT 35.635 0.970 35.805 1.050 ;
        RECT 36.115 0.765 36.285 0.845 ;
        RECT 35.145 0.595 36.285 0.765 ;
        RECT 35.145 0.515 35.315 0.595 ;
        RECT 36.115 0.515 36.285 0.595 ;
        RECT 36.685 0.765 36.855 1.050 ;
        RECT 37.170 1.720 37.825 1.890 ;
        RECT 38.985 1.815 39.155 1.895 ;
        RECT 39.955 1.815 40.125 1.895 ;
        RECT 40.925 1.815 41.095 1.895 ;
        RECT 37.170 0.985 37.340 1.720 ;
        RECT 38.985 1.645 41.095 1.815 ;
        RECT 37.655 0.765 37.825 1.535 ;
        RECT 36.685 0.595 37.825 0.765 ;
        RECT 36.685 0.515 36.855 0.595 ;
        RECT 37.655 0.515 37.825 0.595 ;
        RECT 38.985 0.515 39.155 1.645 ;
        RECT 39.955 0.765 40.125 1.645 ;
        RECT 40.925 1.565 41.095 1.645 ;
        RECT 40.445 1.220 40.615 1.300 ;
        RECT 41.495 1.220 41.665 1.895 ;
        RECT 42.465 1.890 42.635 5.300 ;
        RECT 44.315 2.055 44.485 5.095 ;
        RECT 40.445 1.050 41.665 1.220 ;
        RECT 40.445 0.970 40.615 1.050 ;
        RECT 40.925 0.765 41.095 0.845 ;
        RECT 39.955 0.595 41.095 0.765 ;
        RECT 39.955 0.515 40.125 0.595 ;
        RECT 40.925 0.515 41.095 0.595 ;
        RECT 41.495 0.765 41.665 1.050 ;
        RECT 41.980 1.720 42.635 1.890 ;
        RECT 43.795 1.815 43.965 1.895 ;
        RECT 44.765 1.815 44.935 1.895 ;
        RECT 45.735 1.815 45.905 1.895 ;
        RECT 41.980 0.985 42.150 1.720 ;
        RECT 43.795 1.645 45.905 1.815 ;
        RECT 42.465 0.765 42.635 1.535 ;
        RECT 41.495 0.595 42.635 0.765 ;
        RECT 41.495 0.515 41.665 0.595 ;
        RECT 42.465 0.515 42.635 0.595 ;
        RECT 43.795 0.515 43.965 1.645 ;
        RECT 44.765 0.765 44.935 1.645 ;
        RECT 45.735 1.565 45.905 1.645 ;
        RECT 45.255 1.220 45.425 1.300 ;
        RECT 46.305 1.220 46.475 1.895 ;
        RECT 47.275 1.890 47.445 5.300 ;
        RECT 49.125 2.055 49.295 5.095 ;
        RECT 51.345 2.055 51.515 5.095 ;
        RECT 45.255 1.050 46.475 1.220 ;
        RECT 45.255 0.970 45.425 1.050 ;
        RECT 45.735 0.765 45.905 0.845 ;
        RECT 44.765 0.595 45.905 0.765 ;
        RECT 44.765 0.515 44.935 0.595 ;
        RECT 45.735 0.515 45.905 0.595 ;
        RECT 46.305 0.765 46.475 1.050 ;
        RECT 46.790 1.720 47.445 1.890 ;
        RECT 48.605 1.815 48.775 1.895 ;
        RECT 49.575 1.815 49.745 1.895 ;
        RECT 50.545 1.815 50.715 1.895 ;
        RECT 46.790 0.985 46.960 1.720 ;
        RECT 48.605 1.645 50.715 1.815 ;
        RECT 47.275 0.765 47.445 1.535 ;
        RECT 46.305 0.595 47.445 0.765 ;
        RECT 46.305 0.515 46.475 0.595 ;
        RECT 47.275 0.515 47.445 0.595 ;
        RECT 48.605 0.515 48.775 1.645 ;
        RECT 49.575 0.765 49.745 1.645 ;
        RECT 50.545 1.565 50.715 1.645 ;
        RECT 50.065 1.220 50.235 1.300 ;
        RECT 51.115 1.220 51.285 1.895 ;
        RECT 52.085 1.890 52.255 5.300 ;
        RECT 53.935 2.055 54.105 5.095 ;
        RECT 56.155 2.055 56.325 5.095 ;
        RECT 50.065 1.050 51.285 1.220 ;
        RECT 50.065 0.970 50.235 1.050 ;
        RECT 50.545 0.765 50.715 0.845 ;
        RECT 49.575 0.595 50.715 0.765 ;
        RECT 49.575 0.515 49.745 0.595 ;
        RECT 50.545 0.515 50.715 0.595 ;
        RECT 51.115 0.765 51.285 1.050 ;
        RECT 51.600 1.720 52.255 1.890 ;
        RECT 53.415 1.815 53.585 1.895 ;
        RECT 54.385 1.815 54.555 1.895 ;
        RECT 55.355 1.815 55.525 1.895 ;
        RECT 51.600 0.985 51.770 1.720 ;
        RECT 53.415 1.645 55.525 1.815 ;
        RECT 52.085 0.765 52.255 1.535 ;
        RECT 51.115 0.595 52.255 0.765 ;
        RECT 51.115 0.515 51.285 0.595 ;
        RECT 52.085 0.515 52.255 0.595 ;
        RECT 53.415 0.515 53.585 1.645 ;
        RECT 54.385 0.765 54.555 1.645 ;
        RECT 55.355 1.565 55.525 1.645 ;
        RECT 54.875 1.220 55.045 1.300 ;
        RECT 55.925 1.220 56.095 1.895 ;
        RECT 56.895 1.890 57.065 5.300 ;
        RECT 60.965 2.055 61.135 5.095 ;
        RECT 54.875 1.050 56.095 1.220 ;
        RECT 54.875 0.970 55.045 1.050 ;
        RECT 55.355 0.765 55.525 0.845 ;
        RECT 54.385 0.595 55.525 0.765 ;
        RECT 54.385 0.515 54.555 0.595 ;
        RECT 55.355 0.515 55.525 0.595 ;
        RECT 55.925 0.765 56.095 1.050 ;
        RECT 56.410 1.720 57.065 1.890 ;
        RECT 58.225 1.815 58.395 1.895 ;
        RECT 59.195 1.815 59.365 1.895 ;
        RECT 60.165 1.815 60.335 1.895 ;
        RECT 56.410 0.985 56.580 1.720 ;
        RECT 58.225 1.645 60.335 1.815 ;
        RECT 56.895 0.765 57.065 1.535 ;
        RECT 55.925 0.595 57.065 0.765 ;
        RECT 55.925 0.515 56.095 0.595 ;
        RECT 56.895 0.515 57.065 0.595 ;
        RECT 58.225 0.515 58.395 1.645 ;
        RECT 59.195 0.765 59.365 1.645 ;
        RECT 60.165 1.565 60.335 1.645 ;
        RECT 59.685 1.220 59.855 1.300 ;
        RECT 60.735 1.220 60.905 1.895 ;
        RECT 61.705 1.890 61.875 5.300 ;
        RECT 63.555 2.055 63.725 5.095 ;
        RECT 65.775 4.235 65.945 5.095 ;
        RECT 65.770 3.905 65.945 4.235 ;
        RECT 65.775 2.055 65.945 3.905 ;
        RECT 59.685 1.050 60.905 1.220 ;
        RECT 59.685 0.970 59.855 1.050 ;
        RECT 60.165 0.765 60.335 0.845 ;
        RECT 59.195 0.595 60.335 0.765 ;
        RECT 59.195 0.515 59.365 0.595 ;
        RECT 60.165 0.515 60.335 0.595 ;
        RECT 60.735 0.765 60.905 1.050 ;
        RECT 61.220 1.720 61.875 1.890 ;
        RECT 63.035 1.815 63.205 1.895 ;
        RECT 64.005 1.815 64.175 1.895 ;
        RECT 64.975 1.815 65.145 1.895 ;
        RECT 61.220 0.985 61.390 1.720 ;
        RECT 63.035 1.645 65.145 1.815 ;
        RECT 61.705 0.765 61.875 1.535 ;
        RECT 60.735 0.595 61.875 0.765 ;
        RECT 60.735 0.515 60.905 0.595 ;
        RECT 61.705 0.515 61.875 0.595 ;
        RECT 63.035 0.515 63.205 1.645 ;
        RECT 64.005 0.765 64.175 1.645 ;
        RECT 64.975 1.565 65.145 1.645 ;
        RECT 64.495 1.220 64.665 1.300 ;
        RECT 65.545 1.220 65.715 1.895 ;
        RECT 66.515 1.890 66.685 5.300 ;
        RECT 68.365 2.055 68.535 5.095 ;
        RECT 70.585 2.055 70.755 5.095 ;
        RECT 64.495 1.050 65.715 1.220 ;
        RECT 64.495 0.970 64.665 1.050 ;
        RECT 64.975 0.765 65.145 0.845 ;
        RECT 64.005 0.595 65.145 0.765 ;
        RECT 64.005 0.515 64.175 0.595 ;
        RECT 64.975 0.515 65.145 0.595 ;
        RECT 65.545 0.765 65.715 1.050 ;
        RECT 66.030 1.720 66.685 1.890 ;
        RECT 67.845 1.815 68.015 1.895 ;
        RECT 68.815 1.815 68.985 1.895 ;
        RECT 69.785 1.815 69.955 1.895 ;
        RECT 66.030 0.985 66.200 1.720 ;
        RECT 67.845 1.645 69.955 1.815 ;
        RECT 66.515 0.765 66.685 1.535 ;
        RECT 65.545 0.595 66.685 0.765 ;
        RECT 65.545 0.515 65.715 0.595 ;
        RECT 66.515 0.515 66.685 0.595 ;
        RECT 67.845 0.515 68.015 1.645 ;
        RECT 68.815 0.765 68.985 1.645 ;
        RECT 69.785 1.565 69.955 1.645 ;
        RECT 69.305 1.220 69.475 1.300 ;
        RECT 70.355 1.220 70.525 1.895 ;
        RECT 71.325 1.890 71.495 5.300 ;
        RECT 73.175 2.055 73.345 5.095 ;
        RECT 69.305 1.050 70.525 1.220 ;
        RECT 69.305 0.970 69.475 1.050 ;
        RECT 69.785 0.765 69.955 0.845 ;
        RECT 68.815 0.595 69.955 0.765 ;
        RECT 68.815 0.515 68.985 0.595 ;
        RECT 69.785 0.515 69.955 0.595 ;
        RECT 70.355 0.765 70.525 1.050 ;
        RECT 70.840 1.720 71.495 1.890 ;
        RECT 72.655 1.815 72.825 1.895 ;
        RECT 73.625 1.815 73.795 1.895 ;
        RECT 74.595 1.815 74.765 1.895 ;
        RECT 70.840 0.985 71.010 1.720 ;
        RECT 72.655 1.645 74.765 1.815 ;
        RECT 71.325 0.765 71.495 1.535 ;
        RECT 70.355 0.595 71.495 0.765 ;
        RECT 70.355 0.515 70.525 0.595 ;
        RECT 71.325 0.515 71.495 0.595 ;
        RECT 72.655 0.515 72.825 1.645 ;
        RECT 73.625 0.765 73.795 1.645 ;
        RECT 74.595 1.565 74.765 1.645 ;
        RECT 74.115 1.220 74.285 1.300 ;
        RECT 75.165 1.220 75.335 1.895 ;
        RECT 76.135 1.890 76.305 5.300 ;
        RECT 77.985 2.055 78.155 5.095 ;
        RECT 80.205 2.055 80.375 5.095 ;
        RECT 74.115 1.050 75.335 1.220 ;
        RECT 74.115 0.970 74.285 1.050 ;
        RECT 74.595 0.765 74.765 0.845 ;
        RECT 73.625 0.595 74.765 0.765 ;
        RECT 73.625 0.515 73.795 0.595 ;
        RECT 74.595 0.515 74.765 0.595 ;
        RECT 75.165 0.765 75.335 1.050 ;
        RECT 75.650 1.720 76.305 1.890 ;
        RECT 77.465 1.815 77.635 1.895 ;
        RECT 78.435 1.815 78.605 1.895 ;
        RECT 79.405 1.815 79.575 1.895 ;
        RECT 75.650 0.985 75.820 1.720 ;
        RECT 77.465 1.645 79.575 1.815 ;
        RECT 76.135 0.765 76.305 1.535 ;
        RECT 75.165 0.595 76.305 0.765 ;
        RECT 75.165 0.515 75.335 0.595 ;
        RECT 76.135 0.515 76.305 0.595 ;
        RECT 77.465 0.515 77.635 1.645 ;
        RECT 78.435 0.765 78.605 1.645 ;
        RECT 79.405 1.565 79.575 1.645 ;
        RECT 78.925 1.220 79.095 1.300 ;
        RECT 79.975 1.220 80.145 1.895 ;
        RECT 80.945 1.890 81.115 5.300 ;
        RECT 82.795 2.055 82.965 5.095 ;
        RECT 85.015 2.055 85.185 5.095 ;
        RECT 78.925 1.050 80.145 1.220 ;
        RECT 78.925 0.970 79.095 1.050 ;
        RECT 79.405 0.765 79.575 0.845 ;
        RECT 78.435 0.595 79.575 0.765 ;
        RECT 78.435 0.515 78.605 0.595 ;
        RECT 79.405 0.515 79.575 0.595 ;
        RECT 79.975 0.765 80.145 1.050 ;
        RECT 80.460 1.720 81.115 1.890 ;
        RECT 82.275 1.815 82.445 1.895 ;
        RECT 83.245 1.815 83.415 1.895 ;
        RECT 84.215 1.815 84.385 1.895 ;
        RECT 80.460 0.985 80.630 1.720 ;
        RECT 82.275 1.645 84.385 1.815 ;
        RECT 80.945 0.765 81.115 1.535 ;
        RECT 79.975 0.595 81.115 0.765 ;
        RECT 79.975 0.515 80.145 0.595 ;
        RECT 80.945 0.515 81.115 0.595 ;
        RECT 82.275 0.515 82.445 1.645 ;
        RECT 83.245 0.765 83.415 1.645 ;
        RECT 84.215 1.565 84.385 1.645 ;
        RECT 83.735 1.220 83.905 1.300 ;
        RECT 84.785 1.220 84.955 1.895 ;
        RECT 85.755 1.890 85.925 5.300 ;
        RECT 88.605 5.275 88.775 5.355 ;
        RECT 90.605 7.055 92.535 7.225 ;
        RECT 90.605 5.275 90.775 7.055 ;
        RECT 91.045 5.525 91.215 6.795 ;
        RECT 91.485 5.785 91.655 7.055 ;
        RECT 91.925 5.525 92.095 6.795 ;
        RECT 92.365 5.605 92.535 7.055 ;
        RECT 93.945 7.055 95.875 7.225 ;
        RECT 91.045 5.355 92.095 5.525 ;
        RECT 91.925 5.275 92.095 5.355 ;
        RECT 93.945 5.275 94.115 7.055 ;
        RECT 94.385 5.525 94.555 6.795 ;
        RECT 94.825 5.785 94.995 7.055 ;
        RECT 95.265 5.525 95.435 6.795 ;
        RECT 95.705 5.785 95.875 7.055 ;
        RECT 94.385 5.355 95.915 5.525 ;
        RECT 87.235 2.055 87.405 5.100 ;
        RECT 88.385 4.940 88.555 5.100 ;
        RECT 88.345 4.770 88.555 4.940 ;
        RECT 88.345 2.055 88.515 4.770 ;
        RECT 90.935 2.055 91.105 5.100 ;
        RECT 92.415 2.055 92.585 5.100 ;
        RECT 93.895 2.055 94.065 5.100 ;
        RECT 95.005 4.770 95.195 5.100 ;
        RECT 95.005 2.055 95.175 4.770 ;
        RECT 83.735 1.050 84.955 1.220 ;
        RECT 83.735 0.970 83.905 1.050 ;
        RECT 84.215 0.765 84.385 0.845 ;
        RECT 83.245 0.595 84.385 0.765 ;
        RECT 83.245 0.515 83.415 0.595 ;
        RECT 84.215 0.515 84.385 0.595 ;
        RECT 84.785 0.765 84.955 1.050 ;
        RECT 85.270 1.720 85.925 1.890 ;
        RECT 87.190 1.805 87.360 1.885 ;
        RECT 88.160 1.805 88.330 1.885 ;
        RECT 85.270 0.985 85.440 1.720 ;
        RECT 87.190 1.635 88.330 1.805 ;
        RECT 85.755 0.765 85.925 1.535 ;
        RECT 84.785 0.595 85.925 0.765 ;
        RECT 84.785 0.515 84.955 0.595 ;
        RECT 85.755 0.515 85.925 0.595 ;
        RECT 87.190 0.505 87.360 1.635 ;
        RECT 88.160 0.755 88.330 1.635 ;
        RECT 88.645 1.310 88.815 1.485 ;
        RECT 88.640 1.155 88.815 1.310 ;
        RECT 88.640 0.975 88.810 1.155 ;
        RECT 89.130 0.755 89.300 1.885 ;
        RECT 88.160 0.585 89.300 0.755 ;
        RECT 88.160 0.505 88.330 0.585 ;
        RECT 89.130 0.505 89.300 0.585 ;
        RECT 90.520 1.805 90.690 1.885 ;
        RECT 91.490 1.805 91.660 1.885 ;
        RECT 90.520 1.635 91.660 1.805 ;
        RECT 90.520 0.505 90.690 1.635 ;
        RECT 91.490 0.755 91.660 1.635 ;
        RECT 91.975 0.975 92.145 1.485 ;
        RECT 92.460 0.755 92.630 1.885 ;
        RECT 91.490 0.585 92.630 0.755 ;
        RECT 91.490 0.505 91.660 0.585 ;
        RECT 92.460 0.505 92.630 0.585 ;
        RECT 93.850 1.805 94.020 1.885 ;
        RECT 94.820 1.805 94.990 1.885 ;
        RECT 95.745 1.870 95.915 5.355 ;
        RECT 97.225 2.055 97.395 5.095 ;
        RECT 93.850 1.635 94.990 1.805 ;
        RECT 93.850 0.505 94.020 1.635 ;
        RECT 94.820 0.755 94.990 1.635 ;
        RECT 95.305 1.700 95.915 1.870 ;
        RECT 95.305 0.975 95.475 1.700 ;
        RECT 95.790 0.755 95.960 1.530 ;
        RECT 94.820 0.585 95.960 0.755 ;
        RECT 94.820 0.505 94.990 0.585 ;
        RECT 95.790 0.505 95.960 0.585 ;
      LAYER mcon ;
        RECT 88.605 5.355 88.775 5.525 ;
        RECT 3.245 3.615 3.415 3.785 ;
        RECT 3.985 2.880 4.155 3.050 ;
        RECT 8.050 3.985 8.220 4.155 ;
        RECT 5.835 2.880 6.005 3.050 ;
        RECT 8.795 3.615 8.965 3.785 ;
        RECT 10.645 2.880 10.815 3.050 ;
        RECT 12.865 3.985 13.035 4.155 ;
        RECT 13.605 2.875 13.775 3.045 ;
        RECT 15.455 2.875 15.625 3.045 ;
        RECT 18.415 3.985 18.585 4.155 ;
        RECT 20.265 3.615 20.435 3.785 ;
        RECT 22.485 3.245 22.655 3.415 ;
        RECT 23.225 3.615 23.395 3.785 ;
        RECT 25.075 3.615 25.245 3.785 ;
        RECT 27.295 3.985 27.465 4.155 ;
        RECT 28.035 3.245 28.205 3.415 ;
        RECT 32.105 3.615 32.275 3.785 ;
        RECT 32.845 2.880 33.015 3.050 ;
        RECT 36.910 3.985 37.080 4.155 ;
        RECT 34.695 2.880 34.865 3.050 ;
        RECT 37.655 3.615 37.825 3.785 ;
        RECT 39.505 2.880 39.675 3.050 ;
        RECT 41.725 3.985 41.895 4.155 ;
        RECT 42.465 2.875 42.635 3.045 ;
        RECT 44.315 2.875 44.485 3.045 ;
        RECT 47.275 3.985 47.445 4.155 ;
        RECT 49.125 3.615 49.295 3.785 ;
        RECT 51.345 2.875 51.515 3.045 ;
        RECT 52.085 3.615 52.255 3.785 ;
        RECT 53.935 3.615 54.105 3.785 ;
        RECT 56.155 3.985 56.325 4.155 ;
        RECT 56.895 3.985 57.065 4.155 ;
        RECT 56.895 2.875 57.065 3.045 ;
        RECT 60.965 3.615 61.135 3.785 ;
        RECT 61.705 2.880 61.875 3.050 ;
        RECT 65.770 3.985 65.940 4.155 ;
        RECT 63.555 2.880 63.725 3.050 ;
        RECT 66.515 3.615 66.685 3.785 ;
        RECT 68.365 2.880 68.535 3.050 ;
        RECT 70.585 3.985 70.755 4.155 ;
        RECT 71.325 2.875 71.495 3.045 ;
        RECT 73.175 2.875 73.345 3.045 ;
        RECT 76.135 3.985 76.305 4.155 ;
        RECT 77.985 3.615 78.155 3.785 ;
        RECT 80.205 2.875 80.375 3.045 ;
        RECT 80.945 3.615 81.115 3.785 ;
        RECT 82.795 3.615 82.965 3.785 ;
        RECT 85.015 3.985 85.185 4.155 ;
        RECT 90.605 5.355 90.775 5.525 ;
        RECT 91.925 5.355 92.095 5.525 ;
        RECT 93.945 5.355 94.115 5.525 ;
        RECT 85.755 3.985 85.925 4.155 ;
        RECT 85.755 2.875 85.925 3.045 ;
        RECT 87.235 4.725 87.405 4.895 ;
        RECT 87.235 3.985 87.405 4.155 ;
        RECT 88.345 4.355 88.515 4.525 ;
        RECT 90.935 4.725 91.105 4.895 ;
        RECT 92.415 3.245 92.585 3.415 ;
        RECT 92.415 2.135 92.585 2.305 ;
        RECT 93.895 2.135 94.065 2.305 ;
        RECT 95.005 4.355 95.175 4.525 ;
        RECT 95.745 3.985 95.915 4.155 ;
        RECT 88.645 1.235 88.815 1.405 ;
        RECT 91.975 1.235 92.145 1.405 ;
        RECT 97.225 3.985 97.395 4.155 ;
        RECT 95.305 1.235 95.475 1.405 ;
      LAYER met1 ;
        RECT 88.575 5.525 88.805 5.555 ;
        RECT 90.575 5.525 90.805 5.555 ;
        RECT 91.895 5.525 92.125 5.555 ;
        RECT 93.915 5.525 94.145 5.555 ;
        RECT 88.545 5.355 90.835 5.525 ;
        RECT 91.865 5.355 94.175 5.525 ;
        RECT 88.575 5.325 88.805 5.355 ;
        RECT 90.575 5.325 90.805 5.355 ;
        RECT 91.895 5.325 92.125 5.355 ;
        RECT 93.915 5.325 94.145 5.355 ;
        RECT 87.205 4.895 87.435 4.925 ;
        RECT 90.905 4.895 91.135 4.925 ;
        RECT 87.175 4.725 91.165 4.895 ;
        RECT 87.205 4.695 87.435 4.725 ;
        RECT 90.905 4.695 91.135 4.725 ;
        RECT 88.315 4.525 88.545 4.555 ;
        RECT 94.975 4.525 95.205 4.555 ;
        RECT 59.855 4.355 95.235 4.525 ;
        RECT 8.020 4.155 8.250 4.185 ;
        RECT 12.835 4.155 13.065 4.185 ;
        RECT 18.385 4.155 18.615 4.185 ;
        RECT 27.265 4.155 27.495 4.185 ;
        RECT 36.880 4.155 37.110 4.185 ;
        RECT 41.695 4.155 41.925 4.185 ;
        RECT 47.245 4.155 47.475 4.185 ;
        RECT 56.125 4.155 56.355 4.185 ;
        RECT 56.865 4.155 57.095 4.185 ;
        RECT 59.855 4.155 60.025 4.355 ;
        RECT 88.315 4.325 88.545 4.355 ;
        RECT 94.975 4.325 95.205 4.355 ;
        RECT 65.740 4.155 65.970 4.185 ;
        RECT 70.555 4.155 70.785 4.185 ;
        RECT 76.105 4.155 76.335 4.185 ;
        RECT 84.985 4.155 85.215 4.185 ;
        RECT 85.725 4.155 85.955 4.185 ;
        RECT 87.205 4.155 87.435 4.185 ;
        RECT 95.715 4.155 95.945 4.185 ;
        RECT 97.195 4.155 97.425 4.185 ;
        RECT 7.990 3.985 27.525 4.155 ;
        RECT 36.850 3.985 56.385 4.155 ;
        RECT 56.835 3.985 60.025 4.155 ;
        RECT 65.710 3.985 85.245 4.155 ;
        RECT 85.695 3.985 87.465 4.155 ;
        RECT 95.685 3.985 97.455 4.155 ;
        RECT 8.020 3.955 8.250 3.985 ;
        RECT 12.835 3.955 13.065 3.985 ;
        RECT 18.385 3.955 18.615 3.985 ;
        RECT 27.265 3.955 27.495 3.985 ;
        RECT 36.880 3.955 37.110 3.985 ;
        RECT 41.695 3.955 41.925 3.985 ;
        RECT 47.245 3.955 47.475 3.985 ;
        RECT 56.125 3.955 56.355 3.985 ;
        RECT 56.865 3.955 57.095 3.985 ;
        RECT 65.740 3.955 65.970 3.985 ;
        RECT 70.555 3.955 70.785 3.985 ;
        RECT 76.105 3.955 76.335 3.985 ;
        RECT 84.985 3.955 85.215 3.985 ;
        RECT 85.725 3.955 85.955 3.985 ;
        RECT 87.205 3.955 87.435 3.985 ;
        RECT 95.715 3.955 95.945 3.985 ;
        RECT 97.195 3.955 97.425 3.985 ;
        RECT 3.215 3.785 3.445 3.815 ;
        RECT 8.765 3.785 8.995 3.815 ;
        RECT 20.235 3.785 20.465 3.815 ;
        RECT 23.195 3.785 23.425 3.815 ;
        RECT 25.045 3.785 25.275 3.815 ;
        RECT 32.075 3.785 32.305 3.815 ;
        RECT 37.625 3.785 37.855 3.815 ;
        RECT 49.095 3.785 49.325 3.815 ;
        RECT 52.055 3.785 52.285 3.815 ;
        RECT 53.905 3.785 54.135 3.815 ;
        RECT 60.935 3.785 61.165 3.815 ;
        RECT 66.485 3.785 66.715 3.815 ;
        RECT 77.955 3.785 78.185 3.815 ;
        RECT 80.915 3.785 81.145 3.815 ;
        RECT 82.765 3.785 82.995 3.815 ;
        RECT 3.185 3.615 20.495 3.785 ;
        RECT 23.165 3.615 25.305 3.785 ;
        RECT 32.045 3.615 49.355 3.785 ;
        RECT 52.025 3.615 54.165 3.785 ;
        RECT 60.905 3.615 78.215 3.785 ;
        RECT 80.885 3.615 83.025 3.785 ;
        RECT 3.215 3.585 3.445 3.615 ;
        RECT 8.765 3.585 8.995 3.615 ;
        RECT 20.235 3.585 20.465 3.615 ;
        RECT 23.195 3.585 23.425 3.615 ;
        RECT 25.045 3.585 25.275 3.615 ;
        RECT 32.075 3.585 32.305 3.615 ;
        RECT 37.625 3.585 37.855 3.615 ;
        RECT 49.095 3.585 49.325 3.615 ;
        RECT 52.055 3.585 52.285 3.615 ;
        RECT 53.905 3.585 54.135 3.615 ;
        RECT 60.935 3.585 61.165 3.615 ;
        RECT 66.485 3.585 66.715 3.615 ;
        RECT 77.955 3.585 78.185 3.615 ;
        RECT 80.915 3.585 81.145 3.615 ;
        RECT 82.765 3.585 82.995 3.615 ;
        RECT 22.455 3.415 22.685 3.445 ;
        RECT 28.005 3.415 28.235 3.445 ;
        RECT 92.385 3.415 92.615 3.445 ;
        RECT 22.425 3.245 92.645 3.415 ;
        RECT 22.455 3.215 22.685 3.245 ;
        RECT 28.005 3.215 28.235 3.245 ;
        RECT 92.385 3.215 92.615 3.245 ;
        RECT 3.955 3.050 4.185 3.080 ;
        RECT 5.805 3.050 6.035 3.080 ;
        RECT 10.615 3.050 10.845 3.080 ;
        RECT 3.925 2.880 10.875 3.050 ;
        RECT 13.575 3.045 13.805 3.075 ;
        RECT 15.425 3.045 15.655 3.075 ;
        RECT 32.815 3.050 33.045 3.080 ;
        RECT 34.665 3.050 34.895 3.080 ;
        RECT 39.475 3.050 39.705 3.080 ;
        RECT 3.955 2.850 4.185 2.880 ;
        RECT 5.805 2.850 6.035 2.880 ;
        RECT 10.615 2.850 10.845 2.880 ;
        RECT 13.545 2.875 15.685 3.045 ;
        RECT 32.785 2.880 39.735 3.050 ;
        RECT 42.435 3.045 42.665 3.075 ;
        RECT 44.285 3.045 44.515 3.075 ;
        RECT 51.315 3.045 51.545 3.075 ;
        RECT 56.865 3.045 57.095 3.075 ;
        RECT 61.675 3.050 61.905 3.080 ;
        RECT 63.525 3.050 63.755 3.080 ;
        RECT 68.335 3.050 68.565 3.080 ;
        RECT 13.575 2.845 13.805 2.875 ;
        RECT 15.425 2.845 15.655 2.875 ;
        RECT 32.815 2.850 33.045 2.880 ;
        RECT 34.665 2.850 34.895 2.880 ;
        RECT 39.475 2.850 39.705 2.880 ;
        RECT 42.405 2.875 44.545 3.045 ;
        RECT 51.285 2.875 57.125 3.045 ;
        RECT 61.645 2.880 68.595 3.050 ;
        RECT 71.295 3.045 71.525 3.075 ;
        RECT 73.145 3.045 73.375 3.075 ;
        RECT 80.175 3.045 80.405 3.075 ;
        RECT 85.725 3.045 85.955 3.075 ;
        RECT 42.435 2.845 42.665 2.875 ;
        RECT 44.285 2.845 44.515 2.875 ;
        RECT 51.315 2.845 51.545 2.875 ;
        RECT 56.865 2.845 57.095 2.875 ;
        RECT 61.675 2.850 61.905 2.880 ;
        RECT 63.525 2.850 63.755 2.880 ;
        RECT 68.335 2.850 68.565 2.880 ;
        RECT 71.265 2.875 73.405 3.045 ;
        RECT 80.145 2.875 85.985 3.045 ;
        RECT 71.295 2.845 71.525 2.875 ;
        RECT 73.145 2.845 73.375 2.875 ;
        RECT 80.175 2.845 80.405 2.875 ;
        RECT 85.725 2.845 85.955 2.875 ;
        RECT 92.385 2.305 92.615 2.335 ;
        RECT 93.865 2.305 94.095 2.335 ;
        RECT 92.355 2.135 94.125 2.305 ;
        RECT 92.385 2.105 92.615 2.135 ;
        RECT 93.865 2.105 94.095 2.135 ;
        RECT 88.615 1.405 88.845 1.435 ;
        RECT 91.945 1.405 92.175 1.435 ;
        RECT 95.275 1.405 95.505 1.435 ;
        RECT 88.585 1.235 95.535 1.405 ;
        RECT 88.615 1.205 88.845 1.235 ;
        RECT 91.945 1.205 92.175 1.235 ;
        RECT 95.275 1.205 95.505 1.235 ;
  END
END TMRDFFSNRNQX1






MACRO VOTER3X1
  CLASS BLOCK ;
  FOREIGN VOTER3X1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 13.050 BY 7.950 ;
  PIN Y
    ANTENNADIFFAREA 0.771900 ;
    PORT
      LAYER li1 ;
        RECT 11.015 4.895 11.185 7.250 ;
        RECT 11.015 4.725 11.555 4.895 ;
        RECT 11.385 2.305 11.555 4.725 ;
        RECT 11.015 2.135 11.555 2.305 ;
        RECT 11.015 0.975 11.185 2.135 ;
      LAYER mcon ;
        RECT 11.385 3.990 11.555 4.160 ;
      LAYER met1 ;
        RECT 11.355 4.160 11.585 4.190 ;
        RECT 11.325 3.990 11.735 4.160 ;
        RECT 11.355 3.960 11.585 3.990 ;
    END
  END Y
  PIN A
    ANTENNAGATEAREA 2.053700 ;
    PORT
      LAYER li1 ;
        RECT 1.805 4.940 1.975 5.100 ;
        RECT 1.765 4.770 1.975 4.940 ;
        RECT 8.425 4.770 8.615 5.100 ;
        RECT 1.765 2.055 1.935 4.770 ;
        RECT 8.425 2.055 8.595 4.770 ;
      LAYER mcon ;
        RECT 1.765 4.355 1.935 4.525 ;
        RECT 8.425 4.355 8.595 4.525 ;
      LAYER met1 ;
        RECT 1.735 4.525 1.965 4.555 ;
        RECT 8.395 4.525 8.625 4.555 ;
        RECT 1.705 4.355 8.655 4.525 ;
        RECT 1.735 4.325 1.965 4.355 ;
        RECT 8.395 4.325 8.625 4.355 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 2.066500 ;
    PORT
      LAYER li1 ;
        RECT 0.655 2.055 0.825 5.100 ;
        RECT 4.355 2.055 4.525 5.100 ;
      LAYER mcon ;
        RECT 0.655 4.725 0.825 4.895 ;
        RECT 4.355 4.725 4.525 4.895 ;
      LAYER met1 ;
        RECT 0.625 4.895 0.855 4.925 ;
        RECT 4.325 4.895 4.555 4.925 ;
        RECT 0.595 4.725 4.585 4.895 ;
        RECT 0.625 4.695 0.855 4.725 ;
        RECT 4.325 4.695 4.555 4.725 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA 2.060500 ;
    PORT
      LAYER li1 ;
        RECT 5.835 2.055 6.005 5.100 ;
        RECT 7.315 2.055 7.485 5.100 ;
      LAYER mcon ;
        RECT 5.835 2.135 6.005 2.305 ;
        RECT 7.315 2.135 7.485 2.305 ;
      LAYER met1 ;
        RECT 5.805 2.305 6.035 2.335 ;
        RECT 7.285 2.305 7.515 2.335 ;
        RECT 5.775 2.135 7.545 2.305 ;
        RECT 5.805 2.105 6.035 2.135 ;
        RECT 7.285 2.105 7.515 2.135 ;
    END
  END C
  PIN VDD
    ANTENNADIFFAREA 13.245850 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 12.630 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 12.365 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 0.705 5.355 0.875 7.460 ;
        RECT 1.585 5.785 1.755 7.460 ;
        RECT 2.465 5.355 2.635 7.460 ;
        RECT 3.175 4.340 3.485 7.460 ;
        RECT 6.505 4.340 6.815 7.460 ;
        RECT 9.835 4.340 10.145 7.460 ;
        RECT 10.575 5.415 10.745 7.460 ;
        RECT 11.455 5.415 11.625 7.460 ;
        RECT 12.055 4.340 12.365 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 0.995 7.525 1.165 7.695 ;
        RECT 1.355 7.525 1.525 7.695 ;
        RECT 1.805 7.525 1.975 7.695 ;
        RECT 2.165 7.525 2.335 7.695 ;
        RECT 2.525 7.525 2.695 7.695 ;
        RECT 2.885 7.525 3.055 7.695 ;
        RECT 3.605 7.525 3.775 7.695 ;
        RECT 3.965 7.525 4.135 7.695 ;
        RECT 4.325 7.525 4.495 7.695 ;
        RECT 4.685 7.525 4.855 7.695 ;
        RECT 5.135 7.525 5.305 7.695 ;
        RECT 5.495 7.525 5.665 7.695 ;
        RECT 5.855 7.525 6.025 7.695 ;
        RECT 6.215 7.525 6.385 7.695 ;
        RECT 6.935 7.525 7.105 7.695 ;
        RECT 7.295 7.525 7.465 7.695 ;
        RECT 7.655 7.525 7.825 7.695 ;
        RECT 8.015 7.525 8.185 7.695 ;
        RECT 8.465 7.525 8.635 7.695 ;
        RECT 8.825 7.525 8.995 7.695 ;
        RECT 9.185 7.525 9.355 7.695 ;
        RECT 9.545 7.525 9.715 7.695 ;
        RECT 10.265 7.525 10.435 7.695 ;
        RECT 10.625 7.525 10.795 7.695 ;
        RECT 11.015 7.525 11.185 7.695 ;
        RECT 11.405 7.525 11.575 7.695 ;
        RECT 11.765 7.525 11.935 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 12.365 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 11.366799 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 12.495 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 3.045 -0.075 3.615 -0.065 ;
        RECT 6.375 -0.075 6.945 -0.065 ;
        RECT 9.705 -0.075 10.275 -0.065 ;
        RECT 11.925 -0.075 12.495 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 1.095 0.310 1.265 1.260 ;
        RECT 3.175 0.310 3.485 2.860 ;
        RECT 4.425 0.310 4.595 1.260 ;
        RECT 6.505 0.310 6.815 2.860 ;
        RECT 7.755 0.310 7.925 1.260 ;
        RECT 9.835 0.310 10.145 2.860 ;
        RECT 10.535 0.755 10.705 1.885 ;
        RECT 11.505 0.755 11.675 1.885 ;
        RECT 10.535 0.585 11.675 0.755 ;
        RECT 10.535 0.310 10.705 0.585 ;
        RECT 11.020 0.310 11.190 0.585 ;
        RECT 11.505 0.310 11.675 0.585 ;
        RECT 12.055 0.310 12.365 2.860 ;
        RECT -0.155 0.235 5.395 0.310 ;
        RECT 5.565 0.235 12.365 0.310 ;
        RECT -0.155 0.000 12.365 0.235 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 0.995 0.065 1.165 0.235 ;
        RECT 1.355 0.065 1.525 0.235 ;
        RECT 1.805 0.065 1.975 0.235 ;
        RECT 2.165 0.065 2.335 0.235 ;
        RECT 2.525 0.065 2.695 0.235 ;
        RECT 2.885 0.065 3.055 0.235 ;
        RECT 3.605 0.065 3.775 0.235 ;
        RECT 3.965 0.065 4.135 0.235 ;
        RECT 4.325 0.065 4.495 0.235 ;
        RECT 4.685 0.065 4.855 0.235 ;
        RECT 5.135 0.065 5.305 0.235 ;
        RECT 5.495 0.065 5.665 0.235 ;
        RECT 5.855 0.065 6.025 0.235 ;
        RECT 6.215 0.065 6.385 0.235 ;
        RECT 6.935 0.065 7.105 0.235 ;
        RECT 7.295 0.065 7.465 0.235 ;
        RECT 7.655 0.065 7.825 0.235 ;
        RECT 8.015 0.065 8.185 0.235 ;
        RECT 8.465 0.065 8.635 0.235 ;
        RECT 8.825 0.065 8.995 0.235 ;
        RECT 9.185 0.065 9.355 0.235 ;
        RECT 9.545 0.065 9.715 0.235 ;
        RECT 10.265 0.065 10.435 0.235 ;
        RECT 10.625 0.065 10.795 0.235 ;
        RECT 11.015 0.065 11.185 0.235 ;
        RECT 11.405 0.065 11.575 0.235 ;
        RECT 11.765 0.065 11.935 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 12.365 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 1.145 7.055 1.325 7.225 ;
        RECT 1.145 5.525 1.315 7.055 ;
        RECT 2.025 5.525 2.195 7.225 ;
        RECT 1.145 5.355 2.195 5.525 ;
        RECT 2.025 5.275 2.195 5.355 ;
        RECT 4.025 7.055 5.955 7.225 ;
        RECT 4.025 5.275 4.195 7.055 ;
        RECT 4.465 5.525 4.635 6.795 ;
        RECT 4.905 5.785 5.075 7.055 ;
        RECT 5.345 5.525 5.515 6.795 ;
        RECT 5.785 5.605 5.955 7.055 ;
        RECT 7.365 7.055 9.295 7.225 ;
        RECT 4.465 5.355 5.515 5.525 ;
        RECT 5.345 5.275 5.515 5.355 ;
        RECT 7.365 5.275 7.535 7.055 ;
        RECT 7.805 5.525 7.975 6.795 ;
        RECT 8.245 5.785 8.415 7.055 ;
        RECT 8.685 5.525 8.855 6.795 ;
        RECT 9.125 5.785 9.295 7.055 ;
        RECT 7.805 5.355 9.335 5.525 ;
        RECT 0.610 1.805 0.780 1.885 ;
        RECT 1.580 1.805 1.750 1.885 ;
        RECT 0.610 1.635 1.750 1.805 ;
        RECT 0.610 0.505 0.780 1.635 ;
        RECT 1.580 0.755 1.750 1.635 ;
        RECT 2.065 1.310 2.235 1.485 ;
        RECT 2.060 1.155 2.235 1.310 ;
        RECT 2.060 0.975 2.230 1.155 ;
        RECT 2.550 0.755 2.720 1.885 ;
        RECT 1.580 0.585 2.720 0.755 ;
        RECT 1.580 0.505 1.750 0.585 ;
        RECT 2.550 0.505 2.720 0.585 ;
        RECT 3.940 1.805 4.110 1.885 ;
        RECT 4.910 1.805 5.080 1.885 ;
        RECT 3.940 1.635 5.080 1.805 ;
        RECT 3.940 0.505 4.110 1.635 ;
        RECT 4.910 0.755 5.080 1.635 ;
        RECT 5.395 0.975 5.565 1.485 ;
        RECT 5.880 0.755 6.050 1.885 ;
        RECT 4.910 0.585 6.050 0.755 ;
        RECT 4.910 0.505 5.080 0.585 ;
        RECT 5.880 0.505 6.050 0.585 ;
        RECT 7.270 1.805 7.440 1.885 ;
        RECT 8.240 1.805 8.410 1.885 ;
        RECT 9.165 1.870 9.335 5.355 ;
        RECT 10.645 2.055 10.815 5.095 ;
        RECT 7.270 1.635 8.410 1.805 ;
        RECT 7.270 0.505 7.440 1.635 ;
        RECT 8.240 0.755 8.410 1.635 ;
        RECT 8.725 1.700 9.335 1.870 ;
        RECT 8.725 0.975 8.895 1.700 ;
        RECT 9.210 0.755 9.380 1.530 ;
        RECT 8.240 0.585 9.380 0.755 ;
        RECT 8.240 0.505 8.410 0.585 ;
        RECT 9.210 0.505 9.380 0.585 ;
      LAYER mcon ;
        RECT 2.025 5.355 2.195 5.525 ;
        RECT 4.025 5.355 4.195 5.525 ;
        RECT 5.345 5.355 5.515 5.525 ;
        RECT 7.365 5.355 7.535 5.525 ;
        RECT 9.165 3.985 9.335 4.155 ;
        RECT 2.065 1.235 2.235 1.405 ;
        RECT 5.395 1.235 5.565 1.405 ;
        RECT 10.645 3.985 10.815 4.155 ;
        RECT 8.725 1.235 8.895 1.405 ;
      LAYER met1 ;
        RECT 1.995 5.525 2.225 5.555 ;
        RECT 3.995 5.525 4.225 5.555 ;
        RECT 5.315 5.525 5.545 5.555 ;
        RECT 7.335 5.525 7.565 5.555 ;
        RECT 1.965 5.355 4.255 5.525 ;
        RECT 5.285 5.355 7.595 5.525 ;
        RECT 1.995 5.325 2.225 5.355 ;
        RECT 3.995 5.325 4.225 5.355 ;
        RECT 5.315 5.325 5.545 5.355 ;
        RECT 7.335 5.325 7.565 5.355 ;
        RECT 9.135 4.155 9.365 4.185 ;
        RECT 10.615 4.155 10.845 4.185 ;
        RECT 9.105 3.985 10.875 4.155 ;
        RECT 9.135 3.955 9.365 3.985 ;
        RECT 10.615 3.955 10.845 3.985 ;
        RECT 2.035 1.405 2.265 1.435 ;
        RECT 5.365 1.405 5.595 1.435 ;
        RECT 8.695 1.405 8.925 1.435 ;
        RECT 2.005 1.235 8.955 1.405 ;
        RECT 2.035 1.205 2.265 1.235 ;
        RECT 5.365 1.205 5.595 1.235 ;
        RECT 8.695 1.205 8.925 1.235 ;
  END
END VOTER3X1






MACRO VOTERN3X1
  CLASS BLOCK ;
  FOREIGN VOTERN3X1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 10.830 BY 7.950 ;
  PIN YN
    ANTENNADIFFAREA 1.734950 ;
    PORT
      LAYER li1 ;
        RECT 7.805 5.525 7.975 6.795 ;
        RECT 8.685 5.525 8.855 6.795 ;
        RECT 7.805 5.355 9.335 5.525 ;
        RECT 9.165 1.870 9.335 5.355 ;
        RECT 8.725 1.700 9.335 1.870 ;
        RECT 2.065 1.310 2.235 1.485 ;
        RECT 2.060 1.155 2.235 1.310 ;
        RECT 2.060 0.975 2.230 1.155 ;
        RECT 5.395 0.975 5.565 1.485 ;
        RECT 8.725 0.975 8.895 1.700 ;
      LAYER mcon ;
        RECT 9.165 3.985 9.335 4.155 ;
        RECT 2.065 1.235 2.235 1.405 ;
        RECT 5.395 1.235 5.565 1.405 ;
        RECT 8.725 1.235 8.895 1.405 ;
      LAYER met1 ;
        RECT 9.135 4.155 9.365 4.185 ;
        RECT 9.105 3.985 9.515 4.155 ;
        RECT 9.135 3.955 9.365 3.985 ;
        RECT 2.035 1.405 2.265 1.435 ;
        RECT 5.365 1.405 5.595 1.435 ;
        RECT 8.695 1.405 8.925 1.435 ;
        RECT 2.005 1.235 8.955 1.405 ;
        RECT 2.035 1.205 2.265 1.235 ;
        RECT 5.365 1.205 5.595 1.235 ;
        RECT 8.695 1.205 8.925 1.235 ;
    END
  END YN
  PIN A
    ANTENNAGATEAREA 2.053700 ;
    PORT
      LAYER li1 ;
        RECT 1.805 4.940 1.975 5.100 ;
        RECT 1.765 4.770 1.975 4.940 ;
        RECT 8.425 4.770 8.615 5.100 ;
        RECT 1.765 2.055 1.935 4.770 ;
        RECT 8.425 2.055 8.595 4.770 ;
      LAYER mcon ;
        RECT 1.765 4.355 1.935 4.525 ;
        RECT 8.425 4.355 8.595 4.525 ;
      LAYER met1 ;
        RECT 1.735 4.525 1.965 4.555 ;
        RECT 8.395 4.525 8.625 4.555 ;
        RECT 1.705 4.355 8.655 4.525 ;
        RECT 1.735 4.325 1.965 4.355 ;
        RECT 8.395 4.325 8.625 4.355 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 2.066500 ;
    PORT
      LAYER li1 ;
        RECT 0.655 2.055 0.825 5.100 ;
        RECT 4.355 2.055 4.525 5.100 ;
      LAYER mcon ;
        RECT 0.655 4.725 0.825 4.895 ;
        RECT 4.355 4.725 4.525 4.895 ;
      LAYER met1 ;
        RECT 0.625 4.895 0.855 4.925 ;
        RECT 4.325 4.895 4.555 4.925 ;
        RECT 0.595 4.725 4.585 4.895 ;
        RECT 0.625 4.695 0.855 4.725 ;
        RECT 4.325 4.695 4.555 4.725 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA 2.060500 ;
    PORT
      LAYER li1 ;
        RECT 5.835 2.055 6.005 5.100 ;
        RECT 7.315 2.055 7.485 5.100 ;
      LAYER mcon ;
        RECT 5.835 2.135 6.005 2.305 ;
        RECT 7.315 2.135 7.485 2.305 ;
      LAYER met1 ;
        RECT 5.805 2.305 6.035 2.335 ;
        RECT 7.285 2.305 7.515 2.335 ;
        RECT 5.775 2.135 7.545 2.305 ;
        RECT 5.805 2.105 6.035 2.135 ;
        RECT 7.285 2.105 7.515 2.135 ;
    END
  END C
  PIN VDD
    ANTENNADIFFAREA 10.189000 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 10.410 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 10.145 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 0.705 5.355 0.875 7.460 ;
        RECT 1.585 5.785 1.755 7.460 ;
        RECT 2.465 5.355 2.635 7.460 ;
        RECT 3.175 4.340 3.485 7.460 ;
        RECT 6.505 4.340 6.815 7.460 ;
        RECT 9.835 4.340 10.145 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 0.995 7.525 1.165 7.695 ;
        RECT 1.355 7.525 1.525 7.695 ;
        RECT 1.805 7.525 1.975 7.695 ;
        RECT 2.165 7.525 2.335 7.695 ;
        RECT 2.525 7.525 2.695 7.695 ;
        RECT 2.885 7.525 3.055 7.695 ;
        RECT 3.605 7.525 3.775 7.695 ;
        RECT 3.965 7.525 4.135 7.695 ;
        RECT 4.325 7.525 4.495 7.695 ;
        RECT 4.685 7.525 4.855 7.695 ;
        RECT 5.135 7.525 5.305 7.695 ;
        RECT 5.495 7.525 5.665 7.695 ;
        RECT 5.855 7.525 6.025 7.695 ;
        RECT 6.215 7.525 6.385 7.695 ;
        RECT 6.935 7.525 7.105 7.695 ;
        RECT 7.295 7.525 7.465 7.695 ;
        RECT 7.655 7.525 7.825 7.695 ;
        RECT 8.015 7.525 8.185 7.695 ;
        RECT 8.465 7.525 8.635 7.695 ;
        RECT 8.825 7.525 8.995 7.695 ;
        RECT 9.185 7.525 9.355 7.695 ;
        RECT 9.545 7.525 9.715 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 10.145 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 8.402699 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 10.275 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 3.045 -0.075 3.615 -0.065 ;
        RECT 6.375 -0.075 6.945 -0.065 ;
        RECT 9.705 -0.075 10.275 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 1.095 0.310 1.265 1.260 ;
        RECT 3.175 0.310 3.485 2.860 ;
        RECT 4.425 0.310 4.595 1.260 ;
        RECT 6.505 0.310 6.815 2.860 ;
        RECT 7.755 0.310 7.925 1.260 ;
        RECT 9.835 0.310 10.145 2.860 ;
        RECT -0.155 0.235 5.395 0.310 ;
        RECT 5.565 0.235 10.145 0.310 ;
        RECT -0.155 0.000 10.145 0.235 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 0.995 0.065 1.165 0.235 ;
        RECT 1.355 0.065 1.525 0.235 ;
        RECT 1.805 0.065 1.975 0.235 ;
        RECT 2.165 0.065 2.335 0.235 ;
        RECT 2.525 0.065 2.695 0.235 ;
        RECT 2.885 0.065 3.055 0.235 ;
        RECT 3.605 0.065 3.775 0.235 ;
        RECT 3.965 0.065 4.135 0.235 ;
        RECT 4.325 0.065 4.495 0.235 ;
        RECT 4.685 0.065 4.855 0.235 ;
        RECT 5.135 0.065 5.305 0.235 ;
        RECT 5.495 0.065 5.665 0.235 ;
        RECT 5.855 0.065 6.025 0.235 ;
        RECT 6.215 0.065 6.385 0.235 ;
        RECT 6.935 0.065 7.105 0.235 ;
        RECT 7.295 0.065 7.465 0.235 ;
        RECT 7.655 0.065 7.825 0.235 ;
        RECT 8.015 0.065 8.185 0.235 ;
        RECT 8.465 0.065 8.635 0.235 ;
        RECT 8.825 0.065 8.995 0.235 ;
        RECT 9.185 0.065 9.355 0.235 ;
        RECT 9.545 0.065 9.715 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 10.145 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 1.145 7.055 1.325 7.225 ;
        RECT 1.145 5.525 1.315 7.055 ;
        RECT 2.025 5.525 2.195 7.225 ;
        RECT 1.145 5.355 2.195 5.525 ;
        RECT 2.025 5.275 2.195 5.355 ;
        RECT 4.025 7.055 5.955 7.225 ;
        RECT 4.025 5.275 4.195 7.055 ;
        RECT 4.465 5.525 4.635 6.795 ;
        RECT 4.905 5.785 5.075 7.055 ;
        RECT 5.345 5.525 5.515 6.795 ;
        RECT 5.785 5.605 5.955 7.055 ;
        RECT 7.365 7.055 9.295 7.225 ;
        RECT 4.465 5.355 5.515 5.525 ;
        RECT 5.345 5.275 5.515 5.355 ;
        RECT 7.365 5.275 7.535 7.055 ;
        RECT 8.245 5.785 8.415 7.055 ;
        RECT 9.125 5.785 9.295 7.055 ;
        RECT 0.610 1.805 0.780 1.885 ;
        RECT 1.580 1.805 1.750 1.885 ;
        RECT 0.610 1.635 1.750 1.805 ;
        RECT 0.610 0.505 0.780 1.635 ;
        RECT 1.580 0.755 1.750 1.635 ;
        RECT 2.550 0.755 2.720 1.885 ;
        RECT 1.580 0.585 2.720 0.755 ;
        RECT 1.580 0.505 1.750 0.585 ;
        RECT 2.550 0.505 2.720 0.585 ;
        RECT 3.940 1.805 4.110 1.885 ;
        RECT 4.910 1.805 5.080 1.885 ;
        RECT 3.940 1.635 5.080 1.805 ;
        RECT 3.940 0.505 4.110 1.635 ;
        RECT 4.910 0.755 5.080 1.635 ;
        RECT 5.880 0.755 6.050 1.885 ;
        RECT 4.910 0.585 6.050 0.755 ;
        RECT 4.910 0.505 5.080 0.585 ;
        RECT 5.880 0.505 6.050 0.585 ;
        RECT 7.270 1.805 7.440 1.885 ;
        RECT 8.240 1.805 8.410 1.885 ;
        RECT 7.270 1.635 8.410 1.805 ;
        RECT 7.270 0.505 7.440 1.635 ;
        RECT 8.240 0.755 8.410 1.635 ;
        RECT 9.210 0.755 9.380 1.530 ;
        RECT 8.240 0.585 9.380 0.755 ;
        RECT 8.240 0.505 8.410 0.585 ;
        RECT 9.210 0.505 9.380 0.585 ;
      LAYER mcon ;
        RECT 2.025 5.355 2.195 5.525 ;
        RECT 4.025 5.355 4.195 5.525 ;
        RECT 5.345 5.355 5.515 5.525 ;
        RECT 7.365 5.355 7.535 5.525 ;
      LAYER met1 ;
        RECT 1.995 5.525 2.225 5.555 ;
        RECT 3.995 5.525 4.225 5.555 ;
        RECT 5.315 5.525 5.545 5.555 ;
        RECT 7.335 5.525 7.565 5.555 ;
        RECT 1.965 5.355 4.255 5.525 ;
        RECT 5.285 5.355 7.595 5.525 ;
        RECT 1.995 5.325 2.225 5.355 ;
        RECT 3.995 5.325 4.225 5.355 ;
        RECT 5.315 5.325 5.545 5.355 ;
        RECT 7.335 5.325 7.565 5.355 ;
  END
END VOTERN3X1






MACRO XNOR2X1
  CLASS BLOCK ;
  FOREIGN XNOR2X1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 11.940 BY 7.950 ;
  PIN Y
    ANTENNADIFFAREA 1.543800 ;
    PORT
      LAYER li1 ;
        RECT 4.245 5.525 4.415 6.795 ;
        RECT 7.575 5.525 7.745 6.795 ;
        RECT 4.245 5.355 4.895 5.525 ;
        RECT 7.575 5.355 8.225 5.525 ;
        RECT 4.725 1.875 4.895 5.355 ;
        RECT 8.055 1.875 8.225 5.355 ;
        RECT 4.285 1.705 4.895 1.875 ;
        RECT 7.615 1.705 8.225 1.875 ;
        RECT 4.285 0.975 4.455 1.705 ;
        RECT 7.615 0.975 7.785 1.705 ;
      LAYER mcon ;
        RECT 4.725 3.615 4.895 3.785 ;
        RECT 8.055 3.615 8.225 3.785 ;
      LAYER met1 ;
        RECT 4.695 3.785 4.925 3.815 ;
        RECT 8.025 3.785 8.255 3.815 ;
        RECT 4.665 3.615 8.285 3.785 ;
        RECT 4.695 3.585 4.925 3.615 ;
        RECT 8.025 3.585 8.255 3.615 ;
    END
  END Y
  PIN A
    ANTENNAGATEAREA 2.060500 ;
    PORT
      LAYER li1 ;
        RECT 0.655 2.055 0.825 5.095 ;
        RECT 3.245 2.055 3.415 5.100 ;
      LAYER mcon ;
        RECT 0.655 4.355 0.825 4.525 ;
        RECT 3.245 4.355 3.415 4.525 ;
      LAYER met1 ;
        RECT 0.625 4.525 0.855 4.555 ;
        RECT 3.215 4.525 3.445 4.555 ;
        RECT 0.595 4.355 3.475 4.525 ;
        RECT 0.625 4.325 0.855 4.355 ;
        RECT 3.215 4.325 3.445 4.355 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 2.060500 ;
    PORT
      LAYER li1 ;
        RECT 4.355 3.905 4.525 5.100 ;
        RECT 6.575 2.055 6.745 3.495 ;
        RECT 10.275 2.055 10.445 5.095 ;
      LAYER mcon ;
        RECT 4.355 3.985 4.525 4.155 ;
        RECT 10.275 3.985 10.445 4.155 ;
        RECT 6.575 3.245 6.745 3.415 ;
        RECT 10.275 3.245 10.445 3.415 ;
        RECT 10.275 2.875 10.445 3.045 ;
      LAYER met1 ;
        RECT 4.325 4.155 4.555 4.185 ;
        RECT 10.245 4.155 10.475 4.185 ;
        RECT 4.295 3.985 10.505 4.155 ;
        RECT 4.325 3.955 4.555 3.985 ;
        RECT 10.245 3.955 10.475 3.985 ;
        RECT 6.545 3.415 6.775 3.445 ;
        RECT 10.245 3.415 10.475 3.445 ;
        RECT 6.515 3.245 10.505 3.415 ;
        RECT 6.545 3.215 6.775 3.245 ;
        RECT 10.245 3.215 10.475 3.245 ;
        RECT 10.245 3.045 10.475 3.075 ;
        RECT 10.095 2.875 10.505 3.045 ;
        RECT 10.245 2.845 10.475 2.875 ;
    END
  END B
  PIN VDD
    ANTENNADIFFAREA 13.293050 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 11.520 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 11.255 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 0.585 5.415 0.755 7.460 ;
        RECT 1.465 5.415 1.635 7.460 ;
        RECT 2.065 4.340 2.375 7.460 ;
        RECT 3.365 5.785 3.535 7.460 ;
        RECT 5.395 4.340 5.705 7.460 ;
        RECT 6.695 5.785 6.865 7.460 ;
        RECT 8.725 4.340 9.035 7.460 ;
        RECT 9.465 5.415 9.635 7.460 ;
        RECT 10.345 5.415 10.515 7.460 ;
        RECT 10.945 4.340 11.255 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 1.025 7.525 1.195 7.695 ;
        RECT 1.415 7.525 1.585 7.695 ;
        RECT 1.775 7.525 1.945 7.695 ;
        RECT 2.495 7.525 2.665 7.695 ;
        RECT 2.855 7.525 3.025 7.695 ;
        RECT 3.215 7.525 3.385 7.695 ;
        RECT 3.575 7.525 3.745 7.695 ;
        RECT 4.025 7.525 4.195 7.695 ;
        RECT 4.385 7.525 4.555 7.695 ;
        RECT 4.745 7.525 4.915 7.695 ;
        RECT 5.105 7.525 5.275 7.695 ;
        RECT 5.825 7.525 5.995 7.695 ;
        RECT 6.185 7.525 6.355 7.695 ;
        RECT 6.545 7.525 6.715 7.695 ;
        RECT 6.905 7.525 7.075 7.695 ;
        RECT 7.355 7.525 7.525 7.695 ;
        RECT 7.715 7.525 7.885 7.695 ;
        RECT 8.075 7.525 8.245 7.695 ;
        RECT 8.435 7.525 8.605 7.695 ;
        RECT 9.155 7.525 9.325 7.695 ;
        RECT 9.515 7.525 9.685 7.695 ;
        RECT 9.905 7.525 10.075 7.695 ;
        RECT 10.295 7.525 10.465 7.695 ;
        RECT 10.655 7.525 10.825 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 11.255 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 11.819850 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 11.385 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 1.935 -0.075 2.505 -0.065 ;
        RECT 5.265 -0.075 5.835 -0.065 ;
        RECT 8.595 -0.075 9.165 -0.065 ;
        RECT 10.815 -0.075 11.385 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 0.545 0.755 0.715 1.885 ;
        RECT 1.515 0.755 1.685 1.885 ;
        RECT 0.545 0.585 1.685 0.755 ;
        RECT 0.545 0.310 0.715 0.585 ;
        RECT 1.030 0.310 1.200 0.585 ;
        RECT 1.515 0.310 1.685 0.585 ;
        RECT 2.065 0.310 2.375 2.860 ;
        RECT 3.315 0.310 3.485 1.260 ;
        RECT 5.395 0.310 5.705 2.860 ;
        RECT 6.645 0.310 6.815 1.260 ;
        RECT 8.725 0.310 9.035 2.860 ;
        RECT 9.415 0.755 9.585 1.885 ;
        RECT 10.385 0.755 10.555 1.885 ;
        RECT 9.415 0.585 10.555 0.755 ;
        RECT 9.415 0.310 9.585 0.585 ;
        RECT 9.900 0.310 10.070 0.585 ;
        RECT 10.385 0.310 10.555 0.585 ;
        RECT 10.945 0.310 11.255 2.860 ;
        RECT -0.155 0.000 11.255 0.310 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 1.025 0.065 1.195 0.235 ;
        RECT 1.415 0.065 1.585 0.235 ;
        RECT 1.775 0.065 1.945 0.235 ;
        RECT 2.495 0.065 2.665 0.235 ;
        RECT 2.855 0.065 3.025 0.235 ;
        RECT 3.215 0.065 3.385 0.235 ;
        RECT 3.575 0.065 3.745 0.235 ;
        RECT 4.025 0.065 4.195 0.235 ;
        RECT 4.385 0.065 4.555 0.235 ;
        RECT 4.745 0.065 4.915 0.235 ;
        RECT 5.105 0.065 5.275 0.235 ;
        RECT 5.825 0.065 5.995 0.235 ;
        RECT 6.185 0.065 6.355 0.235 ;
        RECT 6.545 0.065 6.715 0.235 ;
        RECT 6.905 0.065 7.075 0.235 ;
        RECT 7.355 0.065 7.525 0.235 ;
        RECT 7.715 0.065 7.885 0.235 ;
        RECT 8.075 0.065 8.245 0.235 ;
        RECT 8.435 0.065 8.605 0.235 ;
        RECT 9.155 0.065 9.325 0.235 ;
        RECT 9.515 0.065 9.685 0.235 ;
        RECT 9.905 0.065 10.075 0.235 ;
        RECT 10.295 0.065 10.465 0.235 ;
        RECT 10.655 0.065 10.825 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 11.255 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 1.025 4.895 1.195 7.250 ;
        RECT 2.925 5.525 3.095 7.135 ;
        RECT 3.805 7.055 4.855 7.225 ;
        RECT 3.805 5.525 3.975 7.055 ;
        RECT 4.685 5.785 4.855 7.055 ;
        RECT 2.925 5.355 3.975 5.525 ;
        RECT 6.255 5.525 6.425 7.135 ;
        RECT 7.135 7.055 8.185 7.225 ;
        RECT 7.135 5.525 7.305 7.055 ;
        RECT 8.015 5.785 8.185 7.055 ;
        RECT 6.255 5.355 7.305 5.525 ;
        RECT 1.025 4.725 1.565 4.895 ;
        RECT 1.395 2.305 1.565 4.725 ;
        RECT 6.575 4.275 6.745 5.100 ;
        RECT 1.025 2.135 1.565 2.305 ;
        RECT 1.025 0.975 1.195 2.135 ;
        RECT 4.355 2.055 4.525 3.125 ;
        RECT 7.685 2.055 7.855 5.100 ;
        RECT 9.905 4.895 10.075 7.250 ;
        RECT 9.535 4.725 10.075 4.895 ;
        RECT 9.535 2.305 9.705 4.725 ;
        RECT 9.535 2.135 10.075 2.305 ;
        RECT 2.830 1.805 3.000 1.885 ;
        RECT 3.800 1.805 3.970 1.885 ;
        RECT 2.830 1.635 3.970 1.805 ;
        RECT 2.830 0.505 3.000 1.635 ;
        RECT 3.800 0.755 3.970 1.635 ;
        RECT 6.160 1.805 6.330 1.885 ;
        RECT 7.130 1.805 7.300 1.885 ;
        RECT 6.160 1.635 7.300 1.805 ;
        RECT 4.770 0.755 4.940 1.525 ;
        RECT 3.800 0.585 4.940 0.755 ;
        RECT 3.800 0.505 3.970 0.585 ;
        RECT 4.770 0.505 4.940 0.585 ;
        RECT 6.160 0.505 6.330 1.635 ;
        RECT 7.130 0.755 7.300 1.635 ;
        RECT 8.100 0.755 8.270 1.525 ;
        RECT 9.905 0.975 10.075 2.135 ;
        RECT 7.130 0.585 8.270 0.755 ;
        RECT 7.130 0.505 7.300 0.585 ;
        RECT 8.100 0.505 8.270 0.585 ;
      LAYER mcon ;
        RECT 6.575 4.355 6.745 4.525 ;
        RECT 1.395 2.505 1.565 2.675 ;
        RECT 4.355 2.875 4.525 3.045 ;
        RECT 7.685 2.505 7.855 2.675 ;
        RECT 9.535 4.355 9.705 4.525 ;
        RECT 9.535 2.875 9.705 3.045 ;
      LAYER met1 ;
        RECT 6.545 4.525 6.775 4.555 ;
        RECT 9.505 4.525 9.735 4.555 ;
        RECT 6.515 4.355 9.765 4.525 ;
        RECT 6.545 4.325 6.775 4.355 ;
        RECT 9.505 4.325 9.735 4.355 ;
        RECT 4.325 3.045 4.555 3.075 ;
        RECT 9.505 3.045 9.735 3.075 ;
        RECT 4.295 2.875 9.765 3.045 ;
        RECT 4.325 2.845 4.555 2.875 ;
        RECT 9.505 2.845 9.735 2.875 ;
        RECT 1.365 2.675 1.595 2.705 ;
        RECT 7.655 2.675 7.885 2.705 ;
        RECT 1.335 2.505 7.915 2.675 ;
        RECT 1.365 2.475 1.595 2.505 ;
        RECT 7.655 2.475 7.885 2.505 ;
  END
END XNOR2X1






MACRO XOR2X1
  CLASS BLOCK ;
  FOREIGN XOR2X1 ;
  ORIGIN 0.420 0.075 ;
  SIZE 11.940 BY 7.950 ;
  PIN Y
    ANTENNADIFFAREA 1.543800 ;
    PORT
      LAYER li1 ;
        RECT 4.245 5.525 4.415 6.795 ;
        RECT 7.575 5.525 7.745 6.795 ;
        RECT 4.245 5.355 4.895 5.525 ;
        RECT 7.575 5.355 8.225 5.525 ;
        RECT 4.725 1.875 4.895 5.355 ;
        RECT 8.055 1.875 8.225 5.355 ;
        RECT 4.285 1.705 4.895 1.875 ;
        RECT 7.615 1.705 8.225 1.875 ;
        RECT 4.285 0.975 4.455 1.705 ;
        RECT 7.615 0.975 7.785 1.705 ;
      LAYER mcon ;
        RECT 4.725 3.615 4.895 3.785 ;
        RECT 8.055 3.615 8.225 3.785 ;
      LAYER met1 ;
        RECT 4.695 3.785 4.925 3.815 ;
        RECT 8.025 3.785 8.255 3.815 ;
        RECT 4.665 3.615 8.285 3.785 ;
        RECT 4.695 3.585 4.925 3.615 ;
        RECT 8.025 3.585 8.255 3.615 ;
    END
  END Y
  PIN A
    ANTENNAGATEAREA 2.060500 ;
    PORT
      LAYER li1 ;
        RECT 0.655 2.055 0.825 5.095 ;
        RECT 3.245 2.055 3.415 5.100 ;
      LAYER mcon ;
        RECT 0.655 4.355 0.825 4.525 ;
        RECT 3.245 4.355 3.415 4.525 ;
      LAYER met1 ;
        RECT 0.625 4.525 0.855 4.555 ;
        RECT 3.215 4.525 3.445 4.555 ;
        RECT 0.595 4.355 3.475 4.525 ;
        RECT 0.625 4.325 0.855 4.355 ;
        RECT 3.215 4.325 3.445 4.355 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 2.054500 ;
    PORT
      LAYER li1 ;
        RECT 6.575 4.275 6.745 5.100 ;
        RECT 4.355 2.055 4.525 2.755 ;
        RECT 10.275 2.055 10.445 5.095 ;
      LAYER mcon ;
        RECT 6.575 4.355 6.745 4.525 ;
        RECT 10.275 4.355 10.445 4.525 ;
        RECT 4.355 2.505 4.525 2.675 ;
        RECT 10.275 2.505 10.445 2.675 ;
      LAYER met1 ;
        RECT 6.545 4.525 6.775 4.555 ;
        RECT 10.245 4.525 10.475 4.555 ;
        RECT 6.515 4.355 10.505 4.525 ;
        RECT 6.545 4.325 6.775 4.355 ;
        RECT 10.245 4.325 10.475 4.355 ;
        RECT 4.325 2.675 4.555 2.705 ;
        RECT 10.245 2.675 10.475 2.705 ;
        RECT 4.295 2.505 10.505 2.675 ;
        RECT 4.325 2.475 4.555 2.505 ;
        RECT 10.245 2.475 10.475 2.505 ;
    END
  END B
  PIN VDD
    ANTENNADIFFAREA 13.293050 ;
    PORT
      LAYER nwell ;
        RECT -0.420 4.160 11.520 7.875 ;
      LAYER li1 ;
        RECT -0.155 7.460 11.255 7.770 ;
        RECT -0.155 4.340 0.155 7.460 ;
        RECT 0.585 5.415 0.755 7.460 ;
        RECT 1.465 5.415 1.635 7.460 ;
        RECT 2.065 4.340 2.375 7.460 ;
        RECT 3.365 5.785 3.535 7.460 ;
        RECT 5.395 4.340 5.705 7.460 ;
        RECT 6.695 5.785 6.865 7.460 ;
        RECT 8.725 4.340 9.035 7.460 ;
        RECT 9.465 5.415 9.635 7.460 ;
        RECT 10.345 5.415 10.515 7.460 ;
        RECT 10.945 4.340 11.255 7.460 ;
      LAYER mcon ;
        RECT 0.275 7.525 0.445 7.695 ;
        RECT 0.635 7.525 0.805 7.695 ;
        RECT 1.025 7.525 1.195 7.695 ;
        RECT 1.415 7.525 1.585 7.695 ;
        RECT 1.775 7.525 1.945 7.695 ;
        RECT 2.495 7.525 2.665 7.695 ;
        RECT 2.855 7.525 3.025 7.695 ;
        RECT 3.215 7.525 3.385 7.695 ;
        RECT 3.575 7.525 3.745 7.695 ;
        RECT 4.025 7.525 4.195 7.695 ;
        RECT 4.385 7.525 4.555 7.695 ;
        RECT 4.745 7.525 4.915 7.695 ;
        RECT 5.105 7.525 5.275 7.695 ;
        RECT 5.825 7.525 5.995 7.695 ;
        RECT 6.185 7.525 6.355 7.695 ;
        RECT 6.545 7.525 6.715 7.695 ;
        RECT 6.905 7.525 7.075 7.695 ;
        RECT 7.355 7.525 7.525 7.695 ;
        RECT 7.715 7.525 7.885 7.695 ;
        RECT 8.075 7.525 8.245 7.695 ;
        RECT 8.435 7.525 8.605 7.695 ;
        RECT 9.155 7.525 9.325 7.695 ;
        RECT 9.515 7.525 9.685 7.695 ;
        RECT 9.905 7.525 10.075 7.695 ;
        RECT 10.295 7.525 10.465 7.695 ;
        RECT 10.655 7.525 10.825 7.695 ;
      LAYER met1 ;
        RECT -0.155 7.460 11.255 7.770 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 11.819850 ;
    PORT
      LAYER pwell ;
        RECT -0.285 -0.065 11.385 2.990 ;
        RECT -0.285 -0.075 0.285 -0.065 ;
        RECT 1.935 -0.075 2.505 -0.065 ;
        RECT 5.265 -0.075 5.835 -0.065 ;
        RECT 8.595 -0.075 9.165 -0.065 ;
        RECT 10.815 -0.075 11.385 -0.065 ;
      LAYER li1 ;
        RECT -0.155 0.310 0.155 2.860 ;
        RECT 0.545 0.755 0.715 1.885 ;
        RECT 1.515 0.755 1.685 1.885 ;
        RECT 0.545 0.585 1.685 0.755 ;
        RECT 0.545 0.310 0.715 0.585 ;
        RECT 1.030 0.310 1.200 0.585 ;
        RECT 1.515 0.310 1.685 0.585 ;
        RECT 2.065 0.310 2.375 2.860 ;
        RECT 3.315 0.310 3.485 1.260 ;
        RECT 5.395 0.310 5.705 2.860 ;
        RECT 6.645 0.310 6.815 1.260 ;
        RECT 8.725 0.310 9.035 2.860 ;
        RECT 9.415 0.755 9.585 1.885 ;
        RECT 10.385 0.755 10.555 1.885 ;
        RECT 9.415 0.585 10.555 0.755 ;
        RECT 9.415 0.310 9.585 0.585 ;
        RECT 9.900 0.310 10.070 0.585 ;
        RECT 10.385 0.310 10.555 0.585 ;
        RECT 10.945 0.310 11.255 2.860 ;
        RECT -0.155 0.000 11.255 0.310 ;
      LAYER mcon ;
        RECT 0.275 0.065 0.445 0.235 ;
        RECT 0.635 0.065 0.805 0.235 ;
        RECT 1.025 0.065 1.195 0.235 ;
        RECT 1.415 0.065 1.585 0.235 ;
        RECT 1.775 0.065 1.945 0.235 ;
        RECT 2.495 0.065 2.665 0.235 ;
        RECT 2.855 0.065 3.025 0.235 ;
        RECT 3.215 0.065 3.385 0.235 ;
        RECT 3.575 0.065 3.745 0.235 ;
        RECT 4.025 0.065 4.195 0.235 ;
        RECT 4.385 0.065 4.555 0.235 ;
        RECT 4.745 0.065 4.915 0.235 ;
        RECT 5.105 0.065 5.275 0.235 ;
        RECT 5.825 0.065 5.995 0.235 ;
        RECT 6.185 0.065 6.355 0.235 ;
        RECT 6.545 0.065 6.715 0.235 ;
        RECT 6.905 0.065 7.075 0.235 ;
        RECT 7.355 0.065 7.525 0.235 ;
        RECT 7.715 0.065 7.885 0.235 ;
        RECT 8.075 0.065 8.245 0.235 ;
        RECT 8.435 0.065 8.605 0.235 ;
        RECT 9.155 0.065 9.325 0.235 ;
        RECT 9.515 0.065 9.685 0.235 ;
        RECT 9.905 0.065 10.075 0.235 ;
        RECT 10.295 0.065 10.465 0.235 ;
        RECT 10.655 0.065 10.825 0.235 ;
      LAYER met1 ;
        RECT -0.155 0.000 11.255 0.310 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 1.025 4.895 1.195 7.250 ;
        RECT 2.925 5.525 3.095 7.135 ;
        RECT 3.805 7.055 4.855 7.225 ;
        RECT 3.805 5.525 3.975 7.055 ;
        RECT 4.685 5.785 4.855 7.055 ;
        RECT 2.925 5.355 3.975 5.525 ;
        RECT 6.255 5.525 6.425 7.135 ;
        RECT 7.135 7.055 8.185 7.225 ;
        RECT 7.135 5.525 7.305 7.055 ;
        RECT 8.015 5.785 8.185 7.055 ;
        RECT 6.255 5.355 7.305 5.525 ;
        RECT 1.025 4.725 1.565 4.895 ;
        RECT 1.395 2.305 1.565 4.725 ;
        RECT 4.355 3.905 4.525 5.100 ;
        RECT 1.025 2.135 1.565 2.305 ;
        RECT 1.025 0.975 1.195 2.135 ;
        RECT 6.575 2.055 6.745 3.125 ;
        RECT 7.685 2.055 7.855 5.100 ;
        RECT 9.905 4.895 10.075 7.250 ;
        RECT 9.535 4.725 10.075 4.895 ;
        RECT 9.535 2.305 9.705 4.725 ;
        RECT 9.535 2.135 10.075 2.305 ;
        RECT 2.830 1.805 3.000 1.885 ;
        RECT 3.800 1.805 3.970 1.885 ;
        RECT 2.830 1.635 3.970 1.805 ;
        RECT 2.830 0.505 3.000 1.635 ;
        RECT 3.800 0.755 3.970 1.635 ;
        RECT 6.160 1.805 6.330 1.885 ;
        RECT 7.130 1.805 7.300 1.885 ;
        RECT 6.160 1.635 7.300 1.805 ;
        RECT 4.770 0.755 4.940 1.525 ;
        RECT 3.800 0.585 4.940 0.755 ;
        RECT 3.800 0.505 3.970 0.585 ;
        RECT 4.770 0.505 4.940 0.585 ;
        RECT 6.160 0.505 6.330 1.635 ;
        RECT 7.130 0.755 7.300 1.635 ;
        RECT 8.100 0.755 8.270 1.525 ;
        RECT 9.905 0.975 10.075 2.135 ;
        RECT 7.130 0.585 8.270 0.755 ;
        RECT 7.130 0.505 7.300 0.585 ;
        RECT 8.100 0.505 8.270 0.585 ;
      LAYER mcon ;
        RECT 4.355 3.985 4.525 4.155 ;
        RECT 1.395 3.245 1.565 3.415 ;
        RECT 7.685 3.245 7.855 3.415 ;
        RECT 6.575 2.875 6.745 3.045 ;
        RECT 9.535 3.985 9.705 4.155 ;
        RECT 9.535 2.875 9.705 3.045 ;
      LAYER met1 ;
        RECT 4.325 4.155 4.555 4.185 ;
        RECT 9.505 4.155 9.735 4.185 ;
        RECT 4.295 3.985 9.765 4.155 ;
        RECT 4.325 3.955 4.555 3.985 ;
        RECT 9.505 3.955 9.735 3.985 ;
        RECT 1.365 3.415 1.595 3.445 ;
        RECT 7.655 3.415 7.885 3.445 ;
        RECT 1.335 3.245 7.915 3.415 ;
        RECT 1.365 3.215 1.595 3.245 ;
        RECT 7.655 3.215 7.885 3.245 ;
        RECT 6.545 3.045 6.775 3.075 ;
        RECT 9.505 3.045 9.735 3.075 ;
        RECT 6.515 2.875 9.765 3.045 ;
        RECT 6.545 2.845 6.775 2.875 ;
        RECT 9.505 2.845 9.735 2.875 ;
  END
END XOR2X1


