magic
tech sky130A
magscale 1 2
timestamp 1642971615
<< error_p >>
rect 799 313 800 314
rect 983 313 984 314
rect 800 312 801 313
rect 984 312 985 313
rect 85 310 86 311
rect 86 309 87 310
rect 815 282 816 283
rect 850 282 851 283
rect 999 282 1000 283
rect 1034 282 1035 283
rect 101 279 102 280
rect 136 279 137 280
rect 101 188 102 189
rect 136 188 137 189
rect 815 179 816 180
rect 850 179 851 180
rect 999 179 1000 180
rect 1034 179 1035 180
<< nmos >>
rect 56 310 86 360
rect 56 280 152 310
tri 152 280 182 310 sw
rect 56 196 86 280
tri 86 264 102 280 nw
tri 136 264 152 280 ne
tri 86 196 94 204 sw
tri 144 196 152 204 se
rect 152 196 182 280
rect 56 193 94 196
tri 94 193 97 196 sw
rect 56 188 97 193
tri 97 188 102 193 sw
tri 140 192 144 196 se
rect 144 192 182 196
tri 136 188 140 192 se
rect 140 188 182 192
tri 56 158 86 188 ne
rect 86 158 152 188
tri 152 158 182 188 nw
rect 770 313 800 363
rect 954 313 984 363
rect 770 283 866 313
tri 866 283 896 313 sw
rect 770 179 800 283
tri 800 267 816 283 nw
tri 850 267 866 283 ne
tri 800 179 816 195 sw
tri 850 179 866 195 se
rect 866 179 896 283
rect 954 283 1050 313
tri 1050 283 1080 313 sw
tri 770 149 800 179 ne
rect 800 149 866 179
tri 866 149 896 179 nw
rect 954 179 984 283
tri 984 267 1000 283 nw
tri 1034 267 1050 283 ne
tri 984 179 1000 195 sw
tri 1034 179 1050 195 se
rect 1050 179 1080 283
tri 954 149 984 179 ne
rect 984 149 1050 179
tri 1050 149 1080 179 nw
<< ndiff >>
rect 0 304 56 360
rect 86 310 238 360
rect 0 270 10 304
rect 44 270 56 304
tri 152 280 182 310 ne
rect 182 306 238 310
rect 0 215 56 270
rect 0 181 10 215
rect 44 181 56 215
tri 86 264 102 280 se
rect 102 264 136 280
tri 136 264 152 280 sw
rect 86 242 152 264
rect 86 208 98 242
rect 132 208 152 242
rect 86 204 152 208
tri 86 196 94 204 ne
rect 94 196 144 204
tri 144 196 152 204 nw
rect 182 272 194 306
rect 228 272 238 306
rect 182 215 238 272
tri 94 193 97 196 ne
rect 97 193 140 196
tri 97 188 102 193 ne
rect 102 192 140 193
tri 140 192 144 196 nw
rect 102 188 136 192
tri 136 188 140 192 nw
rect 0 158 56 181
tri 56 158 86 188 sw
tri 152 158 182 188 se
rect 182 181 194 215
rect 228 181 238 215
rect 182 158 238 181
rect 0 147 238 158
rect 0 113 10 147
rect 44 113 98 147
rect 132 113 194 147
rect 228 113 238 147
rect 0 101 238 113
rect 714 307 770 363
rect 800 313 954 363
rect 984 313 1134 363
rect 714 273 724 307
rect 758 273 770 307
tri 866 283 896 313 ne
rect 896 309 954 313
rect 714 206 770 273
rect 714 172 724 206
rect 758 172 770 206
tri 800 267 816 283 se
rect 816 267 850 283
tri 850 267 866 283 sw
rect 800 233 866 267
rect 800 199 812 233
rect 846 199 866 233
rect 800 195 866 199
tri 800 179 816 195 ne
rect 816 179 850 195
tri 850 179 866 195 nw
rect 896 275 908 309
rect 942 275 954 309
tri 1050 283 1080 313 ne
rect 896 206 954 275
rect 714 149 770 172
tri 770 149 800 179 sw
tri 866 149 896 179 se
rect 896 172 908 206
rect 942 172 954 206
tri 984 267 1000 283 se
rect 1000 267 1034 283
tri 1034 267 1050 283 sw
rect 984 233 1050 267
rect 984 199 996 233
rect 1030 199 1050 233
rect 984 195 1050 199
tri 984 179 1000 195 ne
rect 1000 179 1034 195
tri 1034 179 1050 195 nw
rect 1080 279 1092 313
rect 1126 279 1134 313
rect 1080 206 1134 279
rect 896 149 954 172
tri 954 149 984 179 sw
tri 1050 149 1080 179 se
rect 1080 172 1092 206
rect 1126 172 1134 206
rect 1080 149 1134 172
rect 714 138 1134 149
rect 714 104 724 138
rect 758 104 812 138
rect 846 104 908 138
rect 942 104 996 138
rect 1030 104 1092 138
rect 1126 104 1134 138
rect 714 92 1134 104
<< ndiffc >>
rect 10 270 44 304
rect 10 181 44 215
rect 98 208 132 242
rect 194 272 228 306
rect 194 181 228 215
rect 10 113 44 147
rect 98 113 132 147
rect 194 113 228 147
rect 724 273 758 307
rect 724 172 758 206
rect 812 199 846 233
rect 908 275 942 309
rect 908 172 942 206
rect 996 199 1030 233
rect 1092 279 1126 313
rect 1092 172 1126 206
rect 724 104 758 138
rect 812 104 846 138
rect 908 104 942 138
rect 996 104 1030 138
rect 1092 104 1126 138
<< psubdiff >>
rect -116 429 354 491
rect -116 47 -54 429
rect 292 47 354 429
rect -116 13 24 47
rect 58 13 92 47
rect 126 13 160 47
rect 194 13 354 47
rect -116 0 354 13
rect 598 420 1250 482
rect 598 38 660 420
rect 1188 38 1250 420
rect 598 4 738 38
rect 772 4 806 38
rect 840 4 874 38
rect 908 4 942 38
rect 976 4 1010 38
rect 1044 4 1078 38
rect 1112 4 1250 38
rect 598 -9 1250 4
<< psubdiffcont >>
rect 24 13 58 47
rect 92 13 126 47
rect 160 13 194 47
rect 738 4 772 38
rect 806 4 840 38
rect 874 4 908 38
rect 942 4 976 38
rect 1010 4 1044 38
rect 1078 4 1112 38
<< poly >>
rect 56 360 86 402
rect 770 363 800 405
rect 954 363 984 405
<< locali >>
rect -116 62 -54 491
rect 10 304 44 331
rect 10 215 44 270
rect 194 306 228 331
rect 98 242 132 258
rect 98 192 132 208
rect 194 215 228 272
rect 10 147 44 181
rect 194 147 228 181
rect 44 113 98 147
rect 132 113 194 147
rect 228 113 238 147
rect 10 62 44 113
rect 194 62 228 113
rect 292 62 354 491
rect -116 47 354 62
rect -116 13 24 47
rect 58 13 92 47
rect 126 13 160 47
rect 194 13 354 47
rect -116 0 354 13
rect 598 53 660 482
rect 724 307 758 334
rect 908 309 942 334
rect 724 206 758 273
rect 812 269 846 278
rect 812 233 846 235
rect 812 183 846 199
rect 1092 313 1126 334
rect 908 206 942 275
rect 724 138 758 172
rect 996 269 1030 279
rect 996 233 1030 235
rect 996 183 1030 199
rect 1092 206 1126 279
rect 908 138 942 172
rect 1092 138 1126 172
rect 758 104 812 138
rect 846 104 908 138
rect 942 104 996 138
rect 1030 104 1092 138
rect 724 53 758 104
rect 908 53 942 104
rect 1092 53 1126 104
rect 1188 53 1250 482
rect 598 38 1250 53
rect 598 4 738 38
rect 772 4 806 38
rect 840 4 874 38
rect 908 4 942 38
rect 976 4 1010 38
rect 1044 4 1078 38
rect 1112 4 1250 38
rect 598 -9 1250 4
<< viali >>
rect 24 13 58 47
rect 92 13 126 47
rect 160 13 194 47
rect 812 235 846 269
rect 996 235 1030 269
rect 738 4 772 38
rect 806 4 840 38
rect 874 4 908 38
rect 942 4 976 38
rect 1010 4 1044 38
rect 1078 4 1112 38
<< metal1 >>
rect -116 62 -54 491
rect 292 62 354 491
rect -116 47 354 62
rect -116 13 24 47
rect 58 13 92 47
rect 126 13 160 47
rect 194 13 354 47
rect -116 0 354 13
rect 598 53 660 482
rect 812 276 846 281
rect 996 276 1030 281
rect 806 269 852 276
rect 990 269 1036 276
rect 806 235 812 269
rect 846 235 996 269
rect 1030 235 1036 269
rect 806 228 852 235
rect 990 228 1036 235
rect 812 223 846 228
rect 996 223 1030 228
rect 1188 53 1250 482
rect 598 38 1250 53
rect 598 4 738 38
rect 772 4 806 38
rect 840 4 874 38
rect 908 4 942 38
rect 976 4 1010 38
rect 1044 4 1078 38
rect 1112 4 1250 38
rect 598 -9 1250 4
<< labels >>
rlabel metal1 992 17 992 17 1 VSS
port 1 n
rlabel metal1 812 235 846 269 1 A
port 2 n
<< end >>
