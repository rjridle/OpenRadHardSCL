* SPICE3 file created from INVX1.ext - technology: sky130A

.subckt INVX1 VDD VSS
M1000 VDD a_56_401# a_102_270# VDD pshort w=1.26u l=0.15u
+  ad=0.693p pd=6.14u as=0p ps=0u
M1001 a_102_270# a_56_401# VDD VDD pshort w=1.26u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_102_270# a_56_401# VSS VSS nshort w=3u l=0.15u
+  ad=0p pd=0u as=1.12185p ps=7.97u
.ends
