* SPICE3 file created from AOA4X1.ext - technology: sky130A

.subckt AOA4X1 Y A B C D VDD GND
X0 VDD.t13 A.t0 a_217_1050.t2 ��8V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X1 VDD.t23 a_217_1050.t5 a_797_1051.t3 �&=9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X2 Y.t2 a_1549_1050.t5 VDD.t5  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X3 VDD.t25 B.t0 a_217_1050.t4 VDD.t24 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X4 VDD.t19 a_864_209.t4 a_1549_1050.t4  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X5 GND A.t1 a_112_101.t0 GND sky130_fd_pr__nfet_01v8 ad=3.4356p pd=2.418u as=0p ps=0u w=0u l=0u
X6 GND a_864_209.t5 a_1444_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X7 VDD.t1 a_1549_1050.t6 Y.t1 |�P� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X8 a_797_1051.t0 C.t0 a_864_209.t0  |�P� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X9 a_217_1050.t3 A.t2 VDD.t11 �{�P� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X10 Y a_1549_1050.t7 GND.t3 GND sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=0p ps=0u w=0u l=0u
X11 a_797_1051.t2 a_217_1050.t7 VDD.t21  |�P� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X12 VDD.t15 D.t0 a_1549_1050.t2 �{�P� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X13 a_217_1050.t1 B.t1 VDD.t8  |�P� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X14 a_1549_1050.t3 a_864_209.t6 VDD.t17 �{�P� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X15 a_864_209.t2 C.t1 a_797_1051.t1  |�P� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X16 a_1549_1050.t1 D.t2 VDD.t3 �{�P� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
C0 A B 0.27fF
C1 C VDD 0.32fF
C2 Y VDD 1.07fF
C3 VDD B 0.32fF
C4 A VDD 0.32fF
C5 D VDD 0.33fF
R0 A.n0 A.t0 480.392
R1 A.n0 A.t2 403.272
R2 A.n1 A.t1 301.486
R3 A.n1 A.n0 227.006
R4 A.n2 A.n1 4.65
R5 A.n2 A 0.046
R6 a_217_1050.n3 a_217_1050.t7 486.819
R7 a_217_1050.n3 a_217_1050.t5 384.527
R8 a_217_1050.n4 a_217_1050.t6 267.201
R9 a_217_1050.n4 a_217_1050.n3 262.705
R10 a_217_1050.n5 a_217_1050.n2 243.576
R11 a_217_1050.n7 a_217_1050.n5 228.526
R12 a_217_1050.n2 a_217_1050.n1 157.964
R13 a_217_1050.n2 a_217_1050.n0 91.706
R14 a_217_1050.n7 a_217_1050.n6 15.218
R15 a_217_1050.n0 a_217_1050.t4 14.282
R16 a_217_1050.n0 a_217_1050.t1 14.282
R17 a_217_1050.n1 a_217_1050.t2 14.282
R18 a_217_1050.n1 a_217_1050.t3 14.282
R19 a_217_1050.n8 a_217_1050.n7 12.014
R20 a_217_1050.n5 a_217_1050.n4 10.615
R21 VDD.n123 VDD.n116 144.705
R22 VDD.n204 VDD.n193 144.705
R23 VDD.n66 VDD.n55 144.705
R24 VDD.n171 VDD.t25 143.754
R25 VDD.n69 VDD.t15 143.754
R26 VDD.n149 VDD.t11 135.17
R27 VDD.n91 VDD.t17 135.17
R28 VDD.n35 VDD.t5 135.17
R29 VDD.n24 VDD.t1 135.17
R30 VDD.n212 VDD.n211 129.849
R31 VDD.n163 VDD.n162 129.472
R32 VDD.n79 VDD.n78 129.472
R33 VDD.n51 VDD.n50 92.5
R34 VDD.n49 VDD.n48 92.5
R35 VDD.n47 VDD.n46 92.5
R36 VDD.n45 VDD.n44 92.5
R37 VDD.n53 VDD.n52 92.5
R38 VDD.n112 VDD.n111 92.5
R39 VDD.n110 VDD.n109 92.5
R40 VDD.n108 VDD.n107 92.5
R41 VDD.n106 VDD.n105 92.5
R42 VDD.n114 VDD.n113 92.5
R43 VDD.n189 VDD.n188 92.5
R44 VDD.n187 VDD.n186 92.5
R45 VDD.n185 VDD.n184 92.5
R46 VDD.n183 VDD.n182 92.5
R47 VDD.n191 VDD.n190 92.5
R48 VDD.n137 VDD.n136 92.5
R49 VDD.n135 VDD.n134 92.5
R50 VDD.n133 VDD.n132 92.5
R51 VDD.n131 VDD.n130 92.5
R52 VDD.n139 VDD.n138 92.5
R53 VDD.n14 VDD.n1 92.5
R54 VDD.n5 VDD.n4 92.5
R55 VDD.n7 VDD.n6 92.5
R56 VDD.n9 VDD.n8 92.5
R57 VDD.n11 VDD.n10 92.5
R58 VDD.n13 VDD.n12 92.5
R59 VDD.n21 VDD.n20 92.059
R60 VDD.n65 VDD.n64 92.059
R61 VDD.n122 VDD.n121 92.059
R62 VDD.n203 VDD.n202 92.059
R63 VDD.n145 VDD.n144 92.059
R64 VDD.n20 VDD.n16 67.194
R65 VDD.n20 VDD.n17 67.194
R66 VDD.n20 VDD.n18 67.194
R67 VDD.n20 VDD.n19 67.194
R68 VDD.n129 VDD.n128 44.141
R69 VDD.n104 VDD.n103 44.141
R70 VDD.n5 VDD.n3 44.141
R71 VDD.n103 VDD.n101 44.107
R72 VDD.n128 VDD.n126 44.107
R73 VDD.n3 VDD.n2 44.107
R74 VDD.n25 |�P� 43.472
R75 VDD.n33 �l[9V 43.472
R76 VDD.n20 VDD.n15 41.052
R77 VDD.n59 VDD.n57 39.742
R78 VDD.n59 VDD.n58 39.742
R79 VDD.n61 VDD.n60 39.742
R80 VDD.n118 VDD.n117 39.742
R81 VDD.n141 VDD.n140 39.742
R82 VDD.n201 VDD.n198 39.742
R83 VDD.n201 VDD.n200 39.742
R84 VDD.n197 VDD.n196 39.742
R85 VDD.n103 VDD.n102 38
R86 VDD.n128 VDD.n127 38
R87 VDD.n101 VDD.n100 36.774
R88 VDD.n57 VDD.n56 36.774
R89 VDD.n200 VDD.n199 36.774
R90 VDD.n1 VDD.n0 30.923
R91 VDD.n64 VDD.n62 26.38
R92 VDD.n64 VDD.n61 26.38
R93 VDD.n64 VDD.n59 26.38
R94 VDD.n64 VDD.n63 26.38
R95 VDD.n121 VDD.n119 26.38
R96 VDD.n121 VDD.n118 26.38
R97 VDD.n121 VDD.n120 26.38
R98 VDD.n144 VDD.n142 26.38
R99 VDD.n144 VDD.n141 26.38
R100 VDD.n144 VDD.n143 26.38
R101 VDD.n202 VDD.n201 26.38
R102 VDD.n202 VDD.n197 26.38
R103 VDD.n202 VDD.n195 26.38
R104 VDD.n202 VDD.n194 26.38
R105 VDD.n147 VDD.n139 22.915
R106 VDD.n23 VDD.n14 22.915
R107 VDD.n74 �{�P� 20.457
R108 VDD.n224  |�P� 20.457
R109 VDD.n167 VDD.t24 20.457
R110 VDD.n87 �{�P� 17.9
R111 VDD.n213 �&=9V 17.9
R112 VDD.n154 �{�P� 17.9
R113 VDD.n139 VDD.n137 14.864
R114 VDD.n137 VDD.n135 14.864
R115 VDD.n135 VDD.n133 14.864
R116 VDD.n133 VDD.n131 14.864
R117 VDD.n131 VDD.n129 14.864
R118 VDD.n114 VDD.n112 14.864
R119 VDD.n112 VDD.n110 14.864
R120 VDD.n110 VDD.n108 14.864
R121 VDD.n108 VDD.n106 14.864
R122 VDD.n106 VDD.n104 14.864
R123 VDD.n53 VDD.n51 14.864
R124 VDD.n51 VDD.n49 14.864
R125 VDD.n49 VDD.n47 14.864
R126 VDD.n47 VDD.n45 14.864
R127 VDD.n45 VDD.n43 14.864
R128 VDD.n43 VDD.n42 14.864
R129 VDD.n191 VDD.n189 14.864
R130 VDD.n189 VDD.n187 14.864
R131 VDD.n187 VDD.n185 14.864
R132 VDD.n185 VDD.n183 14.864
R133 VDD.n183 VDD.n181 14.864
R134 VDD.n181 VDD.n180 14.864
R135 VDD.n14 VDD.n13 14.864
R136 VDD.n13 VDD.n11 14.864
R137 VDD.n11 VDD.n9 14.864
R138 VDD.n9 VDD.n7 14.864
R139 VDD.n7 VDD.n5 14.864
R140 VDD.n67 VDD.n54 14.864
R141 VDD.n124 VDD.n115 14.864
R142 VDD.n205 VDD.n192 14.864
R143 VDD.n162 VDD.t8 14.282
R144 VDD.n162 VDD.t13 14.282
R145 VDD.n211 VDD.t21 14.282
R146 VDD.n211 VDD.t23 14.282
R147 VDD.n78 VDD.t3 14.282
R148 VDD.n78 VDD.t19 14.282
R149 VDD.n81 VDD.n79 9.083
R150 VDD.n165 VDD.n163 9.083
R151 VDD.n23 VDD.n22 8.855
R152 VDD.n22 VDD.n21 8.855
R153 VDD.n27 VDD.n26 8.855
R154 VDD.n26 VDD.n25 8.855
R155 VDD.n31 VDD.n30 8.855
R156 VDD.n30 VDD.n29 8.855
R157 VDD.n36 VDD.n34 8.855
R158 VDD.n34 VDD.n33 8.855
R159 VDD.n40 VDD.n39 8.855
R160 VDD.n39 VDD.n38 8.855
R161 VDD.n67 VDD.n66 8.855
R162 VDD.n66 VDD.n65 8.855
R163 VDD.n72 VDD.n71 8.855
R164 VDD.n71 VDD.n70 8.855
R165 VDD.n76 VDD.n75 8.855
R166 VDD.n75 VDD.n74 8.855
R167 VDD.n81 VDD.n80 8.855
R168 VDD.n80 �{�P� 8.855
R169 VDD.n85 VDD.n84 8.855
R170 VDD.n84 VDD.n83 8.855
R171 VDD.n89 VDD.n88 8.855
R172 VDD.n88 VDD.n87 8.855
R173 VDD.n94 VDD.n93 8.855
R174 VDD.n93 VDD.n92 8.855
R175 VDD.n98 VDD.n97 8.855
R176 VDD.n97 VDD.n96 8.855
R177 VDD.n124 VDD.n123 8.855
R178 VDD.n123 VDD.n122 8.855
R179 VDD.n230 VDD.n229 8.855
R180 VDD.n229 VDD.n228 8.855
R181 VDD.n226 VDD.n225 8.855
R182 VDD.n225 VDD.n224 8.855
R183 VDD.n222 VDD.n221 8.855
R184 VDD.n221  |�P� 8.855
R185 VDD.n219 VDD.n218 8.855
R186 VDD.n218 VDD.n217 8.855
R187 VDD.n215 VDD.n214 8.855
R188 VDD.n214 VDD.n213 8.855
R189 VDD.n209 VDD.n208 8.855
R190 VDD.n208 VDD.n207 8.855
R191 VDD.n205 VDD.n204 8.855
R192 VDD.n204 VDD.n203 8.855
R193 VDD.n178 VDD.n177 8.855
R194 VDD.n177 VDD.n176 8.855
R195 VDD.n174 VDD.n173 8.855
R196 VDD.n173 VDD.n172 8.855
R197 VDD.n169 VDD.n168 8.855
R198 VDD.n168 VDD.n167 8.855
R199 VDD.n165 VDD.n164 8.855
R200 VDD.n164  |�P� 8.855
R201 VDD.n160 VDD.n159 8.855
R202 VDD.n159 VDD.n158 8.855
R203 VDD.n156 VDD.n155 8.855
R204 VDD.n155 VDD.n154 8.855
R205 VDD.n152 VDD.n151 8.855
R206 VDD.n151 VDD.n150 8.855
R207 VDD.n147 VDD.n146 8.855
R208 VDD.n146 VDD.n145 8.855
R209 VDD.n115 VDD.n114 8.051
R210 VDD.n54 VDD.n53 8.051
R211 VDD.n192 VDD.n191 8.051
R212 VDD.n215 VDD.n212 6.193
R213 VDD.n28 VDD.n23 4.795
R214 VDD.n28 VDD.n27 4.65
R215 VDD.n32 VDD.n31 4.65
R216 VDD.n37 VDD.n36 4.65
R217 VDD.n41 VDD.n40 4.65
R218 VDD.n68 VDD.n67 4.65
R219 VDD.n73 VDD.n72 4.65
R220 VDD.n77 VDD.n76 4.65
R221 VDD.n82 VDD.n81 4.65
R222 VDD.n86 VDD.n85 4.65
R223 VDD.n90 VDD.n89 4.65
R224 VDD.n95 VDD.n94 4.65
R225 VDD.n99 VDD.n98 4.65
R226 VDD.n125 VDD.n124 4.65
R227 VDD.n231 VDD.n230 4.65
R228 VDD.n227 VDD.n226 4.65
R229 VDD.n223 VDD.n222 4.65
R230 VDD.n220 VDD.n219 4.65
R231 VDD.n216 VDD.n215 4.65
R232 VDD.n210 VDD.n209 4.65
R233 VDD.n206 VDD.n205 4.65
R234 VDD.n179 VDD.n178 4.65
R235 VDD.n175 VDD.n174 4.65
R236 VDD.n170 VDD.n169 4.65
R237 VDD.n166 VDD.n165 4.65
R238 VDD.n161 VDD.n160 4.65
R239 VDD.n157 VDD.n156 4.65
R240 VDD.n153 VDD.n152 4.65
R241 VDD.n148 VDD.n147 4.65
R242 VDD.n94 VDD.n91 2.89
R243 VDD.n152 VDD.n149 2.89
R244 VDD.n83  2.557
R245 VDD.n217  |�P� 2.557
R246 VDD.n158 ��8V 2.557
R247 VDD.n72 VDD.n69 2.477
R248 VDD.n174 VDD.n171 2.477
R249 VDD.n27 VDD.n24 2.064
R250 VDD.n36 VDD.n35 2.064
R251 VDD.n68 VDD.n41 0.29
R252 VDD.n125 VDD.n99 0.29
R253 VDD.n206 VDD.n179 0.29
R254 VDD.n148 VDD 0.207
R255 VDD.n86 VDD.n82 0.181
R256 VDD.n223 VDD.n220 0.181
R257 VDD.n166 VDD.n161 0.181
R258 VDD.n32 VDD.n28 0.157
R259 VDD.n37 VDD.n32 0.157
R260 VDD.n41 VDD.n37 0.145
R261 VDD.n73 VDD.n68 0.145
R262 VDD.n77 VDD.n73 0.145
R263 VDD.n82 VDD.n77 0.145
R264 VDD.n90 VDD.n86 0.145
R265 VDD.n95 VDD.n90 0.145
R266 VDD.n99 VDD.n95 0.145
R267 VDD.n231 VDD.n227 0.145
R268 VDD.n227 VDD.n223 0.145
R269 VDD.n220 VDD.n216 0.145
R270 VDD.n216 VDD.n210 0.145
R271 VDD.n210 VDD.n206 0.145
R272 VDD.n179 VDD.n175 0.145
R273 VDD.n175 VDD.n170 0.145
R274 VDD.n170 VDD.n166 0.145
R275 VDD.n161 VDD.n157 0.145
R276 VDD.n157 VDD.n153 0.145
R277 VDD.n153 VDD.n148 0.145
R278 VDD VDD.n125 0.078
R279 VDD VDD.n231 0.066
R280 a_797_1051.n0 a_797_1051.t0 228.369
R281 a_797_1051.n0 a_797_1051.t3 219.778
R282 a_797_1051.n1 a_797_1051.n0 42.29
R283 a_797_1051.n1 a_797_1051.t1 14.282
R284 a_797_1051.t2 a_797_1051.n1 14.282
R285 a_1549_1050.n4 a_1549_1050.t6 512.525
R286 a_1549_1050.n4 a_1549_1050.t5 371.139
R287 a_1549_1050.n5 a_1549_1050.n4 303.065
R288 a_1549_1050.n6 a_1549_1050.n3 243.576
R289 a_1549_1050.n5 a_1549_1050.t7 227.134
R290 a_1549_1050.n8 a_1549_1050.n6 222.004
R291 a_1549_1050.n3 a_1549_1050.n2 157.964
R292 a_1549_1050.n3 a_1549_1050.n1 91.706
R293 a_1549_1050.n8 a_1549_1050.n7 30
R294 a_1549_1050.n9 a_1549_1050.n0 24.383
R295 a_1549_1050.n9 a_1549_1050.n8 23.684
R296 a_1549_1050.n1 a_1549_1050.t2 14.282
R297 a_1549_1050.n1 a_1549_1050.t1 14.282
R298 a_1549_1050.n2 a_1549_1050.t4 14.282
R299 a_1549_1050.n2 a_1549_1050.t3 14.282
R300 a_1549_1050.n6 a_1549_1050.n5 10.343
R301 Y.n5 Y.n0 299.141
R302 Y.n5 Y.n4 244.592
R303 Y.n4 Y.n3 30
R304 Y.n2 Y.n1 24.383
R305 Y.n4 Y.n2 23.684
R306 Y.n0 Y.t1 14.282
R307 Y.n0 Y.t2 14.282
R308 Y.n6 Y.n5 4.65
R309 Y.n6 Y 0.046
R310 B.n0 B.t0 472.359
R311 B.n0 B.t1 384.527
R312 B.n1 B.t2 287.037
R313 B.n1 B.n0 210.673
R314 B.n2 B.n1 4.65
R315 B.n2 B 0.046
R316 a_864_209.n1 a_864_209.t4 480.392
R317 a_864_209.n1 a_864_209.t6 403.272
R318 a_864_209.n3 a_864_209.n0 343.684
R319 a_864_209.n2 a_864_209.t5 273.627
R320 a_864_209.n2 a_864_209.n1 254.865
R321 a_864_209.n8 a_864_209.n7 208.452
R322 a_864_209.n10 a_864_209.n8 142.275
R323 a_864_209.n8 a_864_209.n3 86.587
R324 a_864_209.n7 a_864_209.n6 30
R325 a_864_209.n5 a_864_209.n4 24.383
R326 a_864_209.n7 a_864_209.n5 23.684
R327 a_864_209.n10 a_864_209.n9 15.001
R328 a_864_209.n0 a_864_209.t0 14.282
R329 a_864_209.n0 a_864_209.t2 14.282
R330 a_864_209.n11 a_864_209.n10 12.632
R331 a_864_209.n3 a_864_209.n2 10.615
R332 C.n0 C.t0 470.752
R333 C.n0 C.t1 384.527
R334 C.n1 C.t2 314.896
R335 C.n1 C.n0 182.932
R336 C.n2 C.n1 4.65
R337 C.n2 C 0.046
R338 a_112_101.n10 a_112_101.n9 93.333
R339 a_112_101.n12 a_112_101.n11 68.43
R340 a_112_101.n3 a_112_101.n2 51.907
R341 a_112_101.n3 a_112_101.n1 51.594
R342 a_112_101.t0 a_112_101.n3 38.864
R343 a_112_101.n7 a_112_101.n6 38.626
R344 a_112_101.n6 a_112_101.n5 35.955
R345 a_112_101.t1 a_112_101.n8 8.137
R346 a_112_101.t0 a_112_101.n0 6.109
R347 a_112_101.t1 a_112_101.n7 4.864
R348 a_112_101.t0 a_112_101.n4 3.871
R349 a_112_101.t0 a_112_101.n13 2.535
R350 a_112_101.n13 a_112_101.t1 1.145
R351 a_112_101.t1 a_112_101.n12 0.763
R352 a_112_101.n12 a_112_101.n10 0.185
R353 GND.n65 GND.n64 237.558
R354 GND.n95 GND.n94 237.558
R355 GND.n32 GND.n31 237.558
R356 GND.n29 GND.n28 210.82
R357 GND.n97 GND.n96 210.82
R358 GND.n62 GND.n61 210.82
R359 GND.n75 GND.n74 172.612
R360 GND.n51 GND.n50 151.605
R361 GND.n119 GND.n118 40.431
R362 GND.n130 GND.n129 40.003
R363 GND.n21 GND.n20 37.582
R364 GND.n104 GND.n103 37.582
R365 GND.t3 GND.n18 32.601
R366 GND.n50 GND.n49 28.421
R367 GND.n50 GND.n48 25.263
R368 GND.n48 GND.n47 24.383
R369 GND.n18 GND.n17 21.734
R370 GND.n4 GND.n3 20.705
R371 GND.n10 GND.n9 20.705
R372 GND.n22 GND.n21 20.705
R373 GND.n109 GND.n108 20.705
R374 GND.n120 GND.n119 20.705
R375 GND.n125 GND.n124 20.705
R376 GND.n131 GND.n130 20.705
R377 GND.n105 GND.n104 20.705
R378 GND.n3 GND.n2 19.952
R379 GND.n30 GND.n29 18.953
R380 GND.n98 GND.n97 18.953
R381 GND.n63 GND.n62 18.953
R382 GND.n129 GND.n128 17.258
R383 GND.n20 GND.t3 15.644
R384 GND.n103 GND.t6 15.644
R385 GND.n33 GND.n30 14.864
R386 GND.n66 GND.n63 14.864
R387 GND.n99 GND.n98 14.864
R388 GND.n118 GND.t0 13.654
R389 GND.n20 GND.n19 13.541
R390 GND.n103 GND.n102 13.541
R391 GND.n121 GND.n120 9.29
R392 GND.n72 GND.n71 9.154
R393 GND.n77 GND.n76 9.154
R394 GND.n80 GND.n79 9.154
R395 GND.n83 GND.n82 9.154
R396 GND.n86 GND.n85 9.154
R397 GND.n89 GND.n88 9.154
R398 GND.n92 GND.n91 9.154
R399 GND.n99 GND.n95 9.154
R400 GND.n106 GND.n101 9.154
R401 GND.n111 GND.n110 9.154
R402 GND.n114 GND.n113 9.154
R403 GND.n121 GND.n116 9.154
R404 GND.n126 GND.n123 9.154
R405 GND.n133 GND.n132 9.154
R406 GND.n66 GND.n65 9.154
R407 GND.n59 GND.n58 9.154
R408 GND.n56 GND.n55 9.154
R409 GND.n53 GND.n52 9.154
R410 GND.n45 GND.n44 9.154
R411 GND.n42 GND.n41 9.154
R412 GND.n39 GND.n38 9.154
R413 GND.n36 GND.n35 9.154
R414 GND.n33 GND.n32 9.154
R415 GND.n26 GND.n25 9.154
R416 GND.n23 GND.n14 9.154
R417 GND.n12 GND.n11 9.154
R418 GND.n6 GND.n5 9.154
R419 GND.t0 GND.n117 7.04
R420 GND.n7 GND.n1 4.795
R421 GND.n70 GND.n69 4.65
R422 GND.n7 GND.n6 4.65
R423 GND.n13 GND.n12 4.65
R424 GND.n24 GND.n23 4.65
R425 GND.n27 GND.n26 4.65
R426 GND.n34 GND.n33 4.65
R427 GND.n37 GND.n36 4.65
R428 GND.n40 GND.n39 4.65
R429 GND.n43 GND.n42 4.65
R430 GND.n46 GND.n45 4.65
R431 GND.n54 GND.n53 4.65
R432 GND.n57 GND.n56 4.65
R433 GND.n60 GND.n59 4.65
R434 GND.n67 GND.n66 4.65
R435 GND.n134 GND.n133 4.65
R436 GND.n127 GND.n126 4.65
R437 GND.n122 GND.n121 4.65
R438 GND.n115 GND.n114 4.65
R439 GND.n112 GND.n111 4.65
R440 GND.n107 GND.n106 4.65
R441 GND.n100 GND.n99 4.65
R442 GND.n93 GND.n92 4.65
R443 GND.n90 GND.n89 4.65
R444 GND.n87 GND.n86 4.65
R445 GND.n84 GND.n83 4.65
R446 GND.n81 GND.n80 4.65
R447 GND.n78 GND.n77 4.65
R448 GND.n73 GND.n72 4.65
R449 GND.n16 GND.n15 4.504
R450 GND.n6 GND.n4 4.129
R451 GND.n53 GND.n51 4.129
R452 GND.n126 GND.n125 4.129
R453 GND.n111 GND.n109 4.129
R454 GND.n77 GND.n75 4.129
R455 GND.n23 GND.n22 3.716
R456 GND.t3 GND.n16 2.452
R457 GND.n133 GND.n131 1.032
R458 GND.n106 GND.n105 1.032
R459 GND.n1 GND.n0 0.474
R460 GND.n69 GND.n68 0.474
R461 GND.n9 GND.n8 0.376
R462 GND.n34 GND.n27 0.29
R463 GND.n67 GND.n60 0.29
R464 GND.n100 GND.n93 0.29
R465 GND.n70 GND 0.207
R466 GND.n12 GND.n10 0.206
R467 GND.n46 GND.n43 0.181
R468 GND.n122 GND.n115 0.181
R469 GND.n84 GND.n81 0.181
R470 GND.n13 GND.n7 0.157
R471 GND.n24 GND.n13 0.157
R472 GND.n27 GND.n24 0.145
R473 GND.n37 GND.n34 0.145
R474 GND.n40 GND.n37 0.145
R475 GND.n43 GND.n40 0.145
R476 GND.n54 GND.n46 0.145
R477 GND.n57 GND.n54 0.145
R478 GND.n60 GND.n57 0.145
R479 GND.n134 GND.n127 0.145
R480 GND.n127 GND.n122 0.145
R481 GND.n115 GND.n112 0.145
R482 GND.n112 GND.n107 0.145
R483 GND.n107 GND.n100 0.145
R484 GND.n93 GND.n90 0.145
R485 GND.n90 GND.n87 0.145
R486 GND.n87 GND.n84 0.145
R487 GND.n81 GND.n78 0.145
R488 GND.n78 GND.n73 0.145
R489 GND.n73 GND.n70 0.145
R490 GND GND.n67 0.078
R491 GND GND.n134 0.066
R492 a_1444_101.n3 a_1444_101.n1 42.788
R493 a_1444_101.t0 a_1444_101.n0 8.137
R494 a_1444_101.n3 a_1444_101.n2 4.665
R495 a_1444_101.t0 a_1444_101.n3 0.06
R496 D.n0 D.t0 472.359
R497 D.n0 D.t2 384.527
R498 D.n1 D.t1 342.755
R499 D.n1 D.n0 154.955
R500 D.n2 D.n1 4.65
R501 D.n2 D 0.046
C6 VDD GND 4.31fF
C7 a_1444_101.n0 GND 0.05fF
C8 a_1444_101.n1 GND 0.12fF
C9 a_1444_101.n2 GND 0.04fF
C10 a_1444_101.n3 GND 0.17fF
C11 a_112_101.n0 GND 0.02fF
C12 a_112_101.n1 GND 0.09fF
C13 a_112_101.n2 GND 0.07fF
C14 a_112_101.n3 GND 0.04fF
C15 a_112_101.n4 GND 0.01fF
C16 a_112_101.n5 GND 0.04fF
C17 a_112_101.n6 GND 0.04fF
C18 a_112_101.n7 GND 0.02fF
C19 a_112_101.n8 GND 0.05fF
C20 a_112_101.n9 GND 0.02fF
C21 a_112_101.n10 GND 0.14fF
C22 a_112_101.n11 GND 0.08fF
C23 a_112_101.n12 GND 0.08fF
C24 a_112_101.t1 GND 0.22fF
C25 a_112_101.n13 GND 0.01fF
C26 a_864_209.n0 GND 0.50fF
C27 a_864_209.n1 GND 0.32fF
C28 a_864_209.n2 GND 0.46fF
C29 a_864_209.n3 GND 0.52fF
C30 a_864_209.n4 GND 0.03fF
C31 a_864_209.n5 GND 0.04fF
C32 a_864_209.n6 GND 0.03fF
C33 a_864_209.n7 GND 0.09fF
C34 a_864_209.n8 GND 0.31fF
C35 a_864_209.n9 GND 0.06fF
C36 a_864_209.n10 GND 0.04fF
C37 a_864_209.n11 GND 0.04fF
C38 Y.n0 GND 0.68fF
C39 Y.n1 GND 0.04fF
C40 Y.n2 GND 0.05fF
C41 Y.n3 GND 0.03fF
C42 Y.n4 GND 0.16fF
C43 Y.n5 GND 0.62fF
C44 Y.n6 GND 0.01fF
C45 a_1549_1050.n0 GND 0.03fF
C46 a_1549_1050.n1 GND 0.29fF
C47 a_1549_1050.n2 GND 0.37fF
C48 a_1549_1050.n3 GND 0.50fF
C49 a_1549_1050.n4 GND 0.30fF
C50 a_1549_1050.n5 GND 0.43fF
C51 a_1549_1050.n6 GND 0.48fF
C52 a_1549_1050.n7 GND 0.03fF
C53 a_1549_1050.n8 GND 0.10fF
C54 a_1549_1050.n9 GND 0.04fF
C55 a_797_1051.n0 GND 0.52fF
C56 a_797_1051.n1 GND 0.22fF
C57 VDD.n1 GND 0.03fF
C58 VDD.n2 GND 0.08fF
C59 VDD.n3 GND 0.02fF
C60 VDD.n4 GND 0.02fF
C61 VDD.n5 GND 0.05fF
C62 VDD.n6 GND 0.02fF
C63 VDD.n7 GND 0.02fF
C64 VDD.n8 GND 0.02fF
C65 VDD.n9 GND 0.02fF
C66 VDD.n10 GND 0.02fF
C67 VDD.n11 GND 0.02fF
C68 VDD.n12 GND 0.02fF
C69 VDD.n13 GND 0.02fF
C70 VDD.n14 GND 0.03fF
C71 VDD.n15 GND 0.01fF
C72 VDD.n20 GND 0.38fF
C73 VDD.n21 GND 0.23fF
C74 VDD.n22 GND 0.02fF
C75 VDD.n23 GND 0.03fF
C76 VDD.n24 GND 0.05fF
C77 VDD.n25 GND 0.17fF
C78 VDD.n26 GND 0.01fF
C79 VDD.n27 GND 0.01fF
C80 VDD.n28 GND 0.06fF
C81 VDD.n29 GND 0.14fF
C82 VDD.n30 GND 0.01fF
C83 VDD.n31 GND 0.02fF
C84 VDD.n32 GND 0.02fF
C85 VDD.n33 GND 0.17fF
C86 VDD.n34 GND 0.01fF
C87 VDD.n35 GND 0.05fF
C88 VDD.n36 GND 0.01fF
C89 VDD.n37 GND 0.02fF
C90 VDD.n38 GND 0.23fF
C91 VDD.n39 GND 0.01fF
C92 VDD.n40 GND 0.02fF
C93 VDD.n41 GND 0.03fF
C94 VDD.n42 GND 0.05fF
C95 VDD.n43 GND 0.02fF
C96 VDD.n44 GND 0.02fF
C97 VDD.n45 GND 0.02fF
C98 VDD.n46 GND 0.02fF
C99 VDD.n47 GND 0.02fF
C100 VDD.n48 GND 0.02fF
C101 VDD.n49 GND 0.02fF
C102 VDD.n50 GND 0.02fF
C103 VDD.n51 GND 0.02fF
C104 VDD.n52 GND 0.02fF
C105 VDD.n53 GND 0.01fF
C106 VDD.n54 GND 0.02fF
C107 VDD.n55 GND 0.02fF
C108 VDD.n56 GND 0.15fF
C109 VDD.n57 GND 0.02fF
C110 VDD.n58 GND 0.02fF
C111 VDD.n60 GND 0.02fF
C112 VDD.n64 GND 0.23fF
C113 VDD.n65 GND 0.23fF
C114 VDD.n66 GND 0.01fF
C115 VDD.n67 GND 0.02fF
C116 VDD.n68 GND 0.03fF
C117 VDD.n69 GND 0.05fF
C118 VDD.n70 GND 0.20fF
C119 VDD.n71 GND 0.01fF
C120 VDD.n72 GND 0.01fF
C121 VDD.n73 GND 0.02fF
C122 VDD.n74 GND 0.14fF
C123 VDD.n75 GND 0.01fF
C124 VDD.n76 GND 0.02fF
C125 VDD.n77 GND 0.02fF
C126 VDD.n78 GND 0.07fF
C127 VDD.n79 GND 0.04fF
C128 VDD.n80 GND 0.01fF
C129 VDD.n81 GND 0.02fF
C130 VDD.n82 GND 0.02fF
C131 VDD.n83 GND 0.12fF
C132 VDD.n84 GND 0.01fF
C133 VDD.n85 GND 0.02fF
C134 VDD.n86 GND 0.02fF
C135 VDD.n87 GND 0.14fF
C136 VDD.n88 GND 0.01fF
C137 VDD.n89 GND 0.02fF
C138 VDD.n90 GND 0.02fF
C139 VDD.n91 GND 0.05fF
C140 VDD.n92 GND 0.20fF
C141 VDD.n93 GND 0.01fF
C142 VDD.n94 GND 0.01fF
C143 VDD.n95 GND 0.02fF
C144 VDD.n96 GND 0.23fF
C145 VDD.n97 GND 0.01fF
C146 VDD.n98 GND 0.02fF
C147 VDD.n99 GND 0.03fF
C148 VDD.n100 GND 0.18fF
C149 VDD.n101 GND 0.02fF
C150 VDD.n102 GND 0.02fF
C151 VDD.n103 GND 0.02fF
C152 VDD.n104 GND 0.05fF
C153 VDD.n105 GND 0.02fF
C154 VDD.n106 GND 0.02fF
C155 VDD.n107 GND 0.02fF
C156 VDD.n108 GND 0.02fF
C157 VDD.n109 GND 0.02fF
C158 VDD.n110 GND 0.02fF
C159 VDD.n111 GND 0.02fF
C160 VDD.n112 GND 0.02fF
C161 VDD.n113 GND 0.02fF
C162 VDD.n114 GND 0.01fF
C163 VDD.n115 GND 0.02fF
C164 VDD.n116 GND 0.02fF
C165 VDD.n117 GND 0.02fF
C166 VDD.n121 GND 0.23fF
C167 VDD.n122 GND 0.23fF
C168