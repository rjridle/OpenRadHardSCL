magic
tech sky130A
magscale 1 2
timestamp 1645052634
<< nmos >>
rect 125 181 155 243
tri 29 151 59 181 se
rect 59 151 155 181
rect 29 59 59 151
tri 59 135 75 151 nw
tri 109 135 125 151 ne
tri 59 59 75 75 sw
tri 109 59 125 75 se
rect 125 59 155 151
tri 29 29 59 59 ne
rect 59 29 125 59
tri 125 29 155 59 nw
<< ndiff >>
rect -27 227 125 243
rect -27 193 -17 227
rect 17 193 125 227
rect -27 181 125 193
rect 155 227 211 243
rect 155 193 167 227
rect 201 193 211 227
rect -27 29 29 181
tri 29 151 59 181 nw
rect 155 156 211 193
tri 59 135 75 151 se
rect 75 135 109 151
tri 109 135 125 151 sw
rect 59 122 125 135
rect 59 88 75 122
rect 109 88 125 122
rect 59 75 125 88
tri 59 59 75 75 ne
rect 75 59 109 75
tri 109 59 125 75 nw
rect 155 122 167 156
rect 201 122 211 156
rect 155 88 211 122
tri 29 29 59 59 sw
tri 125 29 155 59 se
rect 155 54 167 88
rect 201 54 211 88
rect 155 29 211 54
rect -27 17 211 29
rect -27 -17 -17 17
rect 17 -17 71 17
rect 105 -17 167 17
rect 201 -17 211 17
rect -27 -33 211 -17
<< ndiffc >>
rect -17 193 17 227
rect 167 193 201 227
rect 75 88 109 122
rect 167 122 201 156
rect 167 54 201 88
rect -17 -17 17 17
rect 71 -17 105 17
rect 167 -17 201 17
<< poly >>
rect 125 243 155 269
<< locali >>
rect -17 227 17 243
rect 167 227 201 243
rect 17 193 167 227
rect -17 175 17 193
rect 167 156 201 193
rect 75 122 109 138
rect -17 88 75 122
rect 75 72 109 88
rect 167 88 201 122
rect -17 17 17 35
rect 167 17 201 54
rect 17 -17 71 17
rect 105 -17 167 17
rect -17 -33 17 -17
rect 167 -33 201 -17
<< end >>
