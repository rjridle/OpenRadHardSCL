* SPICE3 file created from INVX3.ext - technology: sky130A

.subckt INVX3 VDD A VSS Y
M1000 Y A VDD VDD pshort w=3u l=0.15u
+  ad=1.71p pd=13.14u as=1.71p ps=13.14u
M1001 Y A VSS VSS nshort w=3u l=0.15u
+  ad=0.1588p pd=1.5u as=1.094p ps=7.96u
M1002 Y A VDD VDD pshort w=3u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 VDD A Y VDD pshort w=3u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
.ends
