magic
tech sky130A
magscale 1 2
timestamp 1647338072
<< locali >>
rect 797 551 831 781
rect 1389 551 1423 855
<< metal1 >>
rect 55 1505 89 1539
rect 131 871 165 905
rect 167 871 1358 905
rect 1611 649 1645 683
rect 1351 575 2019 609
rect 2055 575 2089 609
rect 1425 501 1503 535
rect 55 13 89 47
use li1_M1_contact  li1_M1_contact_3 pcells
timestamp 1646004885
transform 1 0 1554 0 1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_2
timestamp 1646004885
transform 1 0 2072 0 1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_7
timestamp 1646004885
transform -1 0 1332 0 -1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_8
timestamp 1646004885
transform 1 0 888 0 1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_6
timestamp 1646004885
transform -1 0 814 0 -1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_5
timestamp 1646004885
transform -1 0 814 0 -1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1646004885
transform -1 0 1406 0 -1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_9
timestamp 1646004885
transform 1 0 1406 0 1 888
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_1
timestamp 1646004885
transform -1 0 148 0 -1 888
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_4
timestamp 1646004885
transform 1 0 888 0 1 888
box -53 -33 29 33
use xor2X1_pcell  xor2X1_pcell_0 pcells
timestamp 1647338052
transform 1 0 0 0 1 0
box -84 0 2304 1575
<< labels >>
rlabel metal1 72 1522 72 1522 1 VDD
port 4 n
rlabel metal1 72 30 72 30 1 VSS
port 5 n
rlabel metal1 55 1505 89 1539 1 VDD
rlabel metal1 55 13 89 47 1 VSS
rlabel metal1 2055 575 2089 609 1 B
rlabel metal1 1611 649 1645 683 1 Y
rlabel metal1 131 871 165 905 1 A
<< end >>
