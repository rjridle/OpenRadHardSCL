* SPICE3 file created from AOAI4X1.ext - technology: sky130A

.subckt AOAI4X1 YN A B C D VDD GND
X0 VDD.t21 A.t0 a_217_1050.t3  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X1 VDD.t17 a_217_1050.t5 a_797_1051.t3 VDD.t16 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X2 VDD.t11 B.t0 a_217_1050.t2 ,O�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X3 VDD.t9 a_864_209.t4 YN.t4  ,O�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X4 GND A.t1 a_112_101.t0 GND sky130_fd_pr__nfet_01v8 ad=2.2948p pd=1.608u as=0p ps=0u w=0u l=0u
X5 GND a_864_209.t5 a_1444_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X6 YN D.t1 a_1444_101.t0 GND sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=0p ps=0u w=0u l=0u
X7 a_797_1051.t0 C.t0 a_864_209.t0 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X8 a_217_1050.t4 A.t2 VDD.t19  ,O�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X9 a_797_1051.t2 a_217_1050.t7 VDD.t15 �+O�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X10 VDD.t13 D.t0 YN.t1  ,O�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X11 a_217_1050.t1 B.t1 VDD.t3 �+O�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X12 YN.t3 a_864_209.t6 VDD.t1  ,O�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X13 a_864_209.t1 C.t1 a_797_1051.t1 �+O�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X14 YN.t0 D.t2 VDD.t5  ,O�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
C0 D VDD 0.33fF
C1 B VDD 0.32fF
C2 C VDD 0.32fF
C3 YN D 0.26fF
C4 B A 0.27fF
C5 YN VDD 1.82fF
C6 VDD A 0.32fF
R0 A.n0 A.t0 480.392
R1 A.n0 A.t2 403.272
R2 A.n1 A.t1 301.486
R3 A.n1 A.n0 227.006
R4 A.n2 A.n1 4.65
R5 A.n2 A 0.046
R6 a_217_1050.n3 a_217_1050.t7 486.819
R7 a_217_1050.n3 a_217_1050.t5 384.527
R8 a_217_1050.n4 a_217_1050.t6 267.201
R9 a_217_1050.n4 a_217_1050.n3 262.705
R10 a_217_1050.n5 a_217_1050.n2 243.576
R11 a_217_1050.n7 a_217_1050.n5 228.526
R12 a_217_1050.n2 a_217_1050.n1 157.964
R13 a_217_1050.n2 a_217_1050.n0 91.706
R14 a_217_1050.n7 a_217_1050.n6 15.218
R15 a_217_1050.n0 a_217_1050.t2 14.282
R16 a_217_1050.n0 a_217_1050.t1 14.282
R17 a_217_1050.n1 a_217_1050.t3 14.282
R18 a_217_1050.n1 a_217_1050.t4 14.282
R19 a_217_1050.n8 a_217_1050.n7 12.014
R20 a_217_1050.n5 a_217_1050.n4 10.615
R21 VDD.n79 VDD.n68 144.705
R22 VDD.n171 VDD.n160 144.705
R23 VDD.n138 VDD.t11 143.754
R24 VDD.n24 VDD.t13 143.754
R25 VDD.n116 VDD.t19 135.17
R26 VDD.n46 VDD.t1 135.17
R27 VDD.n179 VDD.n178 129.849
R28 VDD.n130 VDD.n129 129.472
R29 VDD.n34 VDD.n33 129.472
R30 VDD.n64 VDD.n63 92.5
R31 VDD.n62 VDD.n61 92.5
R32 VDD.n60 VDD.n59 92.5
R33 VDD.n58 VDD.n57 92.5
R34 VDD.n66 VDD.n65 92.5
R35 VDD.n156 VDD.n155 92.5
R36 VDD.n154 VDD.n153 92.5
R37 VDD.n152 VDD.n151 92.5
R38 VDD.n150 VDD.n149 92.5
R39 VDD.n158 VDD.n157 92.5
R40 VDD.n104 VDD.n103 92.5
R41 VDD.n102 VDD.n101 92.5
R42 VDD.n100 VDD.n99 92.5
R43 VDD.n98 VDD.n97 92.5
R44 VDD.n106 VDD.n105 92.5
R45 VDD.n14 VDD.n1 92.5
R46 VDD.n5 VDD.n4 92.5
R47 VDD.n7 VDD.n6 92.5
R48 VDD.n9 VDD.n8 92.5
R49 VDD.n11 VDD.n10 92.5
R50 VDD.n13 VDD.n12 92.5
R51 VDD.n21 VDD.n20 92.059
R52 VDD.n78 VDD.n77 92.059
R53 VDD.n170 VDD.n169 92.059
R54 VDD.n112 VDD.n111 92.059
R55 VDD.n20 VDD.n16 67.194
R56 VDD.n20 VDD.n17 67.194
R57 VDD.n20 VDD.n18 67.194
R58 VDD.n20 VDD.n19 67.194
R59 VDD.n96 VDD.n95 44.141
R60 VDD.n5 VDD.n3 44.141
R61 VDD.n95 VDD.n93 44.107
R62 VDD.n3 VDD.n2 44.107
R63 VDD.n20 VDD.n15 41.052
R64 VDD.n72 VDD.n70 39.742
R65 VDD.n72 VDD.n71 39.742
R66 VDD.n74 VDD.n73 39.742
R67 VDD.n108 VDD.n107 39.742
R68 VDD.n168 VDD.n165 39.742
R69 VDD.n168 VDD.n167 39.742
R70 VDD.n164 VDD.n163 39.742
R71 VDD.n95 VDD.n94 38
R72 VDD.n70 VDD.n69 36.774
R73 VDD.n167 VDD.n166 36.774
R74 VDD.n1 VDD.n0 30.923
R75 VDD.n77 VDD.n75 26.38
R76 VDD.n77 VDD.n74 26.38
R77 VDD.n77 VDD.n72 26.38
R78 VDD.n77 VDD.n76 26.38
R79 VDD.n111 VDD.n109 26.38
R80 VDD.n111 VDD.n108 26.38
R81 VDD.n111 VDD.n110 26.38
R82 VDD.n169 VDD.n168 26.38
R83 VDD.n169 VDD.n164 26.38
R84 VDD.n169 VDD.n162 26.38
R85 VDD.n169 VDD.n161 26.38
R86 VDD.n114 VDD.n106 22.915
R87 VDD.n23 VDD.n14 22.915
R88 VDD.n29  ,O�� 20.457
R89 VDD.n86 VDD.t6 20.457
R90 VDD.n134 ,O�� 20.457
R91 VDD.n42  ,O�� 17.9
R92 VDD.n180 VDD.t16 17.9
R93 VDD.n121  ,O�� 17.9
R94 VDD.n106 VDD.n104 14.864
R95 VDD.n104 VDD.n102 14.864
R96 VDD.n102 VDD.n100 14.864
R97 VDD.n100 VDD.n98 14.864
R98 VDD.n98 VDD.n96 14.864
R99 VDD.n66 VDD.n64 14.864
R100 VDD.n64 VDD.n62 14.864
R101 VDD.n62 VDD.n60 14.864
R102 VDD.n60 VDD.n58 14.864
R103 VDD.n58 VDD.n56 14.864
R104 VDD.n56 VDD.n55 14.864
R105 VDD.n158 VDD.n156 14.864
R106 VDD.n156 VDD.n154 14.864
R107 VDD.n154 VDD.n152 14.864
R108 VDD.n152 VDD.n150 14.864
R109 VDD.n150 VDD.n148 14.864
R110 VDD.n148 VDD.n147 14.864
R111 VDD.n14 VDD.n13 14.864
R112 VDD.n13 VDD.n11 14.864
R113 VDD.n11 VDD.n9 14.864
R114 VDD.n9 VDD.n7 14.864
R115 VDD.n7 VDD.n5 14.864
R116 VDD.n80 VDD.n67 14.864
R117 VDD.n172 VDD.n159 14.864
R118 VDD.n129 VDD.t3 14.282
R119 VDD.n129 VDD.t21 14.282
R120 VDD.n178 VDD.t15 14.282
R121 VDD.n178 VDD.t17 14.282
R122 VDD.n33 VDD.t5 14.282
R123 VDD.n33 VDD.t9 14.282
R124 VDD.n36 VDD.n34 9.083
R125 VDD.n132 VDD.n130 9.083
R126 VDD.n23 VDD.n22 8.855
R127 VDD.n22 VDD.n21 8.855
R128 VDD.n27 VDD.n26 8.855
R129 VDD.n26 VDD.n25 8.855
R130 VDD.n31 VDD.n30 8.855
R131 VDD.n30 VDD.n29 8.855
R132 VDD.n36 VDD.n35 8.855
R133 VDD.n35  ,O�� 8.855
R134 VDD.n40 VDD.n39 8.855
R135 VDD.n39 VDD.n38 8.855
R136 VDD.n44 VDD.n43 8.855
R137 VDD.n43 VDD.n42 8.855
R138 VDD.n49 VDD.n48 8.855
R139 VDD.n48 VDD.n47 8.855
R140 VDD.n53 VDD.n52 8.855
R141 VDD.n52 VDD.n51 8.855
R142 VDD.n80 VDD.n79 8.855
R143 VDD.n79 VDD.n78 8.855
R144 VDD.n84 VDD.n83 8.855
R145 VDD.n83 VDD.n82 8.855
R146 VDD.n88 VDD.n87 8.855
R147 VDD.n87 VDD.n86 8.855
R148 VDD.n91 VDD.n90 8.855
R149 VDD.n90 �+O�� 8.855
R150 VDD.n186 VDD.n185 8.855
R151 VDD.n185 VDD.n184 8.855
R152 VDD.n182 VDD.n181 8.855
R153 VDD.n181 VDD.n180 8.855
R154 VDD.n176 VDD.n175 8.855
R155 VDD.n175 VDD.n174 8.855
R156 VDD.n172 VDD.n171 8.855
R157 VDD.n171 VDD.n170 8.855
R158 VDD.n145 VDD.n144 8.855
R159 VDD.n144 VDD.n143 8.855
R160 VDD.n141 VDD.n140 8.855
R161 VDD.n140 VDD.n139 8.855
R162 VDD.n136 VDD.n135 8.855
R163 VDD.n135 VDD.n134 8.855
R164 VDD.n132 VDD.n131 8.855
R165 VDD.n131 �+O�� 8.855
R166 VDD.n127 VDD.n126 8.855
R167 VDD.n126 VDD.n125 8.855
R168 VDD.n123 VDD.n122 8.855
R169 VDD.n122 VDD.n121 8.855
R170 VDD.n119 VDD.n118 8.855
R171 VDD.n118 VDD.n117 8.855
R172 VDD.n114 VDD.n113 8.855
R173 VDD.n113 VDD.n112 8.855
R174 VDD.n67 VDD.n66 8.051
R175 VDD.n159 VDD.n158 8.051
R176 VDD.n182 VDD.n179 6.193
R177 VDD.n32 VDD.n31 4.65
R178 VDD.n37 VDD.n36 4.65
R179 VDD.n41 VDD.n40 4.65
R180 VDD.n45 VDD.n44 4.65
R181 VDD.n50 VDD.n49 4.65
R182 VDD.n54 VDD.n53 4.65
R183 VDD.n81 VDD.n80 4.65
R184 VDD.n85 VDD.n84 4.65
R185 VDD.n89 VDD.n88 4.65
R186 VDD.n92 VDD.n91 4.65
R187 VDD.n187 VDD.n186 4.65
R188 VDD.n183 VDD.n182 4.65
R189 VDD.n177 VDD.n176 4.65
R190 VDD.n173 VDD.n172 4.65
R191 VDD.n146 VDD.n145 4.65
R192 VDD.n142 VDD.n141 4.65
R193 VDD.n137 VDD.n136 4.65
R194 VDD.n133 VDD.n132 4.65
R195 VDD.n128 VDD.n127 4.65
R196 VDD.n124 VDD.n123 4.65
R197 VDD.n120 VDD.n119 4.65
R198 VDD.n115 VDD.n114 4.65
R199 VDD.n28 VDD.n23 2.933
R200 VDD.n49 VDD.n46 2.89
R201 VDD.n119 VDD.n116 2.89
R202 VDD.n28 VDD.n27 2.844
R203 VDD.n38  ,O�� 2.557
R204 VDD.n184 �+O�� 2.557
R205 VDD.n125 �B�gU 2.557
R206 VDD.n27 VDD.n24 2.477
R207 VDD.n141 VDD.n138 2.477
R208 VDD.n32 VDD.n28 1.063
R209 VDD.n81 VDD.n54 0.29
R210 VDD.n173 VDD.n146 0.29
R211 VDD.n115 VDD 0.207
R212 VDD.n41 VDD.n37 0.181
R213 VDD.n133 VDD.n128 0.181
R214 VDD.n37 VDD.n32 0.145
R215 VDD.n45 VDD.n41 0.145
R216 VDD.n50 VDD.n45 0.145
R217 VDD.n54 VDD.n50 0.145
R218 VDD.n85 VDD.n81 0.145
R219 VDD.n89 VDD.n85 0.145
R220 VDD.n92 VDD.n89 0.145
R221 VDD.n187 VDD.n183 0.145
R222 VDD.n183 VDD.n177 0.145
R223 VDD.n177 VDD.n173 0.145
R224 VDD.n146 VDD.n142 0.145
R225 VDD.n142 VDD.n137 0.145
R226 VDD.n137 VDD.n133 0.145
R227 VDD.n128 VDD.n124 0.145
R228 VDD.n124 VDD.n120 0.145
R229 VDD.n120 VDD.n115 0.145
R230 VDD VDD.n92 0.09
R231 VDD VDD.n187 0.09
R232 a_797_1051.n0 a_797_1051.t0 228.369
R233 a_797_1051.n0 a_797_1051.t3 219.778
R234 a_797_1051.n1 a_797_1051.n0 42.29
R235 a_797_1051.n1 a_797_1051.t1 14.282
R236 a_797_1051.t2 a_797_1051.n1 14.282
R237 B.n0 B.t0 472.359
R238 B.n0 B.t1 384.527
R239 B.n1 B.t2 287.037
R240 B.n1 B.n0 210.673
R241 B.n2 B.n1 4.65
R242 B.n2 B 0.046
R243 a_864_209.n1 a_864_209.t4 480.392
R244 a_864_209.n1 a_864_209.t6 403.272
R245 a_864_209.n3 a_864_209.n0 343.684
R246 a_864_209.n2 a_864_209.t5 273.627
R247 a_864_209.n2 a_864_209.n1 254.865
R248 a_864_209.n8 a_864_209.n7 208.452
R249 a_864_209.n10 a_864_209.n8 142.275
R250 a_864_209.n8 a_864_209.n3 86.587
R251 a_864_209.n7 a_864_209.n6 30
R252 a_864_209.n5 a_864_209.n4 24.383
R253 a_864_209.n7 a_864_209.n5 23.684
R254 a_864_209.n10 a_864_209.n9 15.001
R255 a_864_209.n0 a_864_209.t0 14.282
R256 a_864_209.n0 a_864_209.t1 14.282
R257 a_864_209.n11 a_864_209.n10 12.632
R258 a_864_209.n3 a_864_209.n2 10.615
R259 YN.n7 YN.n6 249.863
R260 YN.n7 YN.n2 215.717
R261 YN.n2 YN.n1 157.964
R262 YN.n2 YN.n0 91.706
R263 YN.n6 YN.n5 30
R264 YN.n4 YN.n3 24.383
R265 YN.n6 YN.n4 23.684
R266 YN.n0 YN.t1 14.282
R267 YN.n0 YN.t0 14.282
R268 YN.n1 YN.t4 14.282
R269 YN.n1 YN.t3 14.282
R270 YN.n8 YN.n7 4.65
R271 YN.n8 YN 0.046
R272 C.n0 C.t0 470.752
R273 C.n0 C.t1 384.527
R274 C.n1 C.t2 314.896
R275 C.n1 C.n0 182.932
R276 C.n2 C.n1 4.65
R277 C.n2 C 0.046
R278 a_112_101.n10 a_112_101.n9 93.333
R279 a_112_101.n12 a_112_101.n11 68.43
R280 a_112_101.n3 a_112_101.n2 51.907
R281 a_112_101.n3 a_112_101.n1 51.594
R282 a_112_101.t0 a_112_101.n3 38.864
R283 a_112_101.n7 a_112_101.n6 38.626
R284 a_112_101.n6 a_112_101.n5 35.955
R285 a_112_101.t1 a_112_101.n8 8.137
R286 a_112_101.t0 a_112_101.n0 6.109
R287 a_112_101.t1 a_112_101.n7 4.864
R288 a_112_101.t0 a_112_101.n4 3.871
R289 a_112_101.t0 a_112_101.n13 2.535
R290 a_112_101.n13 a_112_101.t1 1.145
R291 a_112_101.t1 a_112_101.n12 0.763
R292 a_112_101.n12 a_112_101.n10 0.185
R293 GND.n31 GND.n30 237.558
R294 GND.n80 GND.n79 237.558
R295 GND.n28 GND.n27 210.82
R296 GND.n82 GND.n81 210.82
R297 GND.n60 GND.n59 172.612
R298 GND.n17 GND.n16 151.605
R299 GND.n49 GND.n48 40.431
R300 GND.n36 GND.n35 40.003
R301 GND.n89 GND.n88 37.582
R302 GND.n16 GND.n15 28.421
R303 GND.n16 GND.n14 25.263
R304 GND.n14 GND.n13 24.383
R305 GND.n94 GND.n93 20.705
R306 GND.n50 GND.n49 20.705
R307 GND.n43 GND.n42 20.705
R308 GND.n37 GND.n36 20.705
R309 GND.n90 GND.n89 20.705
R310 GND.n29 GND.n28 18.953
R311 GND.n83 GND.n82 18.953
R312 GND.n35 GND.n34 17.258
R313 GND.n88 GND.t0 15.644
R314 GND.n32 GND.n29 14.864
R315 GND.n84 GND.n83 14.864
R316 GND.n48 GND.t3 13.654
R317 GND.n88 GND.n87 13.541
R318 GND.n51 GND.n50 9.29
R319 GND.n57 GND.n56 9.154
R320 GND.n62 GND.n61 9.154
R321 GND.n65 GND.n64 9.154
R322 GND.n68 GND.n67 9.154
R323 GND.n71 GND.n70 9.154
R324 GND.n74 GND.n73 9.154
R325 GND.n77 GND.n76 9.154
R326 GND.n84 GND.n80 9.154
R327 GND.n91 GND.n86 9.154
R328 GND.n96 GND.n95 9.154
R329 GND.n99 GND.n98 9.154
R330 GND.n51 GND.n46 9.154
R331 GND.n44 GND.n41 9.154
R332 GND.n39 GND.n38 9.154
R333 GND.n32 GND.n31 9.154
R334 GND.n25 GND.n24 9.154
R335 GND.n22 GND.n21 9.154
R336 GND.n19 GND.n18 9.154
R337 GND.n11 GND.n10 9.154
R338 GND.n8 GND.n7 9.154
R339 GND.n5 GND.n4 9.154
R340 GND.n2 GND.n1 9.154
R341 GND.t3 GND.n47 7.04
R342 GND.n55 GND.n54 4.65
R343 GND.n6 GND.n5 4.65
R344 GND.n9 GND.n8 4.65
R345 GND.n12 GND.n11 4.65
R346 GND.n20 GND.n19 4.65
R347 GND.n23 GND.n22 4.65
R348 GND.n26 GND.n25 4.65
R349 GND.n33 GND.n32 4.65
R350 GND.n40 GND.n39 4.65
R351 GND.n45 GND.n44 4.65
R352 GND.n52 GND.n51 4.65
R353 GND.n100 GND.n99 4.65
R354 GND.n97 GND.n96 4.65
R355 GND.n92 GND.n91 4.65
R356 GND.n85 GND.n84 4.65
R357 GND.n78 GND.n77 4.65
R358 GND.n75 GND.n74 4.65
R359 GND.n72 GND.n71 4.65
R360 GND.n69 GND.n68 4.65
R361 GND.n66 GND.n65 4.65
R362 GND.n63 GND.n62 4.65
R363 GND.n58 GND.n57 4.65
R364 GND.n19 GND.n17 4.129
R365 GND.n44 GND.n43 4.129
R366 GND.n96 GND.n94 4.129
R367 GND.n62 GND.n60 4.129
R368 GND.n3 GND.n0 3.407
R369 GND.n3 GND.n2 2.844
R370 GND.n6 GND.n3 1.063
R371 GND.n39 GND.n37 1.032
R372 GND.n91 GND.n90 1.032
R373 GND.n54 GND.n53 0.474
R374 GND.n33 GND.n26 0.29
R375 GND.n85 GND.n78 0.29
R376 GND.n55 GND 0.207
R377 GND.n12 GND.n9 0.181
R378 GND.n69 GND.n66 0.181
R379 GND.n9 GND.n6 0.145
R380 GND.n20 GND.n12 0.145
R381 GND.n23 GND.n20 0.145
R382 GND.n26 GND.n23 0.145
R383 GND.n40 GND.n33 0.145
R384 GND.n45 GND.n40 0.145
R385 GND.n52 GND.n45 0.145
R386 GND.n100 GND.n97 0.145
R387 GND.n97 GND.n92 0.145
R388 GND.n92 GND.n85 0.145
R389 GND.n78 GND.n75 0.145
R390 GND.n75 GND.n72 0.145
R391 GND.n72 GND.n69 0.145
R392 GND.n66 GND.n63 0.145
R393 GND.n63 GND.n58 0.145
R394 GND.n58 GND.n55 0.145
R395 GND GND.n52 0.09
R396 GND GND.n100 0.09
R397 a_1444_101.n3 a_1444_101.n1 42.788
R398 a_1444_101.t0 a_1444_101.n0 8.137
R399 a_1444_101.n3 a_1444_101.n2 4.665
R400 a_1444_101.t0 a_1444_101.n3 0.06
R401 D.n0 D.t0 472.359
R402 D.n0 D.t2 384.527
R403 D.n1 D.t1 342.755
R404 D.n1 D.n0 154.955
R405 D.n2 D.n1 4.65
R406 D.n2 D 0.046
C7 VDD GND 3.70fF
C8 a_1444_101.n0 GND 0.05fF
C9 a_1444_101.n1 GND 0.12fF
C10 a_1444_101.n2 GND 0.04fF
C11 a_1444_101.n3 GND 0.16fF
C12 a_112_101.n0 GND 0.02fF
C13 a_112_101.n1 GND 0.09fF
C14 a_112_101.n2 GND 0.07fF
C15 a_112_101.n3 GND 0.04fF
C16 a_112_101.n4 GND 0.01fF
C17 a_112_101.n5 GND 0.04fF
C18 a_112_101.n6 GND 0.04fF
C19 a_112_101.n7 GND 0.02fF
C20 a_112_101.n8 GND 0.05fF
C21 a_112_101.n9 GND 0.02fF
C22 a_112_101.n10 GND 0.14fF
C23 a_112_101.n11 GND 0.08fF
C24 a_112_101.n12 GND 0.08fF
C25 a_112_101.t1 GND 0.22fF
C26 a_112_101.n13 GND 0.01fF
C27 YN.n0 GND 0.33fF
C28 YN.n1 GND 0.43fF
C29 YN.n2 GND 0.56fF
C30 YN.n3 GND 0.03fF
C31 YN.n4 GND 0.05fF
C32 YN.n5 GND 0.03fF
C33 YN.n6 GND 0.14fF
C34 YN.n7 GND 0.43fF
C35 YN.n8 GND 0.01fF
C36 a_864_209.n0 GND 0.50fF
C37 a_864_209.n1 GND 0.32fF
C38 a_864_209.n2 GND 0.45fF
C39 a_864_209.n3 GND 0.52fF
C40 a_864_209.n4 GND 0.03fF
C41 a_864_209.n5 GND 0.04fF
C42 a_864_209.n6 GND 0.03fF
C43 a_864_209.n7 GND 0.09fF
C44 a_864_209.n8 GND 0.31fF
C45 a_864_209.n9 GND 0.06fF
C46 a_864_209.n10 GND 0.04fF
C47 a_864_209.n11 GND 0.04fF
C48 a_797_1051.n0 GND 0.52fF
C49 a_797_1051.n1 GND 0.22fF
C50 VDD.n1 GND 0.03fF
C51 VDD.n2 GND 0.11fF
C52 VDD.n3 GND 0.02fF
C53 VDD.n4 GND 0.02fF
C54 VDD.n5 GND 0.05fF
C55 VDD.n6 GND 0.02fF
C56 VDD.n7 GND 0.02fF
C57 VDD.n8 GND 0.02fF
C58 VDD.n9 GND 0.02fF
C59 VDD.n10 GND 0.02fF
C60 VDD.n11 GND 0.02fF
C61 VDD.n12 GND 0.02fF
C62 VDD.n13 GND 0.02fF
C63 VDD.n14 GND 0.03fF
C64 VDD.n15 GND 0.01fF
C65 VDD.n20 GND 0.39fF
C66 VDD.n21 GND 0.23fF
C67 VDD.n22 GND 0.02fF
C68 VDD.n23 GND 0.03fF
C69 VDD.n24 GND 0.05fF
C70 VDD.n25 GND 0.21fF
C71 VDD.n26 GND 0.01fF
C72 VDD.n27 GND 0.01fF
C73 VDD.n28 GND 0.01fF
C74 VDD.n29 GND 0.14fF
C75 VDD.n30 GND 0.01fF
C76 VDD.n31 GND 0.02fF
C77 VDD.n32 GND 0.07fF
C78 VDD.n33 GND 0.07fF
C79 VDD.n34 GND 0.04fF
C80 VDD.n35 GND 0.01fF
C81 VDD.n36 GND 0.02fF
C82 VDD.n37 GND 0.02fF
C83 VDD.n38 GND 0.12fF
C84 VDD.n39 GND 0.01fF
C85 VDD.n40 GND 0.02fF
C86 VDD.n41 GND 0.02fF
C87 VDD.n42 GND 0.14fF
C88 VDD.n43 GND 0.01fF
C89 VDD.n44 GND 0.02fF
C90 VDD.n45 GND 0.02fF
C91 VDD.n46 GND 0.05fF
C92 VDD.n47 GND 0.21fF
C93 VDD.n48 GND 0.01fF
C94 VDD.n49 GND 0.01fF
C95 VDD.n50 GND 0.02fF
C96 VDD.n51 GND 0.23fF
C97 VDD.n52 GND 0.01fF
C98 VDD.n53 GND 0.02fF
C99 VDD.n54 GND 0.03fF
C100 VDD.n55 GND 0.05fF
C101 VDD.n56 GND 0.02fF
C102 VDD.n57 GND 0.02fF
C103 VDD.n58 GND 0.02fF
C104 VDD.n59 GND 0.02fF
C105 VDD.n60 GND 0.02fF
C106 VDD.n61 GND 0.02fF
C107 VDD.n62 GND 0.02fF
C108 VDD.n63 GND 0.02fF
C109 VDD.n64 GND 0.02fF
C110 VDD.n65 GND 0.02fF
C111 VDD.n66 GND 0.01fF
C112 VDD.n67 GND 0.02fF
C113 VDD.n68 GND 0.02fF
C114 VDD.n69 GND 0.19fF
C115 VDD.n70 GND 0.02fF
C116 VDD.n71 GND 0.02fF
C117 VDD.n73 GND 0.02fF
C118 VDD.n77 GND 0.23fF
C119 VDD.n78 GND 0.23fF
C120 VDD.n79 GND 0.01fF
C121 VDD.n80 GND 0.02fF
C122 VDD.n81 GND 0.03fF
C123 VDD.n82 GND 0.21fF
C124 VDD.n83 GND 0.01fF
C125 VDD.n84 GND 0.02fF
C126 VDD.n85 GND 0.02fF
C127 VDD.n86 GND 0.14fF
C128 VDD.n87 GND 0.01fF
C129 VDD.n88 GND 0.02fF
C130 VDD.n89 GND 0.02fF
C131 VDD.n90 GND 0.01fF
C132 VDD.n91 GND 0.02fF
C133 VDD.n92 GND 0.02fF
C134 VDD.n93 GND 0.