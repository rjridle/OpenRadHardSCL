magic
tech sky130
magscale 1 2
timestamp 1651259578
<< nwell >>
rect 55 1505 89 1539
<< psubdiffcont >>
rect 55 13 89 47
<< nsubdiffcont >>
rect 55 1505 89 1539
<< viali >>
rect 55 1505 89 1539
rect 55 13 89 47
<< metal1 >>
rect 547 649 761 683
use invx1_pcell  invx1_pcell_0
timestamp 1651259471
transform 1 0 666 0 1 0
box -84 0 528 1575
use nand2x1_pcell  nand2x1_pcell_0
timestamp 1651259477
transform 1 0 0 0 1 0
box -84 0 750 1575
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform -1 0 518 0 -1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform 1 0 814 0 1 666
box -53 -33 29 33
<< end >>
