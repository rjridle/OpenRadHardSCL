magic
tech sky130A
magscale 1 2
timestamp 1645911694
<< nwell >>
rect 84 1554 613 1575
rect 84 1492 635 1554
rect 84 1487 613 1492
rect 84 1139 582 1487
rect 84 1105 205 1139
rect 229 1105 582 1139
rect 84 832 582 1105
<< pdiffc >>
rect 229 1105 263 1139
<< psubdiff >>
rect 31 510 635 572
rect 31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 361 47
rect 395 46 635 47
rect 395 13 433 46
rect 31 12 433 13
rect 467 12 505 46
rect 539 12 577 46
rect 611 12 635 46
<< nsubdiff >>
rect 31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 361 1539
rect 395 1505 433 1539
rect 467 1505 505 1539
rect 539 1505 577 1539
rect 611 1505 635 1539
rect 31 868 635 930
<< psubdiffcont >>
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 361 13 395 47
rect 433 12 467 46
rect 505 12 539 46
rect 577 12 611 46
<< nsubdiffcont >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 361 1505 395 1539
rect 433 1505 467 1539
rect 505 1505 539 1539
rect 577 1505 611 1539
<< poly >>
rect 175 990 187 1020
rect 481 990 491 1020
rect 175 411 198 444
rect 168 403 198 411
rect 468 411 491 444
rect 468 410 498 411
<< locali >>
rect 31 1539 635 1554
rect 31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 361 1539
rect 395 1505 433 1539
rect 467 1505 505 1539
rect 539 1505 577 1539
rect 611 1505 635 1539
rect 31 1492 635 1505
rect 229 1047 263 1087
rect 405 1047 439 1087
rect 229 1013 439 1047
rect 131 461 165 954
rect 353 461 387 1013
rect 501 477 535 954
rect 353 427 447 461
rect 413 261 447 427
rect 219 62 253 195
rect 31 47 635 62
rect 31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 361 47
rect 395 46 635 47
rect 395 13 433 46
rect 31 12 433 13
rect 467 12 505 46
rect 539 12 577 46
rect 611 12 635 46
rect 31 0 635 12
<< viali >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 361 1505 395 1539
rect 433 1505 467 1539
rect 505 1505 539 1539
rect 577 1505 611 1539
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 361 13 395 47
rect 433 12 467 46
rect 505 12 539 46
rect 577 12 611 46
<< metal1 >>
rect 31 1539 635 1554
rect 31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 361 1539
rect 395 1505 433 1539
rect 467 1505 505 1539
rect 539 1505 577 1539
rect 611 1505 635 1539
rect 31 1492 635 1505
rect 131 723 165 757
rect 31 47 635 62
rect 31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 361 47
rect 395 46 635 47
rect 395 13 433 46
rect 31 12 433 13
rect 467 12 505 46
rect 539 12 577 46
rect 611 12 635 46
rect 31 0 635 12
use poly_li1_contact  poly_li1_contact_1 pcells
timestamp 1645652543
transform 0 1 148 -1 0 444
box -33 -27 33 27
use pmos2  pmos2_0 pcells
timestamp 1645909547
transform 1 0 43 0 1 1450
box 52 -460 352 42
use nmos_bottom  nmos_bottom_0 ./pcells
timestamp 1645649939
transform 1 0 149 0 1 105
box -37 -4 211 298
use li1_M1_contact_perp_ext  li1_M1_contact_perp_ext_0 pcells
timestamp 1645050501
transform 0 -1 148 1 0 740
box -23 -53 49 29
use poly_li1_contact  poly_li1_contact_0
timestamp 1645652543
transform 0 1 148 -1 0 987
box -33 -27 33 27
use diff_ring_side  diff_ring_side_1 pcells
timestamp 1645641539
transform 1 0 0 0 1 0
box -84 0 84 1575
use li1_M1_contact_perp_ext  li1_M1_contact_perp_ext_1
timestamp 1645050501
transform 0 -1 518 1 0 740
box -23 -53 49 29
use li1_M1_contact_perp_ext  li1_M1_contact_perp_ext_2
timestamp 1645050501
transform 0 -1 370 1 0 666
box -23 -53 49 29
use nmos_top  nmos_top_0 pcells
timestamp 1645648650
transform 1 0 307 0 1 101
box -1 0 247 309
use poly_li1_contact  poly_li1_contact_2
timestamp 1645652543
transform 0 1 518 -1 0 444
box -33 -27 33 27
use poly_li1_contact  poly_li1_contact_3
timestamp 1645652543
transform 0 1 518 -1 0 987
box -33 -27 33 27
use pmos2  pmos2_1
timestamp 1645909547
transform 1 0 219 0 1 1450
box 52 -460 352 42
use diff_ring_side  diff_ring_side_0
timestamp 1645641539
transform 1 0 666 0 1 0
box -84 0 84 1575
<< labels >>
rlabel metal1 148 740 148 740 1 A
port 1 n
rlabel metal1 72 1522 72 1522 1 VDD
port 2 n
rlabel metal1 72 30 72 30 1 VSS
port 3 n
rlabel metal1 370 666 370 666 1 Y
port 4 n
rlabel metal1 518 740 518 740 1 B
port 5 n
<< end >>
