* SPICE3 file created from TMRDFFQNX1.ext - technology: sky130A

.subckt TMRDFFQNX1 QN D CLK VDD GND
X0 QN a_3303_411.t5 a_13654_101.t0 GND sky130_fd_pr__nfet_01v8 ad=5.373p pd=4.72u as=0p ps=0u w=0u l=0u
X1 GND a_3303_411.t6 a_14320_101.t0 GND sky130_fd_pr__nfet_01v8 ad=3.7611p pd=3.297u as=0p ps=0u w=0u l=0u
X2 VDD.t146 a_8731_187.t5 a_8861_1050.t5 �ϟHwU sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X3 a_3177_1050.t4 a_277_1050.t7 VDD.t165 �BvIwU sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X4 VDD.t79 a_1845_1050.t5 a_147_187.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X5 a_11887_411.t1 a_11761_1050.t5 VDD.t101 VDD.t100 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X6 VDD.t17 D.t0 a_9183_989.t3  <p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X7 VDD.t13 D.t1 a_4891_989.t2 �;p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X8 VDD.t46 a_7469_1050.t5 a_7595_411.t2  <p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X9 GND a_8731_187.t8 a_8675_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X10 VDD.t128 CLK.t0 a_277_1050.t5 �;p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X11 GND a_7469_1050.t6 a_8030_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X12 a_13757_1051.t7 a_7595_411.t6 QN.t1  <p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X13 a_3177_1050.t1 a_3303_411.t7 VDD.t53 �;p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X14 VDD.t126 CLK.t1 a_147_187.t4  <p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X15 a_11887_411.t4 a_8731_187.t7 VDD.t144 �;p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X16 VDD.t97 a_11887_411.t5 a_11761_1050.t4  <p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X17 GND a_1845_1050.t6 a_2406_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X18 VDD.t124 CLK.t2 a_4439_187.t4 �;p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X19 a_9183_989.t2 D.t2 VDD.t40  <p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X20 GND a_8861_1050.t8 a_9658_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X21 a_3303_411.t1 a_3177_1050.t5 VDD.t163 �;p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X22 VDD.t44 a_599_989.t5 a_277_1050.t1  <p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X23 VDD.t167 a_277_1050.t9 a_599_989.t4 �;p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X24 a_8731_187.t1 a_10429_1050.t5 VDD.t71  <p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X25 a_4569_1050.t3 a_4891_989.t6 VDD.t94 �;p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X26 a_13757_1051.t3 a_3303_411.t8 QN.t2  <p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X27 VDD.t5 a_9183_989.t5 a_10429_1050.t1 �;p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X28 VDD.t83 a_147_187.t6 a_3303_411.t4  <p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X29 a_7595_411.t3 a_7469_1050.t7 VDD.t130 �;p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X30 VDD.t161 a_4569_1050.t7 a_7469_1050.t4  <p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X31 a_4439_187.t3 CLK.t3 VDD.t122 �;p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X32 a_1845_1050.t3 a_147_187.t7 VDD.t64  <p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X33 a_8861_1050.t1 a_9183_989.t6 VDD.t106 �;p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X34 VDD.t77 a_4439_187.t5 a_4569_1050.t6  <p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X35 GND a_147_187.t10 a_91_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X36 a_6137_1050.t1 a_4439_187.t6 VDD.t73 �;p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X37 a_9183_989.t1 a_8861_1050.t7 VDD.t36  <p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X38 QN a_7595_411.t10 a_14320_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X39 GND a_8861_1050.t10 a_11656_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X40 a_13093_1051.t5 a_3303_411.t9 a_13757_1051.t5 �;p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X41 a_11761_1050.t0 a_11887_411.t6 VDD.t1  <p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X42 a_3303_411.t3 a_147_187.t8 VDD.t28 �;p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X43 VDD.t153 a_7595_411.t8 a_13093_1051.t7  <p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X44 VDD.t159 D.t4 a_599_989.t2 �;p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X45 GND a_10429_1050.t6 a_10990_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X46 GND a_4439_187.t8 a_4383_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X47 a_13757_1051.t1 a_11887_411.t7 a_13093_1051.t3  <p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X48 a_8731_187.t3 CLK.t4 VDD.t120 �;p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X49 VDD.t142 a_8731_187.t10 a_10429_1050.t3  <p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X50 a_277_1050.t0 a_147_187.t9 VDD.t7 �;p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X51 a_4439_187.t1 a_6137_1050.t6 VDD.t9  <p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X52 VDD.t21 a_7595_411.t9 a_7469_1050.t2 �;p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X53 VDD.t118 CLK.t5 a_4569_1050.t1  <p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X54 VDD.t51 a_599_989.t7 a_1845_1050.t0 �;p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X55 a_11761_1050.t2 a_8861_1050.t9 VDD.t34  <p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X56 GND a_599_989.t8 a_1740_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X57 GND a_4569_1050.t8 a_5366_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X58 VDD.t169 a_11887_411.t8 a_13093_1051.t1 �;p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X59 GND a_11887_411.t9 a_13654_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X60 a_4891_989.t1 D.t5 VDD.t148  <p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X61 a_13757_1051.t4 a_3303_411.t11 a_13093_1051.t4 �;p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X62 GND a_11887_411.t10 a_12988_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X63 a_277_1050.t4 CLK.t8 VDD.t116  <p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X64 VDD.t92 a_4891_989.t8 a_4569_1050.t2 �;p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X65 VDD.t38 a_277_1050.t10 a_3177_1050.t3  <p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X66 a_147_187.t3 CLK.t9 VDD.t114 �;p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X67 VDD.t25 a_11761_1050.t6 a_11887_411.t0  <p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X68 GND a_3177_1050.t6 a_3738_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X69 GND a_4569_1050.t11 a_7364_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X70 a_4891_989.t0 a_4569_1050.t9 VDD.t11 �;p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X71 GND a_9183_989.t8 a_10324_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X72 a_7595_411.t0 a_4439_187.t10 VDD.t3  <p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X73 a_277_1050.t3 a_599_989.t9 VDD.t57 �;p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X74 a_599_989.t3 a_277_1050.t11 VDD.t68  <p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X75 a_8861_1050.t6 a_8731_187.t11 VDD.t140 �;p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X76 QN.t3 a_3303_411.t12 a_13757_1051.t2  <p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X77 VDD.t134 CLK.t12 a_8731_187.t4 �;p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X78 a_10429_1050.t0 a_9183_989.t7 VDD.t99  <p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X79 a_7469_1050.t3 a_4569_1050.t10 VDD.t75 �;p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X80 a_147_187.t0 a_1845_1050.t7 VDD.t66  <p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X81 VDD.t55 a_3303_411.t13 a_3177_1050.t2 �;p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X82 VDD.t138 a_8731_187.t12 a_11887_411.t3  <p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X83 VDD.t112 CLK.t14 a_8861_1050.t3 �;p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X84 GND a_277_1050.t12 a_1074_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X85 a_4569_1050.t5 a_4439_187.t11 VDD.t42  <p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X86 VDD.t90 a_4891_989.t9 a_6137_1050.t3 �;p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X87 VDD.t32 a_8861_1050.t11 a_11761_1050.t1  <p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X88 VDD.t81 a_3177_1050.t7 a_3303_411.t0 �;p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X89 a_13093_1051.t6 a_7595_411.t11 VDD.t171  <p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X90 a_599_989.t1 D.t7 VDD.t15 �;p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X91 VDD.t59 a_10429_1050.t7 a_8731_187.t0  <p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X92 QN.t6 a_7595_411.t12 a_13757_1051.t6 �;p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X93 a_10429_1050.t2 a_8731_187.t13 VDD.t136  <p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X94 GND a_11761_1050.t7 a_12322_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X95 a_7469_1050.t1 a_7595_411.t13 VDD.t19 �;p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X96 VDD.t104 a_9183_989.t10 a_8861_1050.t0 0<p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X97 a_4569_1050.t0 CLK.t16 VDD.t110  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X98 VDD.t150 a_4439_187.t12 a_6137_1050.t4 0<p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X99 VDD.t30 a_8861_1050.t12 a_9183_989.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X100 a_1845_1050.t4 a_599_989.t10 VDD.t157 0<p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X101 a_8861_1050.t2 CLK.t17 VDD.t108  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X102 GND a_6137_1050.t5 a_6698_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X103 a_13093_1051.t0 a_11887_411.t12 VDD.t85 0<p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X104 QN a_7595_411.t5 a_12988_101.t1 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X105 GND a_277_1050.t8 a_3072_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X106 VDD.t62 a_147_187.t11 a_1845_1050.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X107 a_6137_1050.t2 a_4891_989.t10 VDD.t88 0<p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X108 VDD.t132 a_4569_1050.t12 a_4891_989.t4  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X109 a_13093_1051.t2 a_11887_411.t13 a_13757_1051.t0 0<p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X110 VDD.t155 a_4439_187.t13 a_7595_411.t4  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X111 GND a_4891_989.t5 a_6032_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X112 VDD.t49 a_147_187.t13 a_277_1050.t2 0<p} sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X113 VDD.t23 a_6137_1050.t7 a_4439_187.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
C0 VDD CLK 7.71fF
C1 VDD D 0.97fF
C2 CLK D 0.45fF
C3 VDD QN 0.73fF
R0 a_8731_187.n7 a_8731_187.t5 512.525
R1 a_8731_187.n5 a_8731_187.t10 472.359
R2 a_8731_187.n3 a_8731_187.t12 472.359
R3 a_8731_187.n8 a_8731_187.t8 417.109
R4 a_8731_187.n5 a_8731_187.t13 384.527
R5 a_8731_187.n3 a_8731_187.t7 384.527
R6 a_8731_187.n7 a_8731_187.t11 371.139
R7 a_8731_187.n6 a_8731_187.t6 370.613
R8 a_8731_187.n4 a_8731_187.t9 370.613
R9 a_8731_187.n13 a_8731_187.n11 367.82
R10 a_8731_187.n8 a_8731_187.n7 179.837
R11 a_8731_187.n2 a_8731_187.n1 157.964
R12 a_8731_187.n6 a_8731_187.n5 127.096
R13 a_8731_187.n4 a_8731_187.n3 127.096
R14 a_8731_187.n11 a_8731_187.n2 104.282
R15 a_8731_187.n2 a_8731_187.n0 91.706
R16 a_8731_187.n13 a_8731_187.n12 15.218
R17 a_8731_187.n0 a_8731_187.t4 14.282
R18 a_8731_187.n0 a_8731_187.t3 14.282
R19 a_8731_187.n1 a_8731_187.t0 14.282
R20 a_8731_187.n1 a_8731_187.t1 14.282
R21 a_8731_187.n14 a_8731_187.n13 12.014
R22 a_8731_187.n9 a_8731_187.n8 11.134
R23 a_8731_187.n10 a_8731_187.n4 8.957
R24 a_8731_187.n9 a_8731_187.n6 4.65
R25 a_8731_187.n11 a_8731_187.n10 4.65
R26 a_8731_187.n10 a_8731_187.n9 2.947
R27 a_8861_1050.n7 a_8861_1050.t12 480.392
R28 a_8861_1050.n5 a_8861_1050.t11 480.392
R29 a_8861_1050.n7 a_8861_1050.t7 403.272
R30 a_8861_1050.n5 a_8861_1050.t9 403.272
R31 a_8861_1050.n8 a_8861_1050.t8 385.063
R32 a_8861_1050.n6 a_8861_1050.t10 385.063
R33 a_8861_1050.n12 a_8861_1050.n10 342.597
R34 a_8861_1050.n3 a_8861_1050.n2 161.352
R35 a_8861_1050.n10 a_8861_1050.n4 151.34
R36 a_8861_1050.n8 a_8861_1050.n7 143.429
R37 a_8861_1050.n6 a_8861_1050.n5 143.429
R38 a_8861_1050.n4 a_8861_1050.n0 95.095
R39 a_8861_1050.n3 a_8861_1050.n1 95.095
R40 a_8861_1050.n4 a_8861_1050.n3 66.258
R41 a_8861_1050.n12 a_8861_1050.n11 15.218
R42 a_8861_1050.n0 a_8861_1050.t0 14.282
R43 a_8861_1050.n0 a_8861_1050.t1 14.282
R44 a_8861_1050.n1 a_8861_1050.t3 14.282
R45 a_8861_1050.n1 a_8861_1050.t2 14.282
R46 a_8861_1050.n2 a_8861_1050.t5 14.282
R47 a_8861_1050.n2 a_8861_1050.t6 14.282
R48 a_8861_1050.n13 a_8861_1050.n12 12.014
R49 a_8861_1050.n9 a_8861_1050.n6 11.95
R50 a_8861_1050.n10 a_8861_1050.n9 5.965
R51 a_8861_1050.n9 a_8861_1050.n8 4.65
R52 VDD.n723 VDD.n712 144.705
R53 VDD.n780 VDD.n773 144.705
R54 VDD.n837 VDD.n830 144.705
R55 VDD.n894 VDD.n887 144.705
R56 VDD.n951 VDD.n944 144.705
R57 VDD.n1008 VDD.n1001 144.705
R58 VDD.n1083 VDD.n1076 144.705
R59 VDD.n1140 VDD.n1133 144.705
R60 VDD.n1197 VDD.n1190 144.705
R61 VDD.n602 VDD.n595 144.705
R62 VDD.n1254 VDD.n1247 144.705
R63 VDD.n545 VDD.n538 144.705
R64 VDD.n470 VDD.n463 144.705
R65 VDD.n413 VDD.n406 144.705
R66 VDD.n356 VDD.n349 144.705
R67 VDD.n299 VDD.n292 144.705
R68 VDD.n242 VDD.n235 144.705
R69 VDD.n185 VDD.n178 144.705
R70 VDD.n128 VDD.n121 144.705
R71 VDD.n75 VDD.n64 144.705
R72 VDD.n689 VDD.t44 143.754
R73 VDD.n1050 VDD.t92 143.754
R74 VDD.n479 VDD.t104 143.754
R75 VDD.n748 VDD.t159 143.754
R76 VDD.n805 VDD.t62 143.754
R77 VDD.n862 VDD.t126 143.754
R78 VDD.n919 VDD.t55 143.754
R79 VDD.n976 VDD.t83 143.754
R80 VDD.n1108 VDD.t13 143.754
R81 VDD.n1165 VDD.t150 143.754
R82 VDD.n1222 VDD.t124 143.754
R83 VDD.n605 VDD.t21 143.754
R84 VDD.n548 VDD.t155 143.754
R85 VDD.n416 VDD.t17 143.754
R86 VDD.n359 VDD.t142 143.754
R87 VDD.n302 VDD.t134 143.754
R88 VDD.n245 VDD.t97 143.754
R89 VDD.n188 VDD.t138 143.754
R90 VDD.n153 VDD.t85 135.539
R91 VDD.n131 VDD.t153 135.539
R92 VDD.n654 VDD.t7 135.17
R93 VDD.n726 VDD.t68 135.17
R94 VDD.n783 VDD.t157 135.17
R95 VDD.n840 VDD.t66 135.17
R96 VDD.n897 VDD.t165 135.17
R97 VDD.n954 VDD.t163 135.17
R98 VDD.n1015 VDD.t42 135.17
R99 VDD.n1086 VDD.t11 135.17
R100 VDD.n1143 VDD.t88 135.17
R101 VDD.n1200 VDD.t9 135.17
R102 VDD.n1257 VDD.t75 135.17
R103 VDD.n570 VDD.t130 135.17
R104 VDD.n509 VDD.t140 135.17
R105 VDD.n438 VDD.t36 135.17
R106 VDD.n381 VDD.t99 135.17
R107 VDD.n324 VDD.t71 135.17
R108 VDD.n267 VDD.t34 135.17
R109 VDD.n210 VDD.t101 135.17
R110 VDD.n141 VDD.n140 129.849
R111 VDD.n664 VDD.n663 129.472
R112 VDD.n680 VDD.n679 129.472
R113 VDD.n740 VDD.n739 129.472
R114 VDD.n797 VDD.n796 129.472
R115 VDD.n854 VDD.n853 129.472
R116 VDD.n911 VDD.n910 129.472
R117 VDD.n968 VDD.n967 129.472
R118 VDD.n1025 VDD.n1024 129.472
R119 VDD.n1041 VDD.n1040 129.472
R120 VDD.n1100 VDD.n1099 129.472
R121 VDD.n1157 VDD.n1156 129.472
R122 VDD.n1214 VDD.n1213 129.472
R123 VDD.n615 VDD.n614 129.472
R124 VDD.n558 VDD.n557 129.472
R125 VDD.n500 VDD.n499 129.472
R126 VDD.n488 VDD.n487 129.472
R127 VDD.n426 VDD.n425 129.472
R128 VDD.n369 VDD.n368 129.472
R129 VDD.n312 VDD.n311 129.472
R130 VDD.n255 VDD.n254 129.472
R131 VDD.n198 VDD.n197 129.472
R132 VDD.n60 VDD.n59 92.5
R133 VDD.n58 VDD.n57 92.5
R134 VDD.n56 VDD.n55 92.5
R135 VDD.n54 VDD.n53 92.5
R136 VDD.n62 VDD.n61 92.5
R137 VDD.n117 VDD.n116 92.5
R138 VDD.n115 VDD.n114 92.5
R139 VDD.n113 VDD.n112 92.5
R140 VDD.n111 VDD.n110 92.5
R141 VDD.n119 VDD.n118 92.5
R142 VDD.n174 VDD.n173 92.5
R143 VDD.n172 VDD.n171 92.5
R144 VDD.n170 VDD.n169 92.5
R145 VDD.n168 VDD.n167 92.5
R146 VDD.n176 VDD.n175 92.5
R147 VDD.n231 VDD.n230 92.5
R148 VDD.n229 VDD.n228 92.5
R149 VDD.n227 VDD.n226 92.5
R150 VDD.n225 VDD.n224 92.5
R151 VDD.n233 VDD.n232 92.5
R152 VDD.n288 VDD.n287 92.5
R153 VDD.n286 VDD.n285 92.5
R154 VDD.n284 VDD.n283 92.5
R155 VDD.n282 VDD.n281 92.5
R156 VDD.n290 VDD.n289 92.5
R157 VDD.n345 VDD.n344 92.5
R158 VDD.n343 VDD.n342 92.5
R159 VDD.n341 VDD.n340 92.5
R160 VDD.n339 VDD.n338 92.5
R161 VDD.n347 VDD.n346 92.5
R162 VDD.n402 VDD.n401 92.5
R163 VDD.n400 VDD.n399 92.5
R164 VDD.n398 VDD.n397 92.5
R165 VDD.n396 VDD.n395 92.5
R166 VDD.n404 VDD.n403 92.5
R167 VDD.n459 VDD.n458 92.5
R168 VDD.n457 VDD.n456 92.5
R169 VDD.n455 VDD.n454 92.5
R170 VDD.n453 VDD.n452 92.5
R171 VDD.n461 VDD.n460 92.5
R172 VDD.n534 VDD.n533 92.5
R173 VDD.n532 VDD.n531 92.5
R174 VDD.n530 VDD.n529 92.5
R175 VDD.n528 VDD.n527 92.5
R176 VDD.n536 VDD.n535 92.5
R177 VDD.n591 VDD.n590 92.5
R178 VDD.n589 VDD.n588 92.5
R179 VDD.n587 VDD.n586 92.5
R180 VDD.n585 VDD.n584 92.5
R181 VDD.n593 VDD.n592 92.5
R182 VDD.n1243 VDD.n1242 92.5
R183 VDD.n1241 VDD.n1240 92.5
R184 VDD.n1239 VDD.n1238 92.5
R185 VDD.n1237 VDD.n1236 92.5
R186 VDD.n1245 VDD.n1244 92.5
R187 VDD.n1186 VDD.n1185 92.5
R188 VDD.n1184 VDD.n1183 92.5
R189 VDD.n1182 VDD.n1181 92.5
R190 VDD.n1180 VDD.n1179 92.5
R191 VDD.n1188 VDD.n1187 92.5
R192 VDD.n1129 VDD.n1128 92.5
R193 VDD.n1127 VDD.n1126 92.5
R194 VDD.n1125 VDD.n1124 92.5
R195 VDD.n1123 VDD.n1122 92.5
R196 VDD.n1131 VDD.n1130 92.5
R197 VDD.n1072 VDD.n1071 92.5
R198 VDD.n1070 VDD.n1069 92.5
R199 VDD.n1068 VDD.n1067 92.5
R200 VDD.n1066 VDD.n1065 92.5
R201 VDD.n1074 VDD.n1073 92.5
R202 VDD.n997 VDD.n996 92.5
R203 VDD.n995 VDD.n994 92.5
R204 VDD.n993 VDD.n992 92.5
R205 VDD.n991 VDD.n990 92.5
R206 VDD.n999 VDD.n998 92.5
R207 VDD.n940 VDD.n939 92.5
R208 VDD.n938 VDD.n937 92.5
R209 VDD.n936 VDD.n935 92.5
R210 VDD.n934 VDD.n933 92.5
R211 VDD.n942 VDD.n941 92.5
R212 VDD.n883 VDD.n882 92.5
R213 VDD.n881 VDD.n880 92.5
R214 VDD.n879 VDD.n878 92.5
R215 VDD.n877 VDD.n876 92.5
R216 VDD.n885 VDD.n884 92.5
R217 VDD.n826 VDD.n825 92.5
R218 VDD.n824 VDD.n823 92.5
R219 VDD.n822 VDD.n821 92.5
R220 VDD.n820 VDD.n819 92.5
R221 VDD.n828 VDD.n827 92.5
R222 VDD.n769 VDD.n768 92.5
R223 VDD.n767 VDD.n766 92.5
R224 VDD.n765 VDD.n764 92.5
R225 VDD.n763 VDD.n762 92.5
R226 VDD.n771 VDD.n770 92.5
R227 VDD.n708 VDD.n707 92.5
R228 VDD.n706 VDD.n705 92.5
R229 VDD.n704 VDD.n703 92.5
R230 VDD.n702 VDD.n701 92.5
R231 VDD.n710 VDD.n709 92.5
R232 VDD.n638 VDD.n637 92.5
R233 VDD.n636 VDD.n635 92.5
R234 VDD.n634 VDD.n633 92.5
R235 VDD.n632 VDD.n631 92.5
R236 VDD.n640 VDD.n639 92.5
R237 VDD.n14 VDD.n1 92.5
R238 VDD.n5 VDD.n4 92.5
R239 VDD.n7 VDD.n6 92.5
R240 VDD.n9 VDD.n8 92.5
R241 VDD.n11 VDD.n10 92.5
R242 VDD.n13 VDD.n12 92.5
R243 VDD.n21 VDD.n20 92.059
R244 VDD.n74 VDD.n73 92.059
R245 VDD.n127 VDD.n126 92.059
R246 VDD.n184 VDD.n183 92.059
R247 VDD.n241 VDD.n240 92.059
R248 VDD.n298 VDD.n297 92.059
R249 VDD.n355 VDD.n354 92.059
R250 VDD.n412 VDD.n411 92.059
R251 VDD.n469 VDD.n468 92.059
R252 VDD.n544 VDD.n543 92.059
R253 VDD.n601 VDD.n600 92.059
R254 VDD.n1253 VDD.n1252 92.059
R255 VDD.n1196 VDD.n1195 92.059
R256 VDD.n1139 VDD.n1138 92.059
R257 VDD.n1082 VDD.n1081 92.059
R258 VDD.n1007 VDD.n1006 92.059
R259 VDD.n950 VDD.n949 92.059
R260 VDD.n893 VDD.n892 92.059
R261 VDD.n836 VDD.n835 92.059
R262 VDD.n779 VDD.n778 92.059
R263 VDD.n722 VDD.n721 92.059
R264 VDD.n646 VDD.n645 92.059
R265 VDD.n20 VDD.n16 67.194
R266 VDD.n20 VDD.n17 67.194
R267 VDD.n20 VDD.n18 67.194
R268 VDD.n20 VDD.n19 67.194
R269 VDD.n630 VDD.n629 44.141
R270 VDD.n761 VDD.n760 44.141
R271 VDD.n818 VDD.n817 44.141
R272 VDD.n875 VDD.n874 44.141
R273 VDD.n932 VDD.n931 44.141
R274 VDD.n989 VDD.n988 44.141
R275 VDD.n1064 VDD.n1063 44.141
R276 VDD.n1121 VDD.n1120 44.141
R277 VDD.n1178 VDD.n1177 44.141
R278 VDD.n1235 VDD.n1234 44.141
R279 VDD.n583 VDD.n582 44.141
R280 VDD.n526 VDD.n525 44.141
R281 VDD.n451 VDD.n450 44.141
R282 VDD.n394 VDD.n393 44.141
R283 VDD.n337 VDD.n336 44.141
R284 VDD.n280 VDD.n279 44.141
R285 VDD.n223 VDD.n222 44.141
R286 VDD.n166 VDD.n165 44.141
R287 VDD.n109 VDD.n108 44.141
R288 VDD.n5 VDD.n3 44.141
R289 VDD.n760 VDD.n758 44.107
R290 VDD.n817 VDD.n815 44.107
R291 VDD.n874 VDD.n872 44.107
R292 VDD.n931 VDD.n929 44.107
R293 VDD.n988 VDD.n986 44.107
R294 VDD.n1063 VDD.n1061 44.107
R295 VDD.n1120 VDD.n1118 44.107
R296 VDD.n1177 VDD.n1175 44.107
R297 VDD.n1234 VDD.n1232 44.107
R298 VDD.n582 VDD.n580 44.107
R299 VDD.n525 VDD.n523 44.107
R300 VDD.n450 VDD.n448 44.107
R301 VDD.n393 VDD.n391 44.107
R302 VDD.n336 VDD.n334 44.107
R303 VDD.n279 VDD.n277 44.107
R304 VDD.n222 VDD.n220 44.107
R305 VDD.n165 VDD.n163 44.107
R306 VDD.n108 VDD.n106 44.107
R307 VDD.n629 VDD.n627 44.107
R308 VDD.n3 VDD.n2 44.107
R309 VDD.n20 VDD.n15 41.052
R310 VDD.n68 VDD.n66 39.742
R311 VDD.n68 VDD.n67 39.742
R312 VDD.n70 VDD.n69 39.742
R313 VDD.n123 VDD.n122 39.742
R314 VDD.n180 VDD.n179 39.742
R315 VDD.n237 VDD.n236 39.742
R316 VDD.n294 VDD.n293 39.742
R317 VDD.n351 VDD.n350 39.742
R318 VDD.n408 VDD.n407 39.742
R319 VDD.n465 VDD.n464 39.742
R320 VDD.n540 VDD.n539 39.742
R321 VDD.n597 VDD.n596 39.742
R322 VDD.n1249 VDD.n1248 39.742
R323 VDD.n1192 VDD.n1191 39.742
R324 VDD.n1135 VDD.n1134 39.742
R325 VDD.n1078 VDD.n1077 39.742
R326 VDD.n1003 VDD.n1002 39.742
R327 VDD.n946 VDD.n945 39.742
R328 VDD.n889 VDD.n888 39.742
R329 VDD.n832 VDD.n831 39.742
R330 VDD.n775 VDD.n774 39.742
R331 VDD.n642 VDD.n641 39.742
R332 VDD.n720 VDD.n717 39.742
R333 VDD.n720 VDD.n719 39.742
R334 VDD.n716 VDD.n715 39.742
R335 VDD.n108 VDD.n107 38
R336 VDD.n165 VDD.n164 38
R337 VDD.n222 VDD.n221 38
R338 VDD.n279 VDD.n278 38
R339 VDD.n336 VDD.n335 38
R340 VDD.n393 VDD.n392 38
R341 VDD.n450 VDD.n449 38
R342 VDD.n525 VDD.n524 38
R343 VDD.n582 VDD.n581 38
R344 VDD.n1234 VDD.n1233 38
R345 VDD.n1177 VDD.n1176 38
R346 VDD.n1120 VDD.n1119 38
R347 VDD.n1063 VDD.n1062 38
R348 VDD.n988 VDD.n987 38
R349 VDD.n931 VDD.n930 38
R350 VDD.n874 VDD.n873 38
R351 VDD.n817 VDD.n816 38
R352 VDD.n760 VDD.n759 38
R353 VDD.n629 VDD.n628 38
R354 VDD.n758 VDD.n757 36.774
R355 VDD.n815 VDD.n814 36.774
R356 VDD.n872 VDD.n871 36.774
R357 VDD.n929 VDD.n928 36.774
R358 VDD.n986 VDD.n985 36.774
R359 VDD.n1061 VDD.n1060 36.774
R360 VDD.n1118 VDD.n1117 36.774
R361 VDD.n1175 VDD.n1174 36.774
R362 VDD.n1232 VDD.n1231 36.774
R363 VDD.n580 VDD.n579 36.774
R364 VDD.n523 VDD.n522 36.774
R365 VDD.n448 VDD.n447 36.774
R366 VDD.n391 VDD.n390 36.774
R367 VDD.n334 VDD.n333 36.774
R368 VDD.n277 VDD.n276 36.774
R369 VDD.n220 VDD.n219 36.774
R370 VDD.n163 VDD.n162 36.774
R371 VDD.n106 VDD.n105 36.774
R372 VDD.n66 VDD.n65 36.774
R373 VDD.n719 VDD.n718 36.774
R374 VDD.n481 0<p} 35.8
R375 VDD.n1044 �;p} 35.8
R376 VDD.n683  <p} 35.8
R377 VDD.n505  gIwU 33.243
R378 VDD.n1020  <p} 33.243
R379 VDD.n659 �;p} 33.243
R380 VDD.n1 VDD.n0 30.923
R381 VDD.n73 VDD.n71 26.38
R382 VDD.n73 VDD.n70 26.38
R383 VDD.n73 VDD.n68 26.38
R384 VDD.n73 VDD.n72 26.38
R385 VDD.n126 VDD.n124 26.38
R386 VDD.n126 VDD.n123 26.38
R387 VDD.n126 VDD.n125 26.38
R388 VDD.n183 VDD.n181 26.38
R389 VDD.n183 VDD.n180 26.38
R390 VDD.n183 VDD.n182 26.38
R391 VDD.n240 VDD.n238 26.38
R392 VDD.n240 VDD.n237 26.38
R393 VDD.n240 VDD.n239 26.38
R394 VDD.n297 VDD.n295 26.38
R395 VDD.n297 VDD.n294 26.38
R396 VDD.n297 VDD.n296 26.38
R397 VDD.n354 VDD.n352 26.38
R398 VDD.n354 VDD.n351 26.38
R399 VDD.n354 VDD.n353 26.38
R400 VDD.n411 VDD.n409 26.38
R401 VDD.n411 VDD.n408 26.38
R402 VDD.n411 VDD.n410 26.38
R403 VDD.n468 VDD.n466 26.38
R404 VDD.n468 VDD.n465 26.38
R405 VDD.n468 VDD.n467 26.38
R406 VDD.n543 VDD.n541 26.38
R407 VDD.n543 VDD.n540 26.38
R408 VDD.n543 VDD.n542 26.38
R409 VDD.n600 VDD.n598 26.38
R410 VDD.n600 VDD.n597 26.38
R411 VDD.n600 VDD.n599 26.38
R412 VDD.n1252 VDD.n1250 26.38
R413 VDD.n1252 VDD.n1249 26.38
R414 VDD.n1252 VDD.n1251 26.38
R415 VDD.n1195 VDD.n1193 26.38
R416 VDD.n1195 VDD.n1192 26.38
R417 VDD.n1195 VDD.n1194 26.38
R418 VDD.n1138 VDD.n1136 26.38
R419 VDD.n1138 VDD.n1135 26.38
R420 VDD.n1138 VDD.n1137 26.38
R421 VDD.n1081 VDD.n1079 26.38
R422 VDD.n1081 VDD.n1078 26.38
R423 VDD.n1081 VDD.n1080 26.38
R424 VDD.n1006 VDD.n1004 26.38
R425 VDD.n1006 VDD.n1003 26.38
R426 VDD.n1006 VDD.n1005 26.38
R427 VDD.n949 VDD.n947 26.38
R428 VDD.n949 VDD.n946 26.38
R429 VDD.n949 VDD.n948 26.38
R430 VDD.n892 VDD.n890 26.38
R431 VDD.n892 VDD.n889 26.38
R432 VDD.n892 VDD.n891 26.38
R433 VDD.n835 VDD.n833 26.38
R434 VDD.n835 VDD.n832 26.38
R435 VDD.n835 VDD.n834 26.38
R436 VDD.n778 VDD.n776 26.38
R437 VDD.n778 VDD.n775 26.38
R438 VDD.n778 VDD.n777 26.38
R439 VDD.n645 VDD.n643 26.38
R440 VDD.n645 VDD.n642 26.38
R441 VDD.n645 VDD.n644 26.38
R442 VDD.n721 VDD.n720 26.38
R443 VDD.n721 VDD.n716 26.38
R444 VDD.n721 VDD.n714 26.38
R445 VDD.n721 VDD.n713 26.38
R446 VDD.n648 VDD.n640 22.915
R447 VDD.n23 VDD.n14 22.915
R448 VDD.n28  <p} 20.457
R449 VDD.n93  <p} 20.457
R450 VDD.n136  <p} 20.457
R451 VDD.n193  <p} 20.457
R452 VDD.n250  <p} 20.457
R453 VDD.n307 �;p} 20.457
R454 VDD.n364  <p} 20.457
R455 VDD.n421  <p} 20.457
R456 VDD.n553  20.457
R457 VDD.n610 �;p} 20.457
R458 VDD.n1218 �;p} 20.457
R459 VDD.n1161 0<p} 20.457
R460 VDD.n1104 ���IwU 20.457
R461 VDD.n972  <p} 20.457
R462 VDD.n915 �;p} 20.457
R463 VDD.n858  <p} 20.457
R464 VDD.n801  20.457
R465 VDD.n744 �;p} 20.457
R466 VDD.n39  <p} 17.9
R467 VDD.n82 �;p} 17.9
R468 VDD.n149 0<p} 17.9
R469 VDD.n206 VDD.t100 17.9
R470 VDD.n263  <p} 17.9
R471 VDD.n320  <p} 17.9
R472 VDD.n377  <p} 17.9
R473 VDD.n434  <p} 17.9
R474 VDD.n566 �;p} 17.9
R475 VDD.n623 �;p} 17.9
R476 VDD.n1205  <p} 17.9
R477 VDD.n1148 0<p} 17.9
R478 VDD.n1091 �;p} 17.9
R479 VDD.n959 �;p} 17.9
R480 VDD.n902 �BvIwU 17.9
R481 VDD.n845  <p} 17.9
R482 VDD.n788 0<p} 17.9
R483 VDD.n731  <p} 17.9
R484 VDD.n485 0�\IwU 15.343
R485 VDD.n1038 �;p} 15.343
R486 VDD.n677 �;p} 15.343
R487 VDD.n640 VDD.n638 14.864
R488 VDD.n638 VDD.n636 14.864
R489 VDD.n636 VDD.n634 14.864
R490 VDD.n634 VDD.n632 14.864
R491 VDD.n632 VDD.n630 14.864
R492 VDD.n771 VDD.n769 14.864
R493 VDD.n769 VDD.n767 14.864
R494 VDD.n767 VDD.n765 14.864
R495 VDD.n765 VDD.n763 14.864
R496 VDD.n763 VDD.n761 14.864
R497 VDD.n828 VDD.n826 14.864
R498 VDD.n826 VDD.n824 14.864
R499 VDD.n824 VDD.n822 14.864
R500 VDD.n822 VDD.n820 14.864
R501 VDD.n820 VDD.n818 14.864
R502 VDD.n885 VDD.n883 14.864
R503 VDD.n883 VDD.n881 14.864
R504 VDD.n881 VDD.n879 14.864
R505 VDD.n879 VDD.n877 14.864
R506 VDD.n877 VDD.n875 14.864
R507 VDD.n942 VDD.n940 14.864
R508 VDD.n940 VDD.n938 14.864
R509 VDD.n938 VDD.n936 14.864
R510 VDD.n936 VDD.n934 14.864
R511 VDD.n934 VDD.n932 14.864
R512 VDD.n999 VDD.n997 14.864
R513 VDD.n997 VDD.n995 14.864
R514 VDD.n995 VDD.n993 14.864
R515 VDD.n993 VDD.n991 14.864
R516 VDD.n991 VDD.n989 14.864
R517 VDD.n1074 VDD.n1072 14.864
R518 VDD.n1072 VDD.n1070 14.864
R519 VDD.n1070 VDD.n1068 14.864
R520 VDD.n1068 VDD.n1066 14.864
R521 VDD.n1066 VDD.n1064 14.864
R522 VDD.n1131 VDD.n1129 14.864
R523 VDD.n1129 VDD.n1127 14.864
R524 VDD.n1127 VDD.n1125 14.864
R525 VDD.n1125 VDD.n1123 14.864
R526 VDD.n1123 VDD.n1121 14.864
R527 VDD.n1188 VDD.n1186 14.864
R528 VDD.n1186 VDD.n1184 14.864
R529 VDD.n1184 VDD.n1182 14.864
R530 VDD.n1182 VDD.n1180 14.864
R531 VDD.n1180 VDD.n1178 14.864
R532 VDD.n1245 VDD.n1243 14.864
R533 VDD.n1243 VDD.n1241 14.864
R534 VDD.n1241 VDD.n1239 14.864
R535 VDD.n1239 VDD.n1237 14.864
R536 VDD.n1237 VDD.n1235 14.864
R537 VDD.n593 VDD.n591 14.864
R538 VDD.n591 VDD.n589 14.864
R539 VDD.n589 VDD.n587 14.864
R540 VDD.n587 VDD.n585 14.864
R541 VDD.n585 VDD.n583 14.864
R542 VDD.n536 VDD.n534 14.864
R543 VDD.n534 VDD.n532 14.864
R544 VDD.n532 VDD.n530 14.864
R545 VDD.n530 VDD.n528 14.864
R546 VDD.n528 VDD.n526 14.864
R547 VDD.n461 VDD.n459 14.864
R548 VDD.n459 VDD.n457 14.864
R549 VDD.n457 VDD.n455 14.864
R550 VDD.n455 VDD.n453 14.864
R551 VDD.n453 VDD.n451 14.864
R552 VDD.n404 VDD.n402 14.864
R553 VDD.n402 VDD.n400 14.864
R554 VDD.n400 VDD.n398 14.864
R555 VDD.n398 VDD.n396 14.864
R556 VDD.n396 VDD.n394 14.864
R557 VDD.n347 VDD.n345 14.864
R558 VDD.n345 VDD.n343 14.864
R559 VDD.n343 VDD.n341 14.864
R560 VDD.n341 VDD.n339 14.864
R561 VDD.n339 VDD.n337 14.864
R562 VDD.n290 VDD.n288 14.864
R563 VDD.n288 VDD.n286 14.864
R564 VDD.n286 VDD.n284 14.864
R565 VDD.n284 VDD.n282 14.864
R566 VDD.n282 VDD.n280 14.864
R567 VDD.n233 VDD.n231 14.864
R568 VDD.n231 VDD.n229 14.864
R569 VDD.n229 VDD.n227 14.864
R570 VDD.n227 VDD.n225 14.864
R571 VDD.n225 VDD.n223 14.864
R572 VDD.n176 VDD.n174 14.864
R573 VDD.n174 VDD.n172 14.864
R574 VDD.n172 VDD.n170 14.864
R575 VDD.n170 VDD.n168 14.864
R576 VDD.n168 VDD.n166 14.864
R577 VDD.n119 VDD.n117 14.864
R578 VDD.n117 VDD.n115 14.864
R579 VDD.n115 VDD.n113 14.864
R580 VDD.n113 VDD.n111 14.864
R581 VDD.n111 VDD.n109 14.864
R582 VDD.n62 VDD.n60 14.864
R583 VDD.n60 VDD.n58 14.864
R584 VDD.n58 VDD.n56 14.864
R585 VDD.n56 VDD.n54 14.864
R586 VDD.n54 VDD.n52 14.864
R587 VDD.n52 VDD.n51 14.864
R588 VDD.n710 VDD.n708 14.864
R589 VDD.n708 VDD.n706 14.864
R590 VDD.n706 VDD.n704 14.864
R591 VDD.n704 VDD.n702 14.864
R592 VDD.n702 VDD.n700 14.864
R593 VDD.n700 VDD.n699 14.864
R594 VDD.n14 VDD.n13 14.864
R595 VDD.n13 VDD.n11 14.864
R596 VDD.n11 VDD.n9 14.864
R597 VDD.n9 VDD.n7 14.864
R598 VDD.n7 VDD.n5 14.864
R599 VDD.n76 VDD.n63 14.864
R600 VDD.n129 VDD.n120 14.864
R601 VDD.n186 VDD.n177 14.864
R602 VDD.n243 VDD.n234 14.864
R603 VDD.n300 VDD.n291 14.864
R604 VDD.n357 VDD.n348 14.864
R605 VDD.n414 VDD.n405 14.864
R606 VDD.n471 VDD.n462 14.864
R607 VDD.n546 VDD.n537 14.864
R608 VDD.n603 VDD.n594 14.864
R609 VDD.n1255 VDD.n1246 14.864
R610 VDD.n1198 VDD.n1189 14.864
R611 VDD.n1141 VDD.n1132 14.864
R612 VDD.n1084 VDD.n1075 14.864
R613 VDD.n1009 VDD.n1000 14.864
R614 VDD.n952 VDD.n943 14.864
R615 VDD.n895 VDD.n886 14.864
R616 VDD.n838 VDD.n829 14.864
R617 VDD.n781 VDD.n772 14.864
R618 VDD.n724 VDD.n711 14.864
R619 VDD.n663 VDD.t116 14.282
R620 VDD.n663 VDD.t49 14.282
R621 VDD.n679 VDD.t57 14.282
R622 VDD.n679 VDD.t128 14.282
R623 VDD.n739 VDD.t15 14.282
R624 VDD.n739 VDD.t167 14.282
R625 VDD.n796 VDD.t64 14.282
R626 VDD.n796 VDD.t51 14.282
R627 VDD.n853 VDD.t114 14.282
R628 VDD.n853 VDD.t79 14.282
R629 VDD.n910 VDD.t53 14.282
R630 VDD.n910 VDD.t38 14.282
R631 VDD.n967 VDD.t28 14.282
R632 VDD.n967 VDD.t81 14.282
R633 VDD.n1024 VDD.t110 14.282
R634 VDD.n1024 VDD.t77 14.282
R635 VDD.n1040 VDD.t94 14.282
R636 VDD.n1040 VDD.t118 14.282
R637 VDD.n1099 VDD.t148 14.282
R638 VDD.n1099 VDD.t132 14.282
R639 VDD.n1156 VDD.t73 14.282
R640 VDD.n1156 VDD.t90 14.282
R641 VDD.n1213 VDD.t122 14.282
R642 VDD.n1213 VDD.t23 14.282
R643 VDD.n614 VDD.t19 14.282
R644 VDD.n614 VDD.t161 14.282
R645 VDD.n557 VDD.t3 14.282
R646 VDD.n557 VDD.t46 14.282
R647 VDD.n499 VDD.t108 14.282
R648 VDD.n499 VDD.t146 14.282
R649 VDD.n487 VDD.t106 14.282
R650 VDD.n487 VDD.t112 14.282
R651 VDD.n425 VDD.t40 14.282
R652 VDD.n425 VDD.t30 14.282
R653 VDD.n368 VDD.t136 14.282
R654 VDD.n368 VDD.t5 14.282
R655 VDD.n311 VDD.t120 14.282
R656 VDD.n311 VDD.t59 14.282
R657 VDD.n254 VDD.t1 14.282
R658 VDD.n254 VDD.t32 14.282
R659 VDD.n197 VDD.t144 14.282
R660 VDD.n197 VDD.t25 14.282
R661 VDD.n140 VDD.t171 14.282
R662 VDD.n140 VDD.t169 14.282
R663 VDD.n501 �ϟHwU 12.786
R664 VDD.n1026  <p} 12.786
R665 VDD.n665 0<p} 12.786
R666 VDD.n143 VDD.n141 9.083
R667 VDD.n200 VDD.n198 9.083
R668 VDD.n257 VDD.n255 9.083
R669 VDD.n314 VDD.n312 9.083
R670 VDD.n371 VDD.n369 9.083
R671 VDD.n428 VDD.n426 9.083
R672 VDD.n560 VDD.n558 9.083
R673 VDD.n617 VDD.n615 9.083
R674 VDD.n1216 VDD.n1214 9.083
R675 VDD.n1159 VDD.n1157 9.083
R676 VDD.n1102 VDD.n1100 9.083
R677 VDD.n970 VDD.n968 9.083
R678 VDD.n913 VDD.n911 9.083
R679 VDD.n856 VDD.n854 9.083
R680 VDD.n799 VDD.n797 9.083
R681 VDD.n742 VDD.n740 9.083
R682 VDD.n23 VDD.n22 8.855
R683 VDD.n22 VDD.n21 8.855
R684 VDD.n26 VDD.n25 8.855
R685 VDD.n25 VDD.n24 8.855
R686 VDD.n30 VDD.n29 8.855
R687 VDD.n29 VDD.n28 8.855
R688 VDD.n33 VDD.n32 8.855
R689 VDD.n32 �;p} 8.855
R690 VDD.n37 VDD.n36 8.855
R691 VDD.n36 VDD.n35 8.855
R692 VDD.n41 VDD.n40 8.855
R693 VDD.n40 VDD.n39 8.855
R694 VDD.n45 VDD.n44 8.855
R695 VDD.n44 VDD.n43 8.855
R696 VDD.n49 VDD.n48 8.855
R697 VDD.n48 VDD.n47 8.855
R698 VDD.n76 VDD.n75 8.855
R699 VDD.n75 VDD.n74 8.855
R700 VDD.n80 VDD.n79 8.855
R701 VDD.n79 VDD.n78 8.855
R702 VDD.n84 VDD.n83 8.855
R703 VDD.n83 VDD.n82 8.855
R704 VDD.n88 VDD.n87 8.855
R705 VDD.n87 VDD.n86 8.855
R706 VDD.n91 VDD.n90 8.855
R707 VDD.n90 0<p} 8.855
R708 VDD.n95 VDD.n94 8.855
R709 VDD.n94 VDD.n93 8.855
R710 VDD.n99 VDD.n98 8.855
R711 VDD.n98 VDD.n97 8.855
R712 VDD.n103 VDD.n102 8.855
R713 VDD.n102 VDD.n101 8.855
R714 VDD.n129 VDD.n128 8.855
R715 VDD.n128 VDD.n127 8.855
R716 VDD.n134 VDD.n133 8.855
R717 VDD.n133 VDD.n132 8.855
R718 VDD.n138 VDD.n137 8.855
R719 VDD.n137 VDD.n136 8.855
R720 VDD.n143 VDD.n142 8.855
R721 VDD.n142  <p} 8.855
R722 VDD.n147 VDD.n146 8.855
R723 VDD.n146 VDD.n145 8.855
R724 VDD.n151 VDD.n150 8.855
R725 VDD.n150 VDD.n149 8.855
R726 VDD.n156 VDD.n155 8.855
R727 VDD.n155 VDD.n154 8.855
R728 VDD.n160 VDD.n159 8.855
R729 VDD.n159 VDD.n158 8.855
R730 VDD.n186 VDD.n185 8.855
R731 VDD.n185 VDD.n184 8.855
R732 VDD.n191 VDD.n190 8.855
R733 VDD.n190 VDD.n189 8.855
R734 VDD.n195 VDD.n194 8.855
R735 VDD.n194 VDD.n193 8.855
R736 VDD.n200 VDD.n199 8.855
R737 VDD.n199 �;p} 8.855
R738 VDD.n204 VDD.n203 8.855
R739 VDD.n203 VDD.n202 8.855
R740 VDD.n208 VDD.n207 8.855
R741 VDD.n207 VDD.n206 8.855
R742 VDD.n213 VDD.n212 8.855
R743 VDD.n212 VDD.n211 8.855
R744 VDD.n217 VDD.n216 8.855
R745 VDD.n216 VDD.n215 8.855
R746 VDD.n243 VDD.n242 8.855
R747 VDD.n242 VDD.n241 8.855
R748 VDD.n248 VDD.n247 8.855
R749 VDD.n247 VDD.n246 8.855
R750 VDD.n252 VDD.n251 8.855
R751 VDD.n251 VDD.n250 8.855
R752 VDD.n257 VDD.n256 8.855
R753 VDD.n256  <p} 8.855
R754 VDD.n261 VDD.n260 8.855
R755 VDD.n260 VDD.n259 8.855
R756 VDD.n265 VDD.n264 8.855
R757 VDD.n264 VDD.n263 8.855
R758 VDD.n270 VDD.n269 8.855
R759 VDD.n269 VDD.n268 8.855
R760 VDD.n274 VDD.n273 8.855
R761 VDD.n273 VDD.n272 8.855
R762 VDD.n300 VDD.n299 8.855
R763 VDD.n299 VDD.n298 8.855
R764 VDD.n305 VDD.n304 8.855
R765 VDD.n304 VDD.n303 8.855
R766 VDD.n309 VDD.n308 8.855
R767 VDD.n308 VDD.n307 8.855
R768 VDD.n314 VDD.n313 8.855
R769 VDD.n313 �;p} 8.855
R770 VDD.n318 VDD.n317 8.855
R771 VDD.n317 VDD.n316 8.855
R772 VDD.n322 VDD.n321 8.855
R773 VDD.n321 VDD.n320 8.855
R774 VDD.n327 VDD.n326 8.855
R775 VDD.n326 VDD.n325 8.855
R776 VDD.n331 VDD.n330 8.855
R777 VDD.n330 VDD.n329 8.855
R778 VDD.n357 VDD.n356 8.855
R779 VDD.n356 VDD.n355 8.855
R780 VDD.n362 VDD.n361 8.855
R781 VDD.n361 VDD.n360 8.855
R782 VDD.n366 VDD.n365 8.855
R783 VDD.n365 VDD.n364 8.855
R784 VDD.n371 VDD.n370 8.855
R785 VDD.n370  <p} 8.855
R786 VDD.n375 VDD.n374 8.855
R787 VDD.n374 VDD.n373 8.855
R788 VDD.n379 VDD.n378 8.855
R789 VDD.n378 VDD.n377 8.855
R790 VDD.n384 VDD.n383 8.855
R791 VDD.n383 VDD.n382 8.855
R792 VDD.n388 VDD.n387 8.855
R793 VDD.n387 VDD.n386 8.855
R794 VDD.n414 VDD.n413 8.855
R795 VDD.n413 VDD.n412 8.855
R796 VDD.n419 VDD.n418 8.855
R797 VDD.n418 VDD.n417 8.855
R798 VDD.n423 VDD.n422 8.855
R799 VDD.n422 VDD.n421 8.855
R800 VDD.n428 VDD.n427 8.855
R801 VDD.n427  <p} 8.855
R802 VDD.n432 VDD.n431 8.855
R803 VDD.n431 VDD.n430 8.855
R804 VDD.n436 VDD.n435 8.855
R805 VDD.n435 VDD.n434 8.855
R806 VDD.n441 VDD.n440 8.855
R807 VDD.n440 VDD.n439 8.855
R808 VDD.n445 VDD.n444 8.855
R809 VDD.n444 VDD.n443 8.855
R810 VDD.n471 VDD.n470 8.855
R811 VDD.n470 VDD.n469 8.855
R812 VDD.n475 VDD.n474 8.855
R813 VDD.n474 VDD.n473 8.855
R814 VDD.n479 VDD.n478 8.855
R815 VDD.n478 VDD.n477 8.855
R816 VDD.n483 VDD.n482 8.855
R817 VDD.n482 VDD.n481 8.855
R818 VDD.n489 VDD.n486 8.855
R819 VDD.n486 VDD.n485 8.855
R820 VDD.n493 VDD.n492 8.855
R821 VDD.n492 VDD.n491 8.855
R822 VDD.n497 VDD.n496 8.855
R823 VDD.n496 VDD.n495 8.855
R824 VDD.n503 VDD.n502 8.855
R825 VDD.n502 VDD.n501 8.855
R826 VDD.n507 VDD.n506 8.855
R827 VDD.n506 VDD.n505 8.855
R828 VDD.n512 VDD.n511 8.855
R829 VDD.n511 VDD.n510 8.855
R830 VDD.n516 VDD.n515 8.855
R831 VDD.n515 VDD.n514 8.855
R832 VDD.n520 VDD.n519 8.855
R833 VDD.n519 VDD.n518 8.855
R834 VDD.n546 VDD.n545 8.855
R835 VDD.n545 VDD.n544 8.855
R836 VDD.n551 VDD.n550 8.855
R837 VDD.n550 VDD.n549 8.855
R838 VDD.n555 VDD.n554 8.855
R839 VDD.n554 VDD.n553 8.855
R840 VDD.n560 VDD.n559 8.855
R841 VDD.n559  <p} 8.855
R842 VDD.n564 VDD.n563 8.855
R843 VDD.n563 VDD.n562 8.855
R844 VDD.n568 VDD.n567 8.855
R845 VDD.n567 VDD.n566 8.855
R846 VDD.n573 VDD.n572 8.855
R847 VDD.n572 VDD.n571 8.855
R848 VDD.n577 VDD.n576 8.855
R849 VDD.n576 VDD.n575 8.855
R850 VDD.n603 VDD.n602 8.855
R851 VDD.n602 VDD.n601 8.855
R852 VDD.n608 VDD.n607 8.855
R853 VDD.n607 VDD.n606 8.855
R854 VDD.n612 VDD.n611 8.855
R855 VDD.n611 VDD.n610 8.855
R856 VDD.n617 VDD.n616 8.855
R857 VDD.n616 �;p} 8.855
R858 VDD.n621 VDD.n620 8.855
R859 VDD.n620 VDD.n619 8.855
R860 VDD.n625 VDD.n624 8.855
R861 VDD.n624 VDD.n623 8.855
R862 VDD.n1260 VDD.n1259 8.855
R863 VDD.n1259 VDD.n1258 8.855
R864 VDD.n1255 VDD.n1254 8.855
R865 VDD.n1254 VDD.n1253 8.855
R866 VDD.n1229 VDD.n1228 8.855
R867 VDD.n1228 VDD.n1227 8.855
R868 VDD.n1225 VDD.n1224 8.855
R869 VDD.n1224 VDD.n1223 8.855
R870 VDD.n1220 VDD.n1219 8.855
R871 VDD.n1219 VDD.n1218 8.855
R872 VDD.n1216 VDD.n1215 8.855
R873 VDD.n1215 �;p} 8.855
R874 VDD.n1211 VDD.n1210 8.855
R875 VDD.n1210 VDD.n1209 8.855
R876 VDD.n1207 VDD.n1206 8.855
R877 VDD.n1206 VDD.n1205 8.855
R878 VDD.n1203 VDD.n1202 8.855
R879 VDD.n1202 VDD.n1201 8.855
R880 VDD.n1198 VDD.n1197 8.855
R881 VDD.n1197 VDD.n1196 8.855
R882 VDD.n1172 VDD.n1171 8.855
R883 VDD.n1171 VDD.n1170 8.855
R884 VDD.n1168 VDD.n1167 8.855
R885 VDD.n1167 VDD.n1166 8.855
R886 VDD.n1163 VDD.n1162 8.855
R887 VDD.n1162 VDD.n1161 8.855
R888 VDD.n1159 VDD.n1158 8.855
R889 VDD.n1158 �;p} 8.855
R890 VDD.n1154 VDD.n1153 8.855
R891 VDD.n1153 VDD.n1152 8.855
R892 VDD.n1150 VDD.n1149 8.855
R893 VDD.n1149 VDD.n1148 8.855
R894 VDD.n1146 VDD.n1145 8.855
R895 VDD.n1145 VDD.n1144 8.855
R896 VDD.n1141 VDD.n1140 8.855
R897 VDD.n1140 VDD.n1139 8.855
R898 VDD.n1115 VDD.n1114 8.855
R899 VDD.n1114 VDD.n1113 8.855
R900 VDD.n1111 VDD.n1110 8.855
R901 VDD.n1110 VDD.n1109 8.855
R902 VDD.n1106 VDD.n1105 8.855
R903 VDD.n1105 VDD.n1104 8.855
R904 VDD.n1102 VDD.n1101 8.855
R905 VDD.n1101  <p} 8.855
R906 VDD.n1097 VDD.n1096 8.855
R907 VDD.n1096 VDD.n1095 8.855
R908 VDD.n1093 VDD.n1092 8.855
R909 VDD.n1092 VDD.n1091 8.855
R910 VDD.n1089 VDD.n1088 8.855
R911 VDD.n1088 VDD.n1087 8.855
R912 VDD.n1084 VDD.n1083 8.855
R913 VDD.n1083 VDD.n1082 8.855
R914 VDD.n1058 VDD.n1057 8.855
R915 VDD.n1057 VDD.n1056 8.855
R916 VDD.n1054 VDD.n1053 8.855
R917 VDD.n1053 VDD.n1052 8.855
R918 VDD.n1050 VDD.n1049 8.855
R919 VDD.n1049 VDD.n1048 8.855
R920 VDD.n1046 VDD.n1045 8.855
R921 VDD.n1045 VDD.n1044 8.855
R922 VDD.n1042 VDD.n1039 8.855
R923 VDD.n1039 VDD.n1038 8.855
R924 VDD.n1036 VDD.n1035 8.855
R925 VDD.n1035 VDD.n1034 8.855
R926 VDD.n1032 VDD.n1031 8.855
R927 VDD.n1031 VDD.n1030 8.855
R928 VDD.n1028 VDD.n1027 8.855
R929 VDD.n1027 VDD.n1026 8.855
R930 VDD.n1022 VDD.n1021 8.855
R931 VDD.n1021 VDD.n1020 8.855
R932 VDD.n1018 VDD.n1017 8.855
R933 VDD.n1017 VDD.n1016 8.855
R934 VDD.n1013 VDD.n1012 8.855
R935 VDD.n1012 VDD.n1011 8.855
R936 VDD.n1009 VDD.n1008 8.855
R937 VDD.n1008 VDD.n1007 8.855
R938 VDD.n983 VDD.n982 8.855
R939 VDD.n982 VDD.n981 8.855
R940 VDD.n979 VDD.n978 8.855
R941 VDD.n978 VDD.n977 8.855
R942 VDD.n974 VDD.n973 8.855
R943 VDD.n973 VDD.n972 8.855
R944 VDD.n970 VDD.n969 8.855
R945 VDD.n969 �;p} 8.855
R946 VDD.n965 VDD.n964 8.855
R947 VDD.n964 VDD.n963 8.855
R948 VDD.n961 VDD.n960 8.855
R949 VDD.n960 VDD.n959 8.855
R950 VDD.n957 VDD.n956 8.855
R951 VDD.n956 VDD.n955 8.855
R952 VDD.n952 VDD.n951 8.855
R953 VDD.n951 VDD.n950 8.855
R954 VDD.n926 VDD.n925 8.855
R955 VDD.n925 VDD.n924 8.855
R956 VDD.n922 VDD.n921 8.855
R957 VDD.n921 VDD.n920 8.855
R958 VDD.n917 VDD.n916 8.855
R959 VDD.n916 VDD.n915 8.855
R960 VDD.n913 VDD.n912 8.855
R961 VDD.n912 �;p} 8.855
R962 VDD.n908 VDD.n907 8.855
R963 VDD.n907 VDD.n906 8.855
R964 VDD.n904 VDD.n903 8.855
R965 VDD.n903 VDD.n902 8.855
R966 VDD.n900 VDD.n899 8.855
R967 VDD.n899 VDD.n898 8.855
R968 VDD.n895 VDD.n894 8.855
R969 VDD.n894 VDD.n893 8.855
R970 VDD.n869 VDD.n868 8.855
R971 VDD.n868 VDD.n867 8.855
R972 VDD.n865 VDD.n864 8.855
R973 VDD.n864 VDD.n863 8.855
R974 VDD.n860 VDD.n859 8.855
R975 VDD.n859 VDD.n858 8.855
R976 VDD.n856 VDD.n855 8.855
R977 VDD.n855 �;p} 8.855
R978 VDD.n851 VDD.n850 8.855
R979 VDD.n850 VDD.n849 8.855
R980 VDD.n847 VDD.n846 8.855
R981 VDD.n846 VDD.n845 8.855
R982 VDD.n843 VDD.n842 8.855
R983 VDD.n842 VDD.n841 8.855
R984 VDD.n838 VDD.n837 8.855
R985 VDD.n837 VDD.n836 8.855
R986 VDD.n812 VDD.n811 8.855
R987 VDD.n811 VDD.n810 8.855
R988 VDD.n808 VDD.n807 8.855
R989 VDD.n807 VDD.n806 8.855
R990 VDD.n803 VDD.n802 8.855
R991 VDD.n802 VDD.n801 8.855
R992 VDD.n799 VDD.n798 8.855
R993 VDD.n798  <p} 8.855
R994 VDD.n794 VDD.n793 8.855
R995 VDD.n793 VDD.n792 8.855
R996 VDD.n790 VDD.n789 8.855
R997 VDD.n789 VDD.n788 8.855
R998 VDD.n786 VDD.n785 8.855
R999 VDD.n785 VDD.n784 8.855
R1000 VDD.n781 VDD.n780 8.855
R1001 VDD.n780 VDD.n779 8.855
R1002 VDD.n755 VDD.n754 8.855
R1003 VDD.n754 VDD.n753 8.855
R1004 VDD.n751 VDD.n750 8.855
R1005 VDD.n750 VDD.n749 8.855
R1006 VDD.n746 VDD.n745 8.855
R1007 VDD.n745 VDD.n744 8.855
R1008 VDD.n742 VDD.n741 8.855
R1009 VDD.n741 �;p} 8.855
R1010 VDD.n737 VDD.n736 8.855
R1011 VDD.n736 VDD.n735 8.855
R1012 VDD.n733 VDD.n732 8.855
R1013 VDD.n732 VDD.n731 8.855
R1014 VDD.n729 VDD.n728 8.855
R1015 VDD.n728 VDD.n727 8.855
R1016 VDD.n724 VDD.n723 8.855
R1017 VDD.n723 VDD.n722 8.855
R1018 VDD.n697 VDD.n696 8.855
R1019 VDD.n696 VDD.n695 8.855
R1020 VDD.n693 VDD.n692 8.855
R1021 VDD.n692 VDD.n691 8.855
R1022 VDD.n689 VDD.n688 8.855
R1023 VDD.n688 VDD.n687 8.855
R1024 VDD.n685 VDD.n684 8.855
R1025 VDD.n684 VDD.n683 8.855
R1026 VDD.n681 VDD.n678 8.855
R1027 VDD.n678 VDD.n677 8.855
R1028 VDD.n675 VDD.n674 8.855
R1029 VDD.n674 VDD.n673 8.855
R1030 VDD.n671 VDD.n670 8.855
R1031 VDD.n670 VDD.n669 8.855
R1032 VDD.n667 VDD.n666 8.855
R1033 VDD.n666 VDD.n665 8.855
R1034 VDD.n661 VDD.n660 8.855
R1035 VDD.n660 VDD.n659 8.855
R1036 VDD.n657 VDD.n656 8.855
R1037 VDD.n656 VDD.n655 8.855
R1038 VDD.n652 VDD.n651 8.855
R1039 VDD.n651 VDD.n650 8.855
R1040 VDD.n648 VDD.n647 8.855
R1041 VDD.n647 VDD.n646 8.855
R1042 VDD.n772 VDD.n771 8.051
R1043 VDD.n829 VDD.n828 8.051
R1044 VDD.n886 VDD.n885 8.051
R1045 VDD.n943 VDD.n942 8.051
R1046 VDD.n1000 VDD.n999 8.051
R1047 VDD.n1075 VDD.n1074 8.051
R1048 VDD.n1132 VDD.n1131 8.051
R1049 VDD.n1189 VDD.n1188 8.051
R1050 VDD.n1246 VDD.n1245 8.051
R1051 VDD.n594 VDD.n593 8.051
R1052 VDD.n537 VDD.n536 8.051
R1053 VDD.n462 VDD.n461 8.051
R1054 VDD.n405 VDD.n404 8.051
R1055 VDD.n348 VDD.n347 8.051
R1056 VDD.n291 VDD.n290 8.051
R1057 VDD.n234 VDD.n233 8.051
R1058 VDD.n177 VDD.n176 8.051
R1059 VDD.n120 VDD.n119 8.051
R1060 VDD.n63 VDD.n62 8.051
R1061 VDD.n711 VDD.n710 8.051
R1062 VDD.n495  7.671
R1063 VDD.n1030  7.671
R1064 VDD.n669  <p} 7.671
R1065 VDD.n503 VDD.n500 7.019
R1066 VDD.n1028 VDD.n1025 7.019
R1067 VDD.n667 VDD.n664 7.019
R1068 VDD.n489 VDD.n488 6.606
R1069 VDD.n1042 VDD.n1041 6.606
R1070 VDD.n681 VDD.n680 6.606
R1071 VDD.n491 �;p} 5.114
R1072 VDD.n1034  <p} 5.114
R1073 VDD.n673 �;p} 5.114
R1074 VDD.n31 VDD.n30 4.65
R1075 VDD.n34 VDD.n33 4.65
R1076 VDD.n38 VDD.n37 4.65
R1077 VDD.n42 VDD.n41 4.65
R1078 VDD.n46 VDD.n45 4.65
R1079 VDD.n50 VDD.n49 4.65
R1080 VDD.n77 VDD.n76 4.65
R1081 VDD.n81 VDD.n80 4.65
R1082 VDD.n85 VDD.n84 4.65
R1083 VDD.n89 VDD.n88 4.65
R1084 VDD.n92 VDD.n91 4.65
R1085 VDD.n96 VDD.n95 4.65
R1086 VDD.n100 VDD.n99 4.65
R1087 VDD.n104 VDD.n103 4.65
R1088 VDD.n130 VDD.n129 4.65
R1089 VDD.n135 VDD.n134 4.65
R1090 VDD.n139 VDD.n138 4.65
R1091 VDD.n144 VDD.n143 4.65
R1092 VDD.n148 VDD.n147 4.65
R1093 VDD.n152 VDD.n151 4.65
R1094 VDD.n157 VDD.n156 4.65
R1095 VDD.n161 VDD.n160 4.65
R1096 VDD.n187 VDD.n186 4.65
R1097 VDD.n192 VDD.n191 4.65
R1098 VDD.n196 VDD.n195 4.65
R1099 VDD.n201 VDD.n200 4.65
R1100 VDD.n205 VDD.n204 4.65
R1101 VDD.n209 VDD.n208 4.65
R1102 VDD.n214 VDD.n213 4.65
R1103 VDD.n218 VDD.n217 4.65
R1104 VDD.n244 VDD.n243 4.65
R1105 VDD.n249 VDD.n248 4.65
R1106 VDD.n253 VDD.n252 4.65
R1107 VDD.n258 VDD.n257 4.65
R1108 VDD.n262 VDD.n261 4.65
R1109 VDD.n266 VDD.n265 4.65
R1110 VDD.n271 VDD.n270 4.65
R1111 VDD.n275 VDD.n274 4.65
R1112 VDD.n301 VDD.n300 4.65
R1113 VDD.n306 VDD.n305 4.65
R1114 VDD.n310 VDD.n309 4.65
R1115 VDD.n315 VDD.n314 4.65
R1116 VDD.n319 VDD.n318 4.65
R1117 VDD.n323 VDD.n322 4.65
R1118 VDD.n328 VDD.n327 4.65
R1119 VDD.n332 VDD.n331 4.65
R1120 VDD.n358 VDD.n357 4.65
R1121 VDD.n363 VDD.n362 4.65
R1122 VDD.n367 VDD.n366 4.65
R1123 VDD.n372 VDD.n371 4.65
R1124 VDD.n376 VDD.n375 4.65
R1125 VDD.n380 VDD.n379 4.65
R1126 VDD.n385 VDD.n384 4.65
R1127 VDD.n389 VDD.n388 4.65
R1128 VDD.n415 VDD.n414 4.65
R1129 VDD.n420 VDD.n419 4.65
R1130 VDD.n424 VDD.n423 4.65
R1131 VDD.n429 VDD.n428 4.65
R1132 VDD.n433 VDD.n432 4.65
R1133 VDD.n437 VDD.n436 4.65
R1134 VDD.n442 VDD.n441 4.65
R1135 VDD.n446 VDD.n445 4.65
R1136 VDD.n472 VDD.n471 4.65
R1137 VDD.n476 VDD.n475 4.65
R1138 VDD.n480 VDD.n479 4.65
R1139 VDD.n484 VDD.n483 4.65
R1140 VDD.n490 VDD.n489 4.65
R1141 VDD.n494 VDD.n493 4.65
R1142 VDD.n498 VDD.n497 4.65
R1143 VDD.n504 VDD.n503 4.65
R1144 VDD.n508 VDD.n507 4.65
R1145 VDD.n513 VDD.n512 4.65
R1146 VDD.n517 VDD.n516 4.65
R1147 VDD.n521 VDD.n520 4.65
R1148 VDD.n547 VDD.n546 4.65
R1149 VDD.n552 VDD.n551 4.65
R1150 VDD.n556 VDD.n555 4.65
R1151 VDD.n561 VDD.n560 4.65
R1152 VDD.n565 VDD.n564 4.65
R1153 VDD.n569 VDD.n568 4.65
R1154 VDD.n574 VDD.n573 4.65
R1155 VDD.n578 VDD.n577 4.65
R1156 VDD.n604 VDD.n603 4.65
R1157 VDD.n609 VDD.n608 4.65
R1158 VDD.n613 VDD.n612 4.65
R1159 VDD.n618 VDD.n617 4.65
R1160 VDD.n622 VDD.n621 4.65
R1161 VDD.n626 VDD.n625 4.65
R1162 VDD.n1261 VDD.n1260 4.65
R1163 VDD.n1256 VDD.n1255 4.65
R1164 VDD.n1230 VDD.n1229 4.65
R1165 VDD.n1226 VDD.n1225 4.65
R1166 VDD.n1221 VDD.n1220 4.65
R1167 VDD.n1217 VDD.n1216 4.65
R1168 VDD.n1212 VDD.n1211 4.65
R1169 VDD.n1208 VDD.n1207 4.65
R1170 VDD.n1204 VDD.n1203 4.65
R1171 VDD.n1199 VDD.n1198 4.65
R1172 VDD.n1173 VDD.n1172 4.65
R1173 VDD.n1169 VDD.n1168 4.65
R1174 VDD.n1164 VDD.n1163 4.65
R1175 VDD.n1160 VDD.n1159 4.65
R1176 VDD.n1155 VDD.n1154 4.65
R1177 VDD.n1151 VDD.n1150 4.65
R1178 VDD.n1147 VDD.n1146 4.65
R1179 VDD.n1142 VDD.n1141 4.65
R1180 VDD.n1116 VDD.n1115 4.65
R1181 VDD.n1112 VDD.n1111 4.65
R1182 VDD.n1107 VDD.n1106 4.65
R1183 VDD.n1103 VDD.n1102 4.65
R1184 VDD.n1098 VDD.n1097 4.65
R1185 VDD.n1094 VDD.n1093 4.65
R1186 VDD.n1090 VDD.n1089 4.65
R1187 VDD.n1085 VDD.n1084 4.65
R1188 VDD.n1059 VDD.n1058 4.65
R1189 VDD.n1055 VDD.n1054 4.65
R1190 VDD.n1051 VDD.n1050 4.65
R1191 VDD.n1047 VDD.n1046 4.65
R1192 VDD.n1043 VDD.n1042 4.65
R1193 VDD.n1037 VDD.n1036 4.65
R1194 VDD.n1033 VDD.n1032 4.65
R1195 VDD.n1029 VDD.n1028 4.65
R1196 VDD.n1023 VDD.n1022 4.65
R1197 VDD.n1019 VDD.n1018 4.65
R1198 VDD.n1014 VDD.n1013 4.65
R1199 VDD.n1010 VDD.n1009 4.65
R1200 VDD.n984 VDD.n983 4.65
R1201 VDD.n980 VDD.n979 4.65
R1202 VDD.n975 VDD.n974 4.65
R1203 VDD.n971 VDD.n970 4.65
R1204 VDD.n966 VDD.n965 4.65
R1205 VDD.n962 VDD.n961 4.65
R1206 VDD.n958 VDD.n957 4.65
R1207 VDD.n953 VDD.n952 4.65
R1208 VDD.n927 VDD.n926 4.65
R1209 VDD.n923 VDD.n922 4.65
R1210 VDD.n918 VDD.n917 4.65
R1211 VDD.n914 VDD.n913 4.65
R1212 VDD.n909 VDD.n908 4.65
R1213 VDD.n905 VDD.n904 4.65
R1214 VDD.n901 VDD.n900 4.65
R1215 VDD.n896 VDD.n895 4.65
R1216 VDD.n870 VDD.n869 4.65
R1217 VDD.n866 VDD.n865 4.65
R1218 VDD.n861 VDD.n860 4.65
R1219 VDD.n857 VDD.n856 4.65
R1220 VDD.n852 VDD.n851 4.65
R1221 VDD.n848 VDD.n847 4.65
R1222 VDD.n844 VDD.n843 4.65
R1223 VDD.n839 VDD.n838 4.65
R1224 VDD.n813 VDD.n812 4.65
R1225 VDD.n809 VDD.n808 4.65
R1226 VDD.n804 VDD.n803 4.65
R1227 VDD.n800 VDD.n799 4.65
R1228 VDD.n795 VDD.n794 4.65
R1229 VDD.n791 VDD.n790 4.65
R1230 VDD.n787 VDD.n786 4.65
R1231 VDD.n782 VDD.n781 4.65
R1232 VDD.n756 VDD.n755 4.65
R1233 VDD.n752 VDD.n751 4.65
R1234 VDD.n747 VDD.n746 4.65
R1235 VDD.n743 VDD.n742 4.65
R1236 VDD.n738 VDD.n737 4.65
R1237 VDD.n734 VDD.n733 4.65
R1238 VDD.n730 VDD.n729 4.65
R1239 VDD.n725 VDD.n724 4.65
R1240 VDD.n698 VDD.n697 4.65
R1241 VDD.n694 VDD.n693 4.65
R1242 VDD.n690 VDD.n689 4.65
R1243 VDD.n686 VDD.n685 4.65
R1244 VDD.n682 VDD.n681 4.65
R1245 VDD.n676 VDD.n675 4.65
R1246 VDD.n672 VDD.n671 4.65
R1247 VDD.n668 VDD.n667 4.65
R1248 VDD.n662 VDD.n661 4.65
R1249 VDD.n658 VDD.n657 4.65
R1250 VDD.n653 VDD.n652 4.65
R1251 VDD.n649 VDD.n648 4.65
R1252 VDD.n27 VDD.n23 2.933
R1253 VDD.n156 VDD.n153 2.89
R1254 VDD.n213 VDD.n210 2.89
R1255 VDD.n270 VDD.n267 2.89
R1256 VDD.n327 VDD.n324 2.89
R1257 VDD.n384 VDD.n381 2.89
R1258 VDD.n441 VDD.n438 2.89
R1259 VDD.n573 VDD.n570 2.89
R1260 VDD.n1260 VDD.n1257 2.89
R1261 VDD.n1203 VDD.n1200 2.89
R1262 VDD.n1146 VDD.n1143 2.89
R1263 VDD.n1089 VDD.n1086 2.89
R1264 VDD.n957 VDD.n954 2.89
R1265 VDD.n900 VDD.n897 2.89
R1266 VDD.n843 VDD.n840 2.89
R1267 VDD.n786 VDD.n783 2.89
R1268 VDD.n729 VDD.n726 2.89
R1269 VDD.n27 VDD.n26 2.844
R1270 VDD.n35  <p} 2.557
R1271 VDD.n86 �;p} 2.557
R1272 VDD.n145 �;p} 2.557
R1273 VDD.n202  <p} 2.557
R1274 VDD.n259  <p} 2.557
R1275 VDD.n316  <p} 2.557
R1276 VDD.n373 �;p} 2.557
R1277 VDD.n430  2.557
R1278 VDD.n562  <p} 2.557
R1279 VDD.n619  <p} 2.557
R1280 VDD.n1209  2.557
R1281 VDD.n1152 �;p} 2.557
R1282 VDD.n1095  2.557
R1283 VDD.n963 �;p} 2.557
R1284 VDD.n906  <p} 2.557
R1285 VDD.n849 p��IwU 2.557
R1286 VDD.n792 �;p} 2.557
R1287 VDD.n735 �;p} 2.557
R1288 VDD.n134 VDD.n131 2.477
R1289 VDD.n191 VDD.n188 2.477
R1290 VDD.n248 VDD.n245 2.477
R1291 VDD.n305 VDD.n302 2.477
R1292 VDD.n362 VDD.n359 2.477
R1293 VDD.n419 VDD.n416 2.477
R1294 VDD.n551 VDD.n548 2.477
R1295 VDD.n608 VDD.n605 2.477
R1296 VDD.n1225 VDD.n1222 2.477
R1297 VDD.n1168 VDD.n1165 2.477
R1298 VDD.n1111 VDD.n1108 2.477
R1299 VDD.n979 VDD.n976 2.477
R1300 VDD.n922 VDD.n919 2.477
R1301 VDD.n865 VDD.n862 2.477
R1302 VDD.n808 VDD.n805 2.477
R1303 VDD.n751 VDD.n748 2.477
R1304 VDD.n31 VDD.n27 1.063
R1305 VDD.n512 VDD.n509 0.412
R1306 VDD.n1018 VDD.n1015 0.412
R1307 VDD.n657 VDD.n654 0.412
R1308 VDD.n77 VDD.n50 0.29
R1309 VDD.n130 VDD.n104 0.29
R1310 VDD.n187 VDD.n161 0.29
R1311 VDD.n244 VDD.n218 0.29
R1312 VDD.n301 VDD.n275 0.29
R1313 VDD.n358 VDD.n332 0.29
R1314 VDD.n415 VDD.n389 0.29
R1315 VDD.n472 VDD.n446 0.29
R1316 VDD.n547 VDD.n521 0.29
R1317 VDD.n604 VDD.n578 0.29
R1318 VDD.n1256 VDD.n1230 0.29
R1319 VDD.n1199 VDD.n1173 0.29
R1320 VDD.n1142 VDD.n1116 0.29
R1321 VDD.n1085 VDD.n1059 0.29
R1322 VDD.n1010 VDD.n984 0.29
R1323 VDD.n953 VDD.n927 0.29
R1324 VDD.n896 VDD.n870 0.29
R1325 VDD.n839 VDD.n813 0.29
R1326 VDD.n782 VDD.n756 0.29
R1327 VDD.n725 VDD.n698 0.29
R1328 VDD.n649 VDD 0.207
R1329 VDD.n498 VDD.n494 0.197
R1330 VDD.n1037 VDD.n1033 0.197
R1331 VDD.n676 VDD.n672 0.197
R1332 VDD.n38 VDD.n34 0.181
R1333 VDD.n92 VDD.n89 0.181
R1334 VDD.n148 VDD.n144 0.181
R1335 VDD.n205 VDD.n201 0.181
R1336 VDD.n262 VDD.n258 0.181
R1337 VDD.n319 VDD.n315 0.181
R1338 VDD.n376 VDD.n372 0.181
R1339 VDD.n433 VDD.n429 0.181
R1340 VDD.n565 VDD.n561 0.181
R1341 VDD.n622 VDD.n618 0.181
R1342 VDD.n1217 VDD.n1212 0.181
R1343 VDD.n1160 VDD.n1155 0.181
R1344 VDD.n1103 VDD.n1098 0.181
R1345 VDD.n971 VDD.n966 0.181
R1346 VDD.n914 VDD.n909 0.181
R1347 VDD.n857 VDD.n852 0.181
R1348 VDD.n800 VDD.n795 0.181
R1349 VDD.n743 VDD.n738 0.181
R1350 VDD.n34 VDD.n31 0.145
R1351 VDD.n42 VDD.n38 0.145
R1352 VDD.n46 VDD.n42 0.145
R1353 VDD.n50 VDD.n46 0.145
R1354 VDD.n81 VDD.n77 0.145
R1355 VDD.n85 VDD.n81 0.145
R1356 VDD.n89 VDD.n85 0.145
R1357 VDD.n96 VDD.n92 0.145
R1358 VDD.n100 VDD.n96 0.145
R1359 VDD.n104 VDD.n100 0.145
R1360 VDD.n135 VDD.n130 0.145
R1361 VDD.n139 VDD.n135 0.145
R1362 VDD.n144 VDD.n139 0.145
R1363 VDD.n152 VDD.n148 0.145
R1364 VDD.n157 VDD.n152 0.145
R1365 VDD.n161 VDD.n157 0.145
R1366 VDD.n192 VDD.n187 0.145
R1367 VDD.n196 VDD.n192 0.145
R1368 VDD.n201 VDD.n196 0.145
R1369 VDD.n209 VDD.n205 0.145
R1370 VDD.n214 VDD.n209 0.145
R1371 VDD.n218 VDD.n214 0.145
R1372 VDD.n249 VDD.n244 0.145
R1373 VDD.n253 VDD.n249 0.145
R1374 VDD.n258 VDD.n253 0.145
R1375 VDD.n266 VDD.n262 0.145
R1376 VDD.n271 VDD.n266 0.145
R1377 VDD.n275 VDD.n271 0.145
R1378 VDD.n306 VDD.n301 0.145
R1379 VDD.n310 VDD.n306 0.145
R1380 VDD.n315 VDD.n310 0.145
R1381 VDD.n323 VDD.n319 0.145
R1382 VDD.n328 VDD.n323 0.145
R1383 VDD.n332 VDD.n328 0.145
R1384 VDD.n363 VDD.n358 0.145
R1385 VDD.n367 VDD.n363 0.145
R1386 VDD.n372 VDD.n367 0.145
R1387 VDD.n380 VDD.n376 0.145
R1388 VDD.n385 VDD.n380 0.145
R1389 VDD.n389 VDD.n385 0.145
R1390 VDD.n420 VDD.n415 0.145
R1391 VDD.n424 VDD.n420 0.145
R1392 VDD.n429 VDD.n424 0.145
R1393 VDD.n437 VDD.n433 0.145
R1394 VDD.n442 VDD.n437 0.145
R1395 VDD.n446 VDD.n442 0.145
R1396 VDD.n476 VDD.n472 0.145
R1397 VDD.n480 VDD.n476 0.145
R1398 VDD.n484 VDD.n480 0.145
R1399 VDD.n490 VDD.n484 0.145
R1400 VDD.n494 VDD.n490 0.145
R1401 VDD.n504 VDD.n498 0.145
R1402 VDD.n508 VDD.n504 0.145
R1403 VDD.n513 VDD.n508 0.145
R1404 VDD.n517 VDD.n513 0.145
R1405 VDD.n521 VDD.n517 0.145
R1406 VDD.n552 VDD.n547 0.145
R1407 VDD.n556 VDD.n552 0.145
R1408 VDD.n561 VDD.n556 0.145
R1409 VDD.n569 VDD.n565 0.145
R1410 VDD.n574 VDD.n569 0.145
R1411 VDD.n578 VDD.n574 0.145
R1412 VDD.n609 VDD.n604 0.145
R1413 VDD.n613 VDD.n609 0.145
R1414 VDD.n618 VDD.n613 0.145
R1415 VDD.n626 VDD.n622 0.145
R1416 VDD.n1261 VDD.n1256 0.145
R1417 VDD.n1230 VDD.n1226 0.145
R1418 VDD.n1226 VDD.n1221 0.145
R1419 VDD.n1221 VDD.n1217 0.145
R1420 VDD.n1212 VDD.n1208 0.145
R1421 VDD.n1208 VDD.n1204 0.145
R1422 VDD.n1204 VDD.n1199 0.145
R1423 VDD.n1173 VDD.n1169 0.145
R1424 VDD.n1169 VDD.n1164 0.145
R1425 VDD.n1164 VDD.n1160 0.145
R1426 VDD.n1155 VDD.n1151 0.145
R1427 VDD.n1151 VDD.n1147 0.145
R1428 VDD.n1147 VDD.n1142 0.145
R1429 VDD.n1116 VDD.n1112 0.145
R1430 VDD.n1112 VDD.n1107 0.145
R1431 VDD.n1107 VDD.n1103 0.145
R1432 VDD.n1098 VDD.n1094 0.145
R1433 VDD.n1094 VDD.n1090 0.145
R1434 VDD.n1090 VDD.n1085 0.145
R1435 VDD.n1059 VDD.n1055 0.145
R1436 VDD.n1055 VDD.n1051 0.145
R1437 VDD.n1051 VDD.n1047 0.145
R1438 VDD.n1047 VDD.n1043 0.145
R1439 VDD.n1043 VDD.n1037 0.145
R1440 VDD.n1033 VDD.n1029 0.145
R1441 VDD.n1029 VDD.n1023 0.145
R1442 VDD.n1023 VDD.n1019 0.145
R1443 VDD.n1019 VDD.n1014 0.145
R1444 VDD.n1014 VDD.n1010 0.145
R1445 VDD.n984 VDD.n980 0.145
R1446 VDD.n980 VDD.n975 0.145
R1447 VDD.n975 VDD.n971 0.145
R1448 VDD.n966 VDD.n962 0.145
R1449 VDD.n962 VDD.n958 0.145
R1450 VDD.n958 VDD.n953 0.145
R1451 VDD.n927 VDD.n923 0.145
R1452 VDD.n923 VDD.n918 0.145
R1453 VDD.n918 VDD.n914 0.145
R1454 VDD.n909 VDD.n905 0.145
R1455 VDD.n905 VDD.n901 0.145
R1456 VDD.n901 VDD.n896 0.145
R1457 VDD.n870 VDD.n866 0.145
R1458 VDD.n866 VDD.n861 0.145
R1459 VDD.n861 VDD.n857 0.145
R1460 VDD.n852 VDD.n848 0.145
R1461 VDD.n848 VDD.n844 0.145
R1462 VDD.n844 VDD.n839 0.145
R1463 VDD.n813 VDD.n809 0.145
R1464 VDD.n809 VDD.n804 0.145
R1465 VDD.n804 VDD.n800 0.145
R1466 VDD.n795 VDD.n791 0.145
R1467 VDD.n791 VDD.n787 0.145
R1468 VDD.n787 VDD.n782 0.145
R1469 VDD.n756 VDD.n752 0.145
R1470 VDD.n752 VDD.n747 0.145
R1471 VDD.n747 VDD.n743 0.145
R1472 VDD.n738 VDD.n734 0.145
R1473 VDD.n734 VDD.n730 0.145
R1474 VDD.n730 VDD.n725 0.145
R1475 VDD.n698 VDD.n694 0.145
R1476 VDD.n694 VDD.n690 0.145
R1477 VDD.n690 VDD.n686 0.145
R1478 VDD.n686 VDD.n682 0.145
R1479 VDD.n682 VDD.n676 0.145
R1480 VDD.n672 VDD.n668 0.145
R1481 VDD.n668 VDD.n662 0.145
R1482 VDD.n662 VDD.n658 0.145
R1483 VDD.n658 VDD.n653 0.145
R1484 VDD.n653 VDD.n649 0.145
R1485 VDD VDD.n1261 0.082
R1486 VDD VDD.n626 0.062
R1487 a_277_1050.n7 a_277_1050.t9 480.392
R1488 a_277_1050.n5 a_277_1050.t10 480.392
R1489 a_277_1050.n7 a_277_1050.t11 403.272
R1490 a_277_1050.n5 a_277_1050.t7 403.272
R1491 a_277_1050.n8 a_277_1050.t12 385.063
R1492 a_277_1050.n6 a_277_1050.t8 385.063
R1493 a_277_1050.n12 a_277_1050.n10 342.597
R1494 a_277_1050.n3 a_277_1050.n2 161.352
R1495 a_277_1050.n10 a_277_1050.n4 151.34
R1496 a_277_1050.n8 a_277_1050.n7 143.429
R1497 a_277_1050.n6 a_277_1050.n5 143.429
R1498 a_277_1050.n4 a_277_1050.n0 95.095
R1499 a_277_1050.n3 a_277_1050.n1 95.095
R1500 a_277_1050.n4 a_277_1050.n3 66.258
R1501 a_277_1050.n12 a_277_1050.n11 15.218
R1502 a_277_1050.n0 a_277_1050.t1 14.282
R1503 a_277_1050.n0 a_277_1050.t3 14.282
R1504 a_277_1050.n1 a_277_1050.t5 14.282
R1505 a_277_1050.n1 a_277_1050.t4 14.282
R1506 a_277_1050.n2 a_277_1050.t2 14.282
R1507 a_277_1050.n2 a_277_1050.t0 14.282
R1508 a_277_1050.n13 a_277_1050.n12 12.014
R1509 a_277_1050.n9 a_277_1050.n6 11.95
R1510 a_277_1050.n10 a_277_1050.n9 5.965
R1511 a_277_1050.n9 a_277_1050.n8 4.65
R1512 a_3177_1050.n1 a_3177_1050.t7 480.392
R1513 a_3177_1050.n1 a_3177_1050.t5 403.272
R1514 a_3177_1050.n2 a_3177_1050.t6 385.063
R1515 a_3177_1050.n4 a_3177_1050.n3 355.179
R1516 a_3177_1050.n6 a_3177_1050.n5 157.963
R1517 a_3177_1050.n2 a_3177_1050.n1 143.429
R1518 a_3177_1050.n5 a_3177_1050.n4 132.141
R1519 a_3177_1050.n5 a_3177_1050.n0 91.706
R1520 a_3177_1050.n0 a_3177_1050.t2 14.282
R1521 a_3177_1050.n0 a_3177_1050.t1 14.282
R1522 a_3177_1050.n6 a_3177_1050.t3 14.282
R1523 a_3177_1050.t4 a_3177_1050.n6 14.282
R1524 a_3177_1050.n4 a_3177_1050.n2 10.615
R1525 a_1845_1050.n3 a_1845_1050.t5 480.392
R1526 a_1845_1050.n3 a_1845_1050.t7 403.272
R1527 a_1845_1050.n4 a_1845_1050.t6 357.204
R1528 a_1845_1050.n7 a_1845_1050.n5 312.103
R1529 a_1845_1050.n4 a_1845_1050.n3 171.288
R1530 a_1845_1050.n5 a_1845_1050.n2 159.999
R1531 a_1845_1050.n2 a_1845_1050.n1 157.964
R1532 a_1845_1050.n2 a_1845_1050.n0 91.706
R1533 a_1845_1050.n7 a_1845_1050.n6 15.218
R1534 a_1845_1050.n0 a_1845_1050.t1 14.282
R1535 a_1845_1050.n0 a_1845_1050.t3 14.282
R1536 a_1845_1050.n1 a_1845_1050.t0 14.282
R1537 a_1845_1050.n1 a_1845_1050.t4 14.282
R1538 a_1845_1050.n8 a_1845_1050.n7 12.014
R1539 a_1845_1050.n5 a_1845_1050.n4 10.615
R1540 a_147_187.n5 a_147_187.t13 512.525
R1541 a_147_187.n3 a_147_187.t11 472.359
R1542 a_147_187.n1 a_147_187.t6 472.359
R1543 a_147_187.n6 a_147_187.t10 417.109
R1544 a_147_187.n3 a_147_187.t7 384.527
R1545 a_147_187.n1 a_147_187.t8 384.527
R1546 a_147_187.n10 a_147_187.n9 383.037
R1547 a_147_187.n5 a_147_187.t9 371.139
R1548 a_147_187.n4 a_147_187.t12 370.613
R1549 a_147_187.n2 a_147_187.t5 370.613
R1550 a_147_187.n6 a_147_187.n5 179.837
R1551 a_147_187.n12 a_147_187.n11 157.963
R1552 a_147_187.n4 a_147_187.n3 127.096
R1553 a_147_187.n2 a_147_187.n1 127.096
R1554 a_147_187.n11 a_147_187.n10 104.282
R1555 a_147_187.n11 a_147_187.n0 91.706
R1556 a_147_187.n0 a_147_187.t4 14.282
R1557 a_147_187.n0 a_147_187.t3 14.282
R1558 a_147_187.t1 a_147_187.n12 14.282
R1559 a_147_187.n12 a_147_187.t0 14.282
R1560 a_147_187.n7 a_147_187.n6 11.134
R1561 a_147_187.n8 a_147_187.n2 8.957
R1562 a_147_187.n7 a_147_187.n4 4.65
R1563 a_147_187.n10 a_147_187.n8 4.65
R1564 a_147_187.n8 a_147_187.n7 2.947
R1565 a_3303_411.n2 a_3303_411.t8 512.525
R1566 a_3303_411.n1 a_3303_411.t11 512.525
R1567 a_3303_411.n6 a_3303_411.t13 472.359
R1568 a_3303_411.n6 a_3303_411.t7 384.527
R1569 a_3303_411.n2 a_3303_411.t12 371.139
R1570 a_3303_411.n1 a_3303_411.t9 371.139
R1571 a_3303_411.n3 a_3303_411.n2 343.521
R1572 a_3303_411.n7 a_3303_411.t10 287.037
R1573 a_3303_411.n13 a_3303_411.n12 277.722
R1574 a_3303_411.n5 a_3303_411.n1 259.945
R1575 a_3303_411.n7 a_3303_411.n6 210.673
R1576 a_3303_411.n14 a_3303_411.n13 187.858
R1577 a_3303_411.n3 a_3303_411.t6 172.106
R1578 a_3303_411.n4 a_3303_411.t5 165.68
R1579 a_3303_411.n15 a_3303_411.n14 157.963
R1580 a_3303_411.n14 a_3303_411.n0 91.706
R1581 a_3303_411.n5 a_3303_411.n4 83.576
R1582 a_3303_411.n8 a_3303_411.n5 41.06
R1583 a_3303_411.n12 a_3303_411.n11 30
R1584 a_3303_411.n10 a_3303_411.n9 24.383
R1585 a_3303_411.n12 a_3303_411.n10 23.684
R1586 a_3303_411.n0 a_3303_411.t4 14.282
R1587 a_3303_411.n0 a_3303_411.t3 14.282
R1588 a_3303_411.n15 a_3303_411.t0 14.282
R1589 a_3303_411.t1 a_3303_411.n15 14.282
R1590 a_3303_411.n4 a_3303_411.n3 10.343
R1591 a_3303_411.n8 a_3303_411.n7 7.597
R1592 a_3303_411.n13 a_3303_411.n8 4.65
R1593 a_13654_101.t0 a_13654_101.n0 93.333
R1594 a_13654_101.n3 a_13654_101.n1 79.062
R1595 a_13654_101.n3 a_13654_101.n2 2.084
R1596 a_13654_101.t0 a_13654_101.n3 0.182
R1597 QN.n10 QN.n9 227.387
R1598 QN.n2 QN.n1 165.613
R1599 QN.n7 QN.n6 134.51
R1600 QN.n10 QN.n2 132.893
R1601 QN.n9 QN.n8 127.909
R1602 QN.n7 QN.n5 126.225
R1603 QN.n2 QN.n0 99.355
R1604 QN.n5 QN.n4 22.578
R1605 QN.n0 QN.t1 14.282
R1606 QN.n0 QN.t6 14.282
R1607 QN.n1 QN.t2 14.282
R1608 QN.n1 QN.t3 14.282
R1609 QN.n5 QN.n3 8.58
R1610 QN.n9 QN.n7 7.053
R1611 QN.n11 QN.n10 4.65
R1612 QN.n11 QN 0.046
R1613 GND.n31 GND.n30 237.558
R1614 GND.n389 GND.n388 237.558
R1615 GND.n422 GND.n421 237.558
R1616 GND.n452 GND.n451 237.558
R1617 GND.n485 GND.n484 237.558
R1618 GND.n518 GND.n517 237.558
R1619 GND.n551 GND.n550 237.558
R1620 GND.n595 GND.n594 237.558
R1621 GND.n627 GND.n626 237.558
R1622 GND.n659 GND.n658 237.558
R1623 GND.n324 GND.n323 237.558
R1624 GND.n689 GND.n688 237.558
R1625 GND.n294 GND.n293 237.558
R1626 GND.n249 GND.n248 237.558
R1627 GND.n216 GND.n215 237.558
R1628 GND.n186 GND.n185 237.558
R1629 GND.n156 GND.n155 237.558
R1630 GND.n123 GND.n122 237.558
R1631 GND.n93 GND.n92 237.558
R1632 GND.n61 GND.n60 237.558
R1633 GND.n28 GND.n27 210.82
R1634 GND.n58 GND.n57 210.82
R1635 GND.n391 GND.n390 210.82
R1636 GND.n424 GND.n423 210.82
R1637 GND.n454 GND.n453 210.82
R1638 GND.n487 GND.n486 210.82
R1639 GND.n520 GND.n519 210.82
R1640 GND.n553 GND.n552 210.82
R1641 GND.n597 GND.n596 210.82
R1642 GND.n629 GND.n628 210.82
R1643 GND.n661 GND.n660 210.82
R1644 GND.n691 GND.n690 210.82
R1645 GND.n321 GND.n320 210.82
R1646 GND.n291 GND.n290 210.82
R1647 GND.n246 GND.n245 210.82
R1648 GND.n213 GND.n212 210.82
R1649 GND.n183 GND.n182 210.82
R1650 GND.n153 GND.n152 210.82
R1651 GND.n120 GND.n119 210.82
R1652 GND.n90 GND.n89 210.82
R1653 GND.n47 GND.n46 172.612
R1654 GND.n109 GND.n108 172.612
R1655 GND.n172 GND.n171 172.612
R1656 GND.n202 GND.n201 172.612
R1657 GND.n310 GND.n309 172.612
R1658 GND.n669 GND.n668 172.612
R1659 GND.n432 GND.n431 172.612
R1660 GND.n564 GND.n563 167.358
R1661 GND.n79 GND.n78 166.605
R1662 GND.n639 GND.n638 166.605
R1663 GND.n607 GND.n606 166.605
R1664 GND.n281 GND.n280 152.358
R1665 GND.n358 GND.n357 152.358
R1666 GND.n142 GND.n141 151.605
R1667 GND.n235 GND.n234 151.605
R1668 GND.n343 GND.n342 151.605
R1669 GND.n531 GND.n530 151.605
R1670 GND.n498 GND.n497 151.605
R1671 GND.n465 GND.n464 151.605
R1672 GND.n402 GND.n401 151.605
R1673 GND.n17 GND.n16 151.605
R1674 GND.n141 GND.n140 28.421
R1675 GND.n234 GND.n233 28.421
R1676 GND.n280 GND.n279 28.421
R1677 GND.n342 GND.n341 28.421
R1678 GND.n530 GND.n529 28.421
R1679 GND.n497 GND.n496 28.421
R1680 GND.n464 GND.n463 28.421
R1681 GND.n401 GND.n400 28.421
R1682 GND.n357 GND.n356 28.421
R1683 GND.n16 GND.n15 28.421
R1684 GND.n141 GND.n139 25.263
R1685 GND.n234 GND.n232 25.263
R1686 GND.n280 GND.n278 25.263
R1687 GND.n342 GND.n340 25.263
R1688 GND.n530 GND.n528 25.263
R1689 GND.n497 GND.n495 25.263
R1690 GND.n464 GND.n462 25.263
R1691 GND.n401 GND.n399 25.263
R1692 GND.n357 GND.n355 25.263
R1693 GND.n16 GND.n14 25.263
R1694 GND.n139 GND.n138 24.383
R1695 GND.n232 GND.n231 24.383
R1696 GND.n278 GND.n277 24.383
R1697 GND.n340 GND.n339 24.383
R1698 GND.n528 GND.n527 24.383
R1699 GND.n495 GND.n494 24.383
R1700 GND.n462 GND.n461 24.383
R1701 GND.n399 GND.n398 24.383
R1702 GND.n355 GND.n354 24.383
R1703 GND.n14 GND.n13 24.383
R1704 GND.n78 GND.n76 23.03
R1705 GND.n638 GND.n636 23.03
R1706 GND.n606 GND.n604 23.03
R1707 GND.n563 GND.n561 23.03
R1708 GND.n29 GND.n28 18.953
R1709 GND.n59 GND.n58 18.953
R1710 GND.n392 GND.n391 18.953
R1711 GND.n425 GND.n424 18.953
R1712 GND.n455 GND.n454 18.953
R1713 GND.n488 GND.n487 18.953
R1714 GND.n521 GND.n520 18.953
R1715 GND.n554 GND.n553 18.953
R1716 GND.n598 GND.n597 18.953
R1717 GND.n630 GND.n629 18.953
R1718 GND.n662 GND.n661 18.953
R1719 GND.n692 GND.n691 18.953
R1720 GND.n322 GND.n321 18.953
R1721 GND.n292 GND.n291 18.953
R1722 GND.n247 GND.n246 18.953
R1723 GND.n214 GND.n213 18.953
R1724 GND.n184 GND.n183 18.953
R1725 GND.n154 GND.n153 18.953
R1726 GND.n121 GND.n120 18.953
R1727 GND.n91 GND.n90 18.953
R1728 GND.n32 GND.n29 14.864
R1729 GND.n62 GND.n59 14.864
R1730 GND.n94 GND.n91 14.864
R1731 GND.n124 GND.n121 14.864
R1732 GND.n157 GND.n154 14.864
R1733 GND.n187 GND.n184 14.864
R1734 GND.n217 GND.n214 14.864
R1735 GND.n250 GND.n247 14.864
R1736 GND.n295 GND.n292 14.864
R1737 GND.n325 GND.n322 14.864
R1738 GND.n693 GND.n692 14.864
R1739 GND.n663 GND.n662 14.864
R1740 GND.n631 GND.n630 14.864
R1741 GND.n599 GND.n598 14.864
R1742 GND.n555 GND.n554 14.864
R1743 GND.n522 GND.n521 14.864
R1744 GND.n489 GND.n488 14.864
R1745 GND.n456 GND.n455 14.864
R1746 GND.n426 GND.n425 14.864
R1747 GND.n393 GND.n392 14.864
R1748 GND.n351 GND.n350 9.154
R1749 GND.n359 GND.n353 9.154
R1750 GND.n362 GND.n361 9.154
R1751 GND.n365 GND.n364 9.154
R1752 GND.n368 GND.n367 9.154
R1753 GND.n371 GND.n370 9.154
R1754 GND.n374 GND.n373 9.154
R1755 GND.n377 GND.n376 9.154
R1756 GND.n380 GND.n379 9.154
R1757 GND.n383 GND.n382 9.154
R1758 GND.n386 GND.n385 9.154
R1759 GND.n393 GND.n389 9.154
R1760 GND.n396 GND.n395 9.154
R1761 GND.n404 GND.n403 9.154
R1762 GND.n407 GND.n406 9.154
R1763 GND.n410 GND.n409 9.154
R1764 GND.n413 GND.n412 9.154
R1765 GND.n416 GND.n415 9.154
R1766 GND.n419 GND.n418 9.154
R1767 GND.n426 GND.n422 9.154
R1768 GND.n429 GND.n428 9.154
R1769 GND.n434 GND.n433 9.154
R1770 GND.n437 GND.n436 9.154
R1771 GND.n440 GND.n439 9.154
R1772 GND.n443 GND.n442 9.154
R1773 GND.n446 GND.n445 9.154
R1774 GND.n449 GND.n448 9.154
R1775 GND.n456 GND.n452 9.154
R1776 GND.n459 GND.n458 9.154
R1777 GND.n467 GND.n466 9.154
R1778 GND.n470 GND.n469 9.154
R1779 GND.n473 GND.n472 9.154
R1780 GND.n476 GND.n475 9.154
R1781 GND.n479 GND.n478 9.154
R1782 GND.n482 GND.n481 9.154
R1783 GND.n489 GND.n485 9.154
R1784 GND.n492 GND.n491 9.154
R1785 GND.n500 GND.n499 9.154
R1786 GND.n503 GND.n502 9.154
R1787 GND.n506 GND.n505 9.154
R1788 GND.n509 GND.n508 9.154
R1789 GND.n512 GND.n511 9.154
R1790 GND.n515 GND.n514 9.154
R1791 GND.n522 GND.n518 9.154
R1792 GND.n525 GND.n524 9.154
R1793 GND.n533 GND.n532 9.154
R1794 GND.n536 GND.n535 9.154
R1795 GND.n539 GND.n538 9.154
R1796 GND.n542 GND.n541 9.154
R1797 GND.n545 GND.n544 9.154
R1798 GND.n548 GND.n547 9.154
R1799 GND.n555 GND.n551 9.154
R1800 GND.n558 GND.n557 9.154
R1801 GND.n565 GND.n560 9.154
R1802 GND.n568 GND.n567 9.154
R1803 GND.n571 GND.n570 9.154
R1804 GND.n574 GND.n573 9.154
R1805 GND.n577 GND.n576 9.154
R1806 GND.n580 GND.n579 9.154
R1807 GND.n583 GND.n582 9.154
R1808 GND.n586 GND.n585 9.154
R1809 GND.n589 GND.n588 9.154
R1810 GND.n592 GND.n591 9.154
R1811 GND.n599 GND.n595 9.154
R1812 GND.n602 GND.n601 9.154
R1813 GND.n609 GND.n608 9.154
R1814 GND.n612 GND.n611 9.154
R1815 GND.n615 GND.n614 9.154
R1816 GND.n618 GND.n617 9.154
R1817 GND.n621 GND.n620 9.154
R1818 GND.n624 GND.n623 9.154
R1819 GND.n631 GND.n627 9.154
R1820 GND.n634 GND.n633 9.154
R1821 GND.n641 GND.n640 9.154
R1822 GND.n644 GND.n643 9.154
R1823 GND.n647 GND.n646 9.154
R1824 GND.n650 GND.n649 9.154
R1825 GND.n653 GND.n652 9.154
R1826 GND.n656 GND.n655 9.154
R1827 GND.n663 GND.n659 9.154
R1828 GND.n666 GND.n665 9.154
R1829 GND.n671 GND.n670 9.154
R1830 GND.n674 GND.n673 9.154
R1831 GND.n677 GND.n676 9.154
R1832 GND.n680 GND.n679 9.154
R1833 GND.n683 GND.n682 9.154
R1834 GND.n686 GND.n685 9.154
R1835 GND.n693 GND.n689 9.154
R1836 GND.n696 GND.n695 9.154
R1837 GND.n345 GND.n344 9.154
R1838 GND.n337 GND.n336 9.154
R1839 GND.n334 GND.n333 9.154
R1840 GND.n331 GND.n330 9.154
R1841 GND.n328 GND.n327 9.154
R1842 GND.n325 GND.n324 9.154
R1843 GND.n318 GND.n317 9.154
R1844 GND.n315 GND.n314 9.154
R1845 GND.n312 GND.n311 9.154
R1846 GND.n307 GND.n306 9.154
R1847 GND.n304 GND.n303 9.154
R1848 GND.n301 GND.n300 9.154
R1849 GND.n298 GND.n297 9.154
R1850 GND.n295 GND.n294 9.154
R1851 GND.n288 GND.n287 9.154
R1852 GND.n285 GND.n284 9.154
R1853 GND.n282 GND.n276 9.154
R1854 GND.n274 GND.n273 9.154
R1855 GND.n271 GND.n270 9.154
R1856 GND.n268 GND.n267 9.154
R1857 GND.n265 GND.n264 9.154
R1858 GND.n262 GND.n261 9.154
R1859 GND.n259 GND.n258 9.154
R1860 GND.n256 GND.n255 9.154
R1861 GND.n253 GND.n252 9.154
R1862 GND.n250 GND.n249 9.154
R1863 GND.n243 GND.n242 9.154
R1864 GND.n240 GND.n239 9.154
R1865 GND.n237 GND.n236 9.154
R1866 GND.n229 GND.n228 9.154
R1867 GND.n226 GND.n225 9.154
R1868 GND.n223 GND.n222 9.154
R1869 GND.n220 GND.n219 9.154
R1870 GND.n217 GND.n216 9.154
R1871 GND.n210 GND.n209 9.154
R1872 GND.n207 GND.n206 9.154
R1873 GND.n204 GND.n203 9.154
R1874 GND.n199 GND.n198 9.154
R1875 GND.n196 GND.n195 9.154
R1876 GND.n193 GND.n192 9.154
R1877 GND.n190 GND.n189 9.154
R1878 GND.n187 GND.n186 9.154
R1879 GND.n180 GND.n179 9.154
R1880 GND.n177 GND.n176 9.154
R1881 GND.n174 GND.n173 9.154
R1882 GND.n169 GND.n168 9.154
R1883 GND.n166 GND.n165 9.154
R1884 GND.n163 GND.n162 9.154
R1885 GND.n160 GND.n159 9.154
R1886 GND.n157 GND.n156 9.154
R1887 GND.n150 GND.n149 9.154
R1888 GND.n147 GND.n146 9.154
R1889 GND.n144 GND.n143 9.154
R1890 GND.n136 GND.n135 9.154
R1891 GND.n133 GND.n132 9.154
R1892 GND.n130 GND.n129 9.154
R1893 GND.n127 GND.n126 9.154
R1894 GND.n124 GND.n123 9.154
R1895 GND.n117 GND.n116 9.154
R1896 GND.n114 GND.n113 9.154
R1897 GND.n111 GND.n110 9.154
R1898 GND.n106 GND.n105 9.154
R1899 GND.n103 GND.n102 9.154
R1900 GND.n100 GND.n99 9.154
R1901 GND.n97 GND.n96 9.154
R1902 GND.n94 GND.n93 9.154
R1903 GND.n87 GND.n86 9.154
R1904 GND.n84 GND.n83 9.154
R1905 GND.n81 GND.n80 9.154
R1906 GND.n74 GND.n73 9.154
R1907 GND.n71 GND.n70 9.154
R1908 GND.n68 GND.n67 9.154
R1909 GND.n65 GND.n64 9.154
R1910 GND.n62 GND.n61 9.154
R1911 GND.n55 GND.n54 9.154
R1912 GND.n52 GND.n51 9.154
R1913 GND.n49 GND.n48 9.154
R1914 GND.n44 GND.n43 9.154
R1915 GND.n41 GND.n40 9.154
R1916 GND.n1 GND.n0 9.154
R1917 GND.n5 GND.n4 9.154
R1918 GND.n8 GND.n7 9.154
R1919 GND.n11 GND.n10 9.154
R1920 GND.n19 GND.n18 9.154
R1921 GND.n22 GND.n21 9.154
R1922 GND.n25 GND.n24 9.154
R1923 GND.n32 GND.n31 9.154
R1924 GND.n35 GND.n34 9.154
R1925 GND.n38 GND.n37 9.154
R1926 GND.n78 GND.n77 8.128
R1927 GND.n638 GND.n637 8.128
R1928 GND.n606 GND.n605 8.128
R1929 GND.n563 GND.n562 8.128
R1930 GND.n349 GND.n348 4.65
R1931 GND.n42 GND.n41 4.65
R1932 GND.n45 GND.n44 4.65
R1933 GND.n50 GND.n49 4.65
R1934 GND.n53 GND.n52 4.65
R1935 GND.n56 GND.n55 4.65
R1936 GND.n63 GND.n62 4.65
R1937 GND.n66 GND.n65 4.65
R1938 GND.n69 GND.n68 4.65
R1939 GND.n72 GND.n71 4.65
R1940 GND.n75 GND.n74 4.65
R1941 GND.n82 GND.n81 4.65
R1942 GND.n85 GND.n84 4.65
R1943 GND.n88 GND.n87 4.65
R1944 GND.n95 GND.n94 4.65
R1945 GND.n98 GND.n97 4.65
R1946 GND.n101 GND.n100 4.65
R1947 GND.n104 GND.n103 4.65
R1948 GND.n107 GND.n106 4.65
R1949 GND.n112 GND.n111 4.65
R1950 GND.n115 GND.n114 4.65
R1951 GND.n118 GND.n117 4.65
R1952 GND.n125 GND.n124 4.65
R1953 GND.n128 GND.n127 4.65
R1954 GND.n131 GND.n130 4.65
R1955 GND.n134 GND.n133 4.65
R1956 GND.n137 GND.n136 4.65
R1957 GND.n145 GND.n144 4.65
R1958 GND.n148 GND.n147 4.65
R1959 GND.n151 GND.n150 4.65
R1960 GND.n158 GND.n157 4.65
R1961 GND.n161 GND.n160 4.65
R1962 GND.n164 GND.n163 4.65
R1963 GND.n167 GND.n166 4.65
R1964 GND.n170 GND.n169 4.65
R1965 GND.n175 GND.n174 4.65
R1966 GND.n178 GND.n177 4.65
R1967 GND.n181 GND.n180 4.65
R1968 GND.n188 GND.n187 4.65
R1969 GND.n191 GND.n190 4.65
R1970 GND.n194 GND.n193 4.65
R1971 GND.n197 GND.n196 4.65
R1972 GND.n200 GND.n199 4.65
R1973 GND.n205 GND.n204 4.65
R1974 GND.n208 GND.n207 4.65
R1975 GND.n211 GND.n210 4.65
R1976 GND.n218 GND.n217 4.65
R1977 GND.n221 GND.n220 4.65
R1978 GND.n224 GND.n223 4.65
R1979 GND.n227 GND.n226 4.65
R1980 GND.n230 GND.n229 4.65
R1981 GND.n238 GND.n237 4.65
R1982 GND.n241 GND.n240 4.65
R1983 GND.n244 GND.n243 4.65
R1984 GND.n251 GND.n250 4.65
R1985 GND.n254 GND.n253 4.65
R1986 GND.n257 GND.n256 4.65
R1987 GND.n260 GND.n259 4.65
R1988 GND.n263 GND.n262 4.65
R1989 GND.n266 GND.n265 4.65
R1990 GND.n269 GND.n268 4.65
R1991 GND.n272 GND.n271 4.65
R1992 GND.n275 GND.n274 4.65
R1993 GND.n283 GND.n282 4.65
R1994 GND.n286 GND.n285 4.65
R1995 GND.n289 GND.n288 4.65
R1996 GND.n296 GND.n295 4.65
R1997 GND.n299 GND.n298 4.65
R1998 GND.n302 GND.n301 4.65
R1999 GND.n305 GND.n304 4.65
R2000 GND.n308 GND.n307 4.65
R2001 GND.n313 GND.n312 4.65
R2002 GND.n316 GND.n315 4.65
R2003 GND.n319 GND.n318 4.65
R2004 GND.n326 GND.n325 4.65
R2005 GND.n329 GND.n328 4.65
R2006 GND.n332 GND.n331 4.65
R2007 GND.n335 GND.n334 4.65
R2008 GND.n338 GND.n337 4.65
R2009 GND.n346 GND.n345 4.65
R2010 GND.n697 GND.n696 4.65
R2011 GND.n694 GND.n693 4.65
R2012 GND.n687 GND.n686 4.65
R2013 GND.n684 GND.n683 4.65
R2014 GND.n681 GND.n680 4.65
R2015 GND.n678 GND.n677 4.65
R2016 GND.n675 GND.n674 4.65
R2017 GND.n672 GND.n671 4.65
R2018 GND.n667 GND.n666 4.65
R2019 GND.n664 GND.n663 4.65
R2020 GND.n657 GND.n656 4.65
R2021 GND.n654 GND.n653 4.65
R2022 GND.n651 GND.n650 4.65
R2023 GND.n648 GND.n647 4.65
R2024 GND.n645 GND.n644 4.65
R2025 GND.n642 GND.n641 4.65
R2026 GND.n635 GND.n634 4.65
R2027 GND.n632 GND.n631 4.65
R2028 GND.n625 GND.n624 4.65
R2029 GND.n622 GND.n621 4.65
R2030 GND.n619 GND.n618 4.65
R2031 GND.n616 GND.n615 4.65
R2032 GND.n613 GND.n612 4.65
R2033 GND.n610 GND.n609 4.65
R2034 GND.n603 GND.n602 4.65
R2035 GND.n600 GND.n599 4.65
R2036 GND.n593 GND.n592 4.65
R2037 GND.n590 GND.n589 4.65
R2038 GND.n587 GND.n586 4.65
R2039 GND.n584 GND.n583 4.65
R2040 GND.n581 GND.n580 4.65
R2041 GND.n578 GND.n577 4.65
R2042 GND.n575 GND.n574 4.65
R2043 GND.n572 GND.n571 4.65
R2044 GND.n569 GND.n568 4.65
R2045 GND.n566 GND.n565 4.65
R2046 GND.n559 GND.n558 4.65
R2047 GND.n556 GND.n555 4.65
R2048 GND.n549 GND.n548 4.65
R2049 GND.n546 GND.n545 4.65
R2050 GND.n543 GND.n542 4.65
R2051 GND.n540 GND.n539 4.65
R2052 GND.n537 GND.n536 4.65
R2053 GND.n534 GND.n533 4.65
R2054 GND.n526 GND.n525 4.65
R2055 GND.n523 GND.n522 4.65
R2056 GND.n516 GND.n515 4.65
R2057 GND.n513 GND.n512 4.65
R2058 GND.n510 GND.n509 4.65
R2059 GND.n507 GND.n506 4.65
R2060 GND.n504 GND.n503 4.65
R2061 GND.n501 GND.n500 4.65
R2062 GND.n493 GND.n492 4.65
R2063 GND.n490 GND.n489 4.65
R2064 GND.n483 GND.n482 4.65
R2065 GND.n480 GND.n479 4.65
R2066 GND.n477 GND.n476 4.65
R2067 GND.n474 GND.n473 4.65
R2068 GND.n471 GND.n470 4.65
R2069 GND.n468 GND.n467 4.65
R2070 GND.n460 GND.n459 4.65
R2071 GND.n457 GND.n456 4.65
R2072 GND.n450 GND.n449 4.65
R2073 GND.n447 GND.n446 4.65
R2074 GND.n444 GND.n443 4.65
R2075 GND.n441 GND.n440 4.65
R2076 GND.n438 GND.n437 4.65
R2077 GND.n435 GND.n434 4.65
R2078 GND.n430 GND.n429 4.65
R2079 GND.n427 GND.n426 4.65
R2080 GND.n420 GND.n419 4.65
R2081 GND.n417 GND.n416 4.65
R2082 GND.n414 GND.n413 4.65
R2083 GND.n411 GND.n410 4.65
R2084 GND.n408 GND.n407 4.65
R2085 GND.n405 GND.n404 4.65
R2086 GND.n397 GND.n396 4.65
R2087 GND.n394 GND.n393 4.65
R2088 GND.n387 GND.n386 4.65
R2089 GND.n384 GND.n383 4.65
R2090 GND.n381 GND.n380 4.65
R2091 GND.n378 GND.n377 4.65
R2092 GND.n375 GND.n374 4.65
R2093 GND.n372 GND.n371 4.65
R2094 GND.n369 GND.n368 4.65
R2095 GND.n366 GND.n365 4.65
R2096 GND.n363 GND.n362 4.65
R2097 GND.n360 GND.n359 4.65
R2098 GND.n352 GND.n351 4.65
R2099 GND.n6 GND.n5 4.65
R2100 GND.n9 GND.n8 4.65
R2101 GND.n12 GND.n11 4.65
R2102 GND.n20 GND.n19 4.65
R2103 GND.n23 GND.n22 4.65
R2104 GND.n26 GND.n25 4.65
R2105 GND.n33 GND.n32 4.65
R2106 GND.n36 GND.n35 4.65
R2107 GND.n39 GND.n38 4.65
R2108 GND.n19 GND.n17 4.129
R2109 GND.n49 GND.n47 4.129
R2110 GND.n81 GND.n79 4.129
R2111 GND.n111 GND.n109 4.129
R2112 GND.n144 GND.n142 4.129
R2113 GND.n174 GND.n172 4.129
R2114 GND.n204 GND.n202 4.129
R2115 GND.n237 GND.n235 4.129
R2116 GND.n312 GND.n310 4.129
R2117 GND.n345 GND.n343 4.129
R2118 GND.n671 GND.n669 4.129
R2119 GND.n641 GND.n639 4.129
R2120 GND.n609 GND.n607 4.129
R2121 GND.n533 GND.n531 4.129
R2122 GND.n500 GND.n498 4.129
R2123 GND.n467 GND.n465 4.129
R2124 GND.n434 GND.n432 4.129
R2125 GND.n404 GND.n402 4.129
R2126 GND.n3 GND.n2 3.408
R2127 GND.n3 GND.n1 2.844
R2128 GND.n6 GND.n3 1.063
R2129 GND.n348 GND.n347 0.474
R2130 GND.n33 GND.n26 0.29
R2131 GND.n63 GND.n56 0.29
R2132 GND.n95 GND.n88 0.29
R2133 GND.n125 GND.n118 0.29
R2134 GND.n158 GND.n151 0.29
R2135 GND.n188 GND.n181 0.29
R2136 GND.n218 GND.n211 0.29
R2137 GND.n251 GND.n244 0.29
R2138 GND.n296 GND.n289 0.29
R2139 GND.n326 GND.n319 0.29
R2140 GND.n694 GND.n687 0.29
R2141 GND.n664 GND.n657 0.29
R2142 GND.n632 GND.n625 0.29
R2143 GND.n600 GND.n593 0.29
R2144 GND.n556 GND.n549 0.29
R2145 GND.n523 GND.n516 0.29
R2146 GND.n490 GND.n483 0.29
R2147 GND.n457 GND.n450 0.29
R2148 GND.n427 GND.n420 0.29
R2149 GND.n394 GND.n387 0.29
R2150 GND.n349 GND 0.207
R2151 GND.n282 GND.n281 0.206
R2152 GND.n565 GND.n564 0.206
R2153 GND.n359 GND.n358 0.206
R2154 GND.n269 GND.n266 0.197
R2155 GND.n578 GND.n575 0.197
R2156 GND.n372 GND.n369 0.197
R2157 GND.n12 GND.n9 0.181
R2158 GND.n45 GND.n42 0.181
R2159 GND.n75 GND.n72 0.181
R2160 GND.n107 GND.n104 0.181
R2161 GND.n137 GND.n134 0.181
R2162 GND.n170 GND.n167 0.181
R2163 GND.n200 GND.n197 0.181
R2164 GND.n230 GND.n227 0.181
R2165 GND.n308 GND.n305 0.181
R2166 GND.n338 GND.n335 0.181
R2167 GND.n678 GND.n675 0.181
R2168 GND.n648 GND.n645 0.181
R2169 GND.n616 GND.n613 0.181
R2170 GND.n540 GND.n537 0.181
R2171 GND.n507 GND.n504 0.181
R2172 GND.n474 GND.n471 0.181
R2173 GND.n441 GND.n438 0.181
R2174 GND.n411 GND.n408 0.181
R2175 GND.n9 GND.n6 0.145
R2176 GND.n20 GND.n12 0.145
R2177 GND.n23 GND.n20 0.145
R2178 GND.n26 GND.n23 0.145
R2179 GND.n36 GND.n33 0.145
R2180 GND.n39 GND.n36 0.145
R2181 GND.n42 GND.n39 0.145
R2182 GND.n50 GND.n45 0.145
R2183 GND.n53 GND.n50 0.145
R2184 GND.n56 GND.n53 0.145
R2185 GND.n66 GND.n63 0.145
R2186 GND.n69 GND.n66 0.145
R2187 GND.n72 GND.n69 0.145
R2188 GND.n82 GND.n75 0.145
R2189 GND.n85 GND.n82 0.145
R2190 GND.n88 GND.n85 0.145
R2191 GND.n98 GND.n95 0.145
R2192 GND.n101 GND.n98 0.145
R2193 GND.n104 GND.n101 0.145
R2194 GND.n112 GND.n107 0.145
R2195 GND.n115 GND.n112 0.145
R2196 GND.n118 GND.n115 0.145
R2197 GND.n128 GND.n125 0.145
R2198 GND.n131 GND.n128 0.145
R2199 GND.n134 GND.n131 0.145
R2200 GND.n145 GND.n137 0.145
R2201 GND.n148 GND.n145 0.145
R2202 GND.n151 GND.n148 0.145
R2203 GND.n161 GND.n158 0.145
R2204 GND.n164 GND.n161 0.145
R2205 GND.n167 GND.n164 0.145
R2206 GND.n175 GND.n170 0.145
R2207 GND.n178 GND.n175 0.145
R2208 GND.n181 GND.n178 0.145
R2209 GND.n191 GND.n188 0.145
R2210 GND.n194 GND.n191 0.145
R2211 GND.n197 GND.n194 0.145
R2212 GND.n205 GND.n200 0.145
R2213 GND.n208 GND.n205 0.145
R2214 GND.n211 GND.n208 0.145
R2215 GND.n221 GND.n218 0.145
R2216 GND.n224 GND.n221 0.145
R2217 GND.n227 GND.n224 0.145
R2218 GND.n238 GND.n230 0.145
R2219 GND.n241 GND.n238 0.145
R2220 GND.n244 GND.n241 0.145
R2221 GND.n254 GND.n251 0.145
R2222 GND.n257 GND.n254 0.145
R2223 GND.n260 GND.n257 0.145
R2224 GND.n263 GND.n260 0.145
R2225 GND.n266 GND.n263 0.145
R2226 GND.n272 GND.n269 0.145
R2227 GND.n275 GND.n272 0.145
R2228 GND.n283 GND.n275 0.145
R2229 GND.n286 GND.n283 0.145
R2230 GND.n289 GND.n286 0.145
R2231 GND.n299 GND.n296 0.145
R2232 GND.n302 GND.n299 0.145
R2233 GND.n305 GND.n302 0.145
R2234 GND.n313 GND.n308 0.145
R2235 GND.n316 GND.n313 0.145
R2236 GND.n319 GND.n316 0.145
R2237 GND.n329 GND.n326 0.145
R2238 GND.n332 GND.n329 0.145
R2239 GND.n335 GND.n332 0.145
R2240 GND.n346 GND.n338 0.145
R2241 GND.n697 GND.n694 0.145
R2242 GND.n687 GND.n684 0.145
R2243 GND.n684 GND.n681 0.145
R2244 GND.n681 GND.n678 0.145
R2245 GND.n675 GND.n672 0.145
R2246 GND.n672 GND.n667 0.145
R2247 GND.n667 GND.n664 0.145
R2248 GND.n657 GND.n654 0.145
R2249 GND.n654 GND.n651 0.145
R2250 GND.n651 GND.n648 0.145
R2251 GND.n645 GND.n642 0.145
R2252 GND.n642 GND.n635 0.145
R2253 GND.n635 GND.n632 0.145
R2254 GND.n625 GND.n622 0.145
R2255 GND.n622 GND.n619 0.145
R2256 GND.n619 GND.n616 0.145
R2257 GND.n613 GND.n610 0.145
R2258 GND.n610 GND.n603 0.145
R2259 GND.n603 GND.n600 0.145
R2260 GND.n593 GND.n590 0.145
R2261 GND.n590 GND.n587 0.145
R2262 GND.n587 GND.n584 0.145
R2263 GND.n584 GND.n581 0.145
R2264 GND.n581 GND.n578 0.145
R2265 GND.n575 GND.n572 0.145
R2266 GND.n572 GND.n569 0.145
R2267 GND.n569 GND.n566 0.145
R2268 GND.n566 GND.n559 0.145
R2269 GND.n559 GND.n556 0.145
R2270 GND.n549 GND.n546 0.145
R2271 GND.n546 GND.n543 0.145
R2272 GND.n543 GND.n540 0.145
R2273 GND.n537 GND.n534 0.145
R2274 GND.n534 GND.n526 0.145
R2275 GND.n526 GND.n523 0.145
R2276 GND.n516 GND.n513 0.145
R2277 GND.n513 GND.n510 0.145
R2278 GND.n510 GND.n507 0.145
R2279 GND.n504 GND.n501 0.145
R2280 GND.n501 GND.n493 0.145
R2281 GND.n493 GND.n490 0.145
R2282 GND.n483 GND.n480 0.145
R2283 GND.n480 GND.n477 0.145
R2284 GND.n477 GND.n474 0.145
R2285 GND.n471 GND.n468 0.145
R2286 GND.n468 GND.n460 0.145
R2287 GND.n460 GND.n457 0.145
R2288 GND.n450 GND.n447 0.145
R2289 GND.n447 GND.n444 0.145
R2290 GND.n444 GND.n441 0.145
R2291 GND.n438 GND.n435 0.145
R2292 GND.n435 GND.n430 0.145
R2293 GND.n430 GND.n427 0.145
R2294 GND.n420 GND.n417 0.145
R2295 GND.n417 GND.n414 0.145
R2296 GND.n414 GND.n411 0.145
R2297 GND.n408 GND.n405 0.145
R2298 GND.n405 GND.n397 0.145
R2299 GND.n397 GND.n394 0.145
R2300 GND.n387 GND.n384 0.145
R2301 GND.n384 GND.n381 0.145
R2302 GND.n381 GND.n378 0.145
R2303 GND.n378 GND.n375 0.145
R2304 GND.n375 GND.n372 0.145
R2305 GND.n369 GND.n366 0.145
R2306 GND.n366 GND.n363 0.145
R2307 GND.n363 GND.n360 0.145
R2308 GND.n360 GND.n352 0.145
R2309 GND.n352 GND.n349 0.145
R2310 GND GND.n697 0.082
R2311 GND GND.n346 0.062
R2312 a_11761_1050.n1 a_11761_1050.t6 480.392
R2313 a_11761_1050.n2 a_11761_1050.t7 440.954
R2314 a_11761_1050.n4 a_11761_1050.n3 410.896
R2315 a_11761_1050.n1 a_11761_1050.t5 403.272
R2316 a_11761_1050.n6 a_11761_1050.n5 157.963
R2317 a_11761_1050.n5 a_11761_1050.n0 91.706
R2318 a_11761_1050.n5 a_11761_1050.n4 76.423
R2319 a_11761_1050.n2 a_11761_1050.n1 20.835
R2320 a_11761_1050.n0 a_11761_1050.t4 14.282
R2321 a_11761_1050.n0 a_11761_1050.t0 14.282
R2322 a_11761_1050.n6 a_11761_1050.t1 14.282
R2323 a_11761_1050.t2 a_11761_1050.n6 14.282
R2324 a_11761_1050.n4 a_11761_1050.n2 8.044
R2325 a_11887_411.n3 a_11887_411.t8 512.525
R2326 a_11887_411.n1 a_11887_411.t13 477.179
R2327 a_11887_411.n6 a_11887_411.t5 472.359
R2328 a_11887_411.n2 a_11887_411.t9 440.954
R2329 a_11887_411.n1 a_11887_411.t7 406.485
R2330 a_11887_411.n6 a_11887_411.t6 384.527
R2331 a_11887_411.n5 a_11887_411.t10 378.636
R2332 a_11887_411.n3 a_11887_411.t12 371.139
R2333 a_11887_411.n7 a_11887_411.t11 342.755
R2334 a_11887_411.n13 a_11887_411.n12 333.44
R2335 a_11887_411.n15 a_11887_411.n14 157.963
R2336 a_11887_411.n7 a_11887_411.n6 154.955
R2337 a_11887_411.n14 a_11887_411.n13 132.141
R2338 a_11887_411.n14 a_11887_411.n0 91.706
R2339 a_11887_411.n4 a_11887_411.n3 77.972
R2340 a_11887_411.n5 a_11887_411.n4 55.891
R2341 a_11887_411.n12 a_11887_411.n11 30
R2342 a_11887_411.n10 a_11887_411.n9 24.383
R2343 a_11887_411.n12 a_11887_411.n10 23.684
R2344 a_11887_411.n2 a_11887_411.n1 21.4
R2345 a_11887_411.n0 a_11887_411.t3 14.282
R2346 a_11887_411.n0 a_11887_411.t4 14.282
R2347 a_11887_411.n15 a_11887_411.t0 14.282
R2348 a_11887_411.t1 a_11887_411.n15 14.282
R2349 a_11887_411.n8 a_11887_411.n7 7.597
R2350 a_11887_411.n4 a_11887_411.n2 6.833
R2351 a_11887_411.n8 a_11887_411.n5 5.693
R2352 a_11887_411.n13 a_11887_411.n8 4.65
R2353 D.n5 D.t4 472.359
R2354 D.n2 D.t1 472.359
R2355 D.n0 D.t0 472.359
R2356 D.n5 D.t7 384.527
R2357 D.n2 D.t5 384.527
R2358 D.n0 D.t2 384.527
R2359 D.n6 D.n5 294.249
R2360 D.n3 D.n2 294.249
R2361 D.n1 D.n0 294.249
R2362 D.n6 D.t3 136.225
R2363 D.n3 D.t8 136.225
R2364 D.n1 D.t6 136.225
R2365 D.n4 D.n1 20.384
R2366 D.n7 D.n4 15.734
R2367 D.n4 D.n3 4.65
R2368 D.n7 D.n6 4.65
R2369 D.n7 D 0.046
R2370 a_9183_989.n1 a_9183_989.t5 480.392
R2371 a_9183_989.n3 a_9183_989.t6 454.685
R2372 a_9183_989.n3 a_9183_989.t10 428.979
R2373 a_9183_989.n1 a_9183_989.t7 403.272
R2374 a_9183_989.n2 a_9183_989.t8 357.204
R2375 a_9183_989.n4 a_9183_989.t9 311.683
R2376 a_9183_989.n10 a_9183_989.n9 305.581
R2377 a_9183_989.n4 a_9183_989.n3 171.288
R2378 a_9183_989.n2 a_9183_989.n1 171.288
R2379 a_9183_989.n11 a_9183_989.n10 159.999
R2380 a_9183_989.n12 a_9183_989.n11 157.963
R2381 a_9183_989.n11 a_9183_989.n0 91.706
R2382 a_9183_989.n9 a_9183_989.n8 30
R2383 a_9183_989.n7 a_9183_989.n6 24.383
R2384 a_9183_989.n9 a_9183_989.n7 23.684
R2385 a_9183_989.n0 a_9183_989.t3 14.282
R2386 a_9183_989.n0 a_9183_989.t2 14.282
R2387 a_9183_989.n12 a_9183_989.t0 14.282
R2388 a_9183_989.t1 a_9183_989.n12 14.282
R2389 a_9183_989.n5 a_9183_989.n4 7.597
R2390 a_9183_989.n5 a_9183_989.n2 5.965
R2391 a_9183_989.n10 a_9183_989.n5 4.65
R2392 a_6137_1050.n4 a_6137_1050.t7 480.392
R2393 a_6137_1050.n4 a_6137_1050.t6 403.272
R2394 a_6137_1050.n5 a_6137_1050.t5 357.204
R2395 a_6137_1050.n8 a_6137_1050.n6 305.581
R2396 a_6137_1050.n5 a_6137_1050.n4 171.288
R2397 a_6137_1050.n6 a_6137_1050.n3 159.999
R2398 a_6137_1050.n3 a_6137_1050.n2 157.964
R2399 a_6137_1050.n3 a_6137_1050.n1 91.706
R2400 a_6137_1050.n8 a_6137_1050.n7 30
R2401 a_6137_1050.n9 a_6137_1050.n0 24.383
R2402 a_6137_1050.n9 a_6137_1050.n8 23.684
R2403 a_6137_1050.n1 a_6137_1050.t4 14.282
R2404 a_6137_1050.n1 a_6137_1050.t1 14.282
R2405 a_6137_1050.n2 a_6137_1050.t3 14.282
R2406 a_6137_1050.n2 a_6137_1050.t2 14.282
R2407 a_6137_1050.n6 a_6137_1050.n5 10.615
R2408 a_6698_101.n11 a_6698_101.n10 68.43
R2409 a_6698_101.n3 a_6698_101.n2 62.817
R2410 a_6698_101.n7 a_6698_101.n6 38.626
R2411 a_6698_101.n6 a_6698_101.n5 35.955
R2412 a_6698_101.n3 a_6698_101.n1 26.202
R2413 a_6698_101.t0 a_6698_101.n3 19.737
R2414 a_6698_101.t1 a_6698_101.n8 8.137
R2415 a_6698_101.t0 a_6698_101.n4 7.273
R2416 a_6698_101.t0 a_6698_101.n0 6.109
R2417 a_6698_101.t1 a_6698_101.n7 4.864
R2418 a_6698_101.t0 a_6698_101.n12 2.074
R2419 a_6698_101.n12 a_6698_101.t1 0.937
R2420 a_6698_101.t1 a_6698_101.n11 0.763
R2421 a_6698_101.n11 a_6698_101.n9 0.185
R2422 a_7595_411.n4 a_7595_411.t6 475.572
R2423 a_7595_411.n8 a_7595_411.t9 472.359
R2424 a_7595_411.n3 a_7595_411.t8 469.145
R2425 a_7595_411.n8 a_7595_411.t13 384.527
R2426 a_7595_411.n4 a_7595_411.t12 384.527
R2427 a_7595_411.n3 a_7595_411.t11 384.527
R2428 a_7595_411.n5 a_7595_411.t10 370.613
R2429 a_7595_411.n9 a_7595_411.n8 266.39
R2430 a_7595_411.n11 a_7595_411.n2 243.576
R2431 a_7595_411.n9 a_7595_411.t7 231.319
R2432 a_7595_411.n7 a_7595_411.t5 231.319
R2433 a_7595_411.n13 a_7595_411.n11 228.526
R2434 a_7595_411.n2 a_7595_411.n1 157.964
R2435 a_7595_411.n7 a_7595_411.n6 139.294
R2436 a_7595_411.n5 a_7595_411.n4 128.028
R2437 a_7595_411.n6 a_7595_411.n3 126.97
R2438 a_7595_411.n2 a_7595_411.n0 91.706
R2439 a_7595_411.n10 a_7595_411.n7 22.288
R2440 a_7595_411.n13 a_7595_411.n12 15.218
R2441 a_7595_411.n0 a_7595_411.t4 14.282
R2442 a_7595_411.n0 a_7595_411.t0 14.282
R2443 a_7595_411.n1 a_7595_411.t2 14.282
R2444 a_7595_411.n1 a_7595_411.t3 14.282
R2445 a_7595_411.n6 a_7595_411.n5 14.151
R2446 a_7595_411.n14 a_7595_411.n13 12.014
R2447 a_7595_411.n10 a_7595_411.n9 7.597
R2448 a_7595_411.n11 a_7595_411.n10 4.65
R2449 a_12988_101.n3 a_12988_101.n2 62.817
R2450 a_12988_101.n11 a_12988_101.n10 46.054
R2451 a_12988_101.n7 a_12988_101.n6 38.626
R2452 a_12988_101.n6 a_12988_101.n5 35.955
R2453 a_12988_101.n12 a_12988_101.n11 27.923
R2454 a_12988_101.n3 a_12988_101.n1 26.202
R2455 a_12988_101.t0 a_12988_101.n3 19.737
R2456 a_12988_101.t0 a_12988_101.n4 7.273
R2457 a_12988_101.n9 a_12988_101.n8 6.883
R2458 a_12988_101.t0 a_12988_101.n0 6.109
R2459 a_12988_101.t1 a_12988_101.n7 4.864
R2460 a_12988_101.t0 a_12988_101.n13 2.074
R2461 a_12988_101.t1 a_12988_101.n9 1.179
R2462 a_12988_101.t1 a_12988_101.n12 0.958
R2463 a_12988_101.n13 a_12988_101.t1 0.937
R2464 a_3072_101.n3 a_3072_101.n1 42.788
R2465 a_3072_101.t0 a_3072_101.n0 8.137
R2466 a_3072_101.n3 a_3072_101.n2 4.665
R2467 a_3072_101.t0 a_3072_101.n3 0.06
R2468 a_4891_989.n0 a_4891_989.t9 480.392
R2469 a_4891_989.n2 a_4891_989.t6 454.685
R2470 a_4891_989.n2 a_4891_989.t8 428.979
R2471 a_4891_989.n0 a_4891_989.t10 403.272
R2472 a_4891_989.n1 a_4891_989.t5 357.204
R2473 a_4891_989.n3 a_4891_989.t7 311.683
R2474 a_4891_989.n9 a_4891_989.n8 305.581
R2475 a_4891_989.n3 a_4891_989.n2 171.288
R2476 a_4891_989.n1 a_4891_989.n0 171.288
R2477 a_4891_989.n11 a_4891_989.n9 159.999
R2478 a_4891_989.n11 a_4891_989.n10 157.964
R2479 a_4891_989.n12 a_4891_989.n11 91.705
R2480 a_4891_989.n8 a_4891_989.n7 30
R2481 a_4891_989.n6 a_4891_989.n5 24.383
R2482 a_4891_989.n8 a_4891_989.n6 23.684
R2483 a_4891_989.n10 a_4891_989.t4 14.282
R2484 a_4891_989.n10 a_4891_989.t0 14.282
R2485 a_4891_989.t2 a_4891_989.n12 14.282
R2486 a_4891_989.n12 a_4891_989.t1 14.282
R2487 a_4891_989.n4 a_4891_989.n3 7.597
R2488 a_4891_989.n4 a_4891_989.n1 5.965
R2489 a_4891_989.n9 a_4891_989.n4 4.65
R2490 a_7469_1050.n0 a_7469_1050.t5 480.392
R2491 a_7469_1050.n0 a_7469_1050.t7 403.272
R2492 a_7469_1050.n1 a_7469_1050.t6 385.063
R2493 a_7469_1050.n6 a_7469_1050.n5 333.44
R2494 a_7469_1050.n8 a_7469_1050.n7 157.964
R2495 a_7469_1050.n1 a_7469_1050.n0 143.429
R2496 a_7469_1050.n8 a_7469_1050.n6 132.141
R2497 a_7469_1050.n9 a_7469_1050.n8 91.705
R2498 a_7469_1050.n5 a_7469_1050.n4 30
R2499 a_7469_1050.n3 a_7469_1050.n2 24.383
R2500 a_7469_1050.n5 a_7469_1050.n3 23.684
R2501 a_7469_1050.n7 a_7469_1050.t4 14.282
R2502 a_7469_1050.n7 a_7469_1050.t3 14.282
R2503 a_7469_1050.t2 a_7469_1050.n9 14.282
R2504 a_7469_1050.n9 a_7469_1050.t1 14.282
R2505 a_7469_1050.n6 a_7469_1050.n1 10.615
R2506 a_6032_101.n3 a_6032_101.n1 42.788
R2507 a_6032_101.t0 a_6032_101.n0 8.137
R2508 a_6032_101.n3 a_6032_101.n2 4.665
R2509 a_6032_101.t0 a_6032_101.n3 0.06
R2510 CLK.n15 CLK.t1 472.359
R2511 CLK.n6 CLK.t2 472.359
R2512 CLK.n0 CLK.t12 472.359
R2513 CLK.n20 CLK.t0 459.505
R2514 CLK.n11 CLK.t5 459.505
R2515 CLK.n2 CLK.t14 459.505
R2516 CLK.n21 CLK.t10 399.181
R2517 CLK.n12 CLK.t13 399.181
R2518 CLK.n3 CLK.t7 399.181
R2519 CLK.n1 CLK.t15 398.558
R2520 CLK.n17 CLK.t11 397.101
R2521 CLK.n8 CLK.t6 397.101
R2522 CLK.n20 CLK.t8 384.527
R2523 CLK.n15 CLK.t9 384.527
R2524 CLK.n11 CLK.t16 384.527
R2525 CLK.n6 CLK.t3 384.527
R2526 CLK.n2 CLK.t17 384.527
R2527 CLK.n0 CLK.t4 384.527
R2528 CLK.n21 CLK.n20 33.832
R2529 CLK.n3 CLK.n2 33.832
R2530 CLK.n12 CLK.n11 33.832
R2531 CLK.n1 CLK.n0 32.394
R2532 CLK.n16 CLK.n15 30.822
R2533 CLK.n7 CLK.n6 30.822
R2534 CLK.n4 CLK.n1 9.575
R2535 CLK.n13 CLK.n10 8.078
R2536 CLK.n22 CLK.n19 8.078
R2537 CLK.n14 CLK.n13 7.797
R2538 CLK.n5 CLK.n4 7.564
R2539 CLK.n17 CLK.n16 4.577
R2540 CLK.n8 CLK.n7 4.577
R2541 CLK.n9 CLK.n8 4.282
R2542 CLK.n18 CLK.n17 4.282
R2543 CLK.n4 CLK.n3 2.079
R2544 CLK.n13 CLK.n12 2.079
R2545 CLK.n22 CLK.n21 2.079
R2546 CLK.n22 CLK 0.046
R2547 CLK.n10 CLK.n9 0.038
R2548 CLK.n19 CLK.n18 0.038
R2549 CLK.n9 CLK.n5 0.008
R2550 CLK.n18 CLK.n14 0.008
R2551 a_14320_101.n3 a_14320_101.n1 42.788
R2552 a_14320_101.t0 a_14320_101.n0 8.137
R2553 a_14320_101.n3 a_14320_101.n2 4.665
R2554 a_14320_101.t0 a_14320_101.n3 0.06
R2555 a_13757_1051.n4 a_13757_1051.t7 179.895
R2556 a_13757_1051.n2 a_13757_1051.n1 165.613
R2557 a_13757_1051.n2 a_13757_1051.n0 142.653
R2558 a_13757_1051.n4 a_13757_1051.n3 106.183
R2559 a_13757_1051.n5 a_13757_1051.n4 99.358
R2560 a_13757_1051.n3 a_13757_1051.n2 82.665
R2561 a_13757_1051.n3 a_13757_1051.t2 73.712
R2562 a_13757_1051.n0 a_13757_1051.t5 14.282
R2563 a_13757_1051.n0 a_13757_1051.t4 14.282
R2564 a_13757_1051.n1 a_13757_1051.t0 14.282
R2565 a_13757_1051.n1 a_13757_1051.t1 14.282
R2566 a_13757_1051.n5 a_13757_1051.t6 14.282
R2567 a_13757_1051.t3 a_13757_1051.n5 14.282
R2568 a_7364_101.n11 a_7364_101.n10 68.43
R2569 a_7364_101.n3 a_7364_101.n2 62.817
R2570 a_7364_101.n7 a_7364_101.n6 38.626
R2571 a_7364_101.n6 a_7364_101.n5 35.955
R2572 a_7364_101.n3 a_7364_101.n1 26.202
R2573 a_7364_101.t0 a_7364_101.n3 19.737
R2574 a_7364_101.t1 a_7364_101.n8 8.137
R2575 a_7364_101.t0 a_7364_101.n4 7.273
R2576 a_7364_101.t0 a_7364_101.n0 6.109
R2577 a_7364_101.t1 a_7364_101.n7 4.864
R2578 a_7364_101.t0 a_7364_101.n12 2.074
R2579 a_7364_101.n12 a_7364_101.t1 0.937
R2580 a_7364_101.t1 a_7364_101.n11 0.763
R2581 a_7364_101.n11 a_7364_101.n9 0.185
R2582 a_3738_101.n11 a_3738_101.n10 68.43
R2583 a_3738_101.n3 a_3738_101.n2 62.817
R2584 a_3738_101.n7 a_3738_101.n6 38.626
R2585 a_3738_101.n6 a_3738_101.n5 35.955
R2586 a_3738_101.n3 a_3738_101.n1 26.202
R2587 a_3738_101.t0 a_3738_101.n3 19.737
R2588 a_3738_101.t1 a_3738_101.n8 8.137
R2589 a_3738_101.t0 a_3738_101.n4 7.273
R2590 a_3738_101.t0 a_3738_101.n0 6.109
R2591 a_3738_101.t1 a_3738_101.n7 4.864
R2592 a_3738_101.t0 a_3738_101.n12 2.074
R2593 a_3738_101.n12 a_3738_101.t1 0.937
R2594 a_3738_101.t1 a_3738_101.n11 0.763
R2595 a_3738_101.n11 a_3738_101.n9 0.185
R2596 a_10324_101.n5 a_10324_101.n4 62.817
R2597 a_10324_101.n2 a_10324_101.n0 41.528
R2598 a_10324_101.n5 a_10324_101.n3 26.202
R2599 a_10324_101.t0 a_10324_101.n5 19.737
R2600 a_10324_101.t0 a_10324_101.n6 8.137
R2601 a_10324_101.n2 a_10324_101.n1 3.644
R2602 a_10324_101.t0 a_10324_101.n2 1.093
R2603 a_10429_1050.n1 a_10429_1050.t7 480.392
R2604 a_10429_1050.n1 a_10429_1050.t5 403.272
R2605 a_10429_1050.n2 a_10429_1050.t6 357.204
R2606 a_10429_1050.n4 a_10429_1050.n3 327.32
R2607 a_10429_1050.n2 a_10429_1050.n1 171.288
R2608 a_10429_1050.n5 a_10429_1050.n4 159.999
R2609 a_10429_1050.n6 a_10429_1050.n5 157.963
R2610 a_10429_1050.n5 a_10429_1050.n0 91.706
R2611 a_10429_1050.n0 a_10429_1050.t3 14.282
R2612 a_10429_1050.n0 a_10429_1050.t2 14.282
R2613 a_10429_1050.t1 a_10429_1050.n6 14.282
R2614 a_10429_1050.n6 a_10429_1050.t0 14.282
R2615 a_10429_1050.n4 a_10429_1050.n2 10.615
R2616 a_4439_187.n5 a_4439_187.t5 512.525
R2617 a_4439_187.n3 a_4439_187.t12 472.359
R2618 a_4439_187.n1 a_4439_187.t13 472.359
R2619 a_4439_187.n6 a_4439_187.t8 417.109
R2620 a_4439_187.n3 a_4439_187.t6 384.527
R2621 a_4439_187.n1 a_4439_187.t10 384.527
R2622 a_4439_187.n10 a_4439_187.n9 383.037
R2623 a_4439_187.n5 a_4439_187.t11 371.139
R2624 a_4439_187.n4 a_4439_187.t7 370.613
R2625 a_4439_187.n2 a_4439_187.t9 370.613
R2626 a_4439_187.n6 a_4439_187.n5 179.837
R2627 a_4439_187.n12 a_4439_187.n11 157.963
R2628 a_4439_187.n4 a_4439_187.n3 127.096
R2629 a_4439_187.n2 a_4439_187.n1 127.096
R2630 a_4439_187.n11 a_4439_187.n10 104.282
R2631 a_4439_187.n11 a_4439_187.n0 91.706
R2632 a_4439_187.n0 a_4439_187.t4 14.282
R2633 a_4439_187.n0 a_4439_187.t3 14.282
R2634 a_4439_187.n12 a_4439_187.t0 14.282
R2635 a_4439_187.t1 a_4439_187.n12 14.282
R2636 a_4439_187.n7 a_4439_187.n6 11.134
R2637 a_4439_187.n8 a_4439_187.n2 8.957
R2638 a_4439_187.n7 a_4439_187.n4 4.65
R2639 a_4439_187.n10 a_4439_187.n8 4.65
R2640 a_4439_187.n8 a_4439_187.n7 2.947
R2641 a_8675_103.t0 a_8675_103.n7 59.616
R2642 a_8675_103.n4 a_8675_103.n2 54.496
R2643 a_8675_103.n4 a_8675_103.n3 54.496
R2644 a_8675_103.n1 a_8675_103.n0 24.679
R2645 a_8675_103.n6 a_8675_103.n4 7.859
R2646 a_8675_103.t0 a_8675_103.n1 7.505
R2647 a_8675_103.t0 a_8675_103.n6 3.034
R2648 a_8675_103.n6 a_8675_103.n5 0.443
R2649 a_599_989.n0 a_599_989.t7 480.392
R2650 a_599_989.n2 a_599_989.t9 454.685
R2651 a_599_989.n2 a_599_989.t5 428.979
R2652 a_599_989.n0 a_599_989.t10 403.272
R2653 a_599_989.n1 a_599_989.t8 357.204
R2654 a_599_989.n3 a_599_989.t6 311.683
R2655 a_599_989.n9 a_599_989.n8 305.581
R2656 a_599_989.n3 a_599_989.n2 171.288
R2657 a_599_989.n1 a_599_989.n0 171.288
R2658 a_599_989.n11 a_599_989.n9 159.999
R2659 a_599_989.n11 a_599_989.n10 157.964
R2660 a_599_989.n12 a_599_989.n11 91.705
R2661 a_599_989.n8 a_599_989.n7 30
R2662 a_599_989.n6 a_599_989.n5 24.383
R2663 a_599_989.n8 a_599_989.n6 23.684
R2664 a_599_989.n10 a_599_989.t4 14.282
R2665 a_599_989.n10 a_599_989.t3 14.282
R2666 a_599_989.t2 a_599_989.n12 14.282
R2667 a_599_989.n12 a_599_989.t1 14.282
R2668 a_599_989.n4 a_599_989.n3 7.597
R2669 a_599_989.n4 a_599_989.n1 5.965
R2670 a_599_989.n9 a_599_989.n4 4.65
R2671 a_8030_101.n11 a_8030_101.n10 68.43
R2672 a_8030_101.n3 a_8030_101.n2 62.817
R2673 a_8030_101.n7 a_8030_101.n6 38.626
R2674 a_8030_101.n6 a_8030_101.n5 35.955
R2675 a_8030_101.n3 a_8030_101.n1 26.202
R2676 a_8030_101.t0 a_8030_101.n3 19.737
R2677 a_8030_101.t1 a_8030_101.n8 8.137
R2678 a_8030_101.t0 a_8030_101.n4 7.273
R2679 a_8030_101.t0 a_8030_101.n0 6.109
R2680 a_8030_101.t1 a_8030_101.n7 4.864
R2681 a_8030_101.t0 a_8030_101.n12 2.074
R2682 a_8030_101.n12 a_8030_101.t1 0.937
R2683 a_8030_101.t1 a_8030_101.n11 0.763
R2684 a_8030_101.n11 a_8030_101.n9 0.185
R2685 a_1074_101.n3 a_1074_101.n1 42.788
R2686 a_1074_101.t0 a_1074_101.n0 8.137
R2687 a_1074_101.n3 a_1074_101.n2 4.665
R2688 a_1074_101.t0 a_1074_101.n3 0.06
R2689 a_4569_1050.n3 a_4569_1050.t12 480.392
R2690 a_4569_1050.n1 a_4569_1050.t7 480.392
R2691 a_4569_1050.n3 a_4569_1050.t9 403.272
R2692 a_4569_1050.n1 a_4569_1050.t10 403.272
R2693 a_4569_1050.n4 a_4569_1050.t8 385.063
R2694 a_4569_1050.n2 a_4569_1050.t11 385.063
R2695 a_4569_1050.n10 a_4569_1050.n9 336.075
R2696 a_4569_1050.n13 a_4569_1050.n12 161.352
R2697 a_4569_1050.n11 a_4569_1050.n10 151.34
R2698 a_4569_1050.n4 a_4569_1050.n3 143.429
R2699 a_4569_1050.n2 a_4569_1050.n1 143.429
R2700 a_4569_1050.n11 a_4569_1050.n0 95.095
R2701 a_4569_1050.n14 a_4569_1050.n13 95.094
R2702 a_4569_1050.n13 a_4569_1050.n11 66.258
R2703 a_4569_1050.n9 a_4569_1050.n8 30
R2704 a_4569_1050.n7 a_4569_1050.n6 24.383
R2705 a_4569_1050.n9 a_4569_1050.n7 23.684
R2706 a_4569_1050.n0 a_4569_1050.t2 14.282
R2707 a_4569_1050.n0 a_4569_1050.t3 14.282
R2708 a_4569_1050.n12 a_4569_1050.t6 14.282
R2709 a_4569_1050.n12 a_4569_1050.t5 14.282
R2710 a_4569_1050.t1 a_4569_1050.n14 14.282
R2711 a_4569_1050.n14 a_4569_1050.t0 14.282
R2712 a_4569_1050.n5 a_4569_1050.n2 11.95
R2713 a_4569_1050.n10 a_4569_1050.n5 5.965
R2714 a_4569_1050.n5 a_4569_1050.n4 4.65
R2715 a_12322_101.n11 a_12322_101.n10 68.43
R2716 a_12322_101.n3 a_12322_101.n2 62.817
R2717 a_12322_101.n7 a_12322_101.n6 38.626
R2718 a_12322_101.n6 a_12322_101.n5 35.955
R2719 a_12322_101.n3 a_12322_101.n1 26.202
R2720 a_12322_101.t0 a_12322_101.n3 19.737
R2721 a_12322_101.t1 a_12322_101.n8 8.137
R2722 a_12322_101.t0 a_12322_101.n4 7.273
R2723 a_12322_101.t0 a_12322_101.n0 6.109
R2724 a_12322_101.t1 a_12322_101.n7 4.864
R2725 a_12322_101.t0 a_12322_101.n12 2.074
R2726 a_12322_101.n12 a_12322_101.t1 0.937
R2727 a_12322_101.t1 a_12322_101.n11 0.763
R2728 a_12322_101.n11 a_12322_101.n9 0.185
R2729 a_2406_101.n11 a_2406_101.n10 68.43
R2730 a_2406_101.n3 a_2406_101.n2 62.817
R2731 a_2406_101.n7 a_2406_101.n6 38.626
R2732 a_2406_101.n6 a_2406_101.n5 35.955
R2733 a_2406_101.n3 a_2406_101.n1 26.202
R2734 a_2406_101.t0 a_2406_101.n3 19.737
R2735 a_2406_101.t1 a_2406_101.n8 8.137
R2736 a_2406_101.t0 a_2406_101.n4 7.273
R2737 a_2406_101.t0 a_2406_101.n0 6.109
R2738 a_2406_101.t1 a_2406_101.n7 4.864
R2739 a_2406_101.t0 a_2406_101.n12 2.074
R2740 a_2406_101.n12 a_2406_101.t1 0.937
R2741 a_2406_101.t1 a_2406_101.n11 0.763
R2742 a_2406_101.n11 a_2406_101.n9 0.185
R2743 a_372_210.n10 a_372_210.n8 171.558
R2744 a_372_210.n8 a_372_210.t1 75.764
R2745 a_372_210.n3 a_372_210.n2 27.476
R2746 a_372_210.n10 a_372_210.n9 27.2
R2747 a_372_210.n11 a_372_210.n0 23.498
R2748 a_372_210.n11 a_372_210.n10 22.4
R2749 a_372_210.t1 a_372_210.n5 20.241
R2750 a_372_210.n7 a_372_210.n6 19.952
R2751 a_372_210.t1 a_372_210.n3 13.984
R2752 a_372_210.n5 a_372_210.n4 13.494
R2753 a_372_210.t1 a_372_210.n1 7.04
R2754 a_372_210.n8 a_372_210.n7 1.505
R2755 a_9658_101.n11 a_9658_101.n10 68.43
R2756 a_9658_101.n3 a_9658_101.n2 62.817
R2757 a_9658_101.n7 a_9658_101.n6 38.626
R2758 a_9658_101.n6 a_9658_101.n5 35.955
R2759 a_9658_101.n3 a_9658_101.n1 26.202
R2760 a_9658_101.t0 a_9658_101.n3 19.737
R2761 a_9658_101.t1 a_9658_101.n8 8.137
R2762 a_9658_101.t0 a_9658_101.n4 7.273
R2763 a_9658_101.t0 a_9658_101.n0 6.109
R2764 a_9658_101.t1 a_9658_101.n7 4.864
R2765 a_9658_101.t0 a_9658_101.n12 2.074
R2766 a_9658_101.n12 a_9658_101.t1 0.937
R2767 a_9658_101.t1 a_9658_101.n11 0.763
R2768 a_9658_101.n11 a_9658_101.n9 0.185
R2769 a_13093_1051.n2 a_13093_1051.t5 179.895
R2770 a_13093_1051.n5 a_13093_1051.n4 157.021
R2771 a_13093_1051.n4 a_13093_1051.n0 124.955
R2772 a_13093_1051.n3 a_13093_1051.n2 106.183
R2773 a_13093_1051.n2 a_13093_1051.n1 99.355
R2774 a_13093_1051.n4 a_13093_1051.n3 82.65
R2775 a_13093_1051.n3 a_13093_1051.t3 73.712
R2776 a_13093_1051.n0 a_13093_1051.t7 14.282
R2777 a_13093_1051.n0 a_13093_1051.t6 14.282
R2778 a_13093_1051.n1 a_13093_1051.t4 14.282
R2779 a_13093_1051.n1 a_13093_1051.t2 14.282
R2780 a_13093_1051.t1 a_13093_1051.n5 14.282
R2781 a_13093_1051.n5 a_13093_1051.t0 14.282
R2782 a_4664_210.n10 a_4664_210.n8 171.558
R2783 a_4664_210.n8 a_4664_210.t1 75.764
R2784 a_4664_210.n3 a_4664_210.n2 27.476
R2785 a_4664_210.n10 a_4664_210.n9 27.2
R2786 a_4664_210.n11 a_4664_210.n0 23.498
R2787 a_4664_210.n11 a_4664_210.n10 22.4
R2788 a_4664_210.t1 a_4664_210.n5 20.241
R2789 a_4664_210.n7 a_4664_210.n6 19.952
R2790 a_4664_210.t1 a_4664_210.n3 13.984
R2791 a_4664_210.n5 a_4664_210.n4 13.494
R2792 a_4664_210.t1 a_4664_210.n1 7.04
R2793 a_4664_210.n8 a_4664_210.n7 1.505
R2794 a_8956_210.n8 a_8956_210.n6 185.173
R2795 a_8956_210.t0 a_8956_210.n8 75.765
R2796 a_8956_210.n3 a_8956_210.n1 74.827
R2797 a_8956_210.n3 a_8956_210.n2 27.476
R2798 a_8956_210.n6 a_8956_210.n5 22.349
R2799 a_8956_210.t0 a_8956_210.n10 20.241
R2800 a_8956_210.t0 a_8956_210.n3 13.984
R2801 a_8956_210.n10 a_8956_210.n9 13.494
R2802 a_8956_210.n6 a_8956_210.n4 8.443
R2803 a_8956_210.t0 a_8956_210.n0 8.137
R2804 a_8956_210.n8 a_8956_210.n7 1.505
R2805 a_91_103.n5 a_91_103.n4 66.708
R2806 a_91_103.n2 a_91_103.n0 25.439
R2807 a_91_103.n5 a_91_103.n3 19.496
R2808 a_91_103.t0 a_91_103.n5 13.756
R2809 a_91_103.n2 a_91_103.n1 2.455
R2810 a_91_103.t0 a_91_103.n2 0.246
R2811 a_11656_101.n3 a_11656_101.n1 42.788
R2812 a_11656_101.t0 a_11656_101.n0 8.137
R2813 a_11656_101.n3 a_11656_101.n2 4.665
R2814 a_11656_101.t0 a_11656_101.n3 0.06
R2815 a_10990_101.n3 a_10990_101.n1 42.788
R2816 a_10990_101.t0 a_10990_101.n0 8.137
R2817 a_10990_101.n3 a_10990_101.n2 4.665
R2818 a_10990_101.t0 a_10990_101.n3 0.06
R2819 a_4383_103.t0 a_4383_103.n7 59.616
R2820 a_4383_103.n4 a_4383_103.n2 54.496
R2821 a_4383_103.n4 a_4383_103.n3 54.496
R2822 a_4383_103.n1 a_4383_103.n0 24.679
R2823 a_4383_103.t0 a_4383_103.n1 7.505
R2824 a_4383_103.n6 a_4383_103.n5 2.455
R2825 a_4383_103.n6 a_4383_103.n4 0.636
R2826 a_4383_103.t0 a_4383_103.n6 0.246
R2827 a_1740_101.n3 a_1740_101.n1 42.788
R2828 a_1740_101.t0 a_1740_101.n0 8.137
R2829 a_1740_101.n3 a_1740_101.n2 4.665
R2830 a_1740_101.t0 a_1740_101.n3 0.06
R2831 a_5366_101.n3 a_5366_101.n1 42.788
R2832 a_5366_101.t0 a_5366_101.n0 8.137
R2833 a_5366_101.n3 a_5366_101.n2 4.665
R2834 a_5366_101.t0 a_5366_101.n3 0.06
C4 VDD GND 23.90fF
C5 a_5366_101.n0 GND 0.05fF
C6 a_5366_101.n1 GND 0.12fF
C7 a_5366_101.n2 GND 0.04fF
C8 a_5366_101.n3 GND 0.17fF
C9 a_1740_101.n0 GND 0.05fF
C10 a_1740_101.n1 GND 0.12fF
C11 a_1740_101.n2 GND 0.04fF
C12 a_1740_101.n3 GND 0.17fF
C13 a_4383_103.n0 GND 0.08fF
C14 a_4383_103.n1 GND 0.07fF
C15 a_4383_103.n2 GND 0.04fF
C16 a_4383_103.n3 GND 0.06fF
C17 a_4383_103.n4 GND 0.03fF
C18 a_4383_103.n5 GND 0.04fF
C19 a_4383_103.n7 GND 0.08fF
C20 a_10990_101.n0 GND 0.05fF
C21 a_10990_101.n1 GND 0.12fF
C22 a_10990_101.n2 GND 0.04fF
C23 a_10990_101.n3 GND 0.17fF
C24 a_11656_101.n0 GND 0.05fF
C25 a_11656_101.n1 GND 0.12fF
C26 a_11656_101.n2 GND 0.04fF
C27 a_11656_101.n3 GND 0.17fF
C28 a_91_103.n0 GND 0.10fF
C29 a_91_103.n1 GND 0.03fF
C30 a_91_103.n2 GND 0.03fF
C31 a_91_103.n3 GND 0.07fF
C32 a_91_103.n4 GND 0.08fF
C33 a_91_103.n5 GND 0.03fF
C34 a_8956_210.n0 GND 0.07fF
C35 a_8956_210.n1 GND 0.09fF
C36 a_8956_210.n2 GND 0.12fF
C37 a_8956_210.n3 GND 0.08fF
C38 a_8956_210.n4 GND 0.02fF
C39 a_8956_210.n5 GND 0.03fF
C40 a_8956_210.n6 GND 0.05fF
C41 a_8956_210.n7 GND 0.02fF
C42 a_8956_210.n8 GND 0.14fF
C43 a_8956_210.n9 GND 0.08fF
C44 a_8956_210.n10 GND 0.02fF
C45 a_8956_210.t0 GND 0.31fF
C46 a_4664_210.n0 GND 0.02fF
C47 a_4664_210.n1 GND 0.09fF
C48 a_4664_210.n2 GND 0.12fF
C49 a_4664_210.n3 GND 0.08fF
C50 a_4664_210.n4 GND 0.08fF
C51 a_4664_210.n5 GND 0.02fF
C52 a_4664_210.t1 GND 0.29fF
C53 a_4664_210.n6 GND 0.09fF
C54 a_4664_210.n7 GND 0.02fF
C55 a_4664_210.n8 GND 0.13fF
C56 a_4664_210.n9 GND 0.02fF
C57 a_4664_210.n10 GND 0.03fF
C58 a_4664_210.n11 GND 0.03fF
C59 a_13093_1051.n0 GND 0.36fF
C60 a_13093_1051.n1 GND 0.32fF
C61 a_13093_1051.n2 GND 0.53fF
C62 a_13093_1051.n3 GND 0.30fF
C63 a_13093_1051.n4 GND 0.81fF
C64 a_13093_1051.n5 GND 0.43fF
C65 a_9658_101.n0 GND 0.02fF
C66 a_9658_101.n1 GND 0.09fF
C67 a_9658_101.n2 GND 0.08fF
C68 a_9658_101.n3 GND 0.03fF
C69 a_9658_101.n4 GND 0.01fF
C70 a_9658_101.n5 GND 0.04fF
C71 a_9658_101.n6 GND 0.04fF
C72 a_9658_101.n7 GND 0.02fF
C73 a_9658_101.n8 GND 0.05fF
C74 a_9658_101.n9 GND 0.15fF
C75 a_9658_101.n10 GND 0.08fF
C76 a_9658_101.n11 GND 0.08fF
C77 a_9658_101.t1 GND 0.23fF
C78 a_9658_101.n12 GND 0.01fF
C79 a_372_210.n0 GND 0.02fF
C80 a_372_210.n1 GND 0.09fF
C81 a_372_210.n2 GND 0.12fF
C82 a_372_210.n3 GND 0.08fF
C83 a_372_210.n4 GND 0.08fF
C84 a_372_210.n5 GND 0.02fF
C85 a_372_210.t1 GND 0.29fF
C86 a_372_210.n6 GND 0.09fF
C87 a_372_210.n7 GND 0.02fF
C88 a_372_210.n8 GND 0.13fF
C89 a_372_210.n9 GND 0.02fF
C90 a_372_210.n10 GND 0.03fF
C91 a_372_210.n11 GND 0.03fF
C92 a_2406_101.n0 GND 0.02fF
C93 a_2406_101.n1 GND 0.09fF
C94 a_2406_101.n2 GND 0.08fF
C95 a_2406_101.n3 GND 0.03fF
C96 a_2406_101.n4 GND 0.01fF
C97 a_2406_101.n5 GND 0.04fF
C98 a_2406_101.n6 GND 0.04fF
C99 a_2406_101.n7 GND 0.02fF
C100 a_2406_101.n8 GND 0.05fF
C101 a_2406_101.n9 GND 0.15fF
C102 a_2406_101.n10 GND 0.08fF
C103 a_2406_101.n11 GND 0.08fF
C104 a_2406_101.t1 GND 0.23fF
C105 a_2406_101.n12 GND 0.01fF
C106 a_12322_101.n0 GND 0.02fF
C107 a_12322_101.n1 GND 0.09fF
C108 a_12322_101.n2 GND 0.08fF
C109 a_12322_101.n3 GND 0.03fF
C110 a_12322_101.n4 GND 0.01fF
C111 a_12322_101.n5 GND 0.04fF
C112 a_12322_101.n6 GND 0.04fF
C113 a_12322_101.n7 GND 0.02fF
C114 a_12322_101.n8 GND 0.05fF
C115 a_12322_101.n9 GND 0.15fF
C116 a_12322_101.n10 GND 0.08fF
C117 a_12322_101.n11 GND 0.08fF
C118 a_12322_101.t1 GND 0.23fF
C119 a_12322_101.n12 GND 0.01fF
C120 a_4569_1050.n0 GND 0.57fF
C121 a_4569_1050.n1 GND 0.44fF
C122 a_4569_1050.n2 GND 1.38fF
C123 a_4569_1050.n3 GND 0.44fF
C124 a_4569_1050.n4 GND 0.63fF
C125 a_4569_1050.n5 GND 2.09fF
C126 a_4569_1050.n6 GND 0.06fF
C127 a_4569_1050.n7 GND 0.08fF
C128 a_4569_1050.n8 GND 0.05fF
C129 a_4569_1050.n9 GND 0.37fF
C130 a_4569_1050.n10 GND 0.82fF
C131 a_4569_1050.n11 GND 0.61fF
C132 a_4569_1050.n12 GND 0.72fF
C133 a_4569_1050.n13 GND 0.69fF
C134 a_4569_1050.n14 GND 0.57fF
C135 a_1074_101.n0 GND 0.05fF
C136 a_1074_101.n1 GND 0.12fF
C137 a_1074_101.n2 GND 0.04fF
C138 a_1074_101.n3 GND 0.17fF
C139 a_8030_101.n0 GND 0.02fF
C140 a_8030_101.n1 GND 0.09fF
C141 a_8030_101.n2 GND 0.08fF
C142 a_8030_101.n3 GND 0.03fF
C143 a_8030_101.n4 GND 0.01fF
C144 a_8030_101.n5 GND 0.04fF
C145 a_8030_101.n6 GND 0.04fF
C146 a_8030_101.n7 GND 0.02fF
C147 a_8030_101.n8 GND 0.05fF
C148 a_8030_101.n9 GND 0.15fF
C149 a_8030_101.n10 GND 0.08fF
C150 a_8030_101.n11 GND 0.08fF
C151 a_8030_101.t1 GND 0.23fF
C152 a_8030_101.n12 GND 0.01fF
C153 a_599_989.n0 GND 0.34fF
C154 a_599_989.n1 GND 0.49fF
C155 a_599_989.n2 GND 0.34fF
C156 a_599_989.t6 GND 0.55fF
C157 a_599_989.n3 GND 0.57fF
C158 a_599_989.n4 GND 0.89fF
C159 a_599_989.n5 GND 0.04fF
C160 a_599_989.n6 GND 0.06fF
C161 a_599_989.n7 GND 0.04fF
C162 a_599_989.n8 GND 0.23fF
C163 a_599_989.n9 GND 0.52fF
C164 a_599_989.n10 GND 0.52fF
C165 a_599_989.n11 GND 0.60fF
C166 a_599_989.n12 GND 0.40fF
C167 a_8675_103.n0 GND 0.08fF
C168 a_8675_103.n1 GND 0.07fF
C169 a_8675_103.n2 GND 0.04fF
C170 a_8675_103.n3 GND 0.06fF
C171 a_8675_103.n4 GND 0.11fF
C172 a_8675_103.n5 GND 0.04fF
C173 a_8675_103.n7 GND 0.08fF
C174 a_4439_187.n0 GND 0.65fF
C175 a_4439_187.n1 GND 0.47fF
C176 a_4439_187.t9 GND 0.98fF
C177 a_4439_187.n2 GND 1.08fF
C178 a_4439_187.n3 GND 0.47fF
C179 a_4439_187.t7 GND 0.98fF
C180 a_4439_187.n4 GND 0.66fF
C181 a_4439_187.n5 GND 0.48fF
C182 a_4439_187.n6 GND 1.55fF
C183 a_4439_187.n7 GND 2.34fF
C184 a_4439_187.n8 GND 1.85fF
C185 a_4439_187.n9 GND 0.67fF
C186 a_4439_187.n10 GND 0.88fF
C187 a_4439_187.n11 GND 0.88fF
C188 a_4439_187.n12 GND 0.84fF
C189 a_10429_1050.n0 GND 0.42fF
C190 a_10429_1050.n1 GND 0.36fF
C191 a_10429_1050.n2 GND 0.67fF
C192 a_10429_1050.n3 GND 0.37fF
C193 a_10429_1050.n4 GND 0.76fF
C194 a_10429_1050.n5 GND 0.64fF
C195 a_10429_1050.n6 GND 0.54fF
C196 a_10324_101.n0 GND 0.08fF
C197 a_10324_101.n1 GND 0.02fF
C198 a_10324_101.n2 GND 0.02fF
C199 a_10324_101.n3 GND 0.09fF
C200 a_10324_101.n4 GND 0.08fF
C201 a_10324_101.n5 GND 0.03fF
C202 a_10324_101.n6 GND 0.05fF
C203 a_3738_101.n0 GND 0.02fF
C204 a_3738_101.n1 GND 0.09fF
C205 a_3738_101.n2 GND 0.08fF
C206 a_3738_101.n3 GND 0.03fF
C207 a_3738_101.n4 GND 0.01fF
C208 a_3738_101.n5 GND 0.04fF
C209 a_3738_101.n6 GND 0.04fF
C210 a_3738_101.n7 GND 0.02fF
C211 a_3738_101.n8 GND 0.05fF
C212 a_3738_101.n9 GND 0.15fF
C213 a_3738_101.n10 GND 0.08fF
C214 a_3738_101.n11 GND 0.08fF
C215 a_3738_101.t1 GND 0.23fF
C216 a_3738_101.n12 GND 0.01fF
C217 a_7364_101.n0 GND 0.02fF
C218 a_7364_101.n1 GND 0.09fF
C219 a_7364_101.n2 GND 0.08fF
C220 a_7364_101.n3 GND 0.03fF
C221 a_7364_101.n4 GND 0.01fF
C222 a_7364_101.n5 GND 0.04fF
C223 a_7364_101.n6 GND 0.04fF
C224 a_7364_101.n7 GND 0.02fF
C225 a_7364_101.n8 GND 0.05fF
C226 a_7364_101.n9 GND 0.15fF
C227 a_7364_101.n10 GND 0.08fF
C228 a_7364_101.n11 GND 0.08fF
C229 a_7364_101.t1 GND 0.23fF
C230 a_7364_101.n12 GND 0.01fF
C231 a_13757_1051.n0 GND 0.28fF
C232 a_13757_1051.n1 GND 0.36fF
C233 a_13757_1051.n2 GND 0.70fF
C234 a_13757_1051.n3 GND 0.27fF
C235 a_13757_1051.n4 GND 0.45fF
C236 a_13757_1051.n5 GND 0.28fF
C237 a_14320_101.n0 GND 0.05fF
C238 a_14320_101.n1 GND 0.13fF
C239 a_14320_101.n2 GND 0.04fF
C240 a_14320_101.n3 GND 0.18fF
C241 a_6032_101.n0 GND 0.05fF
C242 a_6032_101.n1 GND 0.12fF
C243 a_6032_101.n2 GND 0.04fF
C244 a_6032_101.n3 GND 0.17fF
C245 a_7469_1050.n0 GND 0.31fF
C246 a_7469_1050.n1 GND 0.63fF
C247 a_7469_1050.n2 GND 0.04fF
C248 a_7469_1050.n3 GND 0.06fF
C249 a_7469_1050.n4 GND 0.04fF
C250 a_7469_1050.n5 GND 0.26fF
C251 a_7469_1050.n6 GND 0.69fF
C252 a_7469_1050.n7 GND 0.51fF
C253 a_7469_1050.n8 GND 0.56fF
C254 a_7469_1050.n9 GND 0.40fF
C255 a_4891_989.n0 GND 0.42fF
C256 a_4891_989.n1 GND 0.60fF
C257 a_4891_989.n2 GND 0.42fF
C258 a_4891_989.t7 GND 0.67fF
C259 a_4891_989.n3 GND 0.70fF
C260 a_4891_989.n4 GND 1.09fF
C261 a_4891_989.n5 GND 0.05fF
C262 a_4891_989.n6 GND 0.07fF
C263 a_4891_989.n7 GND 0.04fF
C264 a_4891_989.n8 GND 0.29fF
C265 a_4891_989.n9 GND 0.63fF
C266 a_4891_989.n10 GND 0.63fF
C267 a_4891_989.n11 GND 0.74fF
C268 a_4891_989.n12 GND 0.49fF
C269 a_3072_101.n0 GND 0.05fF
C270 a_3072_101.n1 GND 0.12fF
C271 a_3072_101.n2 GND 0.04fF
C272 a_3072_101.n3 GND 0.17fF
C273 a_12988_101.n0 GND 0.02fF
C274 a_12988_101.n1 GND 0.09fF
C275 a_12988_101.n2 GND 0.07fF
C276 a_12988_101.n3 GND 0.03fF
C277 a_12988_101.n4 GND 0.01fF
C278 a_12988_101.n5 GND 0.03fF
C279 a_12988_101.n6 GND 0.04fF
C280 a_12988_101.n7 GND 0.02fF
C281 a_12988_101.n8 GND 0.04fF
C282 a_12988_101.n9 GND 0.08fF
C283 a_12988_101.n10 GND 0.04fF
C284 a_12988_101.n11 GND 0.12fF
C285 a_12988_101.n12 GND 0.14fF
C286 a_12988_101.n13 GND 0.01fF
C287 a_7595_411.n0 GND 0.49fF
C288 a_7595_411.n1 GND 0.63fF
C289 a_7595_411.n2 GND 0.86fF
C290 a_7595_411.n3 GND 0.35fF
C291 a_7595_411.n4 GND 0.37fF
C292 a_7595_411.n5 GND 1.27fF
C293 a_7595_411.n6 GND 1.00fF
C294 a_7595_411.n7 GND 2.36fF
C295 a_7595_411.n8 GND 0.50fF
C296 a_7595_411.t7 GND 0.60fF
C297 a_7595_411.n9 GND 0.67fF
C298 a_7595_411.n10 GND 3.74fF
C299 a_7595_411.n11 GND 0.63fF
C300 a_7595_411.n12 GND 0.11fF
C301 a_7595_411.n13 GND 0.17fF
C302 a_7595_411.n14 GND 0.06fF
C303 a_6698_101.n0 GND 0.02fF
C304 a_6698_101.n1 GND 0.09fF
C305 a_6698_101.n2 GND 0.08fF
C306 a_6698_101.n3 GND 0.03fF
C307 a_6698_101.n4 GND 0.01fF
C308 a_6698_101.n5 GND 0.04fF
C309 a_6698_101.n6 GND 0.04fF
C310 a_6698_101.n7 GND 0.02fF
C311 a_6698_101.n8 GND 0.05fF
C312 a_6698_101.n9 GND 0.15fF
C313 a_6698_101.n10 GND 0.08fF
C314 a_6698_101.n11 GND 0.08fF
C315 a_6698_101.t1 GND 0.23fF
C316 a_6698_101.n12 GND 0.01fF
C317 a_6137_1050.n0 GND 0.04fF
C318 a_6137_1050.n1 GND 0.42fF
C319 a_6137_1050.n2 GND 0.54fF
C320 a_6137_1050.n3 GND 0.64fF
C321 a_6137_1050.n4 GND 0.36fF
C322 a_6137_1050.n5 GND 0.67fF
C323 a_6137_1050.n6 GND 0.74fF
C324 a_6137_1050.n7 GND 0.04fF
C325 a_6137_1050.n8 GND 0.25fF
C326 a_6137_1050.n9 GND 0.06fF
C327 a_9183_989.n0 GND 0.50fF
C328 a_9183_989.n1 GND 0.43fF
C329 a_9183_989.n2 GND 0.61fF
C330 a_9183_989.n3 GND 0.43fF
C331 a_9183_989.t9 GND 0.69fF
C332 a_9183_989.n4 GND 0.72fF
C333 a_9183_989.n5 GND 1.11fF
C334 a_9183_989.n6 GND 0.05fF
C335 a_9183_989.n7 GND 0.07fF
C336 a_9183_989.n8 GND 0.04fF
C337 a_9183_989.n9 GND 0.29fF
C338 a_9183_989.n10 GND 0.65fF
C339 a_9183_989.n11 GND 0.76fF
C340 a_9183_989.n12 GND 0.64fF
C341 a_11887_411.n0 GND 0.37fF
C342 a_11887_411.n1 GND 0.24fF
C343 a_11887_411.n2 GND 0.75fF
C344 a_11887_411.n3 GND 0.24fF
C345 a_11887_411.n4 GND 0.49fF
C346 a_11887_411.n5 GND 0.39fF
C347 a_11887_411.n6 GND 0.29fF
C348 a_11887_411.t11 GND 0.54fF
C349 a_11887_411.n7 GND 0.52fF
C350 a_11887_411.n8 GND 0.78fF
C351 a_11887_411.n9 GND 0.04fF
C352 a_11887_411.n10 GND 0.05fF
C353 a_11887_411.n11 GND 0.03fF
C354 a_11887_411.n12 GND 0.25fF
C355 a_11887_411.n13 GND 0.48fF
C356 a_11887_411.n14 GND 0.53fF
C357 a_11887_411.n15 GND 0.48fF
C358 a_11761_1050.n0 GND 0.37fF
C359 a_11761_1050.n1 GND 0.24fF
C360 a_11761_1050.n2 GND 0.65fF
C361 a_11761_1050.n3 GND 0.40fF
C362 a_11761_1050.n4 GND 0.61fF
C363 a_11761_1050.n5 GND 0.46fF
C364 a_11761_1050.n6 GND 0.47fF
C365 QN.n0 GND 0.30fF
C366 QN.n1 GND 0.38fF
C367 QN.n2 GND 0.46fF
C368 QN.n3 GND 0.04fF
C369 QN.n4 GND 0.05fF
C370 QN.n5 GND 0.06fF
C371 QN.n6 GND 0.14fF
C372 QN.n7 GND 1.07fF
C373 QN.n8 GND 0.14fF
C374 QN.n9 GND 0.38fF
C375 QN.n10 GND 0.35fF
C376 QN.n11 GND 0.01fF
C377 a_13654_101.n0 GND 0.02fF
C378 a_13654_101.n1 GND 0.13fF
C379 a_13654_101.n2 GND 0.15fF
C380 a_13654_101.n3 GND 0.16fF
C381 a_3303_411.n0 GND 0.59fF
C382 a_3303_411.n1 GND 0.55fF
C383 a_3303_411.n2 GND 0.67fF
C384 a_3303_411.n3 GND 0.93fF
C385 a_3303_411.n4 GND 0.56fF
C386 a_3303_411.n5 GND 5.97fF
C387 a_3303_411.n6 GND 0.51fF
C388 a_3303_411.t10 GND 0.77fF
C389 a_3303_411.n7 GND 0.82fF
C390 a_3303_411.n8 GND 7.69fF
C391 a_3303_411.n9 GND 0.06fF
C392 a_3303_411.n10 GND 0.08fF
C393 a_3303_411.n11 GND 0.05fF
C394 a_3303_411.n12 GND 0.30fF
C395 a_3303_411.n13 GND 0.75fF
C396 a_3303_411.n14 GND 0.93fF
C397 a_3303_411.n15 GND 0.75fF
C398 a_147_187.n0 GND 0.60fF
C399 a_147_187.n1 GND 0.44fF
C400 a_147_187.t5 GND 0.91fF
C401 a_147_187.n2 GND 0.99fF
C402 a_147_187.n3 GND 0.44fF
C403 a_147_187.t12 GND 0.91fF
C404 a_147_187.n4 GND 0.61fF
C405 a_147_187.n5 GND 0.45fF
C406 a_147_187.n6 GND 1.43fF
C407 a_147_187.n7 GND 2.16fF
C408 a_147_187.n8 GND 1.71fF
C409 a_147_187.n9 GND 0.62fF
C410 a_147_187.n10 GND 0.81fF
C411 a_147_187.n11 GND 0.81fF
C412 a_147_187.n12 GND 0.77fF
C413 a_1845_1050.n0 GND 0.38fF
C414 a_1845_1050.n1 GND 0.49fF
C415 a_1845_1050.n2 GND 0.57fF
C416 a_1845_1050.n3 GND 0.33fF
C417 a_1845_1050.n4 GND 0.60fF
C418 a_1845_1050.n5 GND 0.67fF
C419 a_1845_1050.n6 GND 0.08fF
C420 a_1845_1050.n7 GND 0.22fF
C421 a_1845_1050.n8 GND 0.04fF
C422 a_3177_1050.n0 GND 0.38fF
C423 a_3177_1050.n1 GND 0.30fF
C424 a_3177_1050.n2 GND 0.61fF
C425 a_3177_1050.n3 GND 0.36fF
C426 a_3177_1050.n4 GND 0.69fF
C427 a_3177_1050.n5 GND 0.55fF
C428 a_3177_1050.n6 GND 0.49fF
C429 a_277_1050.n0 GND 0.52fF
C430 a_277_1050.n1 GND 0.52fF
C431 a_277_1050.n2 GND 0.66fF
C432 a_277_1050.n3 GND 0.62fF
C433 a_277_1050.n4 GND 0.55fF
C434 a_277_1050.n5 GND 0.40fF
C435 a_277_1050.n6 GND 1.25fF
C436 a_277_1050.n7 GND 0.40fF
C437 a_277_1050.n8 GND 0.57fF
C438 a_277_1050.n9 GND 1.90fF
C439 a_277_1050.n10 GND 0.75fF
C440 a_277_1050.n11 GND 0.11fF
C441 a_277_1050.n12 GND 0.33fF
C442 a_277_1050.n13 GND 0.06fF
C443 VDD.n1 GND 0.03fF
C444 VDD.n2 GND 0.14fF
C445 VDD.n3 GND 0.03fF
C446 VDD.n4 GND 0.02fF
C447 VDD.n5 GND 0.06fF
C448 VDD.n6 GND 0.02fF
C449 VDD.n7 GND 0.02fF
C450 VDD.n8 GND 0.02fF
C451 VDD.n9 GND 0.02fF
C452 VDD.n10 GND 0.02fF
C453 VDD.n11 GND 0.02fF
C454 VDD.n12 GND 0.02fF
C455 VDD.n13 GND 0.02fF
C456 VDD.n14 GND 0.04fF
C457 VDD.n15 GND 0.01fF
C458 VDD.n20 GND 0.48fF
C459 VDD.n21 GND 0.29fF
C460 VDD.n22 GND 0.02fF
C461 VDD.n23 GND 0.04fF
C462 VDD.n24 GND 0.26fF
C463 VDD.n25 GND 0.01fF
C464 VDD.n26 GND 0.02fF
C465 VDD.n27 GND 0.01fF
C466 VDD.n28 GND 0.18fF
C467 VDD.n29 GND 0.01fF
C468 VDD.n30 GND 0.02fF
C469 VDD.n31 GND 0.08fF
C470 VDD.n32 GND 0.01fF
C471 VDD.n33 GND 0.03fF
C472 VDD.n34 GND 0.03fF
C473 VDD.n35 GND 0.15fF
C474 VDD.n36 GND 0.01fF
C475 VDD.n37 GND 0.03fF
C476 VDD.n38 GND 0.03fF
C477 VDD.n39 GND 0.17fF
C478 VDD.n40 GND 0.01fF
C479 VDD.n41 GND 0.02fF
C480 VDD.n42 GND 0.02fF
C481 VDD.n43 GND 0.26fF
C482 VDD.n44 GND 0.01fF
C483 VDD.n45 GND 0.02fF
C484 VDD.n46 GND 0.02fF
C485 VDD.n47 GND 0.29fF
C486 VDD.n48 GND 0.01fF
C487 VDD.n49 GND 0.02fF
C488 VDD.n50 GND 0.04fF
C489 VDD.n51 GND 0.06fF
C490 VDD.n52 GND 0.02fF
C491 VDD.n53 GND 0.02fF
C492 VDD.n54 GND 0.02fF
C493 VDD.n55 GND 0.02fF
C494 VDD.n56 GND 0.02fF
C495 VDD.n57 GND 0.02fF
C496 VDD.n58 GND 0.02fF
C497 VDD.n59 GND 0.02fF
C498 VDD.n60 GND 0.02fF
C499 VDD.n61 GND 0.02fF
C500 VDD.n62 GND 0.02fF
C501 VDD.n63 GND 0.03fF
C502 VDD.n64 GND 0.02fF
C503 VDD.n65 GND 0.23fF
C504 VDD.n66 GND 0.02fF
C505 VDD.n67 GND 0.02fF
C506 VDD.n69 GND 0.02fF
C507 VDD.n73 GND 0.29fF
C508 VDD.n74 GND 0.29fF
C509 VDD.n75 GND 0.01fF
C510 VDD.n76 GND 0.02fF
C511 VDD.n77 GND 0.04fF
C512 VDD.n78 GND 0.26fF
C513 VDD.n79 GND 0.01fF
C514 VDD.n80 GND 0.02fF
C515 VDD.n81 GND 0.02fF
C516 VDD.n82 GND 0.17fF
C517 VDD.n83 GND 0.01fF
C518 VDD.n84 GND 0.02fF
C519 VDD.n85 GND 0.02fF
C520 VDD.n86 GND 0.15fF
C521 VDD.n87 GND 0.01fF
C522 VDD.n88 GND 0.03fF
C523 VDD.n89 GND 0.03fF
C524 VDD.n90 GND 0.01fF
C525 VDD.n91 GND 0.03fF
C526 VDD.n92 GND 0.03fF
C527 VDD.n93 GND 0.18fF
C528 VDD.n94 GND 0.01fF
C529 VDD.n95 GND 0.02fF
C530 VDD.n96 GND 0.02fF
C531 VDD.n97 GND 0.26fF
C532 VDD.n98 GND 0.01fF
C533 VDD.n99 GND 0.02fF
C534 VDD.n100 GND 0.02fF
C535 VDD.n101 GND 0.29fF
C536 VDD.n102 GND 0.01fF
C537 VDD.n103 GND 0.02fF
C538 VDD.n104 GND 0.04fF
C539 VDD.n105 GND 0.23fF
C540 VDD.n106 GND 0.02fF
C541 VDD.n107 GND 0.02fF
C542 VDD.n108 GND 0.02fF
C543 VDD.n109 GND 0.06fF
C544 VDD.n110 GND 0.02fF
C545 VDD.n111 GND 0.02fF
C546 VDD.n112 GND 0.02fF
C547 VDD.n113 GND 0.02fF
C548 VDD.n114 GND 0.02fF
C549 VDD.n115 GND 0.02fF
C550 VDD.n116 GND 0.02fF
C551 VDD.n117 GND 0.02fF
C552 VDD.n118 GND 0.02fF
C553 VDD.n119 GND 0.02fF
C554 VDD.n120 GND 0.03fF
C555 VDD.n121 GND 0.02fF
C556 VDD.n122 GND 0.02fF
C557 VDD.n126 GND 0.29fF
C558 VDD.n127 GND 0.29fF
C559 VDD.n128 GND 0.01fF
C560 VDD.n129 GND 0.02fF
C561 VDD.n130 GND 0.04fF
C562 VDD.n131 GND 0.07fF
C563 VDD.n132 GND 0.26fF
C564 VDD.n133 GND 0.01fF
C565 VDD.n134 GND 0.01fF
C566 VDD.n135 GND 0.02fF
C567 VDD.n136 GND 0.18fF
C568 VDD.n137 GND 0.01fF
C569 VDD.n138 GND 0.02fF
C570 VDD.n139 GND 0.02fF
C571 VDD.n140 GND 0.09fF
C572 VDD.n141 GND 0.05fF
C573 VDD.n142 GND 0.01fF
C574 VDD.n143 GND 0.02fF
C575 VDD.n144 GND 0.03fF
C576 VDD.n145 GND 0.15fF
C577 VDD.n146 GND 0.01fF
C578 VDD.n147 GND 0.02fF
C579 VDD.n148 GND 0.03fF
C580 VDD.n149 GND 0.17fF
C581 VDD.n150 GND 0.01fF
C582 VDD.n151 GND 0.02fF
C583 VDD.n152 GND 0.02fF
C584 VDD.n153 GND 0.07fF
C585 VDD.n154 GND 0.26fF
C586 VDD.n155 GND 0.01fF
C587 VDD.n156 GND 0.01fF
C588 VDD.n157 GND 0.02fF
C589 VDD.n158 GND 0.29fF
C590 VDD.n159 GND 0.01fF
C591 VDD.n160 GND 0.02fF
C592 VDD.n161 GND 0.04fF
C593 VDD.n162 GND 0.23fF
C594 VDD.n163 GND 0.02fF
C595 VDD.n164 GND 0.02fF
C596 VDD.n165 GND 0.02fF
C597 VDD.n166 GND 0.06fF
C598 VDD.n167 GND 0.02fF
C599 VDD.n168 GND 0.02fF
C600 VDD.n169 GND 0.02fF
C601 VDD.n170 GND 0.02fF
C602 VDD.n171 GND 0.02fF
C603 VDD.n172 GND 0.02fF
C604 VDD.n173 GND 0.02fF
C605 VDD.n174 GND 0.02fF
C606 VDD.n175 GND 0.02fF
C607 VDD.n176 GND 0.02fF
C608 VDD.n177 GND 0.03fF
C609 VDD.n178 GND 0.02fF
C610 VDD.n179 GND 0.02fF
C611 VDD.n183 GND 0.29fF
C612 VDD.n184 GND 0.29fF
C613 VDD.n185 GND 0.01fF
C614 VDD.n186 GND 0.02fF
C615 VDD.n187 GND 0.04fF
C616 VDD.n188 GND 0.06fF
C617 VDD.n189 GND 0.26fF
C618 VDD.n190 GND 0.01fF
C619 VDD.n191 GND 0.01fF
C620 VDD.n192 GND 0.02fF
C621 VDD.n193 GND 0.18fF
C622 VDD.n194 GND 0.01fF
C623 VDD.n195 GND 0.02fF
C624 VDD.n196 GND 0.02fF
C625 VDD.n197 GND 0.09fF
C626 VDD.n198 GND 0.05fF
C627 VDD.n199 GND 0.01fF
C628 VDD.n200 GND 0.02fF
C629 VDD.n201 GND 0.03fF
C630 VDD.n202 GND 0.15fF
C631 VDD.n203 GND 0.01fF
C632 VDD.n204 GND 0.02fF
C633 VDD.n205 GND 0.03fF
C634 VDD.n206 GND 0.17fF
C635 VDD.n207 GND 0.01fF
C636 VDD.n208 GND 0.02fF
C637 VDD.n209 GND 0.02fF
C638 VDD.n210 GND 0.07fF
C639 VDD.n211 GND 0.26fF
C640 VDD.n212 GND 0.01fF
C641 VDD.n213 GND 0.01fF
C642 VDD.n214 GND 0.02fF
C643 VDD.n215 GND 0.29fF
C644 VDD.n216 GND 0.01fF
C645 VDD.n217 GND 0.02fF
C646 VDD.n218 GND 0.04fF
C647 VDD.n219 GND 0.23fF
C648 VDD.n220 GND 0.02fF
C649 VDD.n221 GND 0.02fF
C650 VDD.n222 GND 0.02fF
C651 VDD.n223 GND 0.06fF
C652 VDD.n224 GND 0.02fF
C653 VDD.n225 GND 0.02fF
C654 VDD.n226 GND 0.02fF
C655 VDD.n227 GND 0.02fF
C656 VDD.n228 GND 0.02fF
C657 VDD.n229 GND 0.02fF
C658 VDD.n230 GND 0.02fF
C659 VDD.n231 GND 0.02fF
C660 VDD.n232 GND 0.02fF
C661 VDD.n233 GND 0.02fF
C662 VDD.n234 GND 0.03fF
C663 VDD.n235 GND 0.02fF
C664 VDD.n236 GND 0.02fF
C665 VDD.n240 GND 0.29fF
C666 VDD.n241 GND 0.29fF
C667 VDD.n242 GND 0.01fF
C668 VDD.n243 GND 0.02fF
C669 VDD.n244 GND 0.04fF
C670 VDD.n245 GND 0.06fF
C671 VDD.n246 GND 0.26fF
C672 VDD.n247 GND 0.01fF
C673 VDD.n248 GND 0.01fF
C674 VDD.n249 GND 0.02fF
C675 VDD.n250 GND 0.18fF
C676 VDD.n251 GND 0.01fF
C677 VDD.n252 GND 0.02fF
C678 VDD.n253 GND 0.02fF
C679 VDD.n254 GND 0.09fF
C680 VDD.n255 GND 0.05fF
C681 VDD.n256 GND 0.01fF
C682 VDD.n257 GND 0.02fF
C683 VDD.n258 GND 0.03fF
C684 VDD.n259 GND 0.15fF
C685 VDD.n260 GND 0.01fF
C686 VDD.n261 GND 0.02fF
C687 VDD.n262 GND 0.03fF
C688 VDD.n263 GND 0.17fF
C689 VDD.n264 GND 0.01fF
C690 VDD.n265 GND 0.02fF
C691 VDD.n266 GND 0.02fF
C692 VDD.n267 GND 0.07fF
C693 VDD.n268 GND 0.26fF
C694 VDD.n269 GND 0.01fF
C695 VDD.n270 GND 0.01fF
C696 VDD.n271 GND 0.02fF
C697 VDD.n272 GND 0.29fF
C698 VDD.n273 GND 0.01fF
C699 VDD.n274 GND 0.02fF
C700 VDD.n275 GND 0.04fF
C701 VDD.n276 GND 0.23fF
C702 VDD.n277 GND 0.02fF
C703 VDD.n278 GND 0.02fF
C704 VDD.n279 GND 0.02fF
C705 VDD.n280 GND 0.06fF
C706 VDD.n281 GND 0.02fF
C707 VDD.n282 GND 0.02fF
C708 VDD.n283 GND 0.02fF
C709 VDD.n284 GND 0.02fF
C710 VDD.n285 GND 0.02fF
C711 VDD.n286 GND 0.02fF
C712 VDD.n287 GND 0.02fF
C713 VDD.n288 GND 0.02fF
C714 VDD.n289 GND 0.02fF
C715 VDD.n290 GND 0.02fF
C716 VDD.n291 GND 0.03fF
C717 VDD.n292 GND 0.02fF
C718 VDD.n293 GND 0.02fF
C719 VDD.n297 GND 0.29fF
C720 VDD.n298 GND 0.29fF
C721 VDD.n299 GND 0.01fF
C722 VDD.n300 GND 0.02fF
C723 VDD.n301 GND 0.04fF
C724 VDD.n302 GND 0.06fF
C725 VDD.n303 GND 0.26fF
C726 VDD.n304 GND 0.01fF
C727 VDD.n305 GND 0.01fF
C728 VDD.n306 GND 0.02fF
C729 VDD.n307 GND 0.18fF
C730 VDD.n308 GND 0.01fF
C731 VDD.n309 GND 0.02fF
C732 VDD.n310 GND 0.02fF
C733 VDD.n311 GND 0.09fF
C734 VDD.n312 GND 0.05fF
C735 VDD.n313 GND 0.01fF
C736 VDD.n314 GND 0.02fF
C737 VDD.n315 GND 0.03fF
C738 VDD.n316 GND 0.15fF
C739 VDD.n317 GND 0.01fF
C740 VDD.n318 GND 0.02fF
C741 VDD.n319 GND 0.03fF
C742 VDD.n320 GND 0.17fF
C743 VDD.n321 GND 0.01fF
C744 VDD.n322 GND 0.02fF
C745 VDD.n323 GND 0.02fF
C746 VDD.n324 GND 0.07fF
C747 VDD.n325 GND 0.26fF
C748 VDD.n326 GND 0.01fF
C749 VDD.n327 GND 0.01fF
C750 VDD.n328 GND 0.02fF
C751 VDD.n329 GND 0.29fF
C752 VDD.n330 GND 0.01fF
C753 VDD.n331 GND 0.02fF
C754 VDD.n332 GND 0.04fF
C755 VDD.n333 GND 0.23fF
C756 VDD.n334 GND 0.02fF
C757 VDD.n335 GND 0.02fF
C758 VDD.n336 GND 0.02fF
C759 VDD.n337 GND 0.06fF
C760 VDD.n338 GND 0.02fF
C761 VDD.n339 GND 0.02fF
C762 VDD.n340 GND 0.02fF
C763 VDD.n341 GND 0.02fF
C764 VDD.n342 GND 0.02fF
C765 VDD.n343 GND 0.02fF
C766 VDD.n344 GND 0.02fF
C767 VDD.n345 GND 0.02fF
C768 VDD.n346 GND 0.02fF
C769 VDD.n347 GND 0.02fF
C770 VDD.n348 GND 0.03fF
C771 VDD.n349 GND 0.02fF
C772 VDD.n350 GND 0.02fF
C773 VDD.n354 GND 0.29fF
C774 VDD.n355 GND 0.29fF
C775 VDD.n356 GND 0.01fF
C776 VDD.n357 GND 0.02fF
C777 VDD.n358 GND 0.04fF
C778 VDD.n359 GND 0.06fF
C779 VDD.n360 GND 0.26fF
C780 VDD.n361 GND 0.01fF
C781 VDD.n362 GND 0.01fF
C782 VDD.n363 GND 0.02fF
C783 VDD.n364 GND 0.18fF
C784 VDD.n365 GND 0.01fF
C785 VDD.n366 GND 0.02fF
C786 VDD.n367 GND 0.02fF
C787 VDD.n368 GND 0.09fF
C788 VDD.n369 GND 0.05fF
C789 VDD.n370 GND 0.01fF
C790 VDD.n371 GND 0.02fF
C791 VDD.n372 GND 0.03fF
C792 VDD.n373 GND 0.15fF
C793 VDD.n374 GND 0.01fF
C794 VDD.n375 GND 0.02fF
C795 VDD.n376 GND 0.03fF
C796 VDD.n377 GND 0.17fF
C797 VDD.n378 GND 0.01fF
C798 VDD.n379 GND 0.02fF
C799 VDD.n380 GND 0.02fF
C800 VDD.n381 GND 0.07fF
C801 VDD.n382 GND 0.26fF
C802 VDD.n383 GND 0.01fF
C803 VDD.n384 GND 0.01fF
C804 VDD.n385 GND 0.02fF
C805 VDD.n386 GND 0.29fF
C806 VDD.n387 GND 0.01fF
C807 VDD.n388 GND 0.02fF
C808 VDD.n389 GND 0.04fF
C809 VDD.n390 GND 0.23fF
C810 VDD.n391 GND 0.02fF
C811 VDD.n392 GND 0.02fF
C812 VDD.n393 GND 0.02fF
C813 VDD.n394 GND 0.06fF
C814 VDD.n395 GND 0.02fF
C815 VDD.n396 GND 0.02fF
C816 VDD.n397 GND 0.02fF
C817 VDD.n398 GND 0.02fF
C818 VDD.n399 GND 0.02fF
C819 VDD.n400 GND 0.02fF
C820 VDD.n401 GND 0.02fF
C821 VDD.n402 GND 0.02fF
C822 VDD.n403 GND 0.02fF
C823 VDD.n404 GND 0.02fF
C824 VDD.n405 GND 0.03fF
C825 VDD.n406 GND 0.02fF
C826 VDD.n407 GND 0.02fF
C827 VDD.n411 GND 0.29fF
C828 VDD.n412 GND 0.29fF
C829 VDD.n413 GND 0.01fF
C830 VDD.n414 GND 0.02fF
C831 VDD.n415 GND 0.04fF
C832 VDD.n416 GND 0.06fF
C833 VDD.n417 GND 0.26fF
C834 VDD.n418 GND 0.01fF
C835 VDD.n419 GND 0.01fF
C836 VDD.n420 GND 0.02fF
C837 VDD.n421 GND 0.18fF
C838 VDD.n422 GND 0.01fF
C839 VDD.n423 GND 0.02fF
C840 VDD.n424 GND 0.02fF
C841 VDD.n425 GND 0.09fF
C842 VDD.n426 GND 0.05fF
C843 VDD.n427 GND 0.01fF
C844 VDD.n428 GND 0.02fF
C845 VDD.n429 GND 0.03fF
C846 VDD.n430 GND 0.15fF
C847 VDD.n431 GND 0.01fF
C848 VDD.n432 GND 0.02fF
C849 VDD.n433 GND 0.03fF
C850 VDD.n434 GND 0.17fF
C851 VDD.n435 GND 0.01fF
C852 VDD.n436 GND 0.02fF
C853 VDD.n437 GND 0.02fF
C854 VDD.n438 GND 0.07fF
C855 VDD.n439 GND 0.26fF
C856 VDD.n440 GND 0.01fF
C857 VDD.n441 GND 0.01fF
C858 VDD.n442 GND 0.02fF
C859 VDD.n443 GND 0.29fF
C860 VDD.n444 GND 0.01fF
C861 VDD.n445 GND 0.02fF
C862 VDD.n446 GND 0.04fF
C863 VDD.n447 GND 0.28fF
C864 VDD.n448 GND 0.02fF
C865 VDD.n449 GND 0.02fF
C866 VDD.n450 GND 0.02fF
C867 VDD.n451 GND 0.06fF
C868 VDD.n452 GND 0.02fF
C869 VDD.n453 GND 0.02fF
C870 VDD.n454 GND 0.02fF
C871 VDD.n455 GND 0.02fF
C872 VDD.n456 GND 0.02fF
C873 VDD.n457 GND 0.02fF
C874 VDD.n458 GND 0.02fF
C875 VDD.n459 GND 0.02fF
C876 VDD.n460 GND 0.02fF
C877 VDD.n461 GND 0.02fF
C878 VDD.n462 GND 0.03fF
C879 VDD.n463 GND 0.02fF
C880 VDD.n464 GND 0.02fF
C881 VDD.n468 GND 0.29fF
C882 VDD.n469 GND 0.29fF
C883 VDD.n470 GND 0.01fF
C884 VDD.n471 GND 0.02fF
C885 VDD.n472 GND 0.04fF
C886 VDD.n473 GND 0.29fF
C887 VDD.n474 GND 0.01fF
C888 VDD.n475 GND 0.02fF
C889 VDD.n476 GND 0.02fF
C890 VDD.n477 GND 0.23fF
C891 VDD.n478 GND 0.01fF
C892 VDD.n479 GND 0.07fF
C893 VDD.n480 GND 0.02fF
C894 VDD.n481 GND 0.18fF
C895 VDD.n482 GND 0.01fF
C896 VDD.n483 GND 0.02fF
C897 VDD.n484 GND 0.02fF
C898 VDD.n485 GND 0.17fF
C899 VDD.n486 GND 0.01fF
C900 VDD.n487 GND 0.09fF
C901 VDD.n488 GND 0.05fF
C902 VDD.n489 GND 0.02fF
C903 VDD.n490 GND 0.02fF
C904 VDD.n491 GND 0.15fF
C905 VDD.n492 GND 0.02fF
C906 VDD.n493 GND 0.02fF
C907 VDD.n494 GND 0.03fF
C908 VDD.n495 GND 0.16fF
C909 VDD.n496 GND 0.02fF
C910 VDD.n497 GND 0.02fF
C911 VDD.n498 GND 0.03fF
C912 VDD.n499 GND 0.09fF
C913 VDD.n500 GND 0.05fF
C914 VDD.n501 GND 0.16fF
C915 VDD.n502 GND 0.01fF
C916 VDD.n503 GND 0.02fF
C917 VDD.n504 GND 0.02fF
C918 VDD.n505 GND 0.18fF
C919 VDD.n506 GND 0.01fF
C920 VDD.n507 GND 0.02fF
C921 VDD.n508 GND 0.02fF
C922 VDD.n509 GND 0.07fF
C923 VDD.n510 GND 0.24fF
C924 VDD.n511 GND 0.01fF
C925 VDD.n512 GND 0.01fF
C926 VDD.n513 GND 0.02fF
C927 VDD.n514 GND 0.29fF
C928 VDD.n515 GND 0.01fF
C929 VDD.n516 GND 0.02fF
C930 VDD.n517 GND 0.02fF
C931 VDD.n518 GND 0.29fF
C932 VDD.n519 GND 0.01fF
C933 VDD.n520 GND 0.02fF
C934 VDD.n521 GND 0.04fF
C935 VDD.n522 GND 0.28fF
C936 VDD.n523 GND 0.02fF
C937 VDD.n524 GND 0.02fF
C938 VDD.n525 GND 0.02fF
C939 VDD.n526 GND 0.06fF
C940 VDD.n527 GND 0.02fF
C941 VDD.n528 GND 0.02fF
C942 VDD.n529 GND 0.02fF
C943 VDD.n530 GND 0.02fF
C944 VDD.n531 GND 0.02fF
C945 VDD.n532 GND 0.02fF
C946 VDD.n533 GND 0.02fF
C947 VDD.n534 GND 0.02fF
C948 VDD.n535 GND 0.02fF
C949 VDD.n536 GND 0.02fF
C950 VDD.n537 GND 0.03fF
C951 VDD.n538 GND 0.02fF
C952 VDD.n539 GND 0.02fF
C953 VDD.n543 GND 0.29fF
C954 VDD.n544 GND 0.29fF
C955 VDD.n545 GND 0.01fF
C956 VDD.n546 GND 0.02fF
C957 VDD.n547 GND 0.04fF
C958 VDD.n548 GND 0.06fF
C959 VDD.n549 GND 0.26fF
C960 VDD.n550 GND 0.01fF
C961 VDD.n551 GND 0.01fF
C962 VDD.n552 GND 0.02fF
C963 VDD.n553 GND 0.18fF
C964 VDD.n554 GND 0.01fF
C965 VDD.n555 GND 0.02fF
C966 VDD.n556 GND 0.02fF
C967 VDD.n557 GND 0.09fF
C968 VDD.n558 GND 0.05fF
C969 VDD.n559 GND 0.01fF
C970 VDD.n560 GND 0.02fF
C971 VDD.n561 GND 0.03fF
C972 VDD.n562 GND 0.15fF
C973 VDD.n563 GND 0.01fF
C974 VDD.n564 GND 0.02fF
C975 VDD.n565 GND 0.03fF
C976 VDD.n566 GND 0.17fF
C977 VDD.n567 GND 0.01fF
C978 VDD.n568 GND 0.02fF
C979 VDD.n569 GND 0.02fF
C980 VDD.n570 GND 0.07fF
C981 VDD.n571 GND 0.26fF
C982 VDD.n572 GND 0.01fF
C983 VDD.n573 GND 0.01fF
C984 VDD.n574 GND 0.02fF
C985 VDD.n575 GND 0.29fF
C986 VDD.n576 GND 0.01fF
C987 VDD.n577 GND 0.02fF
C988 VDD.n578 GND 0.04fF
C989 VDD.n579 GND 0.23fF
C990 VDD.n580 GND 0.02fF
C991 VDD.n581 GND 0.02fF
C992 VDD.n582 GND 0.02fF
C993 VDD.n583 GND 0.06fF
C994 VDD.n584 GND 0.02fF
C995 VDD.n585 GND 0.02fF
C996 VDD.n586 GND 0.02fF
C997 VDD.n587 GND 0.02fF
C998 VDD.n588 GND 0.02fF
C999 VDD.n589 GND 0.02fF
C1000 VDD.n590 GND 0.02fF
C1001 VDD.n591 GND 0.02fF
C1002 VDD.n592 GND 0.02fF
C1003 VDD.n593 GND 0.02fF
C1004 VDD.n594 GND 0.03fF
C1005 VDD.n595 GND 0.02fF
C1006 VDD.n596 GND 0.02fF
C1007 VDD.n600 GND 0.29fF
C1008 VDD.n601 GND 0.29fF
C1009 VDD.n602 GND 0.01fF
C1010 VDD.n603 GND 0.02fF
C1011 VDD.n604 GND 0.04fF
C1012 VDD.n605 GND 0.06fF
C1013 VDD.n606 GND 0.26fF
C1014 VDD.n607 GND 0.01fF
C1015 VDD.n608 GND 0.01fF
C1016 VDD.n609 GND 0.02fF
C1017 VDD.n610 GND 0.18fF
C1018 VDD.n611 GND 0.01fF
C1019 VDD.n612 GND 0.02fF
C1020 VDD.n613 GND 0.02fF
C1021 VDD.n614 GND 0.09fF
C1022 VDD.n615 GND 0.05fF
C1023 VDD.n616 GND 0.01fF
C1024 VDD.n617 GND 0.02fF
C1025 VDD.n618 GND 0.03fF
C1026 VDD.n619 GND 0.15fF
C1027 VDD.n620 GND 0.01fF
C1028 VDD.n621 GND 0.02fF
C1029 VDD.n622 GND 0.03fF
C1030 VDD.n623 GND 0.17fF
C1031 VDD.n624 GND 0.01fF
C1032 VDD.n625 GND 0.02fF
C1033 VDD.n626 GND 0.02fF
C1034 VDD.n627 GND 0.19fF
C1035 VDD.n628 GND 0.02fF
C1036 VDD.n629 GND 0.02fF
C1037 VDD.n630 GND 0.06fF
C1038 VDD.n631 GND 0.02fF
C1039 VDD.n632 GND 0.02fF
C1040 VDD.n633 GND 0.02fF
C1041 VDD.n634 GND 0.02fF
C1042 VDD.n635 GND 0.02fF
C1043 VDD.n636 GND 0.02fF
C1044 VDD.n637 GND 0.02fF
C1045 VDD.n638 GND 0.02fF
C1046 VDD.n639 GND 0.03fF
C1047 VDD.n640 GND 0.04fF
C1048 VDD.n641 GND 0.02fF
C1049 VDD.n645 GND 0.48fF
C1050 VDD.n646 GND 0.29fF
C1051 VDD.n647 GND 0.02fF
C1052 VDD.n648 GND 0.03fF
C1053 VDD.n649 GND 0.03fF
C1054 VDD.n650 GND 0.29fF
C1055 VDD.n651 GND 0.01fF
C1056 VDD.n652 GND 0.02fF
C1057 VDD.n653 GND 0.02fF
C1058 VDD.n654 GND 0.07fF
C1059 VDD.n655 GND 0.24fF
C1060 VDD.n656 GND 0.01fF
C1061 VDD.n657 GND 0.01fF
C1062 VDD.n658 GND 0.02fF
C1063 VDD.n659 GND 0.18fF
C1064 VDD.n660 GND 0.01fF
C1065 VDD.n661 GND 0.02fF
C1066 VDD.n662 GND 0.02fF
C1067 VDD.n663 GND 0.09fF
C1068 VDD.n664 GND 0.05fF
C1069 VDD.n665 GND 0.16fF
C1070 VDD.n666 GND 0.01fF
C1071 VDD.n667 GND 0.02fF
C1072 VDD.n668 GND 0.02fF
C1073 VDD.n669 GND 0.16fF
C1074 VDD.n670 GND 0.02fF
C1075 VDD.n671 GND 0.02fF
C1076 VDD.n672 GND 0.03fF
C1077 VDD.n673 GND 0.15fF
C1078 VDD.n674 GND 0.02fF
C1079 VDD.n675 GND 0.02fF
C1080 VDD.n676 GND 0.03fF
C1081 VDD.n677 GND 0.17fF
C1082 VDD.n678 GND 0.01fF
C1083 VDD.n679 GND 0.09fF
C1084 VDD.n680 GND 0.05fF
C1085 VDD.n681 GND 0.02fF
C1086 VDD.n682 GND 0.02fF
C1087 VDD.n683 GND 0.18fF
C1088 VDD.n684 GND 0.01fF
C1089 VDD.n685 GND 0.02fF
C1090 VDD.n686 GND 0.02fF
C1091 VDD.n687 GND 0.23fF
C1092 VDD.n688 GND 0.01fF
C1093 VDD.n689 GND 0.07fF
C1094 VDD.n690 GND 0.02fF
C1095 VDD.n691 GND 0.29fF
C1096 VDD.n692 GND 0.01fF
C1097 VDD.n693 GND 0.02fF
C1098 VDD.n694 GND 0.02fF
C1099 VDD.n695 GND 0.29fF
C1100 VDD.n696 GND 0.01fF
C1101 VDD.n697 GND 0.02fF
C1102 VDD.n698 GND 0.04fF
C1103 VDD.n699 GND 0.06fF
C1104 VDD.n700 GND 0.02fF
C1105 VDD.n701 GND 0.02fF
C1106 VDD.n702 GND 0.02fF
C1107 VDD.n703 GND 0.02fF
C1108 VDD.n704 GND 0.02fF
C1109 VDD.n705 GND 0.02fF
C1110 VDD.n706 GND 0.02fF
C1111 VDD.n707 GND 0.02fF
C1112 VDD.n708 GND 0.02fF
C1113 VDD.n709 GND 0.02fF
C1114 VDD.n710 GND 0.02fF
C1115 VDD.n711 GND 0.03fF
C1116 VDD.n712 GND 0.02fF
C1117 VDD.n715 GND 0.02fF
C1118 VDD.n717 GND 0.02fF
C1119 VDD.n718 GND 0.28fF
C1120 VDD.n719 GND 0.02fF
C1121 VDD.n721 GND 0.29fF
C1122 VDD.n722 GND 0.29fF
C1123 VDD.n723 GND 0.01fF
C1124 VDD.n724 GND 0.02fF
C1125 VDD.n725 GND 0.04fF
C1126 VDD.n726 GND 0.07fF
C1127 VDD.n727 GND 0.26fF
C1128 VDD.n728 GND 0.01fF
C1129 VDD.n729 GND 0.01fF
C1130 VDD.n730 GND 0.02fF
C1131 VDD.n731 GND 0.17fF
C1132 VDD.n732 GND 0.01fF
C1133 VDD.n733 GND 0.02fF
C1134 VDD.n734 GND 0.02fF
C1135 VDD.n735 GND 0.15fF
C1136 VDD.n736 GND 0.01fF
C1137 VDD.n737 GND 0.02fF
C1138 VDD.n738 GND 0.03fF
C1139 VDD.n739 GND 0.09fF
C1140 VDD.n740 GND 0.05fF
C1141 VDD.n741 GND 0.01fF
C1142 VDD.n742 GND 0.02fF
C1143 VDD.n743 GND 0.03fF
C1144 VDD.n744 GND 0.18fF
C1145 VDD.n745 GND 0.01fF
C1146 VDD.n746 GND 0.02fF
C1147 VDD.n747 GND 0.02fF
C1148 VDD.n748 GND 0.06fF
C1149 VDD.n749 GND 0.26fF
C1150 VDD.n750 GND 0.01fF
C1151 VDD.n751 GND 0.01fF
C1152 VDD.n752 GND 0.02fF
C1153 VDD.n753 GND 0.29fF
C1154 VDD.n754 GND 0.01fF
C1155 VDD.n755 GND 0.02fF
C1156 VDD.n756 GND 0.04fF
C1157 VDD.n757 GND 0.23fF
C1158 VDD.n758 GND 0.02fF
C1159 VDD.n759 GND 0.02fF
C1160 VDD.n760 GND 0.02fF
C1161 VDD.n761 GND 0.06fF
C1162 VDD.n762 GND 0.02fF
C1163 VDD.n763 GND 0.02fF
C1164 VDD.n764 GND 0.02fF
C1165 VDD.n765 GND 0.02fF
C1166 VDD.n766 GND 0.02fF
C1167 VDD.n767 GND 0.02fF
C1168 VDD.n768 GND 0.02fF
C1169 VDD.n769 GND 0.02fF
C1170 VDD.n770 GND 0.02fF
C1171 VDD.n771 GND 0.02fF
C1172 VDD.n772 GND 0.03fF
C1173 VDD.n773 GND 0.02fF
C1174 VDD.n774 GND 0.02fF
C1175 VDD.n778 GND 0.29fF
C1176 VDD.n779 GND 0.29fF
C1177 VDD.n780 GND 0.01fF
C1178 VDD.n781 GND 0.02fF
C1179 VDD.n782 GND 0.04fF
C1180 VDD.n783 GND 0.07fF
C1181 VDD.n784 GND 0.26fF
C1182 VDD.n785 GND 0.01fF
C1183 VDD.n786 GND 0.01fF
C1184 VDD.n787 GND 0.02fF
C1185 VDD.n788 GND 0.17fF
C1186 VDD.n789 GND 0.01fF
C1187 VDD.n790 GND 0.02fF
C1188 VDD.n791 GND 0.02fF
C1189 VDD.n792 GND 0.15fF
C1190 VDD.n793 GND 0.01fF
C1191 VDD.n794 GND 0.02fF
C1192 VDD.n795 GND 0.03fF
C1193 VDD.n796 GND 0.09fF
C1194 VDD.n797 GND 0.05fF
C1195 VDD.n798 GND 0.01fF
C1196 VDD.n799 GND 0.02fF
C1197 VDD.n800 GND 0.03fF
C1198 VDD.n801 GND 0.18fF
C1199 VDD.n802 GND 0.01fF
C1200 VDD.n803 GND 0.02fF
C1201 VDD.n804 GND 0.02fF
C1202 VDD.n805 GND 0.06fF
C1203 VDD.n806 GND 0.26fF
C1204 VDD.n807 GND 0.01fF
C1205 VDD.n808 GND 0.01fF
C1206 VDD.n809 GND 0.02fF
C1207 VDD.n810 GND 0.29fF
C1208 VDD.n811 GND 0.01fF
C1209 VDD.n812 GND 0.02fF
C1210 VDD.n813 GND 0.04fF
C1211 VDD.n814 GND 0.23fF
C1212 VDD.n815 GND 0.02fF
C1213 VDD.n816 GND 0.02fF
C1214 VDD.n817 GND 0.02fF
C1215 VDD.n818 GND 0.06fF
C1216 VDD.n819 GND 0.02fF
C1217 VDD.n820 GND 0.02fF
C1218 VDD.n821 GND 0.02fF
C1219 VDD.n822 GND 0.02fF
C1220 VDD.n823 GND 0.02fF
C1221 VDD.n824 GND 0.02fF
C1222 VDD.n825 GND 0.02fF
C1223 VDD.n826 GND 0.02fF
C1224 VDD.n827 GND 0.02fF
C1225 VDD.n828 GND 0.02fF
C1226 VDD.n829 GND 0.03fF
C1227 VDD.n830 GND 0.02fF
C1228 VDD.n831 GND 0.02fF
C1229 VDD.n835 GND 0.29fF
C1230 VDD.n836 GND 0.29fF
C1231 VDD.n837 GND 0.01fF
C1232 VDD.n838 GND 0.02fF
C1233 VDD.n839 GND 0.04fF
C1234 VDD.n840 GND 0.07fF
C1235 VDD.n841 GND 0.26fF
C1236 VDD.n842 GND 0.01fF
C1237 VDD.n843 GND 0.01fF
C1238 VDD.n844 GND 0.02fF
C1239 VDD.n845 GND 0.17fF
C1240 VDD.n846 GND 0.01fF
C1241 VDD.n847 GND 0.02fF
C1242 VDD.n848 GND 0.02fF
C1243 VDD.n849 GND 0.15fF
C1244 VDD.n850 GND 0.01fF
C1245 VDD.n851 GND 0.02fF
C1246 VDD.n852 GND 0.03fF
C1247 VDD.n853 GND 0.09fF
C1248 VDD.n854 GND 0.05fF
C1249 VDD.n855 GND 0.01fF
C1250 VDD.n856 GND 0.02fF
C1251 VDD.n857 GND 0.03fF
C1252 VDD.n858 GND 0.18fF
C1253 VDD.n859 GND 0.01fF
C1254 VDD.n860 GND 0.02fF
C1255 VDD.n861 GND 0.02fF
C1256 VDD.n862 GND 0.06fF
C1257 VDD.n863 GND 0.26fF
C1258 VDD.n864 GND 0.01fF
C1259 VDD.n865 GND 0.01fF
C1260 VDD.n866 GND 0.02fF
C1261 VDD.n867 GND 0.29fF
C1262 VDD.n868 GND 0.01fF
C1263 VDD.n869 GND 0.02fF
C1264 VDD.n870 GND 0.04fF
C1265 VDD.n871 GND 0.23fF
C1266 VDD.n872 GND 0.02fF
C1267 VDD.n873 GND 0.02fF
C1268 VDD.n874 GND 0.02fF
C1269 VDD.n875 GND 0.06fF
C1270 VDD.n876 GND 0.02fF
C1271 VDD.n877 GND 0.02fF
C1272 VDD.n878 GND 0.02fF
C1273 VDD.n879 GND 0.02fF
C1274 VDD.n880 GND 0.02fF
C1275 VDD.n881 GND 0.02fF
C1276 VDD.n882 GND 0.02fF
C1277 VDD.n883 GND 0.02fF
C1278 VDD.n884 GND 0.02fF
C1279 VDD.n885 GND 0.02fF
C1280 VDD.n886 GND 0.03fF
C1281 VDD.n887 GND 0.02fF
C1282 VDD.n888 GND 0.02fF
C1283 VDD.n892 GND 0.29fF
C1284 VDD.n893 GND 0.29fF
C1285 VDD.n894 GND 0.01fF
C1286 VDD.n895 GND 0.02fF
C1287 VDD.n896 GND 0.04fF
C1288 VDD.n897 GND 0.07fF
C1289 VDD.n898 GND 0.26fF
C1290 VDD.n899 GND 0.01fF
C1291 VDD.n900 GND 0.01fF
C1292 VDD.n901 GND 0.02fF
C1293 VDD.n902 GND 0.17fF
C1294 VDD.n903 GND 0.01fF
C1295 VDD.n904 GND 0.02fF
C1296 VDD.n905 GND 0.02fF
C1297 VDD.n906 GND 0.15fF
C1298 VDD.n907 GND 0.01fF
C1299 VDD.n908 GND 0.02fF
C1300 VDD.n909 GND 0.03fF
C1301 VDD.n910 GND 0.09fF
C1302 VDD.n911 GND 0.05fF
C1303 VDD.n912 GND 0.01fF
C1304 VDD.n913 GND 0.02fF
C1305 VDD.n914 GND 0.03fF
C1306 VDD.n915 GND 0.18fF
C1307 VDD.n916 GND 0.01fF
C1308 VDD.n917 GND 0.02fF
C1309 VDD.n918 GND 0.02fF
C1310 VDD.n919 GND 0.06fF
C1311 VDD.n920 GND 0.26fF
C1312 VDD.n921 GND 0.01fF
C1313 VDD.n922 GND 0.01fF
C1314 VDD.n923 GND 0.02fF
C1315 VDD.n924 GND 0.29fF
C1316 VDD.n925 GND 0.01fF
C1317 VDD.n926 GND 0.02fF
C1318 VDD.n927 GND 0.04fF
C1319 VDD.n928 GND 0.23fF
C1320 VDD.n929 GND 0.02fF
C1321 VDD.n930 GND 0.02fF
C1322 VDD.n931 GND 0.02fF
C1323 VDD.n932 GND 0.06fF
C1324 VDD.n933 GND 0.02fF
C1325 VDD.n934 GND 0.02fF
C1326 VDD.n935 GND 0.02fF
C1327 VDD.n936 GND 0.02fF
C1328 VDD.n937 GND 0.02fF
C1329 VDD.n938 GND 0.02fF
C1330 VDD.n939 GND 0.02fF
C1331 VDD.n940 GND 0.02fF
C1332 VDD.n941 GND 0.02fF
C1333 VDD.n942 GND 0.02fF
C1334 VDD.n943 GND 0.03fF
C1335 VDD.n944 GND 0.02fF
C1336 VDD.n945 GND 0.02fF
C1337 VDD.n949 GND 0.29fF
C1338 VDD.n950 GND 0.29fF
C1339 VDD.n951 GND 0.01fF
C1340 VDD.n952 GND 0.02fF
C1341 VDD.n953 GND 0.04fF
C1342 VDD.n954 GND 0.07fF
C1343 VDD.n955 GND 0.26fF
C1344 VDD.n956 GND 0.01fF
C1345 VDD.n957 GND 0.01fF
C1346 VDD.n958 GND 0.02fF
C1347 VDD.n959 GND 0.17fF
C1348 VDD.n960 GND 0.01fF
C1349 VDD.n961 GND 0.02fF
C1350 VDD.n962 GND 0.02fF
C1351 VDD.n963 GND 0.15fF
C1352 VDD.n964 GND 0.01fF
C1353 VDD.n965 GND 0.02fF
C1354 VDD.n966 GND 0.03fF
C1355 VDD.n967 GND 0.09fF
C1356 VDD.n968 GND 0.05fF
C1357 VDD.n969 GND 0.01fF
C1358 VDD.n970 GND 0.02fF
C1359 VDD.n971 GND 0.03fF
C1360 VDD.n972 GND 0.18fF
C1361 VDD.n973 GND 0.01fF
C1362 VDD.n974 GND 0.02fF
C1363 VDD.n975 GND 0.02fF
C1364 VDD.n976 GND 0.06fF
C1365 VDD.n977 GND 0.26fF
C1366 VDD.n978 GND 0.01fF
C1367 VDD.n979 GND 0.01fF
C1368 VDD.n980 GND 0.02fF
C1369 VDD.n981 GND 0.29fF
C1370 VDD.n982 GND 0.01fF
C1371 VDD.n983 GND 0.02fF
C1372 VDD.n984 GND 0.04fF
C1373 VDD.n985 GND 0.28fF
C1374 VDD.n986 GND 0.02fF
C1375 VDD.n987 GND 0.02fF
C1376 VDD.n988 GND 0.02fF
C1377 VDD.n989 GND 0.06fF
C1378 VDD.n990 GND 0.02fF
C1379 VDD.n991 GND 0.02fF
C1380 VDD.n992 GND 0.02fF
C1381 VDD.n993 GND 0.02fF
C1382 VDD.n994 GND 0.02fF
C1383 VDD.n995 GND 0.02fF
C1384 VDD.n996 GND 0.02fF
C1385 VDD.n997 GND 0.02fF
C1386 VDD.n998 GND 0.02fF
C1387 VDD.n999 GND 0.02fF
C1388 VDD.n1000 GND 0.03fF
C1389 VDD.n1001 GND 0.02fF
C1390 VDD.n1002 GND 0.02fF
C1391 VDD.n1006 GND 0.29fF
C1392 VDD.n1007 GND 0.29fF
C1393 VDD.n1008 GND 0.01fF
C1394 VDD.n1009 GND 0.02fF
C1395 VDD.n1010 GND 0.04fF
C1396 VDD.n1011 GND 0.29fF
C1397 VDD.n1012 GND 0.01fF
C1398 VDD.n1013 GND 0.02fF
C1399 VDD.n1014 GND 0.02fF
C1400 VDD.n1015 GND 0.07fF
C1401 VDD.n1016 GND 0.24fF
C1402 VDD.n1017 GND 0.01fF
C1403 VDD.n1018 GND 0.01fF
C1404 VDD.n1019 GND 0.02fF
C1405 VDD.n1020 GND 0.18fF
C1406 VDD.n1021 GND 0.01fF
C1407 VDD.n1022 GND 0.02fF
C1408 VDD.n1023 GND 0.02fF
C1409 VDD.n1024 GND 0.09fF
C1410 VDD.n1025 GND 0.05fF
C1411 VDD.n1026 GND 0.16fF
C1412 VDD.n1027 GND 0.01fF
C1413 VDD.n1028 GND 0.02fF
C1414 VDD.n1029 GND 0.02fF
C1415 VDD.n1030 GND 0.16fF
C1416 VDD.n1031 GND 0.02fF
C1417 VDD.n1032 GND 0.02fF
C1418 VDD.n1033 GND 0.03fF
C1419 VDD.n1034 GND 0.15fF
C1420 VDD.n1035 GND 0.02fF
C1421 VDD.n1036 GND 0.02fF
C1422 VDD.n1037 GND 0.03fF
C1423 VDD.n1038 GND 0.17fF
C1424 VDD.n1039 GND 0.01fF
C1425 VDD.n1040 GND 0.09fF
C1426 VDD.n1041 GND 0.05fF
C1427 VDD.n1042 GND 0.02fF
C1428 VDD.n1043 GND 0.02fF
C1429 VDD.n1044 GND 0.18fF
C1430 VDD.n1045 GND 0.01fF
C1431 VDD.n1046 GND 0.02fF
C1432 VDD.n1047 GND 0.02fF
C1433 VDD.n1048 GND 0.23fF
C1434 VDD.n1049 GND 0.01fF
C1435 VDD.n1050 GND 0.07fF
C1436 VDD.n1051 GND 0.02fF
C1437 VDD.n1052 GND 0.29fF
C1438 VDD.n1053 GND 0.01fF
C1439 VDD.n1054 GND 0.02fF
C1440 VDD.n1055 GND 0.02fF
C1441 VDD.n1056 GND 0.29fF
C1442 VDD.n1057 GND 0.01fF
C1443 VDD.n1058 GND 0.02fF
C1444 VDD.n1059 GND 0.04fF
C1445 VDD.n1060 GND 0.28fF
C1446 VDD.n1061 GND 0.02fF
C1447 VDD.n1062 GND 0.02fF
C1448 VDD.n1063 GND 0.02fF
C1449 VDD.n1064 GND 0.06fF
C1450 VDD.n1065 GND 0.02fF
C1451 VDD.n1066 GND 0.02fF
C1452 VDD.n1067 GND 0.02fF
C1453 VDD.n1068 GND 0.02fF
C1454 VDD.n1069 GND 0.02fF
C1455 VDD.n1070 GND 0.02fF
C1456 VDD.n1071 GND 0.02fF
C1457 VDD.n1072 GND 0.02fF
C1458 VDD.n1073 GND 0.02fF
C1459 VDD.n1074 GND 0.02fF
C1460 VDD.n1075 GND 0.03fF
C1461 VDD.n1076 GND 0.02fF
C1462 VDD.n1077 GND 0.02fF
C1463 VDD.n1081 GND 0.29fF
C1464 VDD.n1082 GND 0.29fF
C1465 VDD.n1083 GND 0.01fF
C1466 VDD.n1084 GND 0.02fF
C1467 VDD.n1085 GND 0.04fF
C1468 VDD.n1086 GND 0.07fF
C1469 VDD.n1087 GND 0.26fF
C1470 VDD.n1088 GND 0.01fF
C1471 VDD.n1089 GND 0.01fF
C1472 VDD.n1090 GND 0.02fF
C1473 VDD.n1091 GND 0.17fF
C1474 VDD.n1092 GND 0.01fF
C1475 VDD.n1093 GND 0.02fF
C1476 VDD.n1094 GND 0.02fF
C1477 VDD.n1095 GND 0.15fF
C1478 VDD.n1096 GND 0.01fF
C1479 VDD.n1097 GND 0.02fF
C1480 VDD.n1098 GND 0.03fF
C1481 VDD.n1099 GND 0.09fF
C1482 VDD.n1100 GND 0.05fF
C1483 VDD.n1101 GND 0.01fF
C1484 VDD.n1102 GND 0.02fF
C1485 VDD.n1103 GND 0.03fF
C1486 VDD.n1104 GND 0.18fF
C1487 VDD.n1105 GND 0.01fF
C1488 VDD.n1106 GND 0.02fF
C1489 VDD.n1107 GND 0.02fF
C1490 VDD.n1108 GND 0.06fF
C1491 VDD.n1109 GND 0.26fF
C1492 VDD.n1110 GND 0.01fF
C1493 VDD.n1111 GND 0.01fF
C1494 VDD.n1112 GND 0.02fF
C1495 VDD.n1113 GND 0.29fF
C1496 VDD.n1114 GND 0.01fF
C1497 VDD.n1115 GND 0.02fF
C1498 VDD.n1116 GND 0.04fF
C1499 VDD.n1117 GND 0.23fF
C1500 VDD.n1118 GND 0.02fF
C1501 VDD.n1119 GND 0.02fF
C1502 VDD.n1120 GND 0.02fF
C1503 VDD.n1121 GND 0.06fF
C1504 VDD.n1122 GND 0.02fF
C1505 VDD.n1123 GND 0.02fF
C1506 VDD.n1124 GND 0.02fF
C1507 VDD.n1125 GND 0.02fF
C1508 VDD.n1126 GND 0.02fF
C1509 VDD.n1127 GND 0.02fF
C1510 VDD.n1128 GND 0.02fF
C1511 VDD.n1129 GND 0.02fF
C1512 VDD.n1130 GND 0.02fF
C1513 VDD.n1131 GND 0.02fF
C1514 VDD.n1132 GND 0.03fF
C1515 VDD.n1133 GND 0.02fF
C1516 VDD.n1134 GND 0.02fF
C1517 VDD.n1138 GND 0.29fF
C1518 VDD.n1139 GND 0.29fF
C1519 VDD.n1140 GND 0.01fF
C1520 VDD.n1141 GND 0.02fF
C1521 VDD.n1142 GND 0.04fF
C1522 VDD.n1143 GND 0.07fF
C1523 VDD.n1144 GND 0.26fF
C1524 VDD.n1145 GND 0.01fF
C1525 VDD.n1146 GND 0.01fF
C1526 VDD.n1147 GND 0.02fF
C1527 VDD.n1148 GND 0.17fF
C1528 VDD.n1149 GND 0.01fF
C1529 VDD.n1150 GND 0.02fF
C1530 VDD.n1151 GND 0.02fF
C1531 VDD.n1152 GND 0.15fF
C1532 VDD.n1153 GND 0.01fF
C1533 VDD.n1154 GND 0.02fF
C1534 VDD.n1155 GND 0.03fF
C1535 VDD.n1156 GND 0.09fF
C1536 VDD.n1157 GND 0.05fF
C1537 VDD.n1158 GND 0.01fF
C1538 VDD.n1159 GND 0.02fF
C1539 VDD.n1160 GND 0.03fF
C1540 VDD.n1161 GND 0.18fF
C1541 VDD.n1162 GND 0.01fF
C1542 VDD.n1163 GND 0.02fF
C1543 VDD.n1164 GND 0.02fF
C1544 VDD.n1165 GND 0.06fF
C1545 VDD.n1166 GND 0.26fF
C1546 VDD.n1167 GND 0.01fF
C1547 VDD.n1168 GND 0.01fF
C1548 VDD.n1169 GND 0.02fF
C1549 VDD.n1170 GND 0.29fF
C1550 VDD.n1171 GND 0.01fF
C1551 VDD.n1172 GND 0.02fF
C1552 VDD.n1173 GND 0.04fF
C1553 VDD.n1174 GND 0.23fF
C1554 VDD.n1175 GND 0.02fF
C1555 VDD.n1176 GND 0.02fF
C1556 VDD.n1177 GND 0.02fF
C1557 VDD.n1178 GND 0.06fF
C1558 VDD.n1179 GND 0.02fF
C1559 VDD.n1180 GND 0.02fF
C1560 VDD.n1181 GND 0.02fF
C1561 VDD.n1182 GND 0.02fF
C1562 VDD.n1183 GND 0.02fF
C1563 VDD.n1184 GND 0.02fF
C1564 VDD.n1185 GND 0.02fF
C1565 VDD.n1186 GND 0.02fF
C1566 VDD.n1187 GND 0.02fF
C1567 VDD.n1188 GND 0.02fF
C1568 VDD.n1189 GND 0.03fF
C1569 VDD.n1190 GND 0.02fF
C1570 VDD.n1191 GND 0.02fF
C1571 VDD.n1195 GND 0.29fF
C1572 VDD.n1196 GND 0.29fF
C1573 VDD.n1197 GND 0.01fF
C1574 VDD.n1198 GND 0.02fF
C1575 VDD.n1199 GND 0.04fF
C1576 VDD.n1200 GND 0.07fF
C1577 VDD.n1201 GND 0.26fF
C1578 VDD.n1202 GND 0.01fF
C1579 VDD.n1203 GND 0.01fF
C1580 VDD.n1204 GND 0.02fF
C1581 VDD.n1205 GND 0.17fF
C1582 VDD.n1206 GND 0.01fF
C1583 VDD.n1207 GND 0.02fF
C1584 VDD.n1208 GND 0.02fF
C1585 VDD.n1209 GND 0.15fF
C1586 VDD.n1210 GND 0.01fF
C1587 VDD.n1211 GND 0.02fF
C1588 VDD.n1212 GND 0.03fF
C1589 VDD.n1213 GND 0.09fF
C1590 VDD.n1214 GND 0.05fF
C1591 VDD.n1215 GND 0.01fF
C1592 VDD.n1216 GND 0.02fF
C1593 VDD.n1217 GND 0.03fF
C1594 VDD.n1218 GND 0.18fF
C1595 VDD.n1219 GND 0.01fF
C1596 VDD.n1220 GND 0.02fF
C1597 VDD.n1221 GND 0.02fF
C1598 VDD.n1222 GND 0.06fF
C1599 VDD.n1223 GND 0.26fF
C1600 VDD.n1224 GND 0.01fF
C1601 VDD.n1225 GND 0.01fF
C1602 VDD.n1226 GND 0.02fF
C1603 VDD.n1227 GND 0.29fF
C1604 VDD.n1228 GND 0.01fF
C1605 VDD.n1229 GND 0.02fF
C1606 VDD.n1230 GND 0.04fF
C1607 VDD.n1231 GND 0.23fF
C1608 VDD.n1232 GND 0.02fF
C1609 VDD.n1233 GND 0.02fF
C1610 VDD.n1234 GND 0.02fF
C1611 VDD.n1235 GND 0.06fF
C1612 VDD.n1236 GND 0.02fF
C1613 VDD.n1237 GND 0.02fF
C1614 VDD.n1238 GND 0.02fF
C1615 VDD.n1239 GND 0.02fF
C1616 VDD.n1240 GND 0.02fF
C1617 VDD.n1241 GND 0.02fF
C1618 VDD.n1242 GND 0.02fF
C1619 VDD.n1243 GND 0.02fF
C1620 VDD.n1244 GND 0.02fF
C1621 VDD.n1245 GND 0.02fF
C1622 VDD.n1246 GND 0.03fF
C1623 VDD.n1247 GND 0.02fF
C1624 VDD.n1248 GND 0.02fF
C1625 VDD.n1252 GND 0.29fF
C1626 VDD.n1253 GND 0.29fF
C1627 VDD.n1254 GND 0.01fF
C1628 VDD.n1255 GND 0.02fF
C