magic
tech sky130A
magscale 1 2
timestamp 1649945909
<< nwell >>
rect -84 832 232 1575
<< psubdiff >>
rect -31 546 179 572
rect -31 512 -17 546
rect 17 512 131 546
rect 165 512 179 546
rect -31 510 179 512
rect -31 474 31 510
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect -31 368 -17 402
rect 17 368 31 402
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect -31 62 31 80
rect 117 474 179 510
rect 117 440 131 474
rect 165 440 179 474
rect 117 402 179 440
rect 117 368 131 402
rect 165 368 179 402
rect 117 330 179 368
rect 117 296 131 330
rect 165 296 179 330
rect 117 258 179 296
rect 117 224 131 258
rect 165 224 179 258
rect 117 186 179 224
rect 117 152 131 186
rect 165 152 179 186
rect 117 114 179 152
rect 117 80 131 114
rect 165 80 179 114
rect 117 62 179 80
rect -31 11 179 62
<< nsubdiff >>
rect -31 1492 179 1539
rect -31 1470 31 1492
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect -31 1038 31 1076
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect -31 930 31 932
rect 117 1470 179 1492
rect 117 1436 131 1470
rect 165 1436 179 1470
rect 117 1398 179 1436
rect 117 1364 131 1398
rect 165 1364 179 1398
rect 117 1326 179 1364
rect 117 1292 131 1326
rect 165 1292 179 1326
rect 117 1254 179 1292
rect 117 1220 131 1254
rect 165 1220 179 1254
rect 117 1182 179 1220
rect 117 1148 131 1182
rect 165 1148 179 1182
rect 117 1110 179 1148
rect 117 1076 131 1110
rect 165 1076 179 1110
rect 117 1038 179 1076
rect 117 1004 131 1038
rect 165 1004 179 1038
rect 117 966 179 1004
rect 117 932 131 966
rect 165 932 179 966
rect 117 930 179 932
rect -31 868 179 930
<< psubdiffcont >>
rect -17 512 17 546
rect 131 512 165 546
rect -17 440 17 474
rect -17 368 17 402
rect -17 296 17 330
rect -17 224 17 258
rect -17 152 17 186
rect -17 80 17 114
rect 131 440 165 474
rect 131 368 165 402
rect 131 296 165 330
rect 131 224 165 258
rect 131 152 165 186
rect 131 80 165 114
<< nsubdiffcont >>
rect -17 1436 17 1470
rect -17 1364 17 1398
rect -17 1292 17 1326
rect -17 1220 17 1254
rect -17 1148 17 1182
rect -17 1076 17 1110
rect -17 1004 17 1038
rect -17 932 17 966
rect 131 1436 165 1470
rect 131 1364 165 1398
rect 131 1292 165 1326
rect 131 1220 165 1254
rect 131 1148 165 1182
rect 131 1076 165 1110
rect 131 1004 165 1038
rect 131 932 165 966
<< locali >>
rect -31 1492 179 1554
rect -31 1470 31 1492
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect -31 1038 31 1076
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect -31 868 31 932
rect 117 1470 179 1492
rect 117 1436 131 1470
rect 165 1436 179 1470
rect 117 1398 179 1436
rect 117 1364 131 1398
rect 165 1364 179 1398
rect 117 1326 179 1364
rect 117 1292 131 1326
rect 165 1292 179 1326
rect 117 1254 179 1292
rect 117 1220 131 1254
rect 165 1220 179 1254
rect 117 1182 179 1220
rect 117 1148 131 1182
rect 165 1148 179 1182
rect 117 1110 179 1148
rect 117 1076 131 1110
rect 165 1076 179 1110
rect 117 1038 179 1076
rect 117 1004 131 1038
rect 165 1004 179 1038
rect 117 966 179 1004
rect 117 932 131 966
rect 165 932 179 966
rect 117 868 179 932
rect -31 546 31 572
rect -31 512 -17 546
rect 17 512 31 546
rect -31 474 31 512
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect -31 368 -17 402
rect 17 368 31 402
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect -31 62 31 80
rect 117 546 179 572
rect 117 512 131 546
rect 165 512 179 546
rect 117 474 179 512
rect 117 440 131 474
rect 165 440 179 474
rect 117 402 179 440
rect 117 368 131 402
rect 165 368 179 402
rect 117 330 179 368
rect 117 296 131 330
rect 165 296 179 330
rect 117 258 179 296
rect 117 224 131 258
rect 165 224 179 258
rect 117 186 179 224
rect 117 152 131 186
rect 165 152 179 186
rect 117 114 179 152
rect 117 80 131 114
rect 165 80 179 114
rect 117 62 179 80
rect -31 0 179 62
<< metal1 >>
rect -31 1492 179 1554
rect -31 0 179 62
<< end >>
