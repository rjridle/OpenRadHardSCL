** sch_path: /home/rjridle/OpenRadHardSCL/lib/xschem/INVX1.sch
.subckt INVX1 A Y
*.PININFO A:I Y:O
M3 Y A VDD VDD pmos w=2u l=0.150u m=1
M2 Y A VDD VDD pmos w=2u l=0.150u m=1
M1 Y A GND GND nmos w=3u l=0.150u m=1
.ends
.GLOBAL GND
.GLOBAL VDD
.end
