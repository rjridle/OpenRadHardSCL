magic
tech sky130
magscale 1 2
timestamp 1645049645
<< poly >>
rect 44 469 110 479
rect 44 435 60 469
rect 94 435 110 469
rect 44 425 110 435
<< polycont >>
rect 60 435 94 469
<< locali >>
rect 44 435 60 469
rect 94 435 110 469
<< viali >>
rect 60 435 94 469
<< metal1 >>
rect 60 475 94 481
rect 54 469 100 475
rect 54 435 60 469
rect 94 435 100 469
rect 54 429 100 435
rect 60 399 94 429
<< end >>
