magic
tech sky130A
magscale 1 2
timestamp 1645051963
<< nmos >>
rect 11 150 41 212
rect 11 120 107 150
tri 107 120 137 150 sw
rect 11 112 49 120
tri 49 112 57 120 nw
tri 91 112 99 120 ne
rect 99 112 137 120
rect 11 31 41 112
tri 41 104 49 112 nw
tri 99 104 107 112 ne
tri 41 31 42 32 sw
tri 106 31 107 32 se
rect 107 31 137 112
rect 11 30 42 31
tri 42 30 43 31 sw
tri 105 30 106 31 se
rect 106 30 137 31
rect 11 29 43 30
tri 43 29 44 30 sw
tri 104 29 105 30 se
rect 105 29 137 30
rect 11 28 44 29
tri 44 28 45 29 sw
tri 103 28 104 29 se
rect 104 28 137 29
rect 11 27 45 28
tri 45 27 46 28 sw
tri 102 27 103 28 se
rect 103 27 137 28
rect 11 26 46 27
tri 46 26 47 27 sw
tri 101 26 102 27 se
rect 102 26 137 27
rect 11 25 47 26
tri 47 25 48 26 sw
tri 100 25 101 26 se
rect 101 25 137 26
rect 11 24 48 25
tri 48 24 49 25 sw
tri 99 24 100 25 se
rect 100 24 137 25
rect 11 23 49 24
tri 49 23 50 24 sw
tri 98 23 99 24 se
rect 99 23 137 24
rect 11 22 50 23
tri 50 22 51 23 sw
tri 97 22 98 23 se
rect 98 22 137 23
rect 11 21 51 22
tri 51 21 52 22 sw
tri 96 21 97 22 se
rect 97 21 137 22
rect 11 16 52 21
tri 52 16 57 21 sw
tri 95 20 96 21 se
rect 96 20 137 21
tri 91 16 95 20 se
rect 95 16 137 20
tri 11 -14 41 16 ne
rect 41 -14 107 16
tri 107 -14 137 16 nw
<< ndiff >>
rect -45 196 11 212
rect -45 162 -35 196
rect -1 162 11 196
rect -45 125 11 162
rect 41 196 193 212
rect 41 162 57 196
rect 91 162 149 196
rect 183 162 193 196
rect 41 150 193 162
rect -45 91 -35 125
rect -1 91 11 125
tri 107 120 137 150 ne
rect 137 125 193 150
tri 49 112 57 120 se
rect 57 112 91 120
tri 91 112 99 120 sw
rect -45 57 11 91
rect -45 23 -35 57
rect -1 23 11 57
tri 41 104 49 112 se
rect 49 104 99 112
tri 99 104 107 112 sw
rect 41 68 107 104
rect 41 34 57 68
rect 91 34 107 68
rect 41 32 107 34
tri 41 31 42 32 ne
rect 42 31 106 32
tri 106 31 107 32 nw
rect 137 91 149 125
rect 183 91 193 125
rect 137 57 193 91
tri 42 30 43 31 ne
rect 43 30 105 31
tri 105 30 106 31 nw
tri 43 29 44 30 ne
rect 44 29 104 30
tri 104 29 105 30 nw
tri 44 28 45 29 ne
rect 45 28 103 29
tri 103 28 104 29 nw
tri 45 27 46 28 ne
rect 46 27 102 28
tri 102 27 103 28 nw
tri 46 26 47 27 ne
rect 47 26 101 27
tri 101 26 102 27 nw
tri 47 25 48 26 ne
rect 48 25 100 26
tri 100 25 101 26 nw
tri 48 24 49 25 ne
rect 49 24 99 25
tri 99 24 100 25 nw
tri 49 23 50 24 ne
rect 50 23 98 24
tri 98 23 99 24 nw
rect 137 23 149 57
rect 183 23 193 57
rect -45 -14 11 23
tri 50 22 51 23 ne
rect 51 22 97 23
tri 97 22 98 23 nw
tri 51 21 52 22 ne
rect 52 21 96 22
tri 96 21 97 22 nw
tri 52 16 57 21 ne
rect 57 20 95 21
tri 95 20 96 21 nw
rect 57 16 91 20
tri 91 16 95 20 nw
tri 11 -14 41 16 sw
tri 107 -14 137 16 se
rect 137 -14 193 23
rect -45 -48 -35 -14
rect -1 -48 149 -14
rect 183 -48 193 -14
rect -45 -64 193 -48
<< ndiffc >>
rect -35 162 -1 196
rect 57 162 91 196
rect 149 162 183 196
rect -35 91 -1 125
rect -35 23 -1 57
rect 57 34 91 68
rect 149 91 183 125
rect 149 23 183 57
rect -35 -48 -1 -14
rect 149 -48 183 -14
<< poly >>
rect 11 212 41 238
<< locali >>
rect -35 196 -1 212
rect 149 196 183 212
rect -1 162 57 196
rect 91 162 149 196
rect -35 125 -1 162
rect -35 57 -1 91
rect 149 125 183 162
rect -35 -14 -1 23
rect -35 -64 -1 -48
rect 57 68 91 84
rect 57 -64 91 34
rect 149 57 183 91
rect 149 -14 183 23
rect 149 -64 183 -48
<< end >>
