* SPICE3 file created from diff_ring_side.ext - technology: sky130A

