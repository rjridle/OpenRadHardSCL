magic
tech sky130A
magscale 1 2
timestamp 1651077508
<< metal1 >>
rect -31 1492 2029 1554
rect 131 945 165 979
rect 353 871 387 905
rect 1833 796 1867 831
rect 1167 427 1201 461
rect -31 0 2029 62
use li1_M1_contact  li1_M1_contact_3 pcells
timestamp 1648061256
transform -1 0 1850 0 -1 814
box -53 -33 29 33
use votern3x1_pcell  votern3x1_pcell_0 pcells
timestamp 1648740297
transform 1 0 0 0 1 0
box -84 0 2082 1575
<< labels >>
rlabel metal1 1833 797 1867 831 1 YN
port 1 n
rlabel metal1 353 871 387 905 1 A
port 2 n
rlabel metal1 131 945 165 979 1 B
port 3 n
rlabel metal1 1167 427 1201 461 1 C
port 4 n
rlabel metal1 -31 1492 2029 1554 1 VDD
rlabel metal1 -31 0 2029 62 1 GND
<< end >>
