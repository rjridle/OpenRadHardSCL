magic
tech sky130A
magscale 1 2
timestamp 1647328248
<< nwell >>
rect 84 1539 360 1575
rect 55 1505 360 1539
rect 84 832 360 1505
<< pdiffc >>
rect 117 1105 151 1139
rect 205 1105 239 1139
rect 293 1105 327 1139
<< psubdiff >>
rect 31 510 413 572
rect 31 13 55 47
rect 89 13 127 47
rect 161 13 205 47
rect 239 13 283 47
rect 317 13 355 47
rect 389 13 413 47
<< nsubdiff >>
rect 31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 205 1539
rect 239 1505 283 1539
rect 317 1505 355 1539
rect 389 1505 413 1539
rect 31 868 413 930
<< psubdiffcont >>
rect 55 13 89 47
rect 127 13 161 47
rect 205 13 239 47
rect 283 13 317 47
rect 355 13 389 47
<< nsubdiffcont >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 205 1505 239 1539
rect 283 1505 317 1539
rect 355 1505 389 1539
<< poly >>
rect 175 411 184 441
rect 154 410 184 411
<< locali >>
rect 31 1539 413 1554
rect 31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 205 1539
rect 239 1505 283 1539
rect 317 1505 355 1539
rect 389 1505 413 1539
rect 31 1492 413 1505
rect 117 1139 151 1157
rect 117 1083 151 1105
rect 205 1139 239 1157
rect 205 979 239 1105
rect 293 1139 327 1157
rect 293 1083 327 1105
rect 131 477 165 954
rect 205 945 313 979
rect 279 461 313 945
rect 205 427 313 461
rect 205 261 239 427
rect 108 62 142 101
rect 205 62 239 117
rect 302 62 336 101
rect 31 47 413 62
rect 31 13 55 47
rect 89 13 127 47
rect 161 13 205 47
rect 239 13 283 47
rect 317 13 355 47
rect 389 13 413 47
rect 31 0 413 13
<< viali >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 205 1505 239 1539
rect 283 1505 317 1539
rect 355 1505 389 1539
rect 55 13 89 47
rect 127 13 161 47
rect 205 13 239 47
rect 283 13 317 47
rect 355 13 389 47
<< metal1 >>
rect 31 1539 413 1554
rect 31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 205 1539
rect 239 1505 283 1539
rect 317 1505 355 1539
rect 389 1505 413 1539
rect 31 1492 413 1505
rect 31 47 413 62
rect 31 13 55 47
rect 89 13 127 47
rect 161 13 205 47
rect 239 13 283 47
rect 317 13 355 47
rect 389 13 413 47
rect 31 0 413 13
use pmos2  pmos2_0
timestamp 1647328240
transform 1 0 19 0 1 1450
box 52 -460 352 42
use poly_li1_contact  poly_li1_contact_0
timestamp 1645652543
transform 0 1 148 -1 0 987
box -33 -27 33 27
use poly_li1_contact  poly_li1_contact_1
timestamp 1645652543
transform 0 -1 148 1 0 444
box -33 -27 33 27
use nmos_top  nmos_top_0
timestamp 1645648650
transform -1 0 345 0 1 101
box -1 0 247 309
use diff_ring_side  diff_ring_side_0
timestamp 1646086970
transform 1 0 444 0 1 0
box -84 0 84 1575
use diff_ring_side  diff_ring_side_1
timestamp 1646086970
transform 1 0 0 0 1 0
box -84 0 84 1575
<< end >>
