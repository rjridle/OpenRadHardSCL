magic
tech sky130A
magscale 1 2
timestamp 1645909608
<< nwell >>
rect 84 832 360 1575
<< ndiff >>
rect 205 195 239 293
<< pdiffc >>
rect 205 1105 239 1139
<< psubdiff >>
rect 31 510 413 572
rect 31 13 55 47
rect 89 13 127 47
rect 161 13 205 47
rect 239 13 283 47
rect 317 13 355 47
rect 389 13 413 47
rect 31 12 413 13
<< nsubdiff >>
rect 31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 205 1539
rect 239 1505 283 1539
rect 317 1505 355 1539
rect 389 1505 413 1539
rect 31 868 413 930
<< psubdiffcont >>
rect 55 13 89 47
rect 127 13 161 47
rect 205 13 239 47
rect 283 13 317 47
rect 355 13 389 47
<< nsubdiffcont >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 205 1505 239 1539
rect 283 1505 317 1539
rect 355 1505 389 1539
<< poly >>
rect 131 470 184 477
rect 121 416 184 470
rect 131 411 184 416
rect 154 410 184 411
<< locali >>
rect 31 1539 413 1554
rect 31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 205 1539
rect 239 1505 283 1539
rect 317 1505 355 1539
rect 389 1505 413 1539
rect 31 1492 413 1505
rect 131 477 165 954
rect 131 461 148 477
rect 131 427 165 461
rect 205 195 239 1090
rect 108 62 142 101
rect 205 62 239 117
rect 302 62 336 101
rect 31 47 413 62
rect 31 13 55 47
rect 89 13 127 47
rect 161 13 205 47
rect 239 13 283 47
rect 317 13 355 47
rect 389 13 413 47
rect 31 0 413 13
<< viali >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 205 1505 239 1539
rect 283 1505 317 1539
rect 355 1505 389 1539
rect 55 13 89 47
rect 127 13 161 47
rect 205 13 239 47
rect 283 13 317 47
rect 355 13 389 47
<< metal1 >>
rect 31 1539 413 1554
rect 31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 205 1539
rect 239 1505 283 1539
rect 317 1505 355 1539
rect 389 1505 413 1539
rect 31 1492 413 1505
rect 131 723 165 757
rect 205 649 239 683
rect 31 47 413 62
rect 31 13 55 47
rect 89 13 127 47
rect 161 13 205 47
rect 239 13 283 47
rect 317 13 355 47
rect 389 13 413 47
rect 31 0 413 13
use pmos2  pmos2_0 pcells
timestamp 1645909547
transform 1 0 19 0 1 1450
box 52 -460 352 42
use diff_ring_side  diff_ring_side_0 pcells
timestamp 1645641539
transform 1 0 444 0 1 0
box -84 0 84 1575
use diff_ring_side  diff_ring_side_1
timestamp 1645641539
transform 1 0 0 0 1 0
box -84 0 84 1575
use nmos_top  nmos_top_0 pcells
timestamp 1645648650
transform -1 0 345 0 1 101
box -1 0 247 309
use poly_li1_contact  poly_li1_contact_0 pcells
timestamp 1645652543
transform 0 1 148 -1 0 987
box -33 -27 33 27
use poly_li1_contact  poly_li1_contact_1
timestamp 1645652543
transform 0 -1 148 1 0 444
box -33 -27 33 27
use li1_M1_contact_perp_ext  li1_M1_contact_perp_ext_0 pcells
timestamp 1645050501
transform 0 -1 148 1 0 740
box -23 -53 49 29
use li1_M1_contact_perp_ext  li1_M1_contact_perp_ext_1
timestamp 1645050501
transform 0 -1 222 1 0 666
box -23 -53 49 29
<< labels >>
rlabel metal1 148 740 148 740 1 A
port 1 n
rlabel metal1 222 666 222 666 1 Y
port 2 n
rlabel metal1 72 1522 72 1522 1 VDD
port 3 n
rlabel metal1 72 30 72 30 1 VSS
port 4 n
<< end >>
