VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO INVX1
  CLASS BLOCK ;
  FOREIGN INVX1 ;
  ORIGIN 0.795 0.000 ;
  SIZE 2.790 BY 6.765 ;
  OBS
      LAYER nwell ;
        RECT -0.795 3.060 1.995 6.765 ;
      LAYER li1 ;
        RECT -0.615 6.350 1.815 6.660 ;
        RECT -0.615 3.240 -0.305 6.350 ;
        RECT 0.050 4.235 0.220 6.350 ;
        RECT -0.010 3.740 0.320 3.910 ;
        RECT -0.615 0.310 -0.305 2.745 ;
        RECT 0.070 1.995 0.240 2.325 ;
        RECT 0.050 0.715 0.220 1.825 ;
        RECT 0.490 0.950 0.660 6.145 ;
        RECT 0.930 4.270 1.100 6.350 ;
        RECT 1.505 3.240 1.815 6.350 ;
        RECT 0.970 0.715 1.140 1.790 ;
        RECT -0.035 0.545 1.225 0.715 ;
        RECT 0.050 0.310 0.220 0.545 ;
        RECT 0.970 0.310 1.140 0.545 ;
        RECT 1.495 0.310 1.805 2.745 ;
        RECT -0.615 0.000 1.805 0.310 ;
      LAYER mcon ;
        RECT -0.220 6.415 -0.050 6.585 ;
        RECT 0.120 6.415 0.290 6.585 ;
        RECT 0.460 6.415 0.630 6.585 ;
        RECT 0.800 6.415 0.975 6.585 ;
        RECT 1.145 6.415 1.320 6.585 ;
        RECT -0.545 6.075 -0.370 6.245 ;
        RECT -0.545 5.735 -0.370 5.905 ;
        RECT -0.545 5.395 -0.370 5.565 ;
        RECT -0.545 5.055 -0.370 5.225 ;
        RECT -0.545 4.715 -0.370 4.885 ;
        RECT -0.545 4.375 -0.370 4.545 ;
        RECT 0.490 4.250 0.660 4.420 ;
        RECT 1.570 6.075 1.745 6.245 ;
        RECT 1.570 5.735 1.745 5.905 ;
        RECT 1.570 5.395 1.745 5.565 ;
        RECT 1.570 5.055 1.745 5.225 ;
        RECT 1.570 4.715 1.745 4.885 ;
        RECT 1.570 4.375 1.745 4.545 ;
        RECT -0.545 4.035 -0.370 4.205 ;
        RECT -0.545 3.695 -0.370 3.865 ;
        RECT 0.070 3.740 0.240 3.910 ;
        RECT -0.540 2.105 -0.370 2.275 ;
        RECT 0.070 2.075 0.240 2.245 ;
        RECT -0.540 1.765 -0.370 1.935 ;
        RECT -0.540 1.425 -0.370 1.595 ;
        RECT -0.540 1.085 -0.370 1.255 ;
        RECT -0.540 0.745 -0.370 0.915 ;
        RECT 1.570 4.035 1.745 4.205 ;
        RECT 1.570 3.695 1.745 3.865 ;
        RECT 1.565 2.105 1.735 2.275 ;
        RECT 1.565 1.765 1.735 1.935 ;
        RECT 1.565 1.425 1.735 1.595 ;
        RECT 1.565 1.085 1.735 1.255 ;
        RECT 1.565 0.745 1.735 0.915 ;
        RECT -0.545 0.405 -0.375 0.575 ;
        RECT 1.565 0.405 1.735 0.575 ;
        RECT -0.220 0.065 -0.050 0.235 ;
        RECT 0.120 0.065 0.290 0.235 ;
        RECT 0.465 0.065 0.635 0.235 ;
        RECT 0.835 0.065 1.005 0.235 ;
        RECT 1.175 0.065 1.345 0.235 ;
      LAYER met1 ;
        RECT -0.615 6.350 1.815 6.660 ;
        RECT -0.615 3.240 -0.305 6.350 ;
        RECT 0.490 4.450 0.660 4.480 ;
        RECT 0.460 4.220 0.690 4.450 ;
        RECT 0.070 3.940 0.240 3.970 ;
        RECT 0.040 3.710 0.270 3.940 ;
        RECT 0.490 3.850 0.660 4.220 ;
        RECT -0.615 0.310 -0.305 2.745 ;
        RECT 0.070 2.280 0.240 3.710 ;
        RECT 1.505 3.240 1.815 6.350 ;
        RECT 0.040 2.040 0.270 2.280 ;
        RECT 0.070 1.960 0.240 2.040 ;
        RECT 1.495 0.310 1.805 2.745 ;
        RECT -0.615 0.000 1.805 0.310 ;
  END
END INVX1
END LIBRARY

