magic
tech sky130A
magscale 1 2
timestamp 1645051859
<< nmos >>
rect 11 162 41 212
rect 11 132 107 162
tri 107 132 137 162 sw
rect 11 28 41 132
tri 41 116 57 132 nw
tri 91 119 104 132 ne
rect 104 119 137 132
tri 104 116 107 119 ne
tri 41 28 57 44 sw
tri 104 41 107 44 se
rect 107 41 137 119
tri 103 40 104 41 se
rect 104 40 137 41
tri 102 39 103 40 se
rect 103 39 137 40
tri 101 38 102 39 se
rect 102 38 137 39
tri 100 37 101 38 se
rect 101 37 137 38
tri 99 36 100 37 se
rect 100 36 137 37
tri 98 35 99 36 se
rect 99 35 137 36
tri 97 34 98 35 se
rect 98 34 137 35
tri 96 33 97 34 se
rect 97 33 137 34
tri 95 32 96 33 se
rect 96 32 137 33
tri 94 31 95 32 se
rect 95 31 137 32
tri 93 30 94 31 se
rect 94 30 137 31
tri 92 29 93 30 se
rect 93 29 137 30
rect 92 28 137 29
tri 11 -2 41 28 ne
rect 41 -2 107 28
tri 107 -2 137 28 nw
<< ndiff >>
rect -45 196 11 212
rect -45 162 -35 196
rect -1 162 11 196
rect 41 196 193 212
rect 41 162 149 196
rect 183 162 193 196
rect -45 125 11 162
tri 107 132 137 162 ne
rect -45 91 -35 125
rect -1 91 11 125
rect -45 57 11 91
rect -45 23 -35 57
rect -1 23 11 57
tri 41 116 57 132 se
rect 57 119 91 132
tri 91 119 104 132 sw
rect 137 125 193 162
rect 57 116 104 119
tri 104 116 107 119 sw
rect 41 80 107 116
rect 41 46 57 80
rect 91 46 107 80
rect 41 44 107 46
tri 41 28 57 44 ne
rect 57 41 104 44
tri 104 41 107 44 nw
rect 137 91 149 125
rect 183 91 193 125
rect 137 57 193 91
rect 57 40 103 41
tri 103 40 104 41 nw
rect 57 39 102 40
tri 102 39 103 40 nw
rect 57 38 101 39
tri 101 38 102 39 nw
rect 57 37 100 38
tri 100 37 101 38 nw
rect 57 36 99 37
tri 99 36 100 37 nw
rect 57 35 98 36
tri 98 35 99 36 nw
rect 57 34 97 35
tri 97 34 98 35 nw
rect 57 33 96 34
tri 96 33 97 34 nw
rect 57 32 95 33
tri 95 32 96 33 nw
rect 57 31 94 32
tri 94 31 95 32 nw
rect 57 30 93 31
tri 93 30 94 31 nw
rect 57 28 92 30
tri 92 29 93 30 nw
rect -45 -2 11 23
tri 11 -2 41 28 sw
tri 107 -2 137 28 se
rect 137 23 149 57
rect 183 23 193 57
rect 137 -2 193 23
rect -45 -14 193 -2
rect -45 -48 -35 -14
rect -1 -48 57 -14
rect 91 -48 149 -14
rect 183 -48 193 -14
rect -45 -64 193 -48
<< ndiffc >>
rect -35 162 -1 196
rect 149 162 183 196
rect -35 91 -1 125
rect -35 23 -1 57
rect 57 46 91 80
rect 149 91 183 125
rect 149 23 183 57
rect -35 -48 -1 -14
rect 57 -48 91 -14
rect 149 -48 183 -14
<< poly >>
rect 11 212 41 238
<< locali >>
rect -35 196 -1 212
rect -35 125 -1 162
rect 149 196 183 212
rect 149 125 183 162
rect -35 57 -1 91
rect 57 80 91 96
rect 57 30 91 46
rect 149 57 183 91
rect -35 -14 -1 23
rect 149 -14 183 23
rect -1 -48 57 -14
rect 91 -48 149 -14
rect -35 -64 -1 -48
rect 149 -64 183 -48
<< end >>
