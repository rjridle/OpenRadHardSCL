magic
tech sky130A
magscale 1 2
timestamp 1643178442
<< nmos >>
rect 107 150 137 212
tri 11 120 41 150 se
rect 41 120 137 150
rect 11 28 41 120
tri 41 104 57 120 nw
tri 91 104 107 120 ne
tri 41 28 57 44 sw
tri 91 28 107 44 se
rect 107 28 137 120
tri 11 -2 41 28 ne
rect 41 -2 107 28
tri 107 -2 137 28 nw
<< ndiff >>
rect -45 196 107 212
rect -45 162 -35 196
rect -1 162 107 196
rect -45 150 107 162
rect 137 196 193 212
rect 137 162 149 196
rect 183 162 193 196
rect -45 125 11 150
rect -45 91 -35 125
rect -1 91 11 125
tri 11 120 41 150 nw
rect -45 57 11 91
rect -45 23 -35 57
rect -1 23 11 57
tri 41 104 57 120 se
rect 57 104 91 120
tri 91 104 107 120 sw
rect 41 91 107 104
rect 41 57 57 91
rect 91 57 107 91
rect 41 44 107 57
tri 41 28 57 44 ne
rect 57 28 91 44
tri 91 28 107 44 nw
rect -45 -2 11 23
tri 11 -2 41 28 sw
tri 107 -2 137 28 se
rect 137 -2 193 162
rect -45 -14 193 -2
rect -45 -48 -35 -14
rect -1 -48 53 -14
rect 87 -48 149 -14
rect 183 -48 193 -14
rect -45 -64 193 -48
<< ndiffc >>
rect -35 162 -1 196
rect 149 162 183 196
rect -35 91 -1 125
rect -35 23 -1 57
rect 57 57 91 91
rect -35 -48 -1 -14
rect 53 -48 87 -14
rect 149 -48 183 -14
<< poly >>
rect 107 212 137 238
<< locali >>
rect -35 196 -1 212
rect 149 196 183 212
rect -1 162 149 196
rect -35 125 -1 162
rect 149 125 183 162
rect -35 57 -1 91
rect 57 91 91 107
rect 91 57 183 91
rect 57 41 91 57
rect -35 -14 -1 23
rect 149 -14 183 17
rect -1 -48 53 -14
rect 87 -48 149 -14
rect -35 -64 -1 -48
rect 149 -64 183 -48
<< end >>
