magic
tech sky130A
magscale 1 2
timestamp 1645917848
<< nmos >>
tri 146 215 162 231 se
rect 162 215 192 276
tri 56 185 86 215 se
rect 86 185 192 215
rect 56 85 86 185
tri 86 169 102 185 nw
tri 146 169 162 185 ne
tri 86 85 102 101 sw
tri 146 85 162 101 se
rect 162 85 192 185
tri 56 55 86 85 ne
rect 86 55 162 85
tri 162 55 192 85 nw
<< ndiff >>
rect 0 260 162 276
rect 0 226 10 260
rect 44 226 107 260
rect 141 231 162 260
rect 141 226 146 231
rect 0 215 146 226
tri 146 215 162 231 nw
rect 192 260 248 276
rect 192 226 204 260
rect 238 226 248 260
rect 0 189 56 215
rect 0 155 10 189
rect 44 155 56 189
tri 56 185 86 215 nw
rect 192 189 248 226
rect 0 121 56 155
rect 0 87 10 121
rect 44 87 56 121
rect 0 55 56 87
tri 86 169 102 185 se
rect 102 169 146 185
tri 146 169 162 185 sw
rect 86 136 162 169
rect 86 102 107 136
rect 141 102 162 136
rect 86 101 162 102
tri 86 85 102 101 ne
rect 102 85 146 101
tri 146 85 162 101 nw
rect 192 155 204 189
rect 238 155 248 189
rect 192 121 248 155
rect 192 87 204 121
rect 238 87 248 121
tri 56 55 86 85 sw
tri 162 55 192 85 se
rect 192 55 248 87
rect 0 50 248 55
rect 0 16 10 50
rect 44 16 204 50
rect 238 16 248 50
rect 0 0 248 16
<< ndiffc >>
rect 10 226 44 260
rect 107 226 141 260
rect 204 226 238 260
rect 10 155 44 189
rect 10 87 44 121
rect 107 102 141 136
rect 204 155 238 189
rect 204 87 238 121
rect 10 16 44 50
rect 204 16 238 50
<< poly >>
rect 162 276 192 302
<< locali >>
rect 10 260 44 276
rect 204 260 238 276
rect 44 226 107 260
rect 141 226 204 260
rect 10 189 44 226
rect 10 121 44 155
rect 204 189 238 226
rect 10 50 44 87
rect 107 136 141 152
rect 107 86 141 102
rect 204 121 238 155
rect 10 0 44 16
rect 204 50 238 87
rect 204 0 238 16
<< end >>
