* SPICE3 file created from TMRDFFSNRNQNX1.ext - technology: sky130A

.subckt TMRDFFSNRNQNX1 QN D CLK SN RN VDD GND
X0 GND a_6049_1050.t8 a_6825_103.t0 GND sky130_fd_pr__nfet_01v8 ad=3.7611p pd=3.297u as=0p ps=0u w=0u l=0u
X1 VDD.t227 RN.t1 a_15669_1050.t5 pV�U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X2 GND a_4125_1050.t7 a_4901_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X3 a_599_989.t5 CLK.t0 VDD.t182 P_��U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X4 VDD.t225 RN.t2 a_9897_1050.t6  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X5 VDD.t67 CLK.t1 a_1561_989.t2 VDD.t66 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X6 a_11821_1050.t4 a_12143_989.t7 VDD.t87 �+���~ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X7 VDD.t163 a_13105_989.t7 a_13745_1050.t5  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X8 VDD.t77 a_277_1050.t7 a_2201_1050.t2  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X9 a_7333_989.t3 CLK.t2 VDD.t24 VDD.t23 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X10 a_10219_989.t1 SN.t0 VDD.t81 �+���~ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X11 VDD.t131 a_7333_989.t7 a_6371_989.t4 �n�U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X12 VDD.t22 CLK.t3 a_12143_989.t3  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X13 GND a_4447_989.t8 a_18760_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X14 GND a_15991_989.t9 a_18094_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X15 a_13105_989.t5 RN.t4 VDD.t223 VDD.t222 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X16 GND D.t0 a_11635_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X17 VDD.t221 RN.t5 a_277_1050.t6 �+���~ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X18 a_6371_989.t1 a_6049_1050.t7 VDD.t29  '8�U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X19 GND a_6049_1050.t9 a_7787_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X20 VDD.t5 a_7973_1050.t7 a_7333_989.t0  HY�U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X21 VDD.t104 a_9897_1050.t7 a_10219_989.t6 ��$�U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X22 a_17533_1051.t4 a_15991_989.t8 VDD.t16  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X23 a_12143_989.t2 CLK.t7 VDD.t123  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X24 GND a_6371_989.t9 a_9711_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X25 QN a_10219_989.t8 a_18760_101.t0 GND sky130_fd_pr__nfet_01v8 ad=5.373p pd=4.72u as=0p ps=0u w=0u l=0u
X26 a_599_989.t3 a_1561_989.t7 VDD.t129 VDD.t128 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X27 a_15991_989.t6 a_15669_1050.t7 VDD.t231 �+���~ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X28 GND D.t1 a_5863_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X29 VDD.t219 RN.t6 a_1561_989.t6 �f�U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X30 a_9897_1050.t4 a_6371_989.t7 VDD.t189 �?�U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X31 a_4125_1050.t4 a_599_989.t8 VDD.t55 @�d�U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X32 VDD.t63 SN.t2 a_2201_1050.t0 @C6�U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X33 a_4125_1050.t0 a_4447_989.t7 VDD.t18 @`
�U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X34 VDD.t89 a_6371_989.t8 a_6049_1050.t4  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X35 a_18197_1051.t1 a_15991_989.t10 a_17533_1051.t2 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X36 a_1561_989.t1 CLK.t8 VDD.t147 �+���~ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X37 GND a_11821_1050.t8 a_12597_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X38 VDD.t135 a_599_989.t9 a_277_1050.t4 0���U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X39 a_13745_1050.t0 SN.t4 VDD.t133 �l��U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X40 GND a_13745_1050.t8 a_14521_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X41 GND a_9897_1050.t8 a_10673_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X42 a_17533_1051.t6 a_10219_989.t7 VDD.t98 ���U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X43 GND a_7973_1050.t9 a_8749_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X44 a_12143_989.t1 a_11821_1050.t7 VDD.t73  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X45 VDD.t110 a_13745_1050.t7 a_13105_989.t3 �`��U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X46 a_15991_989.t1 SN.t5 VDD.t100  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X47 a_15669_1050.t3 a_12143_989.t8 VDD.t125 VDD.t124 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X48 GND D.t4 a_91_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X49 a_4125_1050.t6 RN.t8 VDD.t217 �+���~ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X50 VDD.t151 a_1561_989.t8 a_2201_1050.t5 @r!�U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X51 VDD.t215 RN.t9 a_6049_1050.t6 �,�U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X52 a_7333_989.t1 a_7973_1050.t8 VDD.t139 �̓�U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X53 a_7973_1050.t6 a_7333_989.t8 VDD.t57 ��!�U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X54 a_9897_1050.t3 a_10219_989.t9 VDD.t176 �Q,�U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X55 VDD.t161 a_13105_989.t10 a_15991_989.t4  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X56 a_1561_989.t3 a_2201_1050.t7 VDD.t173 VDD.t172 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X57 a_18197_1051.t5 a_4447_989.t9 a_17533_1051.t7 �+���~ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X58 VDD.t117 a_4125_1050.t8 a_4447_989.t1 ��+�U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X59 GND a_15991_989.t12 a_17428_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X60 a_6371_989.t6 CLK.t10 VDD.t7 �N��U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X61 VDD.t145 CLK.t11 a_7333_989.t2 �!�U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X62 a_6049_1050.t0 D.t2 VDD.t20 ��+�U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X63 GND a_11821_1050.t10 a_13559_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X64 QN.t4 a_10219_989.t10 a_18197_1051.t7 �x��U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X65 GND a_12143_989.t9 a_15483_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X66 QN a_4447_989.t11 a_18094_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X67 a_277_1050.t0 D.t3 VDD.t96  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X68 VDD.t53 CLK.t12 a_13105_989.t2 VDD.t52 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X69 a_15991_989.t3 a_13105_989.t11 VDD.t159 �+���~ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X70 VDD.t137 a_11821_1050.t9 a_13745_1050.t2 ���U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X71 a_10219_989.t4 a_7333_989.t9 VDD.t9 ����U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X72 VDD.t157 a_13105_989.t12 a_12143_989.t6 ���U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X73 a_15669_1050.t6 RN.t10 VDD.t213 �1B�U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X74 VDD.t171 a_277_1050.t8 a_599_989.t6 �xB�U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X75 a_9897_1050.t5 RN.t11 VDD.t211  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X76 VDD.t209 RN.t13 a_11821_1050.t6 VDD.t208 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X77 VDD.t106 a_1561_989.t9 a_599_989.t1 �+���~ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X78 a_13745_1050.t4 a_13105_989.t13 VDD.t155 �>a�U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X79 VDD.t83 SN.t6 a_4447_989.t3 PA�U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X80 a_18197_1051.t2 a_4447_989.t10 QN.t1 @�-�U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X81 VDD.t119 a_15991_989.t11 a_15669_1050.t2 �&��U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X82 a_6371_989.t3 a_7333_989.t10 VDD.t75 �P��U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X83 GND a_15669_1050.t8 a_16445_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X84 VDD.t207 RN.t15 a_7333_989.t6  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X85 VDD.t178 SN.t7 a_7973_1050.t3 VDD.t177 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X86 a_277_1050.t5 RN.t16 VDD.t203 �+���~ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X87 a_11821_1050.t5 RN.t17 VDD.t205 @,�U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X88 VDD.t185 SN.t8 a_13745_1050.t6  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X89 a_10219_989.t5 a_9897_1050.t9 VDD.t61 VDD.t60 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X90 VDD.t180 CLK.t14 a_599_989.t4  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X91 VDD.t108 a_12143_989.t10 a_11821_1050.t3  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X92 a_1561_989.t5 RN.t18 VDD.t201  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X93 VDD.t127 a_1561_989.t10 a_4447_989.t6  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X94 a_2201_1050.t6 SN.t11 VDD.t165  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X95 GND a_277_1050.t11 a_2015_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X96 VDD.t199 RN.t19 a_4125_1050.t5  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X97 a_12143_989.t5 a_13105_989.t14 VDD.t153  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X98 a_599_989.t2 a_277_1050.t9 VDD.t112  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X99 VDD.t51 a_6049_1050.t10 a_7973_1050.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X100 VDD.t197 RN.t21 a_13105_989.t4  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X101 a_277_1050.t3 a_599_989.t11 VDD.t69  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X102 a_11821_1050.t0 D.t5 VDD.t59  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X103 a_13105_989.t0 a_13745_1050.t9 VDD.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X104 VDD.t229 a_15669_1050.t9 a_15991_989.t5  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X105 a_7973_1050.t0 a_6049_1050.t11 VDD.t85  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X106 VDD.t3 a_6371_989.t10 a_9897_1050.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X107 QN a_10219_989.t12 a_17428_101.t1 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X108 a_2201_1050.t1 a_277_1050.t10 VDD.t47  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X109 VDD.t31 a_7333_989.t11 a_10219_989.t3  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X110 a_2201_1050.t4 a_1561_989.t12 VDD.t43  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X111 VDD.t33 a_599_989.t12 a_4125_1050.t3  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X112 GND a_2201_1050.t8 a_2977_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X113 VDD.t191 a_4447_989.t13 a_4125_1050.t2  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X114 a_6049_1050.t5 RN.t23 VDD.t195  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X115 a_17533_1051.t1 a_15991_989.t13 a_18197_1051.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X116 a_4447_989.t0 a_4125_1050.t9 VDD.t115  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X117 VDD.t27 a_6049_1050.t12 a_6371_989.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X118 GND a_277_1050.t12 a_1053_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X119 a_4447_989.t5 a_1561_989.t15 VDD.t41  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X120 a_15669_1050.t0 a_15991_989.t14 VDD.t65  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X121 VDD.t71 a_11821_1050.t11 a_12143_989.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X122 VDD.t187 a_10219_989.t11 a_17533_1051.t5  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X123 a_13105_989.t1 CLK.t16 VDD.t45  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X124 VDD.t13 SN.t13 a_15991_989.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X125 VDD.t39 SN.t14 a_10219_989.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X126 a_13745_1050.t1 a_11821_1050.t12 VDD.t35  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X127 VDD.t149 a_12143_989.t12 a_15669_1050.t4  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X128 GND a_599_989.t7 a_3939_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X129 a_6049_1050.t3 a_6371_989.t12 VDD.t79  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X130 VDD.t37 a_7333_989.t14 a_7973_1050.t5  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X131 VDD.t11 a_10219_989.t14 a_9897_1050.t2  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X132 VDD.t49 a_2201_1050.t9 a_1561_989.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X133 a_4447_989.t2 SN.t15 VDD.t94  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X134 QN.t0 a_4447_989.t14 a_18197_1051.t3  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X135 a_17533_1051.t0 a_4447_989.t15 a_18197_1051.t4  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X136 VDD.t102 CLK.t17 a_6371_989.t5  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X137 a_7333_989.t5 RN.t25 VDD.t193  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X138 VDD.t121 D.t6 a_6049_1050.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X139 a_7973_1050.t2 SN.t16 VDD.t91  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X140 a_18197_1051.t6 a_10219_989.t15 QN.t3  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X141 VDD.t167 a_15991_989.t15 a_17533_1051.t3  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X142 VDD.t143 D.t7 a_277_1050.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X143 VDD.t141 D.t8 a_11821_1050.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
C0 D RN 2.36fF
C1 CLK VDD 8.69fF
C2 CLK D 12.06fF
C3 CLK RN 1.11fF
C4 SN VDD 1.76fF
C5 QN VDD 0.73fF
C6 SN D 0.31fF
C7 SN RN 16.07fF
C8 VDD D 11.48fF
C9 CLK SN 0.63fF
C10 VDD RN 2.65fF
R0 RN.n23 RN.t5 479.223
R1 RN.n17 RN.t19 479.223
R2 RN.n14 RN.t9 479.223
R3 RN.n8 RN.t2 479.223
R4 RN.n5 RN.t13 479.223
R5 RN.n0 RN.t1 479.223
R6 RN.n20 RN.t18 454.685
R7 RN.n11 RN.t25 454.685
R8 RN.n2 RN.t4 454.685
R9 RN.n20 RN.t6 428.979
R10 RN.n11 RN.t15 428.979
R11 RN.n2 RN.t21 428.979
R12 RN.n23 RN.t16 375.52
R13 RN.n17 RN.t8 375.52
R14 RN.n14 RN.t23 375.52
R15 RN.n8 RN.t11 375.52
R16 RN.n5 RN.t17 375.52
R17 RN.n0 RN.t10 375.52
R18 RN.n21 RN.n20 254.865
R19 RN.n12 RN.n11 254.865
R20 RN.n3 RN.n2 254.865
R21 RN.n24 RN.n23 252.188
R22 RN.n18 RN.n17 252.188
R23 RN.n15 RN.n14 252.188
R24 RN.n9 RN.n8 252.188
R25 RN.n6 RN.n5 252.188
R26 RN.n1 RN.n0 252.188
R27 RN.n24 RN.t20 231.854
R28 RN.n18 RN.t26 231.854
R29 RN.n15 RN.t7 231.854
R30 RN.n9 RN.t14 231.854
R31 RN.n6 RN.t12 231.854
R32 RN.n1 RN.t22 231.854
R33 RN.n21 RN.t24 228.106
R34 RN.n12 RN.t3 228.106
R35 RN.n3 RN.t0 228.106
R36 RN.n7 RN.n4 11.381
R37 RN.n16 RN.n13 11.381
R38 RN.n25 RN.n22 11.381
R39 RN.n4 RN.n1 7.325
R40 RN.n10 RN.n7 7.028
R41 RN.n19 RN.n16 7.028
R42 RN.n4 RN.n3 4.65
R43 RN.n7 RN.n6 4.65
R44 RN.n10 RN.n9 4.65
R45 RN.n13 RN.n12 4.65
R46 RN.n16 RN.n15 4.65
R47 RN.n19 RN.n18 4.65
R48 RN.n22 RN.n21 4.65
R49 RN.n25 RN.n24 4.65
R50 RN.n13 RN.n10 2.675
R51 RN.n22 RN.n19 2.675
R52 RN.n25 RN 0.046
R53 a_14802_210.n12 a_14802_210.n10 171.558
R54 a_14802_210.n7 a_14802_210.n6 117.622
R55 a_14802_210.n5 a_14802_210.n4 92.5
R56 a_14802_210.n9 a_14802_210.n8 92.5
R57 a_14802_210.n10 a_14802_210.t1 75.764
R58 a_14802_210.n5 a_14802_210.n3 65.02
R59 a_14802_210.n13 a_14802_210.n0 49.6
R60 a_14802_210.n7 a_14802_210.n5 36.517
R61 a_14802_210.n3 a_14802_210.n2 35.865
R62 a_14802_210.n12 a_14802_210.n11 27.2
R63 a_14802_210.n13 a_14802_210.n12 22.4
R64 a_14802_210.n9 a_14802_210.n7 19.952
R65 a_14802_210.t1 a_14802_210.n1 7.04
R66 a_14802_210.n10 a_14802_210.n9 1.505
R67 a_13105_989.n7 a_13105_989.t13 454.685
R68 a_13105_989.n9 a_13105_989.t14 454.685
R69 a_13105_989.n5 a_13105_989.t11 454.685
R70 a_13105_989.n7 a_13105_989.t7 428.979
R71 a_13105_989.n9 a_13105_989.t12 428.979
R72 a_13105_989.n5 a_13105_989.t10 428.979
R73 a_13105_989.n15 a_13105_989.n13 342.597
R74 a_13105_989.n8 a_13105_989.t8 339.542
R75 a_13105_989.n6 a_13105_989.t9 339.542
R76 a_13105_989.n10 a_13105_989.t15 339.186
R77 a_13105_989.n3 a_13105_989.n2 161.352
R78 a_13105_989.n13 a_13105_989.n4 151.34
R79 a_13105_989.n8 a_13105_989.n7 143.429
R80 a_13105_989.n6 a_13105_989.n5 143.429
R81 a_13105_989.n10 a_13105_989.n9 143.074
R82 a_13105_989.n4 a_13105_989.n0 95.095
R83 a_13105_989.n3 a_13105_989.n1 95.095
R84 a_13105_989.n4 a_13105_989.n3 66.258
R85 a_13105_989.n15 a_13105_989.n14 15.218
R86 a_13105_989.n0 a_13105_989.t4 14.282
R87 a_13105_989.n0 a_13105_989.t5 14.282
R88 a_13105_989.n1 a_13105_989.t2 14.282
R89 a_13105_989.n1 a_13105_989.t1 14.282
R90 a_13105_989.n2 a_13105_989.t3 14.282
R91 a_13105_989.n2 a_13105_989.t0 14.282
R92 a_13105_989.n16 a_13105_989.n15 12.014
R93 a_13105_989.n12 a_13105_989.n6 11.134
R94 a_13105_989.n11 a_13105_989.n10 8.145
R95 a_13105_989.n11 a_13105_989.n8 4.65
R96 a_13105_989.n13 a_13105_989.n12 4.65
R97 a_13105_989.n12 a_13105_989.n11 4.035
R98 GND.n28 GND.n27 237.558
R99 GND.n473 GND.n472 237.558
R100 GND.n517 GND.n516 237.558
R101 GND.n561 GND.n560 237.558
R102 GND.n605 GND.n604 237.558
R103 GND.n647 GND.n646 237.558
R104 GND.n692 GND.n691 237.558
R105 GND.n737 GND.n736 237.558
R106 GND.n782 GND.n781 237.558
R107 GND.n824 GND.n823 237.558
R108 GND.n390 GND.n389 237.558
R109 GND.n428 GND.n427 237.558
R110 GND.n348 GND.n347 237.558
R111 GND.n304 GND.n303 237.558
R112 GND.n260 GND.n259 237.558
R113 GND.n216 GND.n215 237.558
R114 GND.n174 GND.n173 237.558
R115 GND.n130 GND.n129 237.558
R116 GND.n88 GND.n87 237.558
R117 GND.n58 GND.n57 237.558
R118 GND.n25 GND.n24 210.82
R119 GND.n55 GND.n54 210.82
R120 GND.n475 GND.n474 210.82
R121 GND.n519 GND.n518 210.82
R122 GND.n563 GND.n562 210.82
R123 GND.n607 GND.n606 210.82
R124 GND.n649 GND.n648 210.82
R125 GND.n694 GND.n693 210.82
R126 GND.n739 GND.n738 210.82
R127 GND.n784 GND.n783 210.82
R128 GND.n826 GND.n825 210.82
R129 GND.n430 GND.n429 210.82
R130 GND.n387 GND.n386 210.82
R131 GND.n345 GND.n344 210.82
R132 GND.n301 GND.n300 210.82
R133 GND.n257 GND.n256 210.82
R134 GND.n213 GND.n212 210.82
R135 GND.n171 GND.n170 210.82
R136 GND.n127 GND.n126 210.82
R137 GND.n85 GND.n84 210.82
R138 GND.n117 GND.n116 173.365
R139 GND.n203 GND.n202 173.365
R140 GND.n377 GND.n376 173.365
R141 GND.n793 GND.n792 173.365
R142 GND.n616 GND.n615 173.365
R143 GND.n442 GND.n441 173.365
R144 GND.n44 GND.n43 172.612
R145 GND.n74 GND.n73 172.612
R146 GND.n14 GND.n13 172.612
R147 GND.n161 GND.n160 167.358
R148 GND.n247 GND.n246 167.358
R149 GND.n291 GND.n290 167.358
R150 GND.n335 GND.n334 167.358
R151 GND.n421 GND.n420 167.358
R152 GND.n837 GND.n836 167.358
R153 GND.n574 GND.n573 167.358
R154 GND.n530 GND.n529 167.358
R155 GND.n486 GND.n485 167.358
R156 GND.n751 GND.n750 152.358
R157 GND.n706 GND.n705 152.358
R158 GND.n661 GND.n660 152.358
R159 GND.n750 GND.n749 28.421
R160 GND.n705 GND.n704 28.421
R161 GND.n660 GND.n659 28.421
R162 GND.n750 GND.n748 25.263
R163 GND.n705 GND.n703 25.263
R164 GND.n660 GND.n658 25.263
R165 GND.n748 GND.n747 24.383
R166 GND.n703 GND.n702 24.383
R167 GND.n658 GND.n657 24.383
R168 GND.n160 GND.n158 23.03
R169 GND.n246 GND.n244 23.03
R170 GND.n290 GND.n288 23.03
R171 GND.n334 GND.n332 23.03
R172 GND.n420 GND.n418 23.03
R173 GND.n836 GND.n834 23.03
R174 GND.n573 GND.n571 23.03
R175 GND.n529 GND.n527 23.03
R176 GND.n485 GND.n483 23.03
R177 GND.n26 GND.n25 18.953
R178 GND.n56 GND.n55 18.953
R179 GND.n476 GND.n475 18.953
R180 GND.n520 GND.n519 18.953
R181 GND.n564 GND.n563 18.953
R182 GND.n608 GND.n607 18.953
R183 GND.n650 GND.n649 18.953
R184 GND.n695 GND.n694 18.953
R185 GND.n740 GND.n739 18.953
R186 GND.n785 GND.n784 18.953
R187 GND.n827 GND.n826 18.953
R188 GND.n431 GND.n430 18.953
R189 GND.n388 GND.n387 18.953
R190 GND.n346 GND.n345 18.953
R191 GND.n302 GND.n301 18.953
R192 GND.n258 GND.n257 18.953
R193 GND.n214 GND.n213 18.953
R194 GND.n172 GND.n171 18.953
R195 GND.n128 GND.n127 18.953
R196 GND.n86 GND.n85 18.953
R197 GND.n29 GND.n26 14.864
R198 GND.n59 GND.n56 14.864
R199 GND.n89 GND.n86 14.864
R200 GND.n131 GND.n128 14.864
R201 GND.n175 GND.n172 14.864
R202 GND.n217 GND.n214 14.864
R203 GND.n261 GND.n258 14.864
R204 GND.n305 GND.n302 14.864
R205 GND.n349 GND.n346 14.864
R206 GND.n391 GND.n388 14.864
R207 GND.n432 GND.n431 14.864
R208 GND.n828 GND.n827 14.864
R209 GND.n786 GND.n785 14.864
R210 GND.n741 GND.n740 14.864
R211 GND.n696 GND.n695 14.864
R212 GND.n651 GND.n650 14.864
R213 GND.n609 GND.n608 14.864
R214 GND.n565 GND.n564 14.864
R215 GND.n521 GND.n520 14.864
R216 GND.n477 GND.n476 14.864
R217 GND.n438 GND.n437 9.154
R218 GND.n443 GND.n440 9.154
R219 GND.n446 GND.n445 9.154
R220 GND.n449 GND.n448 9.154
R221 GND.n452 GND.n451 9.154
R222 GND.n455 GND.n454 9.154
R223 GND.n458 GND.n457 9.154
R224 GND.n461 GND.n460 9.154
R225 GND.n464 GND.n463 9.154
R226 GND.n467 GND.n466 9.154
R227 GND.n470 GND.n469 9.154
R228 GND.n477 GND.n473 9.154
R229 GND.n480 GND.n479 9.154
R230 GND.n487 GND.n482 9.154
R231 GND.n490 GND.n489 9.154
R232 GND.n493 GND.n492 9.154
R233 GND.n496 GND.n495 9.154
R234 GND.n499 GND.n498 9.154
R235 GND.n502 GND.n501 9.154
R236 GND.n505 GND.n504 9.154
R237 GND.n508 GND.n507 9.154
R238 GND.n511 GND.n510 9.154
R239 GND.n514 GND.n513 9.154
R240 GND.n521 GND.n517 9.154
R241 GND.n524 GND.n523 9.154
R242 GND.n531 GND.n526 9.154
R243 GND.n534 GND.n533 9.154
R244 GND.n537 GND.n536 9.154
R245 GND.n540 GND.n539 9.154
R246 GND.n543 GND.n542 9.154
R247 GND.n546 GND.n545 9.154
R248 GND.n549 GND.n548 9.154
R249 GND.n552 GND.n551 9.154
R250 GND.n555 GND.n554 9.154
R251 GND.n558 GND.n557 9.154
R252 GND.n565 GND.n561 9.154
R253 GND.n568 GND.n567 9.154
R254 GND.n575 GND.n570 9.154
R255 GND.n578 GND.n577 9.154
R256 GND.n581 GND.n580 9.154
R257 GND.n584 GND.n583 9.154
R258 GND.n587 GND.n586 9.154
R259 GND.n590 GND.n589 9.154
R260 GND.n593 GND.n592 9.154
R261 GND.n596 GND.n595 9.154
R262 GND.n599 GND.n598 9.154
R263 GND.n602 GND.n601 9.154
R264 GND.n609 GND.n605 9.154
R265 GND.n612 GND.n611 9.154
R266 GND.n617 GND.n614 9.154
R267 GND.n620 GND.n619 9.154
R268 GND.n623 GND.n622 9.154
R269 GND.n626 GND.n625 9.154
R270 GND.n629 GND.n628 9.154
R271 GND.n632 GND.n631 9.154
R272 GND.n635 GND.n634 9.154
R273 GND.n638 GND.n637 9.154
R274 GND.n641 GND.n640 9.154
R275 GND.n644 GND.n643 9.154
R276 GND.n651 GND.n647 9.154
R277 GND.n654 GND.n653 9.154
R278 GND.n662 GND.n656 9.154
R279 GND.n665 GND.n664 9.154
R280 GND.n668 GND.n667 9.154
R281 GND.n671 GND.n670 9.154
R282 GND.n674 GND.n673 9.154
R283 GND.n677 GND.n676 9.154
R284 GND.n680 GND.n679 9.154
R285 GND.n683 GND.n682 9.154
R286 GND.n686 GND.n685 9.154
R287 GND.n689 GND.n688 9.154
R288 GND.n696 GND.n692 9.154
R289 GND.n699 GND.n698 9.154
R290 GND.n707 GND.n701 9.154
R291 GND.n710 GND.n709 9.154
R292 GND.n713 GND.n712 9.154
R293 GND.n716 GND.n715 9.154
R294 GND.n719 GND.n718 9.154
R295 GND.n722 GND.n721 9.154
R296 GND.n725 GND.n724 9.154
R297 GND.n728 GND.n727 9.154
R298 GND.n731 GND.n730 9.154
R299 GND.n734 GND.n733 9.154
R300 GND.n741 GND.n737 9.154
R301 GND.n744 GND.n743 9.154
R302 GND.n752 GND.n746 9.154
R303 GND.n755 GND.n754 9.154
R304 GND.n758 GND.n757 9.154
R305 GND.n761 GND.n760 9.154
R306 GND.n764 GND.n763 9.154
R307 GND.n767 GND.n766 9.154
R308 GND.n770 GND.n769 9.154
R309 GND.n773 GND.n772 9.154
R310 GND.n776 GND.n775 9.154
R311 GND.n779 GND.n778 9.154
R312 GND.n786 GND.n782 9.154
R313 GND.n789 GND.n788 9.154
R314 GND.n794 GND.n791 9.154
R315 GND.n797 GND.n796 9.154
R316 GND.n800 GND.n799 9.154
R317 GND.n803 GND.n802 9.154
R318 GND.n806 GND.n805 9.154
R319 GND.n809 GND.n808 9.154
R320 GND.n812 GND.n811 9.154
R321 GND.n815 GND.n814 9.154
R322 GND.n818 GND.n817 9.154
R323 GND.n821 GND.n820 9.154
R324 GND.n828 GND.n824 9.154
R325 GND.n831 GND.n830 9.154
R326 GND.n838 GND.n833 9.154
R327 GND.n841 GND.n840 9.154
R328 GND.n844 GND.n843 9.154
R329 GND.n847 GND.n846 9.154
R330 GND.n850 GND.n849 9.154
R331 GND.n853 GND.n852 9.154
R332 GND.n856 GND.n855 9.154
R333 GND.n859 GND.n858 9.154
R334 GND.n862 GND.n861 9.154
R335 GND.n865 GND.n864 9.154
R336 GND.n432 GND.n428 9.154
R337 GND.n425 GND.n424 9.154
R338 GND.n422 GND.n417 9.154
R339 GND.n415 GND.n414 9.154
R340 GND.n412 GND.n411 9.154
R341 GND.n409 GND.n408 9.154
R342 GND.n406 GND.n405 9.154
R343 GND.n403 GND.n402 9.154
R344 GND.n400 GND.n399 9.154
R345 GND.n397 GND.n396 9.154
R346 GND.n394 GND.n393 9.154
R347 GND.n391 GND.n390 9.154
R348 GND.n384 GND.n383 9.154
R349 GND.n381 GND.n380 9.154
R350 GND.n378 GND.n375 9.154
R351 GND.n373 GND.n372 9.154
R352 GND.n370 GND.n369 9.154
R353 GND.n367 GND.n366 9.154
R354 GND.n364 GND.n363 9.154
R355 GND.n361 GND.n360 9.154
R356 GND.n358 GND.n357 9.154
R357 GND.n355 GND.n354 9.154
R358 GND.n352 GND.n351 9.154
R359 GND.n349 GND.n348 9.154
R360 GND.n342 GND.n341 9.154
R361 GND.n339 GND.n338 9.154
R362 GND.n336 GND.n331 9.154
R363 GND.n329 GND.n328 9.154
R364 GND.n326 GND.n325 9.154
R365 GND.n323 GND.n322 9.154
R366 GND.n320 GND.n319 9.154
R367 GND.n317 GND.n316 9.154
R368 GND.n314 GND.n313 9.154
R369 GND.n311 GND.n310 9.154
R370 GND.n308 GND.n307 9.154
R371 GND.n305 GND.n304 9.154
R372 GND.n298 GND.n297 9.154
R373 GND.n295 GND.n294 9.154
R374 GND.n292 GND.n287 9.154
R375 GND.n285 GND.n284 9.154
R376 GND.n282 GND.n281 9.154
R377 GND.n279 GND.n278 9.154
R378 GND.n276 GND.n275 9.154
R379 GND.n273 GND.n272 9.154
R380 GND.n270 GND.n269 9.154
R381 GND.n267 GND.n266 9.154
R382 GND.n264 GND.n263 9.154
R383 GND.n261 GND.n260 9.154
R384 GND.n254 GND.n253 9.154
R385 GND.n251 GND.n250 9.154
R386 GND.n248 GND.n243 9.154
R387 GND.n241 GND.n240 9.154
R388 GND.n238 GND.n237 9.154
R389 GND.n235 GND.n234 9.154
R390 GND.n232 GND.n231 9.154
R391 GND.n229 GND.n228 9.154
R392 GND.n226 GND.n225 9.154
R393 GND.n223 GND.n222 9.154
R394 GND.n220 GND.n219 9.154
R395 GND.n217 GND.n216 9.154
R396 GND.n210 GND.n209 9.154
R397 GND.n207 GND.n206 9.154
R398 GND.n204 GND.n201 9.154
R399 GND.n199 GND.n198 9.154
R400 GND.n196 GND.n195 9.154
R401 GND.n193 GND.n192 9.154
R402 GND.n190 GND.n189 9.154
R403 GND.n187 GND.n186 9.154
R404 GND.n184 GND.n183 9.154
R405 GND.n181 GND.n180 9.154
R406 GND.n178 GND.n177 9.154
R407 GND.n175 GND.n174 9.154
R408 GND.n168 GND.n167 9.154
R409 GND.n165 GND.n164 9.154
R410 GND.n162 GND.n157 9.154
R411 GND.n155 GND.n154 9.154
R412 GND.n152 GND.n151 9.154
R413 GND.n149 GND.n148 9.154
R414 GND.n146 GND.n145 9.154
R415 GND.n143 GND.n142 9.154
R416 GND.n140 GND.n139 9.154
R417 GND.n137 GND.n136 9.154
R418 GND.n134 GND.n133 9.154
R419 GND.n131 GND.n130 9.154
R420 GND.n124 GND.n123 9.154
R421 GND.n121 GND.n120 9.154
R422 GND.n118 GND.n115 9.154
R423 GND.n113 GND.n112 9.154
R424 GND.n110 GND.n109 9.154
R425 GND.n107 GND.n106 9.154
R426 GND.n104 GND.n103 9.154
R427 GND.n101 GND.n100 9.154
R428 GND.n98 GND.n97 9.154
R429 GND.n95 GND.n94 9.154
R430 GND.n92 GND.n91 9.154
R431 GND.n89 GND.n88 9.154
R432 GND.n82 GND.n81 9.154
R433 GND.n79 GND.n78 9.154
R434 GND.n76 GND.n75 9.154
R435 GND.n71 GND.n70 9.154
R436 GND.n68 GND.n67 9.154
R437 GND.n65 GND.n64 9.154
R438 GND.n62 GND.n61 9.154
R439 GND.n59 GND.n58 9.154
R440 GND.n52 GND.n51 9.154
R441 GND.n49 GND.n48 9.154
R442 GND.n46 GND.n45 9.154
R443 GND.n41 GND.n40 9.154
R444 GND.n38 GND.n37 9.154
R445 GND.n1 GND.n0 9.154
R446 GND.n5 GND.n4 9.154
R447 GND.n8 GND.n7 9.154
R448 GND.n11 GND.n10 9.154
R449 GND.n16 GND.n15 9.154
R450 GND.n19 GND.n18 9.154
R451 GND.n22 GND.n21 9.154
R452 GND.n29 GND.n28 9.154
R453 GND.n32 GND.n31 9.154
R454 GND.n35 GND.n34 9.154
R455 GND.n160 GND.n159 8.128
R456 GND.n246 GND.n245 8.128
R457 GND.n290 GND.n289 8.128
R458 GND.n334 GND.n333 8.128
R459 GND.n420 GND.n419 8.128
R460 GND.n836 GND.n835 8.128
R461 GND.n573 GND.n572 8.128
R462 GND.n529 GND.n528 8.128
R463 GND.n485 GND.n484 8.128
R464 GND.n436 GND.n435 4.65
R465 GND.n39 GND.n38 4.65
R466 GND.n42 GND.n41 4.65
R467 GND.n47 GND.n46 4.65
R468 GND.n50 GND.n49 4.65
R469 GND.n53 GND.n52 4.65
R470 GND.n60 GND.n59 4.65
R471 GND.n63 GND.n62 4.65
R472 GND.n66 GND.n65 4.65
R473 GND.n69 GND.n68 4.65
R474 GND.n72 GND.n71 4.65
R475 GND.n77 GND.n76 4.65
R476 GND.n80 GND.n79 4.65
R477 GND.n83 GND.n82 4.65
R478 GND.n90 GND.n89 4.65
R479 GND.n93 GND.n92 4.65
R480 GND.n96 GND.n95 4.65
R481 GND.n99 GND.n98 4.65
R482 GND.n102 GND.n101 4.65
R483 GND.n105 GND.n104 4.65
R484 GND.n108 GND.n107 4.65
R485 GND.n111 GND.n110 4.65
R486 GND.n114 GND.n113 4.65
R487 GND.n119 GND.n118 4.65
R488 GND.n122 GND.n121 4.65
R489 GND.n125 GND.n124 4.65
R490 GND.n132 GND.n131 4.65
R491 GND.n135 GND.n134 4.65
R492 GND.n138 GND.n137 4.65
R493 GND.n141 GND.n140 4.65
R494 GND.n144 GND.n143 4.65
R495 GND.n147 GND.n146 4.65
R496 GND.n150 GND.n149 4.65
R497 GND.n153 GND.n152 4.65
R498 GND.n156 GND.n155 4.65
R499 GND.n163 GND.n162 4.65
R500 GND.n166 GND.n165 4.65
R501 GND.n169 GND.n168 4.65
R502 GND.n176 GND.n175 4.65
R503 GND.n179 GND.n178 4.65
R504 GND.n182 GND.n181 4.65
R505 GND.n185 GND.n184 4.65
R506 GND.n188 GND.n187 4.65
R507 GND.n191 GND.n190 4.65
R508 GND.n194 GND.n193 4.65
R509 GND.n197 GND.n196 4.65
R510 GND.n200 GND.n199 4.65
R511 GND.n205 GND.n204 4.65
R512 GND.n208 GND.n207 4.65
R513 GND.n211 GND.n210 4.65
R514 GND.n218 GND.n217 4.65
R515 GND.n221 GND.n220 4.65
R516 GND.n224 GND.n223 4.65
R517 GND.n227 GND.n226 4.65
R518 GND.n230 GND.n229 4.65
R519 GND.n233 GND.n232 4.65
R520 GND.n236 GND.n235 4.65
R521 GND.n239 GND.n238 4.65
R522 GND.n242 GND.n241 4.65
R523 GND.n249 GND.n248 4.65
R524 GND.n252 GND.n251 4.65
R525 GND.n255 GND.n254 4.65
R526 GND.n262 GND.n261 4.65
R527 GND.n265 GND.n264 4.65
R528 GND.n268 GND.n267 4.65
R529 GND.n271 GND.n270 4.65
R530 GND.n274 GND.n273 4.65
R531 GND.n277 GND.n276 4.65
R532 GND.n280 GND.n279 4.65
R533 GND.n283 GND.n282 4.65
R534 GND.n286 GND.n285 4.65
R535 GND.n293 GND.n292 4.65
R536 GND.n296 GND.n295 4.65
R537 GND.n299 GND.n298 4.65
R538 GND.n306 GND.n305 4.65
R539 GND.n309 GND.n308 4.65
R540 GND.n312 GND.n311 4.65
R541 GND.n315 GND.n314 4.65
R542 GND.n318 GND.n317 4.65
R543 GND.n321 GND.n320 4.65
R544 GND.n324 GND.n323 4.65
R545 GND.n327 GND.n326 4.65
R546 GND.n330 GND.n329 4.65
R547 GND.n337 GND.n336 4.65
R548 GND.n340 GND.n339 4.65
R549 GND.n343 GND.n342 4.65
R550 GND.n350 GND.n349 4.65
R551 GND.n353 GND.n352 4.65
R552 GND.n356 GND.n355 4.65
R553 GND.n359 GND.n358 4.65
R554 GND.n362 GND.n361 4.65
R555 GND.n365 GND.n364 4.65
R556 GND.n368 GND.n367 4.65
R557 GND.n371 GND.n370 4.65
R558 GND.n374 GND.n373 4.65
R559 GND.n379 GND.n378 4.65
R560 GND.n382 GND.n381 4.65
R561 GND.n385 GND.n384 4.65
R562 GND.n392 GND.n391 4.65
R563 GND.n395 GND.n394 4.65
R564 GND.n398 GND.n397 4.65
R565 GND.n401 GND.n400 4.65
R566 GND.n404 GND.n403 4.65
R567 GND.n407 GND.n406 4.65
R568 GND.n410 GND.n409 4.65
R569 GND.n413 GND.n412 4.65
R570 GND.n416 GND.n415 4.65
R571 GND.n423 GND.n422 4.65
R572 GND.n426 GND.n425 4.65
R573 GND.n433 GND.n432 4.65
R574 GND.n866 GND.n865 4.65
R575 GND.n863 GND.n862 4.65
R576 GND.n860 GND.n859 4.65
R577 GND.n857 GND.n856 4.65
R578 GND.n854 GND.n853 4.65
R579 GND.n851 GND.n850 4.65
R580 GND.n848 GND.n847 4.65
R581 GND.n845 GND.n844 4.65
R582 GND.n842 GND.n841 4.65
R583 GND.n839 GND.n838 4.65
R584 GND.n832 GND.n831 4.65
R585 GND.n829 GND.n828 4.65
R586 GND.n822 GND.n821 4.65
R587 GND.n819 GND.n818 4.65
R588 GND.n816 GND.n815 4.65
R589 GND.n813 GND.n812 4.65
R590 GND.n810 GND.n809 4.65
R591 GND.n807 GND.n806 4.65
R592 GND.n804 GND.n803 4.65
R593 GND.n801 GND.n800 4.65
R594 GND.n798 GND.n797 4.65
R595 GND.n795 GND.n794 4.65
R596 GND.n790 GND.n789 4.65
R597 GND.n787 GND.n786 4.65
R598 GND.n780 GND.n779 4.65
R599 GND.n777 GND.n776 4.65
R600 GND.n774 GND.n773 4.65
R601 GND.n771 GND.n770 4.65
R602 GND.n768 GND.n767 4.65
R603 GND.n765 GND.n764 4.65
R604 GND.n762 GND.n761 4.65
R605 GND.n759 GND.n758 4.65
R606 GND.n756 GND.n755 4.65
R607 GND.n753 GND.n752 4.65
R608 GND.n745 GND.n744 4.65
R609 GND.n742 GND.n741 4.65
R610 GND.n735 GND.n734 4.65
R611 GND.n732 GND.n731 4.65
R612 GND.n729 GND.n728 4.65
R613 GND.n726 GND.n725 4.65
R614 GND.n723 GND.n722 4.65
R615 GND.n720 GND.n719 4.65
R616 GND.n717 GND.n716 4.65
R617 GND.n714 GND.n713 4.65
R618 GND.n711 GND.n710 4.65
R619 GND.n708 GND.n707 4.65
R620 GND.n700 GND.n699 4.65
R621 GND.n697 GND.n696 4.65
R622 GND.n690 GND.n689 4.65
R623 GND.n687 GND.n686 4.65
R624 GND.n684 GND.n683 4.65
R625 GND.n681 GND.n680 4.65
R626 GND.n678 GND.n677 4.65
R627 GND.n675 GND.n674 4.65
R628 GND.n672 GND.n671 4.65
R629 GND.n669 GND.n668 4.65
R630 GND.n666 GND.n665 4.65
R631 GND.n663 GND.n662 4.65
R632 GND.n655 GND.n654 4.65
R633 GND.n652 GND.n651 4.65
R634 GND.n645 GND.n644 4.65
R635 GND.n642 GND.n641 4.65
R636 GND.n639 GND.n638 4.65
R637 GND.n636 GND.n635 4.65
R638 GND.n633 GND.n632 4.65
R639 GND.n630 GND.n629 4.65
R640 GND.n627 GND.n626 4.65
R641 GND.n624 GND.n623 4.65
R642 GND.n621 GND.n620 4.65
R643 GND.n618 GND.n617 4.65
R644 GND.n613 GND.n612 4.65
R645 GND.n610 GND.n609 4.65
R646 GND.n603 GND.n602 4.65
R647 GND.n600 GND.n599 4.65
R648 GND.n597 GND.n596 4.65
R649 GND.n594 GND.n593 4.65
R650 GND.n591 GND.n590 4.65
R651 GND.n588 GND.n587 4.65
R652 GND.n585 GND.n584 4.65
R653 GND.n582 GND.n581 4.65
R654 GND.n579 GND.n578 4.65
R655 GND.n576 GND.n575 4.65
R656 GND.n569 GND.n568 4.65
R657 GND.n566 GND.n565 4.65
R658 GND.n559 GND.n558 4.65
R659 GND.n556 GND.n555 4.65
R660 GND.n553 GND.n552 4.65
R661 GND.n550 GND.n549 4.65
R662 GND.n547 GND.n546 4.65
R663 GND.n544 GND.n543 4.65
R664 GND.n541 GND.n540 4.65
R665 GND.n538 GND.n537 4.65
R666 GND.n535 GND.n534 4.65
R667 GND.n532 GND.n531 4.65
R668 GND.n525 GND.n524 4.65
R669 GND.n522 GND.n521 4.65
R670 GND.n515 GND.n514 4.65
R671 GND.n512 GND.n511 4.65
R672 GND.n509 GND.n508 4.65
R673 GND.n506 GND.n505 4.65
R674 GND.n503 GND.n502 4.65
R675 GND.n500 GND.n499 4.65
R676 GND.n497 GND.n496 4.65
R677 GND.n494 GND.n493 4.65
R678 GND.n491 GND.n490 4.65
R679 GND.n488 GND.n487 4.65
R680 GND.n481 GND.n480 4.65
R681 GND.n478 GND.n477 4.65
R682 GND.n471 GND.n470 4.65
R683 GND.n468 GND.n467 4.65
R684 GND.n465 GND.n464 4.65
R685 GND.n462 GND.n461 4.65
R686 GND.n459 GND.n458 4.65
R687 GND.n456 GND.n455 4.65
R688 GND.n453 GND.n452 4.65
R689 GND.n450 GND.n449 4.65
R690 GND.n447 GND.n446 4.65
R691 GND.n444 GND.n443 4.65
R692 GND.n439 GND.n438 4.65
R693 GND.n6 GND.n5 4.65
R694 GND.n9 GND.n8 4.65
R695 GND.n12 GND.n11 4.65
R696 GND.n17 GND.n16 4.65
R697 GND.n20 GND.n19 4.65
R698 GND.n23 GND.n22 4.65
R699 GND.n30 GND.n29 4.65
R700 GND.n33 GND.n32 4.65
R701 GND.n36 GND.n35 4.65
R702 GND.n16 GND.n14 4.129
R703 GND.n46 GND.n44 4.129
R704 GND.n76 GND.n74 4.129
R705 GND.n3 GND.n2 3.408
R706 GND.n3 GND.n1 2.844
R707 GND.n6 GND.n3 1.063
R708 GND.n435 GND.n434 0.474
R709 GND.n30 GND.n23 0.29
R710 GND.n60 GND.n53 0.29
R711 GND.n90 GND.n83 0.29
R712 GND.n132 GND.n125 0.29
R713 GND.n176 GND.n169 0.29
R714 GND.n218 GND.n211 0.29
R715 GND.n262 GND.n255 0.29
R716 GND.n306 GND.n299 0.29
R717 GND.n350 GND.n343 0.29
R718 GND.n392 GND.n385 0.29
R719 GND.n829 GND.n822 0.29
R720 GND.n787 GND.n780 0.29
R721 GND.n742 GND.n735 0.29
R722 GND.n697 GND.n690 0.29
R723 GND.n652 GND.n645 0.29
R724 GND.n610 GND.n603 0.29
R725 GND.n566 GND.n559 0.29
R726 GND.n522 GND.n515 0.29
R727 GND.n478 GND.n471 0.29
R728 GND GND.n866 0.219
R729 GND.n436 GND 0.207
R730 GND.n118 GND.n117 0.206
R731 GND.n162 GND.n161 0.206
R732 GND.n204 GND.n203 0.206
R733 GND.n248 GND.n247 0.206
R734 GND.n292 GND.n291 0.206
R735 GND.n336 GND.n335 0.206
R736 GND.n378 GND.n377 0.206
R737 GND.n422 GND.n421 0.206
R738 GND.n838 GND.n837 0.206
R739 GND.n794 GND.n793 0.206
R740 GND.n752 GND.n751 0.206
R741 GND.n707 GND.n706 0.206
R742 GND.n662 GND.n661 0.206
R743 GND.n617 GND.n616 0.206
R744 GND.n575 GND.n574 0.206
R745 GND.n531 GND.n530 0.206
R746 GND.n487 GND.n486 0.206
R747 GND.n443 GND.n442 0.206
R748 GND.n108 GND.n105 0.197
R749 GND.n150 GND.n147 0.197
R750 GND.n194 GND.n191 0.197
R751 GND.n236 GND.n233 0.197
R752 GND.n280 GND.n277 0.197
R753 GND.n324 GND.n321 0.197
R754 GND.n368 GND.n365 0.197
R755 GND.n410 GND.n407 0.197
R756 GND.n851 GND.n848 0.197
R757 GND.n807 GND.n804 0.197
R758 GND.n765 GND.n762 0.197
R759 GND.n720 GND.n717 0.197
R760 GND.n675 GND.n672 0.197
R761 GND.n630 GND.n627 0.197
R762 GND.n588 GND.n585 0.197
R763 GND.n544 GND.n541 0.197
R764 GND.n500 GND.n497 0.197
R765 GND.n456 GND.n453 0.197
R766 GND.n12 GND.n9 0.181
R767 GND.n42 GND.n39 0.181
R768 GND.n72 GND.n69 0.181
R769 GND.n9 GND.n6 0.145
R770 GND.n17 GND.n12 0.145
R771 GND.n20 GND.n17 0.145
R772 GND.n23 GND.n20 0.145
R773 GND.n33 GND.n30 0.145
R774 GND.n36 GND.n33 0.145
R775 GND.n39 GND.n36 0.145
R776 GND.n47 GND.n42 0.145
R777 GND.n50 GND.n47 0.145
R778 GND.n53 GND.n50 0.145
R779 GND.n63 GND.n60 0.145
R780 GND.n66 GND.n63 0.145
R781 GND.n69 GND.n66 0.145
R782 GND.n77 GND.n72 0.145
R783 GND.n80 GND.n77 0.145
R784 GND.n83 GND.n80 0.145
R785 GND.n93 GND.n90 0.145
R786 GND.n96 GND.n93 0.145
R787 GND.n99 GND.n96 0.145
R788 GND.n102 GND.n99 0.145
R789 GND.n105 GND.n102 0.145
R790 GND.n111 GND.n108 0.145
R791 GND.n114 GND.n111 0.145
R792 GND.n119 GND.n114 0.145
R793 GND.n122 GND.n119 0.145
R794 GND.n125 GND.n122 0.145
R795 GND.n135 GND.n132 0.145
R796 GND.n138 GND.n135 0.145
R797 GND.n141 GND.n138 0.145
R798 GND.n144 GND.n141 0.145
R799 GND.n147 GND.n144 0.145
R800 GND.n153 GND.n150 0.145
R801 GND.n156 GND.n153 0.145
R802 GND.n163 GND.n156 0.145
R803 GND.n166 GND.n163 0.145
R804 GND.n169 GND.n166 0.145
R805 GND.n179 GND.n176 0.145
R806 GND.n182 GND.n179 0.145
R807 GND.n185 GND.n182 0.145
R808 GND.n188 GND.n185 0.145
R809 GND.n191 GND.n188 0.145
R810 GND.n197 GND.n194 0.145
R811 GND.n200 GND.n197 0.145
R812 GND.n205 GND.n200 0.145
R813 GND.n208 GND.n205 0.145
R814 GND.n211 GND.n208 0.145
R815 GND.n221 GND.n218 0.145
R816 GND.n224 GND.n221 0.145
R817 GND.n227 GND.n224 0.145
R818 GND.n230 GND.n227 0.145
R819 GND.n233 GND.n230 0.145
R820 GND.n239 GND.n236 0.145
R821 GND.n242 GND.n239 0.145
R822 GND.n249 GND.n242 0.145
R823 GND.n252 GND.n249 0.145
R824 GND.n255 GND.n252 0.145
R825 GND.n265 GND.n262 0.145
R826 GND.n268 GND.n265 0.145
R827 GND.n271 GND.n268 0.145
R828 GND.n274 GND.n271 0.145
R829 GND.n277 GND.n274 0.145
R830 GND.n283 GND.n280 0.145
R831 GND.n286 GND.n283 0.145
R832 GND.n293 GND.n286 0.145
R833 GND.n296 GND.n293 0.145
R834 GND.n299 GND.n296 0.145
R835 GND.n309 GND.n306 0.145
R836 GND.n312 GND.n309 0.145
R837 GND.n315 GND.n312 0.145
R838 GND.n318 GND.n315 0.145
R839 GND.n321 GND.n318 0.145
R840 GND.n327 GND.n324 0.145
R841 GND.n330 GND.n327 0.145
R842 GND.n337 GND.n330 0.145
R843 GND.n340 GND.n337 0.145
R844 GND.n343 GND.n340 0.145
R845 GND.n353 GND.n350 0.145
R846 GND.n356 GND.n353 0.145
R847 GND.n359 GND.n356 0.145
R848 GND.n362 GND.n359 0.145
R849 GND.n365 GND.n362 0.145
R850 GND.n371 GND.n368 0.145
R851 GND.n374 GND.n371 0.145
R852 GND.n379 GND.n374 0.145
R853 GND.n382 GND.n379 0.145
R854 GND.n385 GND.n382 0.145
R855 GND.n395 GND.n392 0.145
R856 GND.n398 GND.n395 0.145
R857 GND.n401 GND.n398 0.145
R858 GND.n404 GND.n401 0.145
R859 GND.n407 GND.n404 0.145
R860 GND.n413 GND.n410 0.145
R861 GND.n416 GND.n413 0.145
R862 GND.n423 GND.n416 0.145
R863 GND.n426 GND.n423 0.145
R864 GND.n433 GND.n426 0.145
R865 GND.n866 GND.n863 0.145
R866 GND.n863 GND.n860 0.145
R867 GND.n860 GND.n857 0.145
R868 GND.n857 GND.n854 0.145
R869 GND.n854 GND.n851 0.145
R870 GND.n848 GND.n845 0.145
R871 GND.n845 GND.n842 0.145
R872 GND.n842 GND.n839 0.145
R873 GND.n839 GND.n832 0.145
R874 GND.n832 GND.n829 0.145
R875 GND.n822 GND.n819 0.145
R876 GND.n819 GND.n816 0.145
R877 GND.n816 GND.n813 0.145
R878 GND.n813 GND.n810 0.145
R879 GND.n810 GND.n807 0.145
R880 GND.n804 GND.n801 0.145
R881 GND.n801 GND.n798 0.145
R882 GND.n798 GND.n795 0.145
R883 GND.n795 GND.n790 0.145
R884 GND.n790 GND.n787 0.145
R885 GND.n780 GND.n777 0.145
R886 GND.n777 GND.n774 0.145
R887 GND.n774 GND.n771 0.145
R888 GND.n771 GND.n768 0.145
R889 GND.n768 GND.n765 0.145
R890 GND.n762 GND.n759 0.145
R891 GND.n759 GND.n756 0.145
R892 GND.n756 GND.n753 0.145
R893 GND.n753 GND.n745 0.145
R894 GND.n745 GND.n742 0.145
R895 GND.n735 GND.n732 0.145
R896 GND.n732 GND.n729 0.145
R897 GND.n729 GND.n726 0.145
R898 GND.n726 GND.n723 0.145
R899 GND.n723 GND.n720 0.145
R900 GND.n717 GND.n714 0.145
R901 GND.n714 GND.n711 0.145
R902 GND.n711 GND.n708 0.145
R903 GND.n708 GND.n700 0.145
R904 GND.n700 GND.n697 0.145
R905 GND.n690 GND.n687 0.145
R906 GND.n687 GND.n684 0.145
R907 GND.n684 GND.n681 0.145
R908 GND.n681 GND.n678 0.145
R909 GND.n678 GND.n675 0.145
R910 GND.n672 GND.n669 0.145
R911 GND.n669 GND.n666 0.145
R912 GND.n666 GND.n663 0.145
R913 GND.n663 GND.n655 0.145
R914 GND.n655 GND.n652 0.145
R915 GND.n645 GND.n642 0.145
R916 GND.n642 GND.n639 0.145
R917 GND.n639 GND.n636 0.145
R918 GND.n636 GND.n633 0.145
R919 GND.n633 GND.n630 0.145
R920 GND.n627 GND.n624 0.145
R921 GND.n624 GND.n621 0.145
R922 GND.n621 GND.n618 0.145
R923 GND.n618 GND.n613 0.145
R924 GND.n613 GND.n610 0.145
R925 GND.n603 GND.n600 0.145
R926 GND.n600 GND.n597 0.145
R927 GND.n597 GND.n594 0.145
R928 GND.n594 GND.n591 0.145
R929 GND.n591 GND.n588 0.145
R930 GND.n585 GND.n582 0.145
R931 GND.n582 GND.n579 0.145
R932 GND.n579 GND.n576 0.145
R933 GND.n576 GND.n569 0.145
R934 GND.n569 GND.n566 0.145
R935 GND.n559 GND.n556 0.145
R936 GND.n556 GND.n553 0.145
R937 GND.n553 GND.n550 0.145
R938 GND.n550 GND.n547 0.145
R939 GND.n547 GND.n544 0.145
R940 GND.n541 GND.n538 0.145
R941 GND.n538 GND.n535 0.145
R942 GND.n535 GND.n532 0.145
R943 GND.n532 GND.n525 0.145
R944 GND.n525 GND.n522 0.145
R945 GND.n515 GND.n512 0.145
R946 GND.n512 GND.n509 0.145
R947 GND.n509 GND.n506 0.145
R948 GND.n506 GND.n503 0.145
R949 GND.n503 GND.n500 0.145
R950 GND.n497 GND.n494 0.145
R951 GND.n494 GND.n491 0.145
R952 GND.n491 GND.n488 0.145
R953 GND.n488 GND.n481 0.145
R954 GND.n481 GND.n478 0.145
R955 GND.n471 GND.n468 0.145
R956 GND.n468 GND.n465 0.145
R957 GND.n465 GND.n462 0.145
R958 GND.n462 GND.n459 0.145
R959 GND.n459 GND.n456 0.145
R960 GND.n453 GND.n450 0.145
R961 GND.n450 GND.n447 0.145
R962 GND.n447 GND.n444 0.145
R963 GND.n444 GND.n439 0.145
R964 GND.n439 GND.n436 0.145
R965 GND GND.n433 0.07
R966 a_15669_1050.n5 a_15669_1050.t9 512.525
R967 a_15669_1050.n5 a_15669_1050.t7 371.139
R968 a_15669_1050.n6 a_15669_1050.t8 361.392
R969 a_15669_1050.n9 a_15669_1050.n7 314.738
R970 a_15669_1050.n6 a_15669_1050.n5 235.554
R971 a_15669_1050.n7 a_15669_1050.n4 179.199
R972 a_15669_1050.n3 a_15669_1050.n2 161.352
R973 a_15669_1050.n4 a_15669_1050.n0 95.095
R974 a_15669_1050.n3 a_15669_1050.n1 95.095
R975 a_15669_1050.n4 a_15669_1050.n3 66.258
R976 a_15669_1050.n9 a_15669_1050.n8 15.218
R977 a_15669_1050.n0 a_15669_1050.t2 14.282
R978 a_15669_1050.n0 a_15669_1050.t0 14.282
R979 a_15669_1050.n1 a_15669_1050.t5 14.282
R980 a_15669_1050.n1 a_15669_1050.t6 14.282
R981 a_15669_1050.n2 a_15669_1050.t4 14.282
R982 a_15669_1050.n2 a_15669_1050.t3 14.282
R983 a_15669_1050.n10 a_15669_1050.n9 12.014
R984 a_15669_1050.n7 a_15669_1050.n6 10.615
R985 VDD.n880 VDD.n869 144.705
R986 VDD.n955 VDD.n948 144.705
R987 VDD.n1030 VDD.n1023 144.705
R988 VDD.n1105 VDD.n1098 144.705
R989 VDD.n1180 VDD.n1173 144.705
R990 VDD.n1255 VDD.n1248 144.705
R991 VDD.n1330 VDD.n1323 144.705
R992 VDD.n1405 VDD.n1398 144.705
R993 VDD.n1480 VDD.n1473 144.705
R994 VDD.n710 VDD.n703 144.705
R995 VDD.n781 VDD.n774 144.705
R996 VDD.n635 VDD.n628 144.705
R997 VDD.n560 VDD.n553 144.705
R998 VDD.n485 VDD.n478 144.705
R999 VDD.n410 VDD.n403 144.705
R1000 VDD.n335 VDD.n328 144.705
R1001 VDD.n260 VDD.n253 144.705
R1002 VDD.n185 VDD.n178 144.705
R1003 VDD.n128 VDD.n121 144.705
R1004 VDD.n75 VDD.n64 144.705
R1005 VDD.n846 VDD.t135 143.754
R1006 VDD.n922 VDD.t106 143.754
R1007 VDD.n997 VDD.t151 143.754
R1008 VDD.n1072 VDD.t219 143.754
R1009 VDD.n1147 VDD.t191 143.754
R1010 VDD.n1222 VDD.t127 143.754
R1011 VDD.n1297 VDD.t89 143.754
R1012 VDD.n1372 VDD.t131 143.754
R1013 VDD.n1447 VDD.t37 143.754
R1014 VDD.n1522 VDD.t207 143.754
R1015 VDD.n719 VDD.t11 143.754
R1016 VDD.n644 VDD.t31 143.754
R1017 VDD.n569 VDD.t108 143.754
R1018 VDD.n494 VDD.t157 143.754
R1019 VDD.n419 VDD.t163 143.754
R1020 VDD.n344 VDD.t197 143.754
R1021 VDD.n269 VDD.t119 143.754
R1022 VDD.n194 VDD.t161 143.754
R1023 VDD.n153 VDD.t16 135.539
R1024 VDD.n131 VDD.t187 135.539
R1025 VDD.n811 VDD.t96 135.17
R1026 VDD.n887 VDD.t112 135.17
R1027 VDD.n962 VDD.t47 135.17
R1028 VDD.n1037 VDD.t173 135.17
R1029 VDD.n1112 VDD.t55 135.17
R1030 VDD.n1187 VDD.t115 135.17
R1031 VDD.n1262 VDD.t20 135.17
R1032 VDD.n1337 VDD.t29 135.17
R1033 VDD.n1412 VDD.t85 135.17
R1034 VDD.n1487 VDD.t139 135.17
R1035 VDD.n749 VDD.t189 135.17
R1036 VDD.n674 VDD.t61 135.17
R1037 VDD.n599 VDD.t59 135.17
R1038 VDD.n524 VDD.t73 135.17
R1039 VDD.n449 VDD.t35 135.17
R1040 VDD.n374 VDD.t1 135.17
R1041 VDD.n299 VDD.t125 135.17
R1042 VDD.n224 VDD.t231 135.17
R1043 VDD.n141 VDD.n140 129.849
R1044 VDD.n821 VDD.n820 129.472
R1045 VDD.n837 VDD.n836 129.472
R1046 VDD.n897 VDD.n896 129.472
R1047 VDD.n913 VDD.n912 129.472
R1048 VDD.n972 VDD.n971 129.472
R1049 VDD.n988 VDD.n987 129.472
R1050 VDD.n1047 VDD.n1046 129.472
R1051 VDD.n1063 VDD.n1062 129.472
R1052 VDD.n1122 VDD.n1121 129.472
R1053 VDD.n1138 VDD.n1137 129.472
R1054 VDD.n1197 VDD.n1196 129.472
R1055 VDD.n1213 VDD.n1212 129.472
R1056 VDD.n1272 VDD.n1271 129.472
R1057 VDD.n1288 VDD.n1287 129.472
R1058 VDD.n1347 VDD.n1346 129.472
R1059 VDD.n1363 VDD.n1362 129.472
R1060 VDD.n1422 VDD.n1421 129.472
R1061 VDD.n1438 VDD.n1437 129.472
R1062 VDD.n1497 VDD.n1496 129.472
R1063 VDD.n1513 VDD.n1512 129.472
R1064 VDD.n740 VDD.n739 129.472
R1065 VDD.n728 VDD.n727 129.472
R1066 VDD.n665 VDD.n664 129.472
R1067 VDD.n653 VDD.n652 129.472
R1068 VDD.n590 VDD.n589 129.472
R1069 VDD.n578 VDD.n577 129.472
R1070 VDD.n515 VDD.n514 129.472
R1071 VDD.n503 VDD.n502 129.472
R1072 VDD.n440 VDD.n439 129.472
R1073 VDD.n428 VDD.n427 129.472
R1074 VDD.n365 VDD.n364 129.472
R1075 VDD.n353 VDD.n352 129.472
R1076 VDD.n290 VDD.n289 129.472
R1077 VDD.n278 VDD.n277 129.472
R1078 VDD.n215 VDD.n214 129.472
R1079 VDD.n203 VDD.n202 129.472
R1080 VDD.n60 VDD.n59 92.5
R1081 VDD.n58 VDD.n57 92.5
R1082 VDD.n56 VDD.n55 92.5
R1083 VDD.n54 VDD.n53 92.5
R1084 VDD.n62 VDD.n61 92.5
R1085 VDD.n117 VDD.n116 92.5
R1086 VDD.n115 VDD.n114 92.5
R1087 VDD.n113 VDD.n112 92.5
R1088 VDD.n111 VDD.n110 92.5
R1089 VDD.n119 VDD.n118 92.5
R1090 VDD.n174 VDD.n173 92.5
R1091 VDD.n172 VDD.n171 92.5
R1092 VDD.n170 VDD.n169 92.5
R1093 VDD.n168 VDD.n167 92.5
R1094 VDD.n176 VDD.n175 92.5
R1095 VDD.n249 VDD.n248 92.5
R1096 VDD.n247 VDD.n246 92.5
R1097 VDD.n245 VDD.n244 92.5
R1098 VDD.n243 VDD.n242 92.5
R1099 VDD.n251 VDD.n250 92.5
R1100 VDD.n324 VDD.n323 92.5
R1101 VDD.n322 VDD.n321 92.5
R1102 VDD.n320 VDD.n319 92.5
R1103 VDD.n318 VDD.n317 92.5
R1104 VDD.n326 VDD.n325 92.5
R1105 VDD.n399 VDD.n398 92.5
R1106 VDD.n397 VDD.n396 92.5
R1107 VDD.n395 VDD.n394 92.5
R1108 VDD.n393 VDD.n392 92.5
R1109 VDD.n401 VDD.n400 92.5
R1110 VDD.n474 VDD.n473 92.5
R1111 VDD.n472 VDD.n471 92.5
R1112 VDD.n470 VDD.n469 92.5
R1113 VDD.n468 VDD.n467 92.5
R1114 VDD.n476 VDD.n475 92.5
R1115 VDD.n549 VDD.n548 92.5
R1116 VDD.n547 VDD.n546 92.5
R1117 VDD.n545 VDD.n544 92.5
R1118 VDD.n543 VDD.n542 92.5
R1119 VDD.n551 VDD.n550 92.5
R1120 VDD.n624 VDD.n623 92.5
R1121 VDD.n622 VDD.n621 92.5
R1122 VDD.n620 VDD.n619 92.5
R1123 VDD.n618 VDD.n617 92.5
R1124 VDD.n626 VDD.n625 92.5
R1125 VDD.n699 VDD.n698 92.5
R1126 VDD.n697 VDD.n696 92.5
R1127 VDD.n695 VDD.n694 92.5
R1128 VDD.n693 VDD.n692 92.5
R1129 VDD.n701 VDD.n700 92.5
R1130 VDD.n770 VDD.n769 92.5
R1131 VDD.n768 VDD.n767 92.5
R1132 VDD.n766 VDD.n765 92.5
R1133 VDD.n764 VDD.n763 92.5
R1134 VDD.n772 VDD.n771 92.5
R1135 VDD.n1469 VDD.n1468 92.5
R1136 VDD.n1467 VDD.n1466 92.5
R1137 VDD.n1465 VDD.n1464 92.5
R1138 VDD.n1463 VDD.n1462 92.5
R1139 VDD.n1471 VDD.n1470 92.5
R1140 VDD.n1394 VDD.n1393 92.5
R1141 VDD.n1392 VDD.n1391 92.5
R1142 VDD.n1390 VDD.n1389 92.5
R1143 VDD.n1388 VDD.n1387 92.5
R1144 VDD.n1396 VDD.n1395 92.5
R1145 VDD.n1319 VDD.n1318 92.5
R1146 VDD.n1317 VDD.n1316 92.5
R1147 VDD.n1315 VDD.n1314 92.5
R1148 VDD.n1313 VDD.n1312 92.5
R1149 VDD.n1321 VDD.n1320 92.5
R1150 VDD.n1244 VDD.n1243 92.5
R1151 VDD.n1242 VDD.n1241 92.5
R1152 VDD.n1240 VDD.n1239 92.5
R1153 VDD.n1238 VDD.n1237 92.5
R1154 VDD.n1246 VDD.n1245 92.5
R1155 VDD.n1169 VDD.n1168 92.5
R1156 VDD.n1167 VDD.n1166 92.5
R1157 VDD.n1165 VDD.n1164 92.5
R1158 VDD.n1163 VDD.n1162 92.5
R1159 VDD.n1171 VDD.n1170 92.5
R1160 VDD.n1094 VDD.n1093 92.5
R1161 VDD.n1092 VDD.n1091 92.5
R1162 VDD.n1090 VDD.n1089 92.5
R1163 VDD.n1088 VDD.n1087 92.5
R1164 VDD.n1096 VDD.n1095 92.5
R1165 VDD.n1019 VDD.n1018 92.5
R1166 VDD.n1017 VDD.n1016 92.5
R1167 VDD.n1015 VDD.n1014 92.5
R1168 VDD.n1013 VDD.n1012 92.5
R1169 VDD.n1021 VDD.n1020 92.5
R1170 VDD.n944 VDD.n943 92.5
R1171 VDD.n942 VDD.n941 92.5
R1172 VDD.n940 VDD.n939 92.5
R1173 VDD.n938 VDD.n937 92.5
R1174 VDD.n946 VDD.n945 92.5
R1175 VDD.n865 VDD.n864 92.5
R1176 VDD.n863 VDD.n862 92.5
R1177 VDD.n861 VDD.n860 92.5
R1178 VDD.n859 VDD.n858 92.5
R1179 VDD.n867 VDD.n866 92.5
R1180 VDD.n795 VDD.n794 92.5
R1181 VDD.n793 VDD.n792 92.5
R1182 VDD.n791 VDD.n790 92.5
R1183 VDD.n789 VDD.n788 92.5
R1184 VDD.n797 VDD.n796 92.5
R1185 VDD.n14 VDD.n1 92.5
R1186 VDD.n5 VDD.n4 92.5
R1187 VDD.n7 VDD.n6 92.5
R1188 VDD.n9 VDD.n8 92.5
R1189 VDD.n11 VDD.n10 92.5
R1190 VDD.n13 VDD.n12 92.5
R1191 VDD.n21 VDD.n20 92.059
R1192 VDD.n74 VDD.n73 92.059
R1193 VDD.n127 VDD.n126 92.059
R1194 VDD.n184 VDD.n183 92.059
R1195 VDD.n259 VDD.n258 92.059
R1196 VDD.n334 VDD.n333 92.059
R1197 VDD.n409 VDD.n408 92.059
R1198 VDD.n484 VDD.n483 92.059
R1199 VDD.n559 VDD.n558 92.059
R1200 VDD.n634 VDD.n633 92.059
R1201 VDD.n709 VDD.n708 92.059
R1202 VDD.n780 VDD.n779 92.059
R1203 VDD.n1479 VDD.n1478 92.059
R1204 VDD.n1404 VDD.n1403 92.059
R1205 VDD.n1329 VDD.n1328 92.059
R1206 VDD.n1254 VDD.n1253 92.059
R1207 VDD.n1179 VDD.n1178 92.059
R1208 VDD.n1104 VDD.n1103 92.059
R1209 VDD.n1029 VDD.n1028 92.059
R1210 VDD.n954 VDD.n953 92.059
R1211 VDD.n879 VDD.n878 92.059
R1212 VDD.n803 VDD.n802 92.059
R1213 VDD.n20 VDD.n16 67.194
R1214 VDD.n20 VDD.n17 67.194
R1215 VDD.n20 VDD.n18 67.194
R1216 VDD.n20 VDD.n19 67.194
R1217 VDD.n787 VDD.n786 44.141
R1218 VDD.n936 VDD.n935 44.141
R1219 VDD.n1011 VDD.n1010 44.141
R1220 VDD.n1086 VDD.n1085 44.141
R1221 VDD.n1161 VDD.n1160 44.141
R1222 VDD.n1236 VDD.n1235 44.141
R1223 VDD.n1311 VDD.n1310 44.141
R1224 VDD.n1386 VDD.n1385 44.141
R1225 VDD.n1461 VDD.n1460 44.141
R1226 VDD.n762 VDD.n761 44.141
R1227 VDD.n691 VDD.n690 44.141
R1228 VDD.n616 VDD.n615 44.141
R1229 VDD.n541 VDD.n540 44.141
R1230 VDD.n466 VDD.n465 44.141
R1231 VDD.n391 VDD.n390 44.141
R1232 VDD.n316 VDD.n315 44.141
R1233 VDD.n241 VDD.n240 44.141
R1234 VDD.n166 VDD.n165 44.141
R1235 VDD.n109 VDD.n108 44.141
R1236 VDD.n5 VDD.n3 44.141
R1237 VDD.n935 VDD.n933 44.107
R1238 VDD.n1010 VDD.n1008 44.107
R1239 VDD.n1085 VDD.n1083 44.107
R1240 VDD.n1160 VDD.n1158 44.107
R1241 VDD.n1235 VDD.n1233 44.107
R1242 VDD.n1310 VDD.n1308 44.107
R1243 VDD.n1385 VDD.n1383 44.107
R1244 VDD.n1460 VDD.n1458 44.107
R1245 VDD.n761 VDD.n759 44.107
R1246 VDD.n690 VDD.n688 44.107
R1247 VDD.n615 VDD.n613 44.107
R1248 VDD.n540 VDD.n538 44.107
R1249 VDD.n465 VDD.n463 44.107
R1250 VDD.n390 VDD.n388 44.107
R1251 VDD.n315 VDD.n313 44.107
R1252 VDD.n240 VDD.n238 44.107
R1253 VDD.n165 VDD.n163 44.107
R1254 VDD.n108 VDD.n106 44.107
R1255 VDD.n786 VDD.n784 44.107
R1256 VDD.n3 VDD.n2 44.107
R1257 VDD.n20 VDD.n15 41.052
R1258 VDD.n68 VDD.n66 39.742
R1259 VDD.n68 VDD.n67 39.742
R1260 VDD.n70 VDD.n69 39.742
R1261 VDD.n123 VDD.n122 39.742
R1262 VDD.n180 VDD.n179 39.742
R1263 VDD.n255 VDD.n254 39.742
R1264 VDD.n330 VDD.n329 39.742
R1265 VDD.n405 VDD.n404 39.742
R1266 VDD.n480 VDD.n479 39.742
R1267 VDD.n555 VDD.n554 39.742
R1268 VDD.n630 VDD.n629 39.742
R1269 VDD.n705 VDD.n704 39.742
R1270 VDD.n776 VDD.n775 39.742
R1271 VDD.n1475 VDD.n1474 39.742
R1272 VDD.n1400 VDD.n1399 39.742
R1273 VDD.n1325 VDD.n1324 39.742
R1274 VDD.n1250 VDD.n1249 39.742
R1275 VDD.n1175 VDD.n1174 39.742
R1276 VDD.n1100 VDD.n1099 39.742
R1277 VDD.n1025 VDD.n1024 39.742
R1278 VDD.n950 VDD.n949 39.742
R1279 VDD.n799 VDD.n798 39.742
R1280 VDD.n877 VDD.n874 39.742
R1281 VDD.n877 VDD.n876 39.742
R1282 VDD.n873 VDD.n872 39.742
R1283 VDD.n108 VDD.n107 38
R1284 VDD.n165 VDD.n164 38
R1285 VDD.n240 VDD.n239 38
R1286 VDD.n315 VDD.n314 38
R1287 VDD.n390 VDD.n389 38
R1288 VDD.n465 VDD.n464 38
R1289 VDD.n540 VDD.n539 38
R1290 VDD.n615 VDD.n614 38
R1291 VDD.n690 VDD.n689 38
R1292 VDD.n761 VDD.n760 38
R1293 VDD.n1460 VDD.n1459 38
R1294 VDD.n1385 VDD.n1384 38
R1295 VDD.n1310 VDD.n1309 38
R1296 VDD.n1235 VDD.n1234 38
R1297 VDD.n1160 VDD.n1159 38
R1298 VDD.n1085 VDD.n1084 38
R1299 VDD.n1010 VDD.n1009 38
R1300 VDD.n935 VDD.n934 38
R1301 VDD.n786 VDD.n785 38
R1302 VDD.n933 VDD.n932 36.774
R1303 VDD.n1008 VDD.n1007 36.774
R1304 VDD.n1083 VDD.n1082 36.774
R1305 VDD.n1158 VDD.n1157 36.774
R1306 VDD.n1233 VDD.n1232 36.774
R1307 VDD.n1308 VDD.n1307 36.774
R1308 VDD.n1383 VDD.n1382 36.774
R1309 VDD.n1458 VDD.n1457 36.774
R1310 VDD.n759 VDD.n758 36.774
R1311 VDD.n688 VDD.n687 36.774
R1312 VDD.n613 VDD.n612 36.774
R1313 VDD.n538 VDD.n537 36.774
R1314 VDD.n463 VDD.n462 36.774
R1315 VDD.n388 VDD.n387 36.774
R1316 VDD.n313 VDD.n312 36.774
R1317 VDD.n238 VDD.n237 36.774
R1318 VDD.n163 VDD.n162 36.774
R1319 VDD.n106 VDD.n105 36.774
R1320 VDD.n66 VDD.n65 36.774
R1321 VDD.n876 VDD.n875 36.774
R1322 VDD.n196 0A�U 35.8
R1323 VDD.n271 �&��U 35.8
R1324 VDD.n346  35.8
R1325 VDD.n421  35.8
R1326 VDD.n496 ���U 35.8
R1327 VDD.n571  35.8
R1328 VDD.n646  35.8
R1329 VDD.n721  35.8
R1330 VDD.n1516 �`\�U 35.8
R1331 VDD.n1441  35.8
R1332 VDD.n1366 �n�U 35.8
R1333 VDD.n1291  35.8
R1334 VDD.n1216  35.8
R1335 VDD.n1141  35.8
R1336 VDD.n1066 �f�U 35.8
R1337 VDD.n991 @r!�U 35.8
R1338 VDD.n916 `�g�U 35.8
R1339 VDD.n840 0���U 35.8
R1340 VDD.n220 �+���~ 33.243
R1341 VDD.n295 VDD.t124 33.243
R1342 VDD.n370  33.243
R1343 VDD.n445  33.243
R1344 VDD.n520  33.243
R1345 VDD.n595  33.243
R1346 VDD.n670 VDD.t60 33.243
R1347 VDD.n745 �?�U 33.243
R1348 VDD.n1492 �̓�U 33.243
R1349 VDD.n1417  33.243
R1350 VDD.n1342  '8�U 33.243
R1351 VDD.n1267 ��+�U 33.243
R1352 VDD.n1192  33.243
R1353 VDD.n1117 @�d�U 33.243
R1354 VDD.n1042 VDD.t172 33.243
R1355 VDD.n967  33.243
R1356 VDD.n892  33.243
R1357 VDD.n816 ����U 33.243
R1358 VDD.n1 VDD.n0 30.923
R1359 VDD.n73 VDD.n71 26.38
R1360 VDD.n73 VDD.n70 26.38
R1361 VDD.n73 VDD.n68 26.38
R1362 VDD.n73 VDD.n72 26.38
R1363 VDD.n126 VDD.n124 26.38
R1364 VDD.n126 VDD.n123 26.38
R1365 VDD.n126 VDD.n125 26.38
R1366 VDD.n183 VDD.n181 26.38
R1367 VDD.n183 VDD.n180 26.38
R1368 VDD.n183 VDD.n182 26.38
R1369 VDD.n258 VDD.n256 26.38
R1370 VDD.n258 VDD.n255 26.38
R1371 VDD.n258 VDD.n257 26.38
R1372 VDD.n333 VDD.n331 26.38
R1373 VDD.n333 VDD.n330 26.38
R1374 VDD.n333 VDD.n332 26.38
R1375 VDD.n408 VDD.n406 26.38
R1376 VDD.n408 VDD.n405 26.38
R1377 VDD.n408 VDD.n407 26.38
R1378 VDD.n483 VDD.n481 26.38
R1379 VDD.n483 VDD.n480 26.38
R1380 VDD.n483 VDD.n482 26.38
R1381 VDD.n558 VDD.n556 26.38
R1382 VDD.n558 VDD.n555 26.38
R1383 VDD.n558 VDD.n557 26.38
R1384 VDD.n633 VDD.n631 26.38
R1385 VDD.n633 VDD.n630 26.38
R1386 VDD.n633 VDD.n632 26.38
R1387 VDD.n708 VDD.n706 26.38
R1388 VDD.n708 VDD.n705 26.38
R1389 VDD.n708 VDD.n707 26.38
R1390 VDD.n779 VDD.n777 26.38
R1391 VDD.n779 VDD.n776 26.38
R1392 VDD.n779 VDD.n778 26.38
R1393 VDD.n1478 VDD.n1476 26.38
R1394 VDD.n1478 VDD.n1475 26.38
R1395 VDD.n1478 VDD.n1477 26.38
R1396 VDD.n1403 VDD.n1401 26.38
R1397 VDD.n1403 VDD.n1400 26.38
R1398 VDD.n1403 VDD.n1402 26.38
R1399 VDD.n1328 VDD.n1326 26.38
R1400 VDD.n1328 VDD.n1325 26.38
R1401 VDD.n1328 VDD.n1327 26.38
R1402 VDD.n1253 VDD.n1251 26.38
R1403 VDD.n1253 VDD.n1250 26.38
R1404 VDD.n1253 VDD.n1252 26.38
R1405 VDD.n1178 VDD.n1176 26.38
R1406 VDD.n1178 VDD.n1175 26.38
R1407 VDD.n1178 VDD.n1177 26.38
R1408 VDD.n1103 VDD.n1101 26.38
R1409 VDD.n1103 VDD.n1100 26.38
R1410 VDD.n1103 VDD.n1102 26.38
R1411 VDD.n1028 VDD.n1026 26.38
R1412 VDD.n1028 VDD.n1025 26.38
R1413 VDD.n1028 VDD.n1027 26.38
R1414 VDD.n953 VDD.n951 26.38
R1415 VDD.n953 VDD.n950 26.38
R1416 VDD.n953 VDD.n952 26.38
R1417 VDD.n802 VDD.n800 26.38
R1418 VDD.n802 VDD.n799 26.38
R1419 VDD.n802 VDD.n801 26.38
R1420 VDD.n878 VDD.n877 26.38
R1421 VDD.n878 VDD.n873 26.38
R1422 VDD.n878 VDD.n871 26.38
R1423 VDD.n878 VDD.n870 26.38
R1424 VDD.n805 VDD.n797 22.915
R1425 VDD.n23 VDD.n14 22.915
R1426 VDD.n28  20.457
R1427 VDD.n93 VDD.t14 20.457
R1428 VDD.n136  20.457
R1429 VDD.n39  17.9
R1430 VDD.n82  17.9
R1431 VDD.n149  17.9
R1432 VDD.n200 �+���~ 15.343
R1433 VDD.n275  15.343
R1434 VDD.n350 VDD.t222 15.343
R1435 VDD.n425 �>a�U 15.343
R1436 VDD.n500  15.343
R1437 VDD.n575 �+���~ 15.343
R1438 VDD.n650 ����U 15.343
R1439 VDD.n725 �Q,�U 15.343
R1440 VDD.n1510  15.343
R1441 VDD.n1435 ��!�U 15.343
R1442 VDD.n1360 �P��U 15.343
R1443 VDD.n1285  15.343
R1444 VDD.n1210  15.343
R1445 VDD.n1135 @`
�U 15.343
R1446 VDD.n1060  15.343
R1447 VDD.n985  15.343
R1448 VDD.n910 VDD.t128 15.343
R1449 VDD.n834  15.343
R1450 VDD.n797 VDD.n795 14.864
R1451 VDD.n795 VDD.n793 14.864
R1452 VDD.n793 VDD.n791 14.864
R1453 VDD.n791 VDD.n789 14.864
R1454 VDD.n789 VDD.n787 14.864
R1455 VDD.n946 VDD.n944 14.864
R1456 VDD.n944 VDD.n942 14.864
R1457 VDD.n942 VDD.n940 14.864
R1458 VDD.n940 VDD.n938 14.864
R1459 VDD.n938 VDD.n936 14.864
R1460 VDD.n1021 VDD.n1019 14.864
R1461 VDD.n1019 VDD.n1017 14.864
R1462 VDD.n1017 VDD.n1015 14.864
R1463 VDD.n1015 VDD.n1013 14.864
R1464 VDD.n1013 VDD.n1011 14.864
R1465 VDD.n1096 VDD.n1094 14.864
R1466 VDD.n1094 VDD.n1092 14.864
R1467 VDD.n1092 VDD.n1090 14.864
R1468 VDD.n1090 VDD.n1088 14.864
R1469 VDD.n1088 VDD.n1086 14.864
R1470 VDD.n1171 VDD.n1169 14.864
R1471 VDD.n1169 VDD.n1167 14.864
R1472 VDD.n1167 VDD.n1165 14.864
R1473 VDD.n1165 VDD.n1163 14.864
R1474 VDD.n1163 VDD.n1161 14.864
R1475 VDD.n1246 VDD.n1244 14.864
R1476 VDD.n1244 VDD.n1242 14.864
R1477 VDD.n1242 VDD.n1240 14.864
R1478 VDD.n1240 VDD.n1238 14.864
R1479 VDD.n1238 VDD.n1236 14.864
R1480 VDD.n1321 VDD.n1319 14.864
R1481 VDD.n1319 VDD.n1317 14.864
R1482 VDD.n1317 VDD.n1315 14.864
R1483 VDD.n1315 VDD.n1313 14.864
R1484 VDD.n1313 VDD.n1311 14.864
R1485 VDD.n1396 VDD.n1394 14.864
R1486 VDD.n1394 VDD.n1392 14.864
R1487 VDD.n1392 VDD.n1390 14.864
R1488 VDD.n1390 VDD.n1388 14.864
R1489 VDD.n1388 VDD.n1386 14.864
R1490 VDD.n1471 VDD.n1469 14.864
R1491 VDD.n1469 VDD.n1467 14.864
R1492 VDD.n1467 VDD.n1465 14.864
R1493 VDD.n1465 VDD.n1463 14.864
R1494 VDD.n1463 VDD.n1461 14.864
R1495 VDD.n772 VDD.n770 14.864
R1496 VDD.n770 VDD.n768 14.864
R1497 VDD.n768 VDD.n766 14.864
R1498 VDD.n766 VDD.n764 14.864
R1499 VDD.n764 VDD.n762 14.864
R1500 VDD.n701 VDD.n699 14.864
R1501 VDD.n699 VDD.n697 14.864
R1502 VDD.n697 VDD.n695 14.864
R1503 VDD.n695 VDD.n693 14.864
R1504 VDD.n693 VDD.n691 14.864
R1505 VDD.n626 VDD.n624 14.864
R1506 VDD.n624 VDD.n622 14.864
R1507 VDD.n622 VDD.n620 14.864
R1508 VDD.n620 VDD.n618 14.864
R1509 VDD.n618 VDD.n616 14.864
R1510 VDD.n551 VDD.n549 14.864
R1511 VDD.n549 VDD.n547 14.864
R1512 VDD.n547 VDD.n545 14.864
R1513 VDD.n545 VDD.n543 14.864
R1514 VDD.n543 VDD.n541 14.864
R1515 VDD.n476 VDD.n474 14.864
R1516 VDD.n474 VDD.n472 14.864
R1517 VDD.n472 VDD.n470 14.864
R1518 VDD.n470 VDD.n468 14.864
R1519 VDD.n468 VDD.n466 14.864
R1520 VDD.n401 VDD.n399 14.864
R1521 VDD.n399 VDD.n397 14.864
R1522 VDD.n397 VDD.n395 14.864
R1523 VDD.n395 VDD.n393 14.864
R1524 VDD.n393 VDD.n391 14.864
R1525 VDD.n326 VDD.n324 14.864
R1526 VDD.n324 VDD.n322 14.864
R1527 VDD.n322 VDD.n320 14.864
R1528 VDD.n320 VDD.n318 14.864
R1529 VDD.n318 VDD.n316 14.864
R1530 VDD.n251 VDD.n249 14.864
R1531 VDD.n249 VDD.n247 14.864
R1532 VDD.n247 VDD.n245 14.864
R1533 VDD.n245 VDD.n243 14.864
R1534 VDD.n243 VDD.n241 14.864
R1535 VDD.n176 VDD.n174 14.864
R1536 VDD.n174 VDD.n172 14.864
R1537 VDD.n172 VDD.n170 14.864
R1538 VDD.n170 VDD.n168 14.864
R1539 VDD.n168 VDD.n166 14.864
R1540 VDD.n119 VDD.n117 14.864
R1541 VDD.n117 VDD.n115 14.864
R1542 VDD.n115 VDD.n113 14.864
R1543 VDD.n113 VDD.n111 14.864
R1544 VDD.n111 VDD.n109 14.864
R1545 VDD.n62 VDD.n60 14.864
R1546 VDD.n60 VDD.n58 14.864
R1547 VDD.n58 VDD.n56 14.864
R1548 VDD.n56 VDD.n54 14.864
R1549 VDD.n54 VDD.n52 14.864
R1550 VDD.n52 VDD.n51 14.864
R1551 VDD.n867 VDD.n865 14.864
R1552 VDD.n865 VDD.n863 14.864
R1553 VDD.n863 VDD.n861 14.864
R1554 VDD.n861 VDD.n859 14.864
R1555 VDD.n859 VDD.n857 14.864
R1556 VDD.n857 VDD.n856 14.864
R1557 VDD.n14 VDD.n13 14.864
R1558 VDD.n13 VDD.n11 14.864
R1559 VDD.n11 VDD.n9 14.864
R1560 VDD.n9 VDD.n7 14.864
R1561 VDD.n7 VDD.n5 14.864
R1562 VDD.n76 VDD.n63 14.864
R1563 VDD.n129 VDD.n120 14.864
R1564 VDD.n186 VDD.n177 14.864
R1565 VDD.n261 VDD.n252 14.864
R1566 VDD.n336 VDD.n327 14.864
R1567 VDD.n411 VDD.n402 14.864
R1568 VDD.n486 VDD.n477 14.864
R1569 VDD.n561 VDD.n552 14.864
R1570 VDD.n636 VDD.n627 14.864
R1571 VDD.n711 VDD.n702 14.864
R1572 VDD.n782 VDD.n773 14.864
R1573 VDD.n1481 VDD.n1472 14.864
R1574 VDD.n1406 VDD.n1397 14.864
R1575 VDD.n1331 VDD.n1322 14.864
R1576 VDD.n1256 VDD.n1247 14.864
R1577 VDD.n1181 VDD.n1172 14.864
R1578 VDD.n1106 VDD.n1097 14.864
R1579 VDD.n1031 VDD.n1022 14.864
R1580 VDD.n956 VDD.n947 14.864
R1581 VDD.n881 VDD.n868 14.864
R1582 VDD.n820 VDD.t203 14.282
R1583 VDD.n820 VDD.t143 14.282
R1584 VDD.n836 VDD.t69 14.282
R1585 VDD.n836 VDD.t221 14.282
R1586 VDD.n896 VDD.t182 14.282
R1587 VDD.n896 VDD.t171 14.282
R1588 VDD.n912 VDD.t129 14.282
R1589 VDD.n912 VDD.t180 14.282
R1590 VDD.n971 VDD.t165 14.282
R1591 VDD.n971 VDD.t77 14.282
R1592 VDD.n987 VDD.t43 14.282
R1593 VDD.n987 VDD.t63 14.282
R1594 VDD.n1046 VDD.t147 14.282
R1595 VDD.n1046 VDD.t49 14.282
R1596 VDD.n1062 VDD.t201 14.282
R1597 VDD.n1062 VDD.t67 14.282
R1598 VDD.n1121 VDD.t217 14.282
R1599 VDD.n1121 VDD.t33 14.282
R1600 VDD.n1137 VDD.t18 14.282
R1601 VDD.n1137 VDD.t199 14.282
R1602 VDD.n1196 VDD.t94 14.282
R1603 VDD.n1196 VDD.t117 14.282
R1604 VDD.n1212 VDD.t41 14.282
R1605 VDD.n1212 VDD.t83 14.282
R1606 VDD.n1271 VDD.t195 14.282
R1607 VDD.n1271 VDD.t121 14.282
R1608 VDD.n1287 VDD.t79 14.282
R1609 VDD.n1287 VDD.t215 14.282
R1610 VDD.n1346 VDD.t7 14.282
R1611 VDD.n1346 VDD.t27 14.282
R1612 VDD.n1362 VDD.t75 14.282
R1613 VDD.n1362 VDD.t102 14.282
R1614 VDD.n1421 VDD.t91 14.282
R1615 VDD.n1421 VDD.t51 14.282
R1616 VDD.n1437 VDD.t57 14.282
R1617 VDD.n1437 VDD.t178 14.282
R1618 VDD.n1496 VDD.t24 14.282
R1619 VDD.n1496 VDD.t5 14.282
R1620 VDD.n1512 VDD.t193 14.282
R1621 VDD.n1512 VDD.t145 14.282
R1622 VDD.n739 VDD.t211 14.282
R1623 VDD.n739 VDD.t3 14.282
R1624 VDD.n727 VDD.t176 14.282
R1625 VDD.n727 VDD.t225 14.282
R1626 VDD.n664 VDD.t81 14.282
R1627 VDD.n664 VDD.t104 14.282
R1628 VDD.n652 VDD.t9 14.282
R1629 VDD.n652 VDD.t39 14.282
R1630 VDD.n589 VDD.t205 14.282
R1631 VDD.n589 VDD.t141 14.282
R1632 VDD.n577 VDD.t87 14.282
R1633 VDD.n577 VDD.t209 14.282
R1634 VDD.n514 VDD.t123 14.282
R1635 VDD.n514 VDD.t71 14.282
R1636 VDD.n502 VDD.t153 14.282
R1637 VDD.n502 VDD.t22 14.282
R1638 VDD.n439 VDD.t133 14.282
R1639 VDD.n439 VDD.t137 14.282
R1640 VDD.n427 VDD.t155 14.282
R1641 VDD.n427 VDD.t185 14.282
R1642 VDD.n364 VDD.t45 14.282
R1643 VDD.n364 VDD.t110 14.282
R1644 VDD.n352 VDD.t223 14.282
R1645 VDD.n352 VDD.t53 14.282
R1646 VDD.n289 VDD.t213 14.282
R1647 VDD.n289 VDD.t149 14.282
R1648 VDD.n277 VDD.t65 14.282
R1649 VDD.n277 VDD.t227 14.282
R1650 VDD.n214 VDD.t100 14.282
R1651 VDD.n214 VDD.t229 14.282
R1652 VDD.n202 VDD.t159 14.282
R1653 VDD.n202 VDD.t13 14.282
R1654 VDD.n140 VDD.t98 14.282
R1655 VDD.n140 VDD.t167 14.282
R1656 VDD.n216  12.786
R1657 VDD.n291  12.786
R1658 VDD.n366 �`��U 12.786
R1659 VDD.n441 ���U 12.786
R1660 VDD.n516  12.786
R1661 VDD.n591  12.786
R1662 VDD.n666 ��$�U 12.786
R1663 VDD.n741  12.786
R1664 VDD.n1498  HY�U 12.786
R1665 VDD.n1423  12.786
R1666 VDD.n1348  12.786
R1667 VDD.n1273  12.786
R1668 VDD.n1198 ��+�U 12.786
R1669 VDD.n1123  12.786
R1670 VDD.n1048  12.786
R1671 VDD.n973 pe�U 12.786
R1672 VDD.n898 �xB�U 12.786
R1673 VDD.n822  12.786
R1674 VDD.n143 VDD.n141 9.083
R1675 VDD.n23 VDD.n22 8.855
R1676 VDD.n22 VDD.n21 8.855
R1677 VDD.n26 VDD.n25 8.855
R1678 VDD.n25 VDD.n24 8.855
R1679 VDD.n30 VDD.n29 8.855
R1680 VDD.n29 VDD.n28 8.855
R1681 VDD.n33 VDD.n32 8.855
R1682 VDD.n32 �x��U 8.855
R1683 VDD.n37 VDD.n36 8.855
R1684 VDD.n36 VDD.n35 8.855
R1685 VDD.n41 VDD.n40 8.855
R1686 VDD.n40 VDD.n39 8.855
R1687 VDD.n45 VDD.n44 8.855
R1688 VDD.n44 VDD.n43 8.855
R1689 VDD.n49 VDD.n48 8.855
R1690 VDD.n48 VDD.n47 8.855
R1691 VDD.n76 VDD.n75 8.855
R1692 VDD.n75 VDD.n74 8.855
R1693 VDD.n80 VDD.n79 8.855
R1694 VDD.n79 VDD.n78 8.855
R1695 VDD.n84 VDD.n83 8.855
R1696 VDD.n83 VDD.n82 8.855
R1697 VDD.n88 VDD.n87 8.855
R1698 VDD.n87 VDD.n86 8.855
R1699 VDD.n91 VDD.n90 8.855
R1700 VDD.n90  8.855
R1701 VDD.n95 VDD.n94 8.855
R1702 VDD.n94 VDD.n93 8.855
R1703 VDD.n99 VDD.n98 8.855
R1704 VDD.n98 VDD.n97 8.855
R1705 VDD.n103 VDD.n102 8.855
R1706 VDD.n102 VDD.n101 8.855
R1707 VDD.n129 VDD.n128 8.855
R1708 VDD.n128 VDD.n127 8.855
R1709 VDD.n134 VDD.n133 8.855
R1710 VDD.n133 VDD.n132 8.855
R1711 VDD.n138 VDD.n137 8.855
R1712 VDD.n137 VDD.n136 8.855
R1713 VDD.n143 VDD.n142 8.855
R1714 VDD.n142 ���U 8.855
R1715 VDD.n147 VDD.n146 8.855
R1716 VDD.n146 VDD.n145 8.855
R1717 VDD.n151 VDD.n150 8.855
R1718 VDD.n150 VDD.n149 8.855
R1719 VDD.n156 VDD.n155 8.855
R1720 VDD.n155 VDD.n154 8.855
R1721 VDD.n160 VDD.n159 8.855
R1722 VDD.n159 VDD.n158 8.855
R1723 VDD.n186 VDD.n185 8.855
R1724 VDD.n185 VDD.n184 8.855
R1725 VDD.n190 VDD.n189 8.855
R1726 VDD.n189 VDD.n188 8.855
R1727 VDD.n194 VDD.n193 8.855
R1728 VDD.n193 VDD.n192 8.855
R1729 VDD.n198 VDD.n197 8.855
R1730 VDD.n197 VDD.n196 8.855
R1731 VDD.n204 VDD.n201 8.855
R1732 VDD.n201 VDD.n200 8.855
R1733 VDD.n208 VDD.n207 8.855
R1734 VDD.n207 VDD.n206 8.855
R1735 VDD.n212 VDD.n211 8.855
R1736 VDD.n211 VDD.n210 8.855
R1737 VDD.n218 VDD.n217 8.855
R1738 VDD.n217 VDD.n216 8.855
R1739 VDD.n222 VDD.n221 8.855
R1740 VDD.n221 VDD.n220 8.855
R1741 VDD.n227 VDD.n226 8.855
R1742 VDD.n226 VDD.n225 8.855
R1743 VDD.n231 VDD.n230 8.855
R1744 VDD.n230 VDD.n229 8.855
R1745 VDD.n235 VDD.n234 8.855
R1746 VDD.n234 VDD.n233 8.855
R1747 VDD.n261 VDD.n260 8.855
R1748 VDD.n260 VDD.n259 8.855
R1749 VDD.n265 VDD.n264 8.855
R1750 VDD.n264 VDD.n263 8.855
R1751 VDD.n269 VDD.n268 8.855
R1752 VDD.n268 VDD.n267 8.855
R1753 VDD.n273 VDD.n272 8.855
R1754 VDD.n272 VDD.n271 8.855
R1755 VDD.n279 VDD.n276 8.855
R1756 VDD.n276 VDD.n275 8.855
R1757 VDD.n283 VDD.n282 8.855
R1758 VDD.n282 VDD.n281 8.855
R1759 VDD.n287 VDD.n286 8.855
R1760 VDD.n286 VDD.n285 8.855
R1761 VDD.n293 VDD.n292 8.855
R1762 VDD.n292 VDD.n291 8.855
R1763 VDD.n297 VDD.n296 8.855
R1764 VDD.n296 VDD.n295 8.855
R1765 VDD.n302 VDD.n301 8.855
R1766 VDD.n301 VDD.n300 8.855
R1767 VDD.n306 VDD.n305 8.855
R1768 VDD.n305 VDD.n304 8.855
R1769 VDD.n310 VDD.n309 8.855
R1770 VDD.n309 VDD.n308 8.855
R1771 VDD.n336 VDD.n335 8.855
R1772 VDD.n335 VDD.n334 8.855
R1773 VDD.n340 VDD.n339 8.855
R1774 VDD.n339 VDD.n338 8.855
R1775 VDD.n344 VDD.n343 8.855
R1776 VDD.n343 VDD.n342 8.855
R1777 VDD.n348 VDD.n347 8.855
R1778 VDD.n347 VDD.n346 8.855
R1779 VDD.n354 VDD.n351 8.855
R1780 VDD.n351 VDD.n350 8.855
R1781 VDD.n358 VDD.n357 8.855
R1782 VDD.n357 VDD.n356 8.855
R1783 VDD.n362 VDD.n361 8.855
R1784 VDD.n361 VDD.n360 8.855
R1785 VDD.n368 VDD.n367 8.855
R1786 VDD.n367 VDD.n366 8.855
R1787 VDD.n372 VDD.n371 8.855
R1788 VDD.n371 VDD.n370 8.855
R1789 VDD.n377 VDD.n376 8.855
R1790 VDD.n376 VDD.n375 8.855
R1791 VDD.n381 VDD.n380 8.855
R1792 VDD.n380 VDD.n379 8.855
R1793 VDD.n385 VDD.n384 8.855
R1794 VDD.n384 VDD.n383 8.855
R1795 VDD.n411 VDD.n410 8.855
R1796 VDD.n410 VDD.n409 8.855
R1797 VDD.n415 VDD.n414 8.855
R1798 VDD.n414 VDD.n413 8.855
R1799 VDD.n419 VDD.n418 8.855
R1800 VDD.n418 VDD.n417 8.855
R1801 VDD.n423 VDD.n422 8.855
R1802 VDD.n422 VDD.n421 8.855
R1803 VDD.n429 VDD.n426 8.855
R1804 VDD.n426 VDD.n425 8.855
R1805 VDD.n433 VDD.n432 8.855
R1806 VDD.n432 VDD.n431 8.855
R1807 VDD.n437 VDD.n436 8.855
R1808 VDD.n436 VDD.n435 8.855
R1809 VDD.n443 VDD.n442 8.855
R1810 VDD.n442 VDD.n441 8.855
R1811 VDD.n447 VDD.n446 8.855
R1812 VDD.n446 VDD.n445 8.855
R1813 VDD.n452 VDD.n451 8.855
R1814 VDD.n451 VDD.n450 8.855
R1815 VDD.n456 VDD.n455 8.855
R1816 VDD.n455 VDD.n454 8.855
R1817 VDD.n460 VDD.n459 8.855
R1818 VDD.n459 VDD.n458 8.855
R1819 VDD.n486 VDD.n485 8.855
R1820 VDD.n485 VDD.n484 8.855
R1821 VDD.n490 VDD.n489 8.855
R1822 VDD.n489 VDD.n488 8.855
R1823 VDD.n494 VDD.n493 8.855
R1824 VDD.n493 VDD.n492 8.855
R1825 VDD.n498 VDD.n497 8.855
R1826 VDD.n497 VDD.n496 8.855
R1827 VDD.n504 VDD.n501 8.855
R1828 VDD.n501 VDD.n500 8.855
R1829 VDD.n508 VDD.n507 8.855
R1830 VDD.n507 VDD.n506 8.855
R1831 VDD.n512 VDD.n511 8.855
R1832 VDD.n511 VDD.n510 8.855
R1833 VDD.n518 VDD.n517 8.855
R1834 VDD.n517 VDD.n516 8.855
R1835 VDD.n522 VDD.n521 8.855
R1836 VDD.n521 VDD.n520 8.855
R1837 VDD.n527 VDD.n526 8.855
R1838 VDD.n526 VDD.n525 8.855
R1839 VDD.n531 VDD.n530 8.855
R1840 VDD.n530 VDD.n529 8.855
R1841 VDD.n535 VDD.n534 8.855
R1842 VDD.n534 VDD.n533 8.855
R1843 VDD.n561 VDD.n560 8.855
R1844 VDD.n560 VDD.n559 8.855
R1845 VDD.n565 VDD.n564 8.855
R1846 VDD.n564 VDD.n563 8.855
R1847 VDD.n569 VDD.n568 8.855
R1848 VDD.n568 VDD.n567 8.855
R1849 VDD.n573 VDD.n572 8.855
R1850 VDD.n572 VDD.n571 8.855
R1851 VDD.n579 VDD.n576 8.855
R1852 VDD.n576 VDD.n575 8.855
R1853 VDD.n583 VDD.n582 8.855
R1854 VDD.n582 VDD.n581 8.855
R1855 VDD.n587 VDD.n586 8.855
R1856 VDD.n586 VDD.n585 8.855
R1857 VDD.n593 VDD.n592 8.855
R1858 VDD.n592 VDD.n591 8.855
R1859 VDD.n597 VDD.n596 8.855
R1860 VDD.n596 VDD.n595 8.855
R1861 VDD.n602 VDD.n601 8.855
R1862 VDD.n601 VDD.n600 8.855
R1863 VDD.n606 VDD.n605 8.855
R1864 VDD.n605 VDD.n604 8.855
R1865 VDD.n610 VDD.n609 8.855
R1866 VDD.n609 VDD.n608 8.855
R1867 VDD.n636 VDD.n635 8.855
R1868 VDD.n635 VDD.n634 8.855
R1869 VDD.n640 VDD.n639 8.855
R1870 VDD.n639 VDD.n638 8.855
R1871 VDD.n644 VDD.n643 8.855
R1872 VDD.n643 VDD.n642 8.855
R1873 VDD.n648 VDD.n647 8.855
R1874 VDD.n647 VDD.n646 8.855
R1875 VDD.n654 VDD.n651 8.855
R1876 VDD.n651 VDD.n650 8.855
R1877 VDD.n658 VDD.n657 8.855
R1878 VDD.n657 VDD.n656 8.855
R1879 VDD.n662 VDD.n661 8.855
R1880 VDD.n661 VDD.n660 8.855
R1881 VDD.n668 VDD.n667 8.855
R1882 VDD.n667 VDD.n666 8.855
R1883 VDD.n672 VDD.n671 8.855
R1884 VDD.n671 VDD.n670 8.855
R1885 VDD.n677 VDD.n676 8.855
R1886 VDD.n676 VDD.n675 8.855
R1887 VDD.n681 VDD.n680 8.855
R1888 VDD.n680 VDD.n679 8.855
R1889 VDD.n685 VDD.n684 8.855
R1890 VDD.n684 VDD.n683 8.855
R1891 VDD.n711 VDD.n710 8.855
R1892 VDD.n710 VDD.n709 8.855
R1893 VDD.n715 VDD.n714 8.855
R1894 VDD.n714 VDD.n713 8.855
R1895 VDD.n719 VDD.n718 8.855
R1896 VDD.n718 VDD.n717 8.855
R1897 VDD.n723 VDD.n722 8.855
R1898 VDD.n722 VDD.n721 8.855
R1899 VDD.n729 VDD.n726 8.855
R1900 VDD.n726 VDD.n725 8.855
R1901 VDD.n733 VDD.n732 8.855
R1902 VDD.n732 VDD.n731 8.855
R1903 VDD.n737 VDD.n736 8.855
R1904 VDD.n736 VDD.n735 8.855
R1905 VDD.n743 VDD.n742 8.855
R1906 VDD.n742 VDD.n741 8.855
R1907 VDD.n747 VDD.n746 8.855
R1908 VDD.n746 VDD.n745 8.855
R1909 VDD.n752 VDD.n751 8.855
R1910 VDD.n751 VDD.n750 8.855
R1911 VDD.n756 VDD.n755 8.855
R1912 VDD.n755 VDD.n754 8.855
R1913 VDD.n782 VDD.n781 8.855
R1914 VDD.n781 VDD.n780 8.855
R1915 VDD.n1530 VDD.n1529 8.855
R1916 VDD.n1529 VDD.n1528 8.855
R1917 VDD.n1526 VDD.n1525 8.855
R1918 VDD.n1525 VDD.n1524 8.855
R1919 VDD.n1522 VDD.n1521 8.855
R1920 VDD.n1521 VDD.n1520 8.855
R1921 VDD.n1518 VDD.n1517 8.855
R1922 VDD.n1517 VDD.n1516 8.855
R1923 VDD.n1514 VDD.n1511 8.855
R1924 VDD.n1511 VDD.n1510 8.855
R1925 VDD.n1508 VDD.n1507 8.855
R1926 VDD.n1507 VDD.n1506 8.855
R1927 VDD.n1504 VDD.n1503 8.855
R1928 VDD.n1503 VDD.n1502 8.855
R1929 VDD.n1500 VDD.n1499 8.855
R1930 VDD.n1499 VDD.n1498 8.855
R1931 VDD.n1494 VDD.n1493 8.855
R1932 VDD.n1493 VDD.n1492 8.855
R1933 VDD.n1490 VDD.n1489 8.855
R1934 VDD.n1489 VDD.n1488 8.855
R1935 VDD.n1485 VDD.n1484 8.855
R1936 VDD.n1484 VDD.n1483 8.855
R1937 VDD.n1481 VDD.n1480 8.855
R1938 VDD.n1480 VDD.n1479 8.855
R1939 VDD.n1455 VDD.n1454 8.855
R1940 VDD.n1454 VDD.n1453 8.855
R1941 VDD.n1451 VDD.n1450 8.855
R1942 VDD.n1450 VDD.n1449 8.855
R1943 VDD.n1447 VDD.n1446 8.855
R1944 VDD.n1446 VDD.n1445 8.855
R1945 VDD.n1443 VDD.n1442 8.855
R1946 VDD.n1442 VDD.n1441 8.855
R1947 VDD.n1439 VDD.n1436 8.855
R1948 VDD.n1436 VDD.n1435 8.855
R1949 VDD.n1433 VDD.n1432 8.855
R1950 VDD.n1432 VDD.n1431 8.855
R1951 VDD.n1429 VDD.n1428 8.855
R1952 VDD.n1428 VDD.n1427 8.855
R1953 VDD.n1425 VDD.n1424 8.855
R1954 VDD.n1424 VDD.n1423 8.855
R1955 VDD.n1419 VDD.n1418 8.855
R1956 VDD.n1418 VDD.n1417 8.855
R1957 VDD.n1415 VDD.n1414 8.855
R1958 VDD.n1414 VDD.n1413 8.855
R1959 VDD.n1410 VDD.n1409 8.855
R1960 VDD.n1409 VDD.n1408 8.855
R1961 VDD.n1406 VDD.n1405 8.855
R1962 VDD.n1405 VDD.n1404 8.855
R1963 VDD.n1380 VDD.n1379 8.855
R1964 VDD.n1379 VDD.n1378 8.855
R1965 VDD.n1376 VDD.n1375 8.855
R1966 VDD.n1375 VDD.n1374 8.855
R1967 VDD.n1372 VDD.n1371 8.855
R1968 VDD.n1371 VDD.n1370 8.855
R1969 VDD.n1368 VDD.n1367 8.855
R1970 VDD.n1367 VDD.n1366 8.855
R1971 VDD.n1364 VDD.n1361 8.855
R1972 VDD.n1361 VDD.n1360 8.855
R1973 VDD.n1358 VDD.n1357 8.855
R1974 VDD.n1357 VDD.n1356 8.855
R1975 VDD.n1354 VDD.n1353 8.855
R1976 VDD.n1353 VDD.n1352 8.855
R1977 VDD.n1350 VDD.n1349 8.855
R1978 VDD.n1349 VDD.n1348 8.855
R1979 VDD.n1344 VDD.n1343 8.855
R1980 VDD.n1343 VDD.n1342 8.855
R1981 VDD.n1340 VDD.n1339 8.855
R1982 VDD.n1339 VDD.n1338 8.855
R1983 VDD.n1335 VDD.n1334 8.855
R1984 VDD.n1334 VDD.n1333 8.855
R1985 VDD.n1331 VDD.n1330 8.855
R1986 VDD.n1330 VDD.n1329 8.855
R1987 VDD.n1305 VDD.n1304 8.855
R1988 VDD.n1304 VDD.n1303 8.855
R1989 VDD.n1301 VDD.n1300 8.855
R1990 VDD.n1300 VDD.n1299 8.855
R1991 VDD.n1297 VDD.n1296 8.855
R1992 VDD.n1296 VDD.n1295 8.855
R1993 VDD.n1293 VDD.n1292 8.855
R1994 VDD.n1292 VDD.n1291 8.855
R1995 VDD.n1289 VDD.n1286 8.855
R1996 VDD.n1286 VDD.n1285 8.855
R1997 VDD.n1283 VDD.n1282 8.855
R1998 VDD.n1282 VDD.n1281 8.855
R1999 VDD.n1279 VDD.n1278 8.855
R2000 VDD.n1278 VDD.n1277 8.855
R2001 VDD.n1275 VDD.n1274 8.855
R2002 VDD.n1274 VDD.n1273 8.855
R2003 VDD.n1269 VDD.n1268 8.855
R2004 VDD.n1268 VDD.n1267 8.855
R2005 VDD.n1265 VDD.n1264 8.855
R2006 VDD.n1264 VDD.n1263 8.855
R2007 VDD.n1260 VDD.n1259 8.855
R2008 VDD.n1259 VDD.n1258 8.855
R2009 VDD.n1256 VDD.n1255 8.855
R2010 VDD.n1255 VDD.n1254 8.855
R2011 VDD.n1230 VDD.n1229 8.855
R2012 VDD.n1229 VDD.n1228 8.855
R2013 VDD.n1226 VDD.n1225 8.855
R2014 VDD.n1225 VDD.n1224 8.855
R2015 VDD.n1222 VDD.n1221 8.855
R2016 VDD.n1221 VDD.n1220 8.855
R2017 VDD.n1218 VDD.n1217 8.855
R2018 VDD.n1217 VDD.n1216 8.855
R2019 VDD.n1214 VDD.n1211 8.855
R2020 VDD.n1211 VDD.n1210 8.855
R2021 VDD.n1208 VDD.n1207 8.855
R2022 VDD.n1207 VDD.n1206 8.855
R2023 VDD.n1204 VDD.n1203 8.855
R2024 VDD.n1203 VDD.n1202 8.855
R2025 VDD.n1200 VDD.n1199 8.855
R2026 VDD.n1199 VDD.n1198 8.855
R2027 VDD.n1194 VDD.n1193 8.855
R2028 VDD.n1193 VDD.n1192 8.855
R2029 VDD.n1190 VDD.n1189 8.855
R2030 VDD.n1189 VDD.n1188 8.855
R2031 VDD.n1185 VDD.n1184 8.855
R2032 VDD.n1184 VDD.n1183 8.855
R2033 VDD.n1181 VDD.n1180 8.855
R2034 VDD.n1180 VDD.n1179 8.855
R2035 VDD.n1155 VDD.n1154 8.855
R2036 VDD.n1154 VDD.n1153 8.855
R2037 VDD.n1151 VDD.n1150 8.855
R2038 VDD.n1150 VDD.n1149 8.855
R2039 VDD.n1147 VDD.n1146 8.855
R2040 VDD.n1146 VDD.n1145 8.855
R2041 VDD.n1143 VDD.n1142 8.855
R2042 VDD.n1142 VDD.n1141 8.855
R2043 VDD.n1139 VDD.n1136 8.855
R2044 VDD.n1136 VDD.n1135 8.855
R2045 VDD.n1133 VDD.n1132 8.855
R2046 VDD.n1132 VDD.n1131 8.855
R2047 VDD.n1129 VDD.n1128 8.855
R2048 VDD.n1128 VDD.n1127 8.855
R2049 VDD.n1125 VDD.n1124 8.855
R2050 VDD.n1124 VDD.n1123 8.855
R2051 VDD.n1119 VDD.n1118 8.855
R2052 VDD.n1118 VDD.n1117 8.855
R2053 VDD.n1115 VDD.n1114 8.855
R2054 VDD.n1114 VDD.n1113 8.855
R2055 VDD.n1110 VDD.n1109 8.855
R2056 VDD.n1109 VDD.n1108 8.855
R2057 VDD.n1106 VDD.n1105 8.855
R2058 VDD.n1105 VDD.n1104 8.855
R2059 VDD.n1080 VDD.n1079 8.855
R2060 VDD.n1079 VDD.n1078 8.855
R2061 VDD.n1076 VDD.n1075 8.855
R2062 VDD.n1075 VDD.n1074 8.855
R2063 VDD.n1072 VDD.n1071 8.855
R2064 VDD.n1071 VDD.n1070 8.855
R2065 VDD.n1068 VDD.n1067 8.855
R2066 VDD.n1067 VDD.n1066 8.855
R2067 VDD.n1064 VDD.n1061 8.855
R2068 VDD.n1061 VDD.n1060 8.855
R2069 VDD.n1058 VDD.n1057 8.855
R2070 VDD.n1057 VDD.n1056 8.855
R2071 VDD.n1054 VDD.n1053 8.855
R2072 VDD.n1053 VDD.n1052 8.855
R2073 VDD.n1050 VDD.n1049 8.855
R2074 VDD.n1049 VDD.n1048 8.855
R2075 VDD.n1044 VDD.n1043 8.855
R2076 VDD.n1043 VDD.n1042 8.855
R2077 VDD.n1040 VDD.n1039 8.855
R2078 VDD.n1039 VDD.n1038 8.855
R2079 VDD.n1035 VDD.n1034 8.855
R2080 VDD.n1034 VDD.n1033 8.855
R2081 VDD.n1031 VDD.n1030 8.855
R2082 VDD.n1030 VDD.n1029 8.855
R2083 VDD.n1005 VDD.n1004 8.855
R2084 VDD.n1004 VDD.n1003 8.855
R2085 VDD.n1001 VDD.n1000 8.855
R2086 VDD.n1000 VDD.n999 8.855
R2087 VDD.n997 VDD.n996 8.855
R2088 VDD.n996 VDD.n995 8.855
R2089 VDD.n993 VDD.n992 8.855
R2090 VDD.n992 VDD.n991 8.855
R2091 VDD.n989 VDD.n986 8.855
R2092 VDD.n986 VDD.n985 8.855
R2093 VDD.n983 VDD.n982 8.855
R2094 VDD.n982 VDD.n981 8.855
R2095 VDD.n979 VDD.n978 8.855
R2096 VDD.n978 VDD.n977 8.855
R2097 VDD.n975 VDD.n974 8.855
R2098 VDD.n974 VDD.n973 8.855
R2099 VDD.n969 VDD.n968 8.855
R2100 VDD.n968 VDD.n967 8.855
R2101 VDD.n965 VDD.n964 8.855
R2102 VDD.n964 VDD.n963 8.855
R2103 VDD.n960 VDD.n959 8.855
R2104 VDD.n959 VDD.n958 8.855
R2105 VDD.n956 VDD.n955 8.855
R2106 VDD.n955 VDD.n954 8.855
R2107 VDD.n930 VDD.n929 8.855
R2108 VDD.n929 VDD.n928 8.855
R2109 VDD.n926 VDD.n925 8.855
R2110 VDD.n925 VDD.n924 8.855
R2111 VDD.n922 VDD.n921 8.855
R2112 VDD.n921 VDD.n920 8.855
R2113 VDD.n918 VDD.n917 8.855
R2114 VDD.n917 VDD.n916 8.855
R2115 VDD.n914 VDD.n911 8.855
R2116 VDD.n911 VDD.n910 8.855
R2117 VDD.n908 VDD.n907 8.855
R2118 VDD.n907 VDD.n906 8.855
R2119 VDD.n904 VDD.n903 8.855
R2120 VDD.n903 VDD.n902 8.855
R2121 VDD.n900 VDD.n899 8.855
R2122 VDD.n899 VDD.n898 8.855
R2123 VDD.n894 VDD.n893 8.855
R2124 VDD.n893 VDD.n892 8.855
R2125 VDD.n890 VDD.n889 8.855
R2126 VDD.n889 VDD.n888 8.855
R2127 VDD.n885 VDD.n884 8.855
R2128 VDD.n884 VDD.n883 8.855
R2129 VDD.n881 VDD.n880 8.855
R2130 VDD.n880 VDD.n879 8.855
R2131 VDD.n854 VDD.n853 8.855
R2132 VDD.n853 VDD.n852 8.855
R2133 VDD.n850 VDD.n849 8.855
R2134 VDD.n849 VDD.n848 8.855
R2135 VDD.n846 VDD.n845 8.855
R2136 VDD.n845 VDD.n844 8.855
R2137 VDD.n842 VDD.n841 8.855
R2138 VDD.n841 VDD.n840 8.855
R2139 VDD.n838 VDD.n835 8.855
R2140 VDD.n835 VDD.n834 8.855
R2141 VDD.n832 VDD.n831 8.855
R2142 VDD.n831 VDD.n830 8.855
R2143 VDD.n828 VDD.n827 8.855
R2144 VDD.n827 VDD.n826 8.855
R2145 VDD.n824 VDD.n823 8.855
R2146 VDD.n823 VDD.n822 8.855
R2147 VDD.n818 VDD.n817 8.855
R2148 VDD.n817 VDD.n816 8.855
R2149 VDD.n814 VDD.n813 8.855
R2150 VDD.n813 VDD.n812 8.855
R2151 VDD.n809 VDD.n808 8.855
R2152 VDD.n808 VDD.n807 8.855
R2153 VDD.n805 VDD.n804 8.855
R2154 VDD.n804 VDD.n803 8.855
R2155 VDD.n947 VDD.n946 8.051
R2156 VDD.n1022 VDD.n1021 8.051
R2157 VDD.n1097 VDD.n1096 8.051
R2158 VDD.n1172 VDD.n1171 8.051
R2159 VDD.n1247 VDD.n1246 8.051
R2160 VDD.n1322 VDD.n1321 8.051
R2161 VDD.n1397 VDD.n1396 8.051
R2162 VDD.n1472 VDD.n1471 8.051
R2163 VDD.n773 VDD.n772 8.051
R2164 VDD.n702 VDD.n701 8.051
R2165 VDD.n627 VDD.n626 8.051
R2166 VDD.n552 VDD.n551 8.051
R2167 VDD.n477 VDD.n476 8.051
R2168 VDD.n402 VDD.n401 8.051
R2169 VDD.n327 VDD.n326 8.051
R2170 VDD.n252 VDD.n251 8.051
R2171 VDD.n177 VDD.n176 8.051
R2172 VDD.n120 VDD.n119 8.051
R2173 VDD.n63 VDD.n62 8.051
R2174 VDD.n868 VDD.n867 8.051
R2175 VDD.n210 ���U 7.671
R2176 VDD.n285 �1B�U 7.671
R2177 VDD.n360  7.671
R2178 VDD.n435 �l��U 7.671
R2179 VDD.n510 �Nt�U 7.671
R2180 VDD.n585 @,�U 7.671
R2181 VDD.n660 �+���~ 7.671
R2182 VDD.n735 0Ɔ�U 7.671
R2183 VDD.n1502 VDD.t23 7.671
R2184 VDD.n1427  7.671
R2185 VDD.n1352 �N��U 7.671
R2186 VDD.n1277  7.671
R2187 VDD.n1202  7.671
R2188 VDD.n1127 �+���~ 7.671
R2189 VDD.n1052 �+���~ 7.671
R2190 VDD.n977  7.671
R2191 VDD.n902 P_��U 7.671
R2192 VDD.n826 �+���~ 7.671
R2193 VDD.n218 VDD.n215 7.019
R2194 VDD.n293 VDD.n290 7.019
R2195 VDD.n368 VDD.n365 7.019
R2196 VDD.n443 VDD.n440 7.019
R2197 VDD.n518 VDD.n515 7.019
R2198 VDD.n593 VDD.n590 7.019
R2199 VDD.n668 VDD.n665 7.019
R2200 VDD.n743 VDD.n740 7.019
R2201 VDD.n1500 VDD.n1497 7.019
R2202 VDD.n1425 VDD.n1422 7.019
R2203 VDD.n1350 VDD.n1347 7.019
R2204 VDD.n1275 VDD.n1272 7.019
R2205 VDD.n1200 VDD.n1197 7.019
R2206 VDD.n1125 VDD.n1122 7.019
R2207 VDD.n1050 VDD.n1047 7.019
R2208 VDD.n975 VDD.n972 7.019
R2209 VDD.n900 VDD.n897 7.019
R2210 VDD.n824 VDD.n821 7.019
R2211 VDD.n204 VDD.n203 6.606
R2212 VDD.n279 VDD.n278 6.606
R2213 VDD.n354 VDD.n353 6.606
R2214 VDD.n429 VDD.n428 6.606
R2215 VDD.n504 VDD.n503 6.606
R2216 VDD.n579 VDD.n578 6.606
R2217 VDD.n654 VDD.n653 6.606
R2218 VDD.n729 VDD.n728 6.606
R2219 VDD.n1514 VDD.n1513 6.606
R2220 VDD.n1439 VDD.n1438 6.606
R2221 VDD.n1364 VDD.n1363 6.606
R2222 VDD.n1289 VDD.n1288 6.606
R2223 VDD.n1214 VDD.n1213 6.606
R2224 VDD.n1139 VDD.n1138 6.606
R2225 VDD.n1064 VDD.n1063 6.606
R2226 VDD.n989 VDD.n988 6.606
R2227 VDD.n914 VDD.n913 6.606
R2228 VDD.n838 VDD.n837 6.606
R2229 VDD.n206  5.114
R2230 VDD.n281 pV�U 5.114
R2231 VDD.n356 VDD.t52 5.114
R2232 VDD.n431 �B�U 5.114
R2233 VDD.n506 ����U 5.114
R2234 VDD.n581 VDD.t208 5.114
R2235 VDD.n656  5.114
R2236 VDD.n731 �v��U 5.114
R2237 VDD.n1506 �!�U 5.114
R2238 VDD.n1431 VDD.t177 5.114
R2239 VDD.n1356  5.114
R2240 VDD.n1281 �,�U 5.114
R2241 VDD.n1206 PA�U 5.114
R2242 VDD.n1131  5.114
R2243 VDD.n1056 VDD.t66 5.114
R2244 VDD.n981 @C6�U 5.114
R2245 VDD.n906  5.114
R2246 VDD.n830 �+���~ 5.114
R2247 VDD.n31 VDD.n30 4.65
R2248 VDD.n34 VDD.n33 4.65
R2249 VDD.n38 VDD.n37 4.65
R2250 VDD.n42 VDD.n41 4.65
R2251 VDD.n46 VDD.n45 4.65
R2252 VDD.n50 VDD.n49 4.65
R2253 VDD.n77 VDD.n76 4.65
R2254 VDD.n81 VDD.n80 4.65
R2255 VDD.n85 VDD.n84 4.65
R2256 VDD.n89 VDD.n88 4.65
R2257 VDD.n92 VDD.n91 4.65
R2258 VDD.n96 VDD.n95 4.65
R2259 VDD.n100 VDD.n99 4.65
R2260 VDD.n104 VDD.n103 4.65
R2261 VDD.n130 VDD.n129 4.65
R2262 VDD.n135 VDD.n134 4.65
R2263 VDD.n139 VDD.n138 4.65
R2264 VDD.n144 VDD.n143 4.65
R2265 VDD.n148 VDD.n147 4.65
R2266 VDD.n152 VDD.n151 4.65
R2267 VDD.n157 VDD.n156 4.65
R2268 VDD.n161 VDD.n160 4.65
R2269 VDD.n187 VDD.n186 4.65
R2270 VDD.n191 VDD.n190 4.65
R2271 VDD.n195 VDD.n194 4.65
R2272 VDD.n199 VDD.n198 4.65
R2273 VDD.n205 VDD.n204 4.65
R2274 VDD.n209 VDD.n208 4.65
R2275 VDD.n213 VDD.n212 4.65
R2276 VDD.n219 VDD.n218 4.65
R2277 VDD.n223 VDD.n222 4.65
R2278 VDD.n228 VDD.n227 4.65
R2279 VDD.n232 VDD.n231 4.65
R2280 VDD.n236 VDD.n235 4.65
R2281 VDD.n262 VDD.n261 4.65
R2282 VDD.n266 VDD.n265 4.65
R2283 VDD.n270 VDD.n269 4.65
R2284 VDD.n274 VDD.n273 4.65
R2285 VDD.n280 VDD.n279 4.65
R2286 VDD.n284 VDD.n283 4.65
R2287 VDD.n288 VDD.n287 4.65
R2288 VDD.n294 VDD.n293 4.65
R2289 VDD.n298 VDD.n297 4.65
R2290 VDD.n303 VDD.n302 4.65
R2291 VDD.n307 VDD.n306 4.65
R2292 VDD.n311 VDD.n310 4.65
R2293 VDD.n337 VDD.n336 4.65
R2294 VDD.n341 VDD.n340 4.65
R2295 VDD.n345 VDD.n344 4.65
R2296 VDD.n349 VDD.n348 4.65
R2297 VDD.n355 VDD.n354 4.65
R2298 VDD.n359 VDD.n358 4.65
R2299 VDD.n363 VDD.n362 4.65
R2300 VDD.n369 VDD.n368 4.65
R2301 VDD.n373 VDD.n372 4.65
R2302 VDD.n378 VDD.n377 4.65
R2303 VDD.n382 VDD.n381 4.65
R2304 VDD.n386 VDD.n385 4.65
R2305 VDD.n412 VDD.n411 4.65
R2306 VDD.n416 VDD.n415 4.65
R2307 VDD.n420 VDD.n419 4.65
R2308 VDD.n424 VDD.n423 4.65
R2309 VDD.n430 VDD.n429 4.65
R2310 VDD.n434 VDD.n433 4.65
R2311 VDD.n438 VDD.n437 4.65
R2312 VDD.n444 VDD.n443 4.65
R2313 VDD.n448 VDD.n447 4.65
R2314 VDD.n453 VDD.n452 4.65
R2315 VDD.n457 VDD.n456 4.65
R2316 VDD.n461 VDD.n460 4.65
R2317 VDD.n487 VDD.n486 4.65
R2318 VDD.n491 VDD.n490 4.65
R2319 VDD.n495 VDD.n494 4.65
R2320 VDD.n499 VDD.n498 4.65
R2321 VDD.n505 VDD.n504 4.65
R2322 VDD.n509 VDD.n508 4.65
R2323 VDD.n513 VDD.n512 4.65
R2324 VDD.n519 VDD.n518 4.65
R2325 VDD.n523 VDD.n522 4.65
R2326 VDD.n528 VDD.n527 4.65
R2327 VDD.n532 VDD.n531 4.65
R2328 VDD.n536 VDD.n535 4.65
R2329 VDD.n562 VDD.n561 4.65
R2330 VDD.n566 VDD.n565 4.65
R2331 VDD.n570 VDD.n569 4.65
R2332 VDD.n574 VDD.n573 4.65
R2333 VDD.n580 VDD.n579 4.65
R2334 VDD.n584 VDD.n583 4.65
R2335 VDD.n588 VDD.n587 4.65
R2336 VDD.n594 VDD.n593 4.65
R2337 VDD.n598 VDD.n597 4.65
R2338 VDD.n603 VDD.n602 4.65
R2339 VDD.n607 VDD.n606 4.65
R2340 VDD.n611 VDD.n610 4.65
R2341 VDD.n637 VDD.n636 4.65
R2342 VDD.n641 VDD.n640 4.65
R2343 VDD.n645 VDD.n644 4.65
R2344 VDD.n649 VDD.n648 4.65
R2345 VDD.n655 VDD.n654 4.65
R2346 VDD.n659 VDD.n658 4.65
R2347 VDD.n663 VDD.n662 4.65
R2348 VDD.n669 VDD.n668 4.65
R2349 VDD.n673 VDD.n672 4.65
R2350 VDD.n678 VDD.n677 4.65
R2351 VDD.n682 VDD.n681 4.65
R2352 VDD.n686 VDD.n685 4.65
R2353 VDD.n712 VDD.n711 4.65
R2354 VDD.n716 VDD.n715 4.65
R2355 VDD.n720 VDD.n719 4.65
R2356 VDD.n724 VDD.n723 4.65
R2357 VDD.n730 VDD.n729 4.65
R2358 VDD.n734 VDD.n733 4.65
R2359 VDD.n738 VDD.n737 4.65
R2360 VDD.n744 VDD.n743 4.65
R2361 VDD.n748 VDD.n747 4.65
R2362 VDD.n753 VDD.n752 4.65
R2363 VDD.n757 VDD.n756 4.65
R2364 VDD.n783 VDD.n782 4.65
R2365 VDD.n1531 VDD.n1530 4.65
R2366 VDD.n1527 VDD.n1526 4.65
R2367 VDD.n1523 VDD.n1522 4.65
R2368 VDD.n1519 VDD.n1518 4.65
R2369 VDD.n1515 VDD.n1514 4.65
R2370 VDD.n1509 VDD.n1508 4.65
R2371 VDD.n1505 VDD.n1504 4.65
R2372 VDD.n1501 VDD.n1500 4.65
R2373 VDD.n1495 VDD.n1494 4.65
R2374 VDD.n1491 VDD.n1490 4.65
R2375 VDD.n1486 VDD.n1485 4.65
R2376 VDD.n1482 VDD.n1481 4.65
R2377 VDD.n1456 VDD.n1455 4.65
R2378 VDD.n1452 VDD.n1451 4.65
R2379 VDD.n1448 VDD.n1447 4.65
R2380 VDD.n1444 VDD.n1443 4.65
R2381 VDD.n1440 VDD.n1439 4.65
R2382 VDD.n1434 VDD.n1433 4.65
R2383 VDD.n1430 VDD.n1429 4.65
R2384 VDD.n1426 VDD.n1425 4.65
R2385 VDD.n1420 VDD.n1419 4.65
R2386 VDD.n1416 VDD.n1415 4.65
R2387 VDD.n1411 VDD.n1410 4.65
R2388 VDD.n1407 VDD.n1406 4.65
R2389 VDD.n1381 VDD.n1380 4.65
R2390 VDD.n1377 VDD.n1376 4.65
R2391 VDD.n1373 VDD.n1372 4.65
R2392 VDD.n1369 VDD.n1368 4.65
R2393 VDD.n1365 VDD.n1364 4.65
R2394 VDD.n1359 VDD.n1358 4.65
R2395 VDD.n1355 VDD.n1354 4.65
R2396 VDD.n1351 VDD.n1350 4.65
R2397 VDD.n1345 VDD.n1344 4.65
R2398 VDD.n1341 VDD.n1340 4.65
R2399 VDD.n1336 VDD.n1335 4.65
R2400 VDD.n1332 VDD.n1331 4.65
R2401 VDD.n1306 VDD.n1305 4.65
R2402 VDD.n1302 VDD.n1301 4.65
R2403 VDD.n1298 VDD.n1297 4.65
R2404 VDD.n1294 VDD.n1293 4.65
R2405 VDD.n1290 VDD.n1289 4.65
R2406 VDD.n1284 VDD.n1283 4.65
R2407 VDD.n1280 VDD.n1279 4.65
R2408 VDD.n1276 VDD.n1275 4.65
R2409 VDD.n1270 VDD.n1269 4.65
R2410 VDD.n1266 VDD.n1265 4.65
R2411 VDD.n1261 VDD.n1260 4.65
R2412 VDD.n1257 VDD.n1256 4.65
R2413 VDD.n1231 VDD.n1230 4.65
R2414 VDD.n1227 VDD.n1226 4.65
R2415 VDD.n1223 VDD.n1222 4.65
R2416 VDD.n1219 VDD.n1218 4.65
R2417 VDD.n1215 VDD.n1214 4.65
R2418 VDD.n1209 VDD.n1208 4.65
R2419 VDD.n1205 VDD.n1204 4.65
R2420 VDD.n1201 VDD.n1200 4.65
R2421 VDD.n1195 VDD.n1194 4.65
R2422 VDD.n1191 VDD.n1190 4.65
R2423 VDD.n1186 VDD.n1185 4.65
R2424 VDD.n1182 VDD.n1181 4.65
R2425 VDD.n1156 VDD.n1155 4.65
R2426 VDD.n1152 VDD.n1151 4.65
R2427 VDD.n1148 VDD.n1147 4.65
R2428 VDD.n1144 VDD.n1143 4.65
R2429 VDD.n1140 VDD.n1139 4.65
R2430 VDD.n1134 VDD.n1133 4.65
R2431 VDD.n1130 VDD.n1129 4.65
R2432 VDD.n1126 VDD.n1125 4.65
R2433 VDD.n1120 VDD.n1119 4.65
R2434 VDD.n1116 VDD.n1115 4.65
R2435 VDD.n1111 VDD.n1110 4.65
R2436 VDD.n1107 VDD.n1106 4.65
R2437 VDD.n1081 VDD.n1080 4.65
R2438 VDD.n1077 VDD.n1076 4.65
R2439 VDD.n1073 VDD.n1072 4.65
R2440 VDD.n1069 VDD.n1068 4.65
R2441 VDD.n1065 VDD.n1064 4.65
R2442 VDD.n1059 VDD.n1058 4.65
R2443 VDD.n1055 VDD.n1054 4.65
R2444 VDD.n1051 VDD.n1050 4.65
R2445 VDD.n1045 VDD.n1044 4.65
R2446 VDD.n1041 VDD.n1040 4.65
R2447 VDD.n1036 VDD.n1035 4.65
R2448 VDD.n1032 VDD.n1031 4.65
R2449 VDD.n1006 VDD.n1005 4.65
R2450 VDD.n1002 VDD.n1001 4.65
R2451 VDD.n998 VDD.n997 4.65
R2452 VDD.n994 VDD.n993 4.65
R2453 VDD.n990 VDD.n989 4.65
R2454 VDD.n984 VDD.n983 4.65
R2455 VDD.n980 VDD.n979 4.65
R2456 VDD.n976 VDD.n975 4.65
R2457 VDD.n970 VDD.n969 4.65
R2458 VDD.n966 VDD.n965 4.65
R2459 VDD.n961 VDD.n960 4.65
R2460 VDD.n957 VDD.n956 4.65
R2461 VDD.n931 VDD.n930 4.65
R2462 VDD.n927 VDD.n926 4.65
R2463 VDD.n923 VDD.n922 4.65
R2464 VDD.n919 VDD.n918 4.65
R2465 VDD.n915 VDD.n914 4.65
R2466 VDD.n909 VDD.n908 4.65
R2467 VDD.n905 VDD.n904 4.65
R2468 VDD.n901 VDD.n900 4.65
R2469 VDD.n895 VDD.n894 4.65
R2470 VDD.n891 VDD.n890 4.65
R2471 VDD.n886 VDD.n885 4.65
R2472 VDD.n882 VDD.n881 4.65
R2473 VDD.n855 VDD.n854 4.65
R2474 VDD.n851 VDD.n850 4.65
R2475 VDD.n847 VDD.n846 4.65
R2476 VDD.n843 VDD.n842 4.65
R2477 VDD.n839 VDD.n838 4.65
R2478 VDD.n833 VDD.n832 4.65
R2479 VDD.n829 VDD.n828 4.65
R2480 VDD.n825 VDD.n824 4.65
R2481 VDD.n819 VDD.n818 4.65
R2482 VDD.n815 VDD.n814 4.65
R2483 VDD.n810 VDD.n809 4.65
R2484 VDD.n806 VDD.n805 4.65
R2485 VDD.n27 VDD.n23 2.933
R2486 VDD.n156 VDD.n153 2.89
R2487 VDD.n27 VDD.n26 2.844
R2488 VDD.n35 @�-�U 2.557
R2489 VDD.n86 �+���~ 2.557
R2490 VDD.n145  2.557
R2491 VDD.n134 VDD.n131 2.477
R2492 VDD.n31 VDD.n27 1.063
R2493 VDD.n227 VDD.n224 0.412
R2494 VDD.n302 VDD.n299 0.412
R2495 VDD.n377 VDD.n374 0.412
R2496 VDD.n452 VDD.n449 0.412
R2497 VDD.n527 VDD.n524 0.412
R2498 VDD.n602 VDD.n599 0.412
R2499 VDD.n677 VDD.n674 0.412
R2500 VDD.n752 VDD.n749 0.412
R2501 VDD.n1490 VDD.n1487 0.412
R2502 VDD.n1415 VDD.n1412 0.412
R2503 VDD.n1340 VDD.n1337 0.412
R2504 VDD.n1265 VDD.n1262 0.412
R2505 VDD.n1190 VDD.n1187 0.412
R2506 VDD.n1115 VDD.n1112 0.412
R2507 VDD.n1040 VDD.n1037 0.412
R2508 VDD.n965 VDD.n962 0.412
R2509 VDD.n890 VDD.n887 0.412
R2510 VDD.n814 VDD.n811 0.412
R2511 VDD.n77 VDD.n50 0.29
R2512 VDD.n130 VDD.n104 0.29
R2513 VDD.n187 VDD.n161 0.29
R2514 VDD.n262 VDD.n236 0.29
R2515 VDD.n337 VDD.n311 0.29
R2516 VDD.n412 VDD.n386 0.29
R2517 VDD.n487 VDD.n461 0.29
R2518 VDD.n562 VDD.n536 0.29
R2519 VDD.n637 VDD.n611 0.29
R2520 VDD.n712 VDD.n686 0.29
R2521 VDD.n1482 VDD.n1456 0.29
R2522 VDD.n1407 VDD.n1381 0.29
R2523 VDD.n1332 VDD.n1306 0.29
R2524 VDD.n1257 VDD.n1231 0.29
R2525 VDD.n1182 VDD.n1156 0.29
R2526 VDD.n1107 VDD.n1081 0.29
R2527 VDD.n1032 VDD.n1006 0.29
R2528 VDD.n957 VDD.n931 0.29
R2529 VDD.n882 VDD.n855 0.29
R2530 VDD VDD.n1531 0.219
R2531 VDD.n806 VDD 0.207
R2532 VDD.n213 VDD.n209 0.197
R2533 VDD.n288 VDD.n284 0.197
R2534 VDD.n363 VDD.n359 0.197
R2535 VDD.n438 VDD.n434 0.197
R2536 VDD.n513 VDD.n509 0.197
R2537 VDD.n588 VDD.n584 0.197
R2538 VDD.n663 VDD.n659 0.197
R2539 VDD.n738 VDD.n734 0.197
R2540 VDD.n1509 VDD.n1505 0.197
R2541 VDD.n1434 VDD.n1430 0.197
R2542 VDD.n1359 VDD.n1355 0.197
R2543 VDD.n1284 VDD.n1280 0.197
R2544 VDD.n1209 VDD.n1205 0.197
R2545 VDD.n1134 VDD.n1130 0.197
R2546 VDD.n1059 VDD.n1055 0.197
R2547 VDD.n984 VDD.n980 0.197
R2548 VDD.n909 VDD.n905 0.197
R2549 VDD.n833 VDD.n829 0.197
R2550 VDD.n38 VDD.n34 0.181
R2551 VDD.n92 VDD.n89 0.181
R2552 VDD.n148 VDD.n144 0.181
R2553 VDD.n34 VDD.n31 0.145
R2554 VDD.n42 VDD.n38 0.145
R2555 VDD.n46 VDD.n42 0.145
R2556 VDD.n50 VDD.n46 0.145
R2557 VDD.n81 VDD.n77 0.145
R2558 VDD.n85 VDD.n81 0.145
R2559 VDD.n89 VDD.n85 0.145
R2560 VDD.n96 VDD.n92 0.145
R2561 VDD.n100 VDD.n96 0.145
R2562 VDD.n104 VDD.n100 0.145
R2563 VDD.n135 VDD.n130 0.145
R2564 VDD.n139 VDD.n135 0.145
R2565 VDD.n144 VDD.n139 0.145
R2566 VDD.n152 VDD.n148 0.145
R2567 VDD.n157 VDD.n152 0.145
R2568 VDD.n161 VDD.n157 0.145
R2569 VDD.n191 VDD.n187 0.145
R2570 VDD.n195 VDD.n191 0.145
R2571 VDD.n199 VDD.n195 0.145
R2572 VDD.n205 VDD.n199 0.145
R2573 VDD.n209 VDD.n205 0.145
R2574 VDD.n219 VDD.n213 0.145
R2575 VDD.n223 VDD.n219 0.145
R2576 VDD.n228 VDD.n223 0.145
R2577 VDD.n232 VDD.n228 0.145
R2578 VDD.n236 VDD.n232 0.145
R2579 VDD.n266 VDD.n262 0.145
R2580 VDD.n270 VDD.n266 0.145
R2581 VDD.n274 VDD.n270 0.145
R2582 VDD.n280 VDD.n274 0.145
R2583 VDD.n284 VDD.n280 0.145
R2584 VDD.n294 VDD.n288 0.145
R2585 VDD.n298 VDD.n294 0.145
R2586 VDD.n303 VDD.n298 0.145
R2587 VDD.n307 VDD.n303 0.145
R2588 VDD.n311 VDD.n307 0.145
R2589 VDD.n341 VDD.n337 0.145
R2590 VDD.n345 VDD.n341 0.145
R2591 VDD.n349 VDD.n345 0.145
R2592 VDD.n355 VDD.n349 0.145
R2593 VDD.n359 VDD.n355 0.145
R2594 VDD.n369 VDD.n363 0.145
R2595 VDD.n373 VDD.n369 0.145
R2596 VDD.n378 VDD.n373 0.145
R2597 VDD.n382 VDD.n378 0.145
R2598 VDD.n386 VDD.n382 0.145
R2599 VDD.n416 VDD.n412 0.145
R2600 VDD.n420 VDD.n416 0.145
R2601 VDD.n424 VDD.n420 0.145
R2602 VDD.n430 VDD.n424 0.145
R2603 VDD.n434 VDD.n430 0.145
R2604 VDD.n444 VDD.n438 0.145
R2605 VDD.n448 VDD.n444 0.145
R2606 VDD.n453 VDD.n448 0.145
R2607 VDD.n457 VDD.n453 0.145
R2608 VDD.n461 VDD.n457 0.145
R2609 VDD.n491 VDD.n487 0.145
R2610 VDD.n495 VDD.n491 0.145
R2611 VDD.n499 VDD.n495 0.145
R2612 VDD.n505 VDD.n499 0.145
R2613 VDD.n509 VDD.n505 0.145
R2614 VDD.n519 VDD.n513 0.145
R2615 VDD.n523 VDD.n519 0.145
R2616 VDD.n528 VDD.n523 0.145
R2617 VDD.n532 VDD.n528 0.145
R2618 VDD.n536 VDD.n532 0.145
R2619 VDD.n566 VDD.n562 0.145
R2620 VDD.n570 VDD.n566 0.145
R2621 VDD.n574 VDD.n570 0.145
R2622 VDD.n580 VDD.n574 0.145
R2623 VDD.n584 VDD.n580 0.145
R2624 VDD.n594 VDD.n588 0.145
R2625 VDD.n598 VDD.n594 0.145
R2626 VDD.n603 VDD.n598 0.145
R2627 VDD.n607 VDD.n603 0.145
R2628 VDD.n611 VDD.n607 0.145
R2629 VDD.n641 VDD.n637 0.145
R2630 VDD.n645 VDD.n641 0.145
R2631 VDD.n649 VDD.n645 0.145
R2632 VDD.n655 VDD.n649 0.145
R2633 VDD.n659 VDD.n655 0.145
R2634 VDD.n669 VDD.n663 0.145
R2635 VDD.n673 VDD.n669 0.145
R2636 VDD.n678 VDD.n673 0.145
R2637 VDD.n682 VDD.n678 0.145
R2638 VDD.n686 VDD.n682 0.145
R2639 VDD.n716 VDD.n712 0.145
R2640 VDD.n720 VDD.n716 0.145
R2641 VDD.n724 VDD.n720 0.145
R2642 VDD.n730 VDD.n724 0.145
R2643 VDD.n734 VDD.n730 0.145
R2644 VDD.n744 VDD.n738 0.145
R2645 VDD.n748 VDD.n744 0.145
R2646 VDD.n753 VDD.n748 0.145
R2647 VDD.n757 VDD.n753 0.145
R2648 VDD.n783 VDD.n757 0.145
R2649 VDD.n1531 VDD.n1527 0.145
R2650 VDD.n1527 VDD.n1523 0.145
R2651 VDD.n1523 VDD.n1519 0.145
R2652 VDD.n1519 VDD.n1515 0.145
R2653 VDD.n1515 VDD.n1509 0.145
R2654 VDD.n1505 VDD.n1501 0.145
R2655 VDD.n1501 VDD.n1495 0.145
R2656 VDD.n1495 VDD.n1491 0.145
R2657 VDD.n1491 VDD.n1486 0.145
R2658 VDD.n1486 VDD.n1482 0.145
R2659 VDD.n1456 VDD.n1452 0.145
R2660 VDD.n1452 VDD.n1448 0.145
R2661 VDD.n1448 VDD.n1444 0.145
R2662 VDD.n1444 VDD.n1440 0.145
R2663 VDD.n1440 VDD.n1434 0.145
R2664 VDD.n1430 VDD.n1426 0.145
R2665 VDD.n1426 VDD.n1420 0.145
R2666 VDD.n1420 VDD.n1416 0.145
R2667 VDD.n1416 VDD.n1411 0.145
R2668 VDD.n1411 VDD.n1407 0.145
R2669 VDD.n1381 VDD.n1377 0.145
R2670 VDD.n1377 VDD.n1373 0.145
R2671 VDD.n1373 VDD.n1369 0.145
R2672 VDD.n1369 VDD.n1365 0.145
R2673 VDD.n1365 VDD.n1359 0.145
R2674 VDD.n1355 VDD.n1351 0.145
R2675 VDD.n1351 VDD.n1345 0.145
R2676 VDD.n1345 VDD.n1341 0.145
R2677 VDD.n1341 VDD.n1336 0.145
R2678 VDD.n1336 VDD.n1332 0.145
R2679 VDD.n1306 VDD.n1302 0.145
R2680 VDD.n1302 VDD.n1298 0.145
R2681 VDD.n1298 VDD.n1294 0.145
R2682 VDD.n1294 VDD.n1290 0.145
R2683 VDD.n1290 VDD.n1284 0.145
R2684 VDD.n1280 VDD.n1276 0.145
R2685 VDD.n1276 VDD.n1270 0.145
R2686 VDD.n1270 VDD.n1266 0.145
R2687 VDD.n1266 VDD.n1261 0.145
R2688 VDD.n1261 VDD.n1257 0.145
R2689 VDD.n1231 VDD.n1227 0.145
R2690 VDD.n1227 VDD.n1223 0.145
R2691 VDD.n1223 VDD.n1219 0.145
R2692 VDD.n1219 VDD.n1215 0.145
R2693 VDD.n1215 VDD.n1209 0.145
R2694 VDD.n1205 VDD.n1201 0.145
R2695 VDD.n1201 VDD.n1195 0.145
R2696 VDD.n1195 VDD.n1191 0.145
R2697 VDD.n1191 VDD.n1186 0.145
R2698 VDD.n1186 VDD.n1182 0.145
R2699 VDD.n1156 VDD.n1152 0.145
R2700 VDD.n1152 VDD.n1148 0.145
R2701 VDD.n1148 VDD.n1144 0.145
R2702 VDD.n1144 VDD.n1140 0.145
R2703 VDD.n1140 VDD.n1134 0.145
R2704 VDD.n1130 VDD.n1126 0.145
R2705 VDD.n1126 VDD.n1120 0.145
R2706 VDD.n1120 VDD.n1116 0.145
R2707 VDD.n1116 VDD.n1111 0.145
R2708 VDD.n1111 VDD.n1107 0.145
R2709 VDD.n1081 VDD.n1077 0.145
R2710 VDD.n1077 VDD.n1073 0.145
R2711 VDD.n1073 VDD.n1069 0.145
R2712 VDD.n1069 VDD.n1065 0.145
R2713 VDD.n1065 VDD.n1059 0.145
R2714 VDD.n1055 VDD.n1051 0.145
R2715 VDD.n1051 VDD.n1045 0.145
R2716 VDD.n1045 VDD.n1041 0.145
R2717 VDD.n1041 VDD.n1036 0.145
R2718 VDD.n1036 VDD.n1032 0.145
R2719 VDD.n1006 VDD.n1002 0.145
R2720 VDD.n1002 VDD.n998 0.145
R2721 VDD.n998 VDD.n994 0.145
R2722 VDD.n994 VDD.n990 0.145
R2723 VDD.n990 VDD.n984 0.145
R2724 VDD.n980 VDD.n976 0.145
R2725 VDD.n976 VDD.n970 0.145
R2726 VDD.n970 VDD.n966 0.145
R2727 VDD.n966 VDD.n961 0.145
R2728 VDD.n961 VDD.n957 0.145
R2729 VDD.n931 VDD.n927 0.145
R2730 VDD.n927 VDD.n923 0.145
R2731 VDD.n923 VDD.n919 0.145
R2732 VDD.n919 VDD.n915 0.145
R2733 VDD.n915 VDD.n909 0.145
R2734 VDD.n905 VDD.n901 0.145
R2735 VDD.n901 VDD.n895 0.145
R2736 VDD.n895 VDD.n891 0.145
R2737 VDD.n891 VDD.n886 0.145
R2738 VDD.n886 VDD.n882 0.145
R2739 VDD.n855 VDD.n851 0.145
R2740 VDD.n851 VDD.n847 0.145
R2741 VDD.n847 VDD.n843 0.145
R2742 VDD.n843 VDD.n839 0.145
R2743 VDD.n839 VDD.n833 0.145
R2744 VDD.n829 VDD.n825 0.145
R2745 VDD.n825 VDD.n819 0.145
R2746 VDD.n819 VDD.n815 0.145
R2747 VDD.n815 VDD.n810 0.145
R2748 VDD.n810 VDD.n806 0.145
R2749 VDD VDD.n783 0.07
R2750 CLK.n18 CLK.t14 459.505
R2751 CLK.n15 CLK.t1 459.505
R2752 CLK.n12 CLK.t17 459.505
R2753 CLK.n7 CLK.t11 459.505
R2754 CLK.n4 CLK.t3 459.505
R2755 CLK.n0 CLK.t12 459.505
R2756 CLK.n16 CLK.t6 399.181
R2757 CLK.n8 CLK.t9 399.181
R2758 CLK.n1 CLK.t13 399.181
R2759 CLK.n20 CLK.t5 398.835
R2760 CLK.n10 CLK.t4 397.657
R2761 CLK.n2 CLK.t15 397.657
R2762 CLK.n18 CLK.t0 384.527
R2763 CLK.n15 CLK.t8 384.527
R2764 CLK.n12 CLK.t10 384.527
R2765 CLK.n7 CLK.t2 384.527
R2766 CLK.n4 CLK.t7 384.527
R2767 CLK.n0 CLK.t16 384.527
R2768 CLK.n1 CLK.n0 33.832
R2769 CLK.n8 CLK.n7 33.832
R2770 CLK.n16 CLK.n15 33.832
R2771 CLK.n19 CLK.n18 30.851
R2772 CLK.n13 CLK.n12 30.851
R2773 CLK.n5 CLK.n4 30.851
R2774 CLK.n9 CLK.n6 14.075
R2775 CLK.n17 CLK.n14 14.075
R2776 CLK.n19 CLK 9.3
R2777 CLK.n3 CLK.n1 9.111
R2778 CLK.n11 CLK.n9 7.032
R2779 CLK.n21 CLK.n17 7.032
R2780 CLK.n6 CLK.n5 4.639
R2781 CLK.n14 CLK.n13 4.639
R2782 CLK.n3 CLK.n2 4.234
R2783 CLK.n11 CLK.n10 4.234
R2784 CLK.n20 CLK.n19 2.59
R2785 CLK.n21 CLK.n20 2.1
R2786 CLK.n9 CLK.n8 2.079
R2787 CLK.n17 CLK.n16 2.079
R2788 CLK.n21 CLK 0.046
R2789 CLK.n6 CLK.n3 0.023
R2790 CLK.n14 CLK.n11 0.023
R2791 a_599_989.n1 a_599_989.t12 512.525
R2792 a_599_989.n3 a_599_989.t11 454.685
R2793 a_599_989.n3 a_599_989.t9 428.979
R2794 a_599_989.n1 a_599_989.t8 371.139
R2795 a_599_989.n2 a_599_989.t7 361.392
R2796 a_599_989.n7 a_599_989.n6 329.955
R2797 a_599_989.n4 a_599_989.t10 311.683
R2798 a_599_989.n2 a_599_989.n1 235.554
R2799 a_599_989.n8 a_599_989.n7 179.199
R2800 a_599_989.n4 a_599_989.n3 171.288
R2801 a_599_989.n10 a_599_989.n9 161.352
R2802 a_599_989.n8 a_599_989.n0 95.095
R2803 a_599_989.n11 a_599_989.n10 95.094
R2804 a_599_989.n10 a_599_989.n8 66.258
R2805 a_599_989.n0 a_599_989.t1 14.282
R2806 a_599_989.n0 a_599_989.t3 14.282
R2807 a_599_989.n9 a_599_989.t6 14.282
R2808 a_599_989.n9 a_599_989.t2 14.282
R2809 a_599_989.n11 a_599_989.t4 14.282
R2810 a_599_989.t5 a_599_989.n11 14.282
R2811 a_599_989.n5 a_599_989.n2 13.038
R2812 a_599_989.n5 a_599_989.n4 8.685
R2813 a_599_989.n7 a_599_989.n5 4.65
R2814 a_9897_1050.n1 a_9897_1050.t7 512.525
R2815 a_9897_1050.n1 a_9897_1050.t9 371.139
R2816 a_9897_1050.n2 a_9897_1050.t8 361.392
R2817 a_9897_1050.n4 a_9897_1050.n3 329.955
R2818 a_9897_1050.n2 a_9897_1050.n1 235.554
R2819 a_9897_1050.n5 a_9897_1050.n4 179.199
R2820 a_9897_1050.n7 a_9897_1050.n6 161.352
R2821 a_9897_1050.n5 a_9897_1050.n0 95.095
R2822 a_9897_1050.n8 a_9897_1050.n7 95.094
R2823 a_9897_1050.n7 a_9897_1050.n5 66.258
R2824 a_9897_1050.n0 a_9897_1050.t2 14.282
R2825 a_9897_1050.n0 a_9897_1050.t3 14.282
R2826 a_9897_1050.n6 a_9897_1050.t0 14.282
R2827 a_9897_1050.n6 a_9897_1050.t4 14.282
R2828 a_9897_1050.t6 a_9897_1050.n8 14.282
R2829 a_9897_1050.n8 a_9897_1050.t5 14.282
R2830 a_9897_1050.n4 a_9897_1050.n2 10.615
R2831 a_3939_103.n5 a_3939_103.n4 66.708
R2832 a_3939_103.n2 a_3939_103.n0 32.662
R2833 a_3939_103.n5 a_3939_103.n3 19.496
R2834 a_3939_103.t0 a_3939_103.n5 13.756
R2835 a_3939_103.t0 a_3939_103.n2 3.034
R2836 a_3939_103.n2 a_3939_103.n1 0.443
R2837 a_1561_989.n3 a_1561_989.t12 454.685
R2838 a_1561_989.n5 a_1561_989.t7 454.685
R2839 a_1561_989.n1 a_1561_989.t15 454.685
R2840 a_1561_989.n3 a_1561_989.t8 428.979
R2841 a_1561_989.n5 a_1561_989.t9 428.979
R2842 a_1561_989.n1 a_1561_989.t10 428.979
R2843 a_1561_989.n4 a_1561_989.t11 339.542
R2844 a_1561_989.n2 a_1561_989.t14 339.542
R2845 a_1561_989.n6 a_1561_989.t13 339.186
R2846 a_1561_989.n13 a_1561_989.n12 336.075
R2847 a_1561_989.n16 a_1561_989.n15 161.352
R2848 a_1561_989.n14 a_1561_989.n13 151.34
R2849 a_1561_989.n4 a_1561_989.n3 143.429
R2850 a_1561_989.n2 a_1561_989.n1 143.429
R2851 a_1561_989.n6 a_1561_989.n5 143.074
R2852 a_1561_989.n14 a_1561_989.n0 95.095
R2853 a_1561_989.n17 a_1561_989.n16 95.094
R2854 a_1561_989.n16 a_1561_989.n14 66.258
R2855 a_1561_989.n12 a_1561_989.n11 30
R2856 a_1561_989.n10 a_1561_989.n9 24.383
R2857 a_1561_989.n12 a_1561_989.n10 23.684
R2858 a_1561_989.n0 a_1561_989.t6 14.282
R2859 a_1561_989.n0 a_1561_989.t5 14.282
R2860 a_1561_989.n15 a_1561_989.t0 14.282
R2861 a_1561_989.n15 a_1561_989.t3 14.282
R2862 a_1561_989.t2 a_1561_989.n17 14.282
R2863 a_1561_989.n17 a_1561_989.t1 14.282
R2864 a_1561_989.n8 a_1561_989.n2 11.134
R2865 a_1561_989.n7 a_1561_989.n6 8.145
R2866 a_1561_989.n7 a_1561_989.n4 4.65
R2867 a_1561_989.n13 a_1561_989.n8 4.65
R2868 a_1561_989.n8 a_1561_989.n7 4.035
R2869 a_12143_989.n1 a_12143_989.t12 512.525
R2870 a_12143_989.n3 a_12143_989.t7 454.685
R2871 a_12143_989.n3 a_12143_989.t10 428.979
R2872 a_12143_989.n1 a_12143_989.t8 371.139
R2873 a_12143_989.n2 a_12143_989.t9 361.392
R2874 a_12143_989.n4 a_12143_989.t11 311.683
R2875 a_12143_989.n10 a_12143_989.n9 308.216
R2876 a_12143_989.n2 a_12143_989.n1 235.554
R2877 a_12143_989.n11 a_12143_989.n10 179.199
R2878 a_12143_989.n4 a_12143_989.n3 171.288
R2879 a_12143_989.n13 a_12143_989.n12 161.352
R2880 a_12143_989.n11 a_12143_989.n0 95.095
R2881 a_12143_989.n14 a_12143_989.n13 95.094
R2882 a_12143_989.n13 a_12143_989.n11 66.258
R2883 a_12143_989.n9 a_12143_989.n8 30
R2884 a_12143_989.n7 a_12143_989.n6 24.383
R2885 a_12143_989.n9 a_12143_989.n7 23.684
R2886 a_12143_989.n0 a_12143_989.t6 14.282
R2887 a_12143_989.n0 a_12143_989.t5 14.282
R2888 a_12143_989.n12 a_12143_989.t0 14.282
R2889 a_12143_989.n12 a_12143_989.t1 14.282
R2890 a_12143_989.t3 a_12143_989.n14 14.282
R2891 a_12143_989.n14 a_12143_989.t2 14.282
R2892 a_12143_989.n5 a_12143_989.n2 13.038
R2893 a_12143_989.n5 a_12143_989.n4 8.685
R2894 a_12143_989.n10 a_12143_989.n5 4.65
R2895 a_11821_1050.n2 a_11821_1050.t11 512.525
R2896 a_11821_1050.n0 a_11821_1050.t9 512.525
R2897 a_11821_1050.n2 a_11821_1050.t7 371.139
R2898 a_11821_1050.n0 a_11821_1050.t12 371.139
R2899 a_11821_1050.n3 a_11821_1050.t8 306.051
R2900 a_11821_1050.n1 a_11821_1050.t10 306.051
R2901 a_11821_1050.n3 a_11821_1050.n2 290.895
R2902 a_11821_1050.n1 a_11821_1050.n0 290.895
R2903 a_11821_1050.n9 a_11821_1050.n8 252.875
R2904 a_11821_1050.n13 a_11821_1050.n9 234.54
R2905 a_11821_1050.n12 a_11821_1050.n11 161.352
R2906 a_11821_1050.n12 a_11821_1050.n10 95.095
R2907 a_11821_1050.n14 a_11821_1050.n13 95.094
R2908 a_11821_1050.n13 a_11821_1050.n12 66.258
R2909 a_11821_1050.n8 a_11821_1050.n7 30
R2910 a_11821_1050.n6 a_11821_1050.n5 24.383
R2911 a_11821_1050.n8 a_11821_1050.n6 23.684
R2912 a_11821_1050.n10 a_11821_1050.t6 14.282
R2913 a_11821_1050.n10 a_11821_1050.t5 14.282
R2914 a_11821_1050.n11 a_11821_1050.t1 14.282
R2915 a_11821_1050.n11 a_11821_1050.t0 14.282
R2916 a_11821_1050.n14 a_11821_1050.t3 14.282
R2917 a_11821_1050.t4 a_11821_1050.n14 14.282
R2918 a_11821_1050.n4 a_11821_1050.n1 8.141
R2919 a_11821_1050.n9 a_11821_1050.n4 5.965
R2920 a_11821_1050.n4 a_11821_1050.n3 4.65
R2921 a_9030_210.n12 a_9030_210.n10 171.558
R2922 a_9030_210.n7 a_9030_210.n6 117.622
R2923 a_9030_210.n5 a_9030_210.n4 92.5
R2924 a_9030_210.n9 a_9030_210.n8 92.5
R2925 a_9030_210.n10 a_9030_210.t1 75.764
R2926 a_9030_210.n5 a_9030_210.n3 65.02
R2927 a_9030_210.n7 a_9030_210.n5 36.517
R2928 a_9030_210.n3 a_9030_210.n2 35.865
R2929 a_9030_210.n12 a_9030_210.n11 27.2
R2930 a_9030_210.n13 a_9030_210.n0 23.498
R2931 a_9030_210.n13 a_9030_210.n12 22.4
R2932 a_9030_210.n9 a_9030_210.n7 19.952
R2933 a_9030_210.t1 a_9030_210.n1 7.04
R2934 a_9030_210.n10 a_9030_210.n9 1.505
R2935 a_7333_989.n3 a_7333_989.t8 454.685
R2936 a_7333_989.n5 a_7333_989.t10 454.685
R2937 a_7333_989.n1 a_7333_989.t9 454.685
R2938 a_7333_989.n3 a_7333_989.t14 428.979
R2939 a_7333_989.n5 a_7333_989.t7 428.979
R2940 a_7333_989.n1 a_7333_989.t11 428.979
R2941 a_7333_989.n10 a_7333_989.n9 357.814
R2942 a_7333_989.n4 a_7333_989.t13 339.542
R2943 a_7333_989.n2 a_7333_989.t15 339.542
R2944 a_7333_989.n6 a_7333_989.t12 339.186
R2945 a_7333_989.n13 a_7333_989.n12 161.352
R2946 a_7333_989.n11 a_7333_989.n10 151.34
R2947 a_7333_989.n4 a_7333_989.n3 143.429
R2948 a_7333_989.n2 a_7333_989.n1 143.429
R2949 a_7333_989.n6 a_7333_989.n5 143.074
R2950 a_7333_989.n11 a_7333_989.n0 95.095
R2951 a_7333_989.n14 a_7333_989.n13 95.094
R2952 a_7333_989.n13 a_7333_989.n11 66.258
R2953 a_7333_989.n0 a_7333_989.t6 14.282
R2954 a_7333_989.n0 a_7333_989.t5 14.282
R2955 a_7333_989.n12 a_7333_989.t0 14.282
R2956 a_7333_989.n12 a_7333_989.t1 14.282
R2957 a_7333_989.n14 a_7333_989.t2 14.282
R2958 a_7333_989.t3 a_7333_989.n14 14.282
R2959 a_7333_989.n8 a_7333_989.n2 11.134
R2960 a_7333_989.n7 a_7333_989.n6 8.145
R2961 a_7333_989.n7 a_7333_989.n4 4.65
R2962 a_7333_989.n10 a_7333_989.n8 4.65
R2963 a_7333_989.n8 a_7333_989.n7 4.035
R2964 a_13745_1050.n2 a_13745_1050.t7 512.525
R2965 a_13745_1050.n2 a_13745_1050.t9 371.139
R2966 a_13745_1050.n3 a_13745_1050.t8 305.674
R2967 a_13745_1050.n3 a_13745_1050.n2 291.272
R2968 a_13745_1050.n8 a_13745_1050.n7 252.498
R2969 a_13745_1050.n9 a_13745_1050.n8 234.917
R2970 a_13745_1050.n11 a_13745_1050.n10 161.352
R2971 a_13745_1050.n9 a_13745_1050.n1 95.095
R2972 a_13745_1050.n10 a_13745_1050.n0 95.095
R2973 a_13745_1050.n10 a_13745_1050.n9 66.258
R2974 a_13745_1050.n7 a_13745_1050.n6 30
R2975 a_13745_1050.n5 a_13745_1050.n4 24.383
R2976 a_13745_1050.n7 a_13745_1050.n5 23.684
R2977 a_13745_1050.n1 a_13745_1050.t5 14.282
R2978 a_13745_1050.n1 a_13745_1050.t4 14.282
R2979 a_13745_1050.n0 a_13745_1050.t6 14.282
R2980 a_13745_1050.n0 a_13745_1050.t0 14.282
R2981 a_13745_1050.t2 a_13745_1050.n11 14.282
R2982 a_13745_1050.n11 a_13745_1050.t1 14.282
R2983 a_13745_1050.n8 a_13745_1050.n3 10.615
R2984 a_277_1050.n2 a_277_1050.t8 512.525
R2985 a_277_1050.n0 a_277_1050.t7 512.525
R2986 a_277_1050.n2 a_277_1050.t9 371.139
R2987 a_277_1050.n0 a_277_1050.t10 371.139
R2988 a_277_1050.n3 a_277_1050.t12 306.051
R2989 a_277_1050.n1 a_277_1050.t11 306.051
R2990 a_277_1050.n3 a_277_1050.n2 290.895
R2991 a_277_1050.n1 a_277_1050.n0 290.895
R2992 a_277_1050.n9 a_277_1050.n8 252.875
R2993 a_277_1050.n13 a_277_1050.n9 234.54
R2994 a_277_1050.n12 a_277_1050.n11 161.352
R2995 a_277_1050.n12 a_277_1050.n10 95.095
R2996 a_277_1050.n14 a_277_1050.n13 95.094
R2997 a_277_1050.n13 a_277_1050.n12 66.258
R2998 a_277_1050.n8 a_277_1050.n7 30
R2999 a_277_1050.n6 a_277_1050.n5 24.383
R3000 a_277_1050.n8 a_277_1050.n6 23.684
R3001 a_277_1050.n10 a_277_1050.t6 14.282
R3002 a_277_1050.n10 a_277_1050.t5 14.282
R3003 a_277_1050.n11 a_277_1050.t1 14.282
R3004 a_277_1050.n11 a_277_1050.t0 14.282
R3005 a_277_1050.t4 a_277_1050.n14 14.282
R3006 a_277_1050.n14 a_277_1050.t3 14.282
R3007 a_277_1050.n4 a_277_1050.n1 8.141
R3008 a_277_1050.n9 a_277_1050.n4 5.965
R3009 a_277_1050.n4 a_277_1050.n3 4.65
R3010 a_2201_1050.n2 a_2201_1050.t9 512.525
R3011 a_2201_1050.n2 a_2201_1050.t7 371.139
R3012 a_2201_1050.n3 a_2201_1050.t8 305.674
R3013 a_2201_1050.n3 a_2201_1050.n2 291.272
R3014 a_2201_1050.n8 a_2201_1050.n7 252.498
R3015 a_2201_1050.n9 a_2201_1050.n8 234.917
R3016 a_2201_1050.n11 a_2201_1050.n10 161.352
R3017 a_2201_1050.n9 a_2201_1050.n1 95.095
R3018 a_2201_1050.n10 a_2201_1050.n0 95.095
R3019 a_2201_1050.n10 a_2201_1050.n9 66.258
R3020 a_2201_1050.n7 a_2201_1050.n6 30
R3021 a_2201_1050.n5 a_2201_1050.n4 24.383
R3022 a_2201_1050.n7 a_2201_1050.n5 23.684
R3023 a_2201_1050.n1 a_2201_1050.t5 14.282
R3024 a_2201_1050.n1 a_2201_1050.t4 14.282
R3025 a_2201_1050.n0 a_2201_1050.t0 14.282
R3026 a_2201_1050.n0 a_2201_1050.t6 14.282
R3027 a_2201_1050.t2 a_2201_1050.n11 14.282
R3028 a_2201_1050.n11 a_2201_1050.t1 14.282
R3029 a_2201_1050.n8 a_2201_1050.n3 10.615
R3030 SN.n14 SN.t2 479.223
R3031 SN.n11 SN.t6 479.223
R3032 SN.n8 SN.t7 479.223
R3033 SN.n5 SN.t14 479.223
R3034 SN.n2 SN.t8 479.223
R3035 SN.n0 SN.t13 479.223
R3036 SN.n14 SN.t11 375.52
R3037 SN.n11 SN.t15 375.52
R3038 SN.n8 SN.t16 375.52
R3039 SN.n5 SN.t0 375.52
R3040 SN.n2 SN.t4 375.52
R3041 SN.n0 SN.t5 375.52
R3042 SN.n12 SN.n11 280.047
R3043 SN.n6 SN.n5 280.047
R3044 SN.n1 SN.n0 280.047
R3045 SN.n3 SN.n2 276.525
R3046 SN.n9 SN.n8 276.525
R3047 SN.n15 SN.n14 276.525
R3048 SN.n12 SN.t1 136.76
R3049 SN.n6 SN.t9 136.76
R3050 SN.n1 SN.t10 136.76
R3051 SN.n15 SN.t17 135.513
R3052 SN.n9 SN.t3 135.513
R3053 SN.n3 SN.t12 135.513
R3054 SN.n4 SN.n1 15.211
R3055 SN.n7 SN.n4 10.564
R3056 SN.n13 SN.n10 10.564
R3057 SN.n10 SN.n7 10.561
R3058 SN.n16 SN.n13 10.561
R3059 SN.n7 SN.n6 4.65
R3060 SN.n13 SN.n12 4.65
R3061 SN.n4 SN.n3 2.113
R3062 SN.n10 SN.n9 2.113
R3063 SN.n16 SN.n15 2.113
R3064 SN.n16 SN 0.046
R3065 a_10219_989.n1 a_10219_989.t15 475.572
R3066 a_10219_989.n3 a_10219_989.t11 469.145
R3067 a_10219_989.n6 a_10219_989.t9 454.685
R3068 a_10219_989.n6 a_10219_989.t14 428.979
R3069 a_10219_989.n3 a_10219_989.t7 384.527
R3070 a_10219_989.n1 a_10219_989.t10 384.527
R3071 a_10219_989.n4 a_10219_989.t12 370.613
R3072 a_10219_989.n2 a_10219_989.t8 370.613
R3073 a_10219_989.n7 a_10219_989.t13 255.965
R3074 a_10219_989.n12 a_10219_989.n11 252.498
R3075 a_10219_989.n7 a_10219_989.n6 227.006
R3076 a_10219_989.n16 a_10219_989.n15 161.352
R3077 a_10219_989.n14 a_10219_989.n13 151.34
R3078 a_10219_989.n2 a_10219_989.n1 128.028
R3079 a_10219_989.n4 a_10219_989.n3 126.97
R3080 a_10219_989.n14 a_10219_989.n0 95.095
R3081 a_10219_989.n17 a_10219_989.n16 95.094
R3082 a_10219_989.n13 a_10219_989.n12 83.576
R3083 a_10219_989.n16 a_10219_989.n14 66.258
R3084 a_10219_989.n11 a_10219_989.n10 30
R3085 a_10219_989.n13 a_10219_989.n5 27.875
R3086 a_10219_989.n9 a_10219_989.n8 24.383
R3087 a_10219_989.n11 a_10219_989.n9 23.684
R3088 a_10219_989.n0 a_10219_989.t3 14.282
R3089 a_10219_989.n0 a_10219_989.t4 14.282
R3090 a_10219_989.n15 a_10219_989.t6 14.282
R3091 a_10219_989.n15 a_10219_989.t5 14.282
R3092 a_10219_989.n17 a_10219_989.t0 14.282
R3093 a_10219_989.t1 a_10219_989.n17 14.282
R3094 a_10219_989.n12 a_10219_989.n7 13.335
R3095 a_10219_989.n5 a_10219_989.n2 9.501
R3096 a_10219_989.n5 a_10219_989.n4 4.65
R3097 a_6371_989.n0 a_6371_989.t10 512.525
R3098 a_6371_989.n2 a_6371_989.t12 454.685
R3099 a_6371_989.n2 a_6371_989.t8 428.979
R3100 a_6371_989.n0 a_6371_989.t7 371.139
R3101 a_6371_989.n1 a_6371_989.t9 361.392
R3102 a_6371_989.n3 a_6371_989.t11 311.683
R3103 a_6371_989.n9 a_6371_989.n8 308.216
R3104 a_6371_989.n1 a_6371_989.n0 235.554
R3105 a_6371_989.n13 a_6371_989.n9 179.199
R3106 a_6371_989.n3 a_6371_989.n2 171.288
R3107 a_6371_989.n12 a_6371_989.n11 161.352
R3108 a_6371_989.n12 a_6371_989.n10 95.095
R3109 a_6371_989.n14 a_6371_989.n13 95.094
R3110 a_6371_989.n13 a_6371_989.n12 66.258
R3111 a_6371_989.n8 a_6371_989.n7 30
R3112 a_6371_989.n6 a_6371_989.n5 24.383
R3113 a_6371_989.n8 a_6371_989.n6 23.684
R3114 a_6371_989.n10 a_6371_989.t5 14.282
R3115 a_6371_989.n10 a_6371_989.t6 14.282
R3116 a_6371_989.n11 a_6371_989.t0 14.282
R3117 a_6371_989.n11 a_6371_989.t1 14.282
R3118 a_6371_989.t4 a_6371_989.n14 14.282
R3119 a_6371_989.n14 a_6371_989.t3 14.282
R3120 a_6371_989.n4 a_6371_989.n1 13.038
R3121 a_6371_989.n4 a_6371_989.n3 8.685
R3122 a_6371_989.n9 a_6371_989.n4 4.65
R3123 a_4901_103.n5 a_4901_103.n4 66.708
R3124 a_4901_103.n2 a_4901_103.n0 32.662
R3125 a_4901_103.n5 a_4901_103.n3 19.496
R3126 a_4901_103.t0 a_4901_103.n5 13.756
R3127 a_4901_103.t0 a_4901_103.n2 3.034
R3128 a_4901_103.n2 a_4901_103.n1 0.443
R3129 a_5182_210.n12 a_5182_210.n10 171.558
R3130 a_5182_210.n7 a_5182_210.n6 117.622
R3131 a_5182_210.n5 a_5182_210.n4 92.5
R3132 a_5182_210.n9 a_5182_210.n8 92.5
R3133 a_5182_210.n10 a_5182_210.t1 75.764
R3134 a_5182_210.n5 a_5182_210.n3 65.02
R3135 a_5182_210.n13 a_5182_210.n0 49.6
R3136 a_5182_210.n7 a_5182_210.n5 36.517
R3137 a_5182_210.n3 a_5182_210.n2 35.865
R3138 a_5182_210.n12 a_5182_210.n11 27.2
R3139 a_5182_210.n13 a_5182_210.n12 22.4
R3140 a_5182_210.n9 a_5182_210.n7 19.952
R3141 a_5182_210.t1 a_5182_210.n1 7.04
R3142 a_5182_210.n10 a_5182_210.n9 1.505
R3143 a_6825_103.n5 a_6825_103.n4 66.708
R3144 a_6825_103.n2 a_6825_103.n0 32.662
R3145 a_6825_103.n5 a_6825_103.n3 19.496
R3146 a_6825_103.t0 a_6825_103.n5 13.756
R3147 a_6825_103.t0 a_6825_103.n2 3.034
R3148 a_6825_103.n2 a_6825_103.n1 0.443
R3149 a_7106_210.n8 a_7106_210.n6 185.173
R3150 a_7106_210.t0 a_7106_210.n8 75.765
R3151 a_7106_210.n3 a_7106_210.n1 74.827
R3152 a_7106_210.n3 a_7106_210.n2 27.476
R3153 a_7106_210.n6 a_7106_210.n5 22.349
R3154 a_7106_210.t0 a_7106_210.n10 20.241
R3155 a_7106_210.t0 a_7106_210.n3 13.984
R3156 a_7106_210.n10 a_7106_210.n9 13.494
R3157 a_7106_210.n6 a_7106_210.n4 8.443
R3158 a_7106_210.t0 a_7106_210.n0 8.137
R3159 a_7106_210.n8 a_7106_210.n7 1.505
R3160 a_1053_103.n5 a_1053_103.n4 66.708
R3161 a_1053_103.n2 a_1053_103.n0 32.662
R3162 a_1053_103.n5 a_1053_103.n3 19.496
R3163 a_1053_103.t0 a_1053_103.n5 13.756
R3164 a_1053_103.t0 a_1053_103.n2 3.034
R3165 a_1053_103.n2 a_1053_103.n1 0.443
R3166 a_1334_210.n8 a_1334_210.n6 185.173
R3167 a_1334_210.t0 a_1334_210.n8 75.765
R3168 a_1334_210.n3 a_1334_210.n1 74.827
R3169 a_1334_210.n3 a_1334_210.n2 27.476
R3170 a_1334_210.n6 a_1334_210.n5 22.349
R3171 a_1334_210.t0 a_1334_210.n10 20.241
R3172 a_1334_210.t0 a_1334_210.n3 13.984
R3173 a_1334_210.n10 a_1334_210.n9 13.494
R3174 a_1334_210.n6 a_1334_210.n4 8.443
R3175 a_1334_210.t0 a_1334_210.n0 8.137
R3176 a_1334_210.n8 a_1334_210.n7 1.505
R3177 a_15991_989.n3 a_15991_989.t15 512.525
R3178 a_15991_989.n1 a_15991_989.t13 477.179
R3179 a_15991_989.n6 a_15991_989.t14 454.685
R3180 a_15991_989.n2 a_15991_989.t9 440.954
R3181 a_15991_989.n6 a_15991_989.t11 428.979
R3182 a_15991_989.n1 a_15991_989.t10 406.485
R3183 a_15991_989.n5 a_15991_989.t12 378.636
R3184 a_15991_989.n3 a_15991_989.t8 371.139
R3185 a_15991_989.n7 a_15991_989.t7 255.965
R3186 a_15991_989.n12 a_15991_989.n11 252.498
R3187 a_15991_989.n7 a_15991_989.n6 227.006
R3188 a_15991_989.n16 a_15991_989.n15 161.352
R3189 a_15991_989.n14 a_15991_989.n13 151.34
R3190 a_15991_989.n14 a_15991_989.n0 95.095
R3191 a_15991_989.n17 a_15991_989.n16 95.094
R3192 a_15991_989.n13 a_15991_989.n12 83.576
R3193 a_15991_989.n4 a_15991_989.n3 77.972
R3194 a_15991_989.n16 a_15991_989.n14 66.258
R3195 a_15991_989.n5 a_15991_989.n4 55.891
R3196 a_15991_989.n11 a_15991_989.n10 30
R3197 a_15991_989.n9 a_15991_989.n8 24.383
R3198 a_15991_989.n11 a_15991_989.n9 23.684
R3199 a_15991_989.n2 a_15991_989.n1 21.4
R3200 a_15991_989.n0 a_15991_989.t4 14.282
R3201 a_15991_989.n0 a_15991_989.t3 14.282
R3202 a_15991_989.n15 a_15991_989.t5 14.282
R3203 a_15991_989.n15 a_15991_989.t6 14.282
R3204 a_15991_989.n17 a_15991_989.t0 14.282
R3205 a_15991_989.t1 a_15991_989.n17 14.282
R3206 a_15991_989.n12 a_15991_989.n7 13.335
R3207 a_15991_989.n13 a_15991_989.n5 10.343
R3208 a_15991_989.n4 a_15991_989.n2 6.833
R3209 a_15764_210.n9 a_15764_210.n7 171.558
R3210 a_15764_210.t0 a_15764_210.n9 75.765
R3211 a_15764_210.n3 a_15764_210.n1 74.827
R3212 a_15764_210.n3 a_15764_210.n2 27.476
R3213 a_15764_210.n7 a_15764_210.n6 27.2
R3214 a_15764_210.n5 a_15764_210.n4 23.498
R3215 a_15764_210.n7 a_15764_210.n5 22.4
R3216 a_15764_210.t0 a_15764_210.n11 20.241
R3217 a_15764_210.t0 a_15764_210.n3 13.984
R3218 a_15764_210.n11 a_15764_210.n10 13.494
R3219 a_15764_210.t0 a_15764_210.n0 8.137
R3220 a_15764_210.n9 a_15764_210.n8 1.505
R3221 a_2977_103.n5 a_2977_103.n4 66.708
R3222 a_2977_103.n2 a_2977_103.n0 32.662
R3223 a_2977_103.n5 a_2977_103.n3 19.496
R3224 a_2977_103.t0 a_2977_103.n5 13.756
R3225 a_2977_103.t0 a_2977_103.n2 3.034
R3226 a_2977_103.n2 a_2977_103.n1 0.443
R3227 a_3258_210.n10 a_3258_210.n8 171.558
R3228 a_3258_210.n8 a_3258_210.t1 75.764
R3229 a_3258_210.n11 a_3258_210.n0 49.6
R3230 a_3258_210.n3 a_3258_210.n2 27.476
R3231 a_3258_210.n10 a_3258_210.n9 27.2
R3232 a_3258_210.n11 a_3258_210.n10 22.4
R3233 a_3258_210.t1 a_3258_210.n5 20.241
R3234 a_3258_210.n7 a_3258_210.n6 19.952
R3235 a_3258_210.t1 a_3258_210.n3 13.984
R3236 a_3258_210.n5 a_3258_210.n4 13.494
R3237 a_3258_210.t1 a_3258_210.n1 7.04
R3238 a_3258_210.n8 a_3258_210.n7 1.505
R3239 a_6049_1050.n2 a_6049_1050.t12 512.525
R3240 a_6049_1050.n0 a_6049_1050.t10 512.525
R3241 a_6049_1050.n2 a_6049_1050.t7 371.139
R3242 a_6049_1050.n0 a_6049_1050.t11 371.139
R3243 a_6049_1050.n3 a_6049_1050.t8 306.051
R3244 a_6049_1050.n1 a_6049_1050.t9 306.051
R3245 a_6049_1050.n3 a_6049_1050.n2 290.895
R3246 a_6049_1050.n1 a_6049_1050.n0 290.895
R3247 a_6049_1050.n9 a_6049_1050.n8 252.875
R3248 a_6049_1050.n13 a_6049_1050.n9 234.54
R3249 a_6049_1050.n12 a_6049_1050.n11 161.352
R3250 a_6049_1050.n12 a_6049_1050.n10 95.095
R3251 a_6049_1050.n14 a_6049_1050.n13 95.094
R3252 a_6049_1050.n13 a_6049_1050.n12 66.258
R3253 a_6049_1050.n8 a_6049_1050.n7 30
R3254 a_6049_1050.n6 a_6049_1050.n5 24.383
R3255 a_6049_1050.n8 a_6049_1050.n6 23.684
R3256 a_6049_1050.n10 a_6049_1050.t6 14.282
R3257 a_6049_1050.n10 a_6049_1050.t5 14.282
R3258 a_6049_1050.n11 a_6049_1050.t1 14.282
R3259 a_6049_1050.n11 a_6049_1050.t0 14.282
R3260 a_6049_1050.t4 a_6049_1050.n14 14.282
R3261 a_6049_1050.n14 a_6049_1050.t3 14.282
R3262 a_6049_1050.n4 a_6049_1050.n1 8.141
R3263 a_6049_1050.n9 a_6049_1050.n4 5.965
R3264 a_6049_1050.n4 a_6049_1050.n3 4.65
R3265 a_13840_210.n10 a_13840_210.n8 171.558
R3266 a_13840_210.n8 a_13840_210.t1 75.764
R3267 a_13840_210.n3 a_13840_210.n2 27.476
R3268 a_13840_210.n10 a_13840_210.n9 27.2
R3269 a_13840_210.n11 a_13840_210.n0 23.498
R3270 a_13840_210.n11 a_13840_210.n10 22.4
R3271 a_13840_210.t1 a_13840_210.n5 20.241
R3272 a_13840_210.n7 a_13840_210.n6 19.952
R3273 a_13840_210.t1 a_13840_210.n3 13.984
R3274 a_13840_210.n5 a_13840_210.n4 13.494
R3275 a_13840_210.t1 a_13840_210.n1 7.04
R3276 a_13840_210.n8 a_13840_210.n7 1.505
R3277 a_7973_1050.n2 a_7973_1050.t7 512.525
R3278 a_7973_1050.n2 a_7973_1050.t8 371.139
R3279 a_7973_1050.n3 a_7973_1050.t9 305.674
R3280 a_7973_1050.n3 a_7973_1050.n2 291.272
R3281 a_7973_1050.n8 a_7973_1050.n7 252.498
R3282 a_7973_1050.n9 a_7973_1050.n8 234.917
R3283 a_7973_1050.n11 a_7973_1050.n10 161.352
R3284 a_7973_1050.n9 a_7973_1050.n1 95.095
R3285 a_7973_1050.n10 a_7973_1050.n0 95.095
R3286 a_7973_1050.n10 a_7973_1050.n9 66.258
R3287 a_7973_1050.n7 a_7973_1050.n6 30
R3288 a_7973_1050.n5 a_7973_1050.n4 24.383
R3289 a_7973_1050.n7 a_7973_1050.n5 23.684
R3290 a_7973_1050.n1 a_7973_1050.t5 14.282
R3291 a_7973_1050.n1 a_7973_1050.t6 14.282
R3292 a_7973_1050.n0 a_7973_1050.t3 14.282
R3293 a_7973_1050.n0 a_7973_1050.t2 14.282
R3294 a_7973_1050.t1 a_7973_1050.n11 14.282
R3295 a_7973_1050.n11 a_7973_1050.t0 14.282
R3296 a_7973_1050.n8 a_7973_1050.n3 10.615
R3297 a_17533_1051.n2 a_17533_1051.t0 179.895
R3298 a_17533_1051.n5 a_17533_1051.n4 157.021
R3299 a_17533_1051.n4 a_17533_1051.n0 124.955
R3300 a_17533_1051.n3 a_17533_1051.n2 106.183
R3301 a_17533_1051.n2 a_17533_1051.n1 99.355
R3302 a_17533_1051.n4 a_17533_1051.n3 82.65
R3303 a_17533_1051.n3 a_17533_1051.t2 73.712
R3304 a_17533_1051.n0 a_17533_1051.t5 14.282
R3305 a_17533_1051.n0 a_17533_1051.t6 14.282
R3306 a_17533_1051.n1 a_17533_1051.t7 14.282
R3307 a_17533_1051.n1 a_17533_1051.t1 14.282
R3308 a_17533_1051.n5 a_17533_1051.t3 14.282
R3309 a_17533_1051.t4 a_17533_1051.n5 14.282
R3310 a_4125_1050.n2 a_4125_1050.t8 512.525
R3311 a_4125_1050.n2 a_4125_1050.t9 371.139
R3312 a_4125_1050.n3 a_4125_1050.t7 361.392
R3313 a_4125_1050.n5 a_4125_1050.n4 329.955
R3314 a_4125_1050.n3 a_4125_1050.n2 235.554
R3315 a_4125_1050.n6 a_4125_1050.n5 179.199
R3316 a_4125_1050.n8 a_4125_1050.n7 161.352
R3317 a_4125_1050.n6 a_4125_1050.n1 95.095
R3318 a_4125_1050.n7 a_4125_1050.n0 95.095
R3319 a_4125_1050.n7 a_4125_1050.n6 66.258
R3320 a_4125_1050.n1 a_4125_1050.t2 14.282
R3321 a_4125_1050.n1 a_4125_1050.t0 14.282
R3322 a_4125_1050.n0 a_4125_1050.t5 14.282
R3323 a_4125_1050.n0 a_4125_1050.t6 14.282
R3324 a_4125_1050.n8 a_4125_1050.t3 14.282
R3325 a_4125_1050.t4 a_4125_1050.n8 14.282
R3326 a_4125_1050.n5 a_4125_1050.n3 10.615
R3327 a_4447_989.n3 a_4447_989.t10 512.525
R3328 a_4447_989.n2 a_4447_989.t9 512.525
R3329 a_4447_989.n7 a_4447_989.t7 454.685
R3330 a_4447_989.n7 a_4447_989.t13 428.979
R3331 a_4447_989.n3 a_4447_989.t14 371.139
R3332 a_4447_989.n2 a_4447_989.t15 371.139
R3333 a_4447_989.n4 a_4447_989.n3 343.521
R3334 a_4447_989.n13 a_4447_989.n12 295.88
R3335 a_4447_989.n8 a_4447_989.t12 272.577
R3336 a_4447_989.n6 a_4447_989.n2 259.945
R3337 a_4447_989.n14 a_4447_989.n13 207.058
R3338 a_4447_989.n8 a_4447_989.n7 199.147
R3339 a_4447_989.n4 a_4447_989.t8 172.106
R3340 a_4447_989.n5 a_4447_989.t11 165.68
R3341 a_4447_989.n16 a_4447_989.n15 161.352
R3342 a_4447_989.n14 a_4447_989.n1 95.095
R3343 a_4447_989.n15 a_4447_989.n0 95.095
R3344 a_4447_989.n6 a_4447_989.n5 83.576
R3345 a_4447_989.n15 a_4447_989.n14 66.258
R3346 a_4447_989.n9 a_4447_989.n6 51.943
R3347 a_4447_989.n12 a_4447_989.n11 22.578
R3348 a_4447_989.n1 a_4447_989.t6 14.282
R3349 a_4447_989.n1 a_4447_989.t5 14.282
R3350 a_4447_989.n0 a_4447_989.t3 14.282
R3351 a_4447_989.n0 a_4447_989.t2 14.282
R3352 a_4447_989.t1 a_4447_989.n16 14.282
R3353 a_4447_989.n16 a_4447_989.t0 14.282
R3354 a_4447_989.n5 a_4447_989.n4 10.343
R3355 a_4447_989.n9 a_4447_989.n8 8.685
R3356 a_4447_989.n12 a_4447_989.n10 8.58
R3357 a_4447_989.n13 a_4447_989.n9 4.65
R3358 a_18760_101.n3 a_18760_101.n1 42.788
R3359 a_18760_101.t0 a_18760_101.n0 8.137
R3360 a_18760_101.n3 a_18760_101.n2 4.665
R3361 a_18760_101.t0 a_18760_101.n3 0.06
R3362 a_18094_101.n2 a_18094_101.n0 42.761
R3363 a_18094_101.n2 a_18094_101.n1 2.167
R3364 a_18094_101.t0 a_18094_101.n2 0.099
R3365 a_18197_1051.n2 a_18197_1051.t6 179.895
R3366 a_18197_1051.n5 a_18197_1051.n4 165.613
R3367 a_18197_1051.n4 a_18197_1051.n0 142.653
R3368 a_18197_1051.n3 a_18197_1051.n2 106.183
R3369 a_18197_1051.n2 a_18197_1051.n1 99.355
R3370 a_18197_1051.n4 a_18197_1051.n3 82.665
R3371 a_18197_1051.n3 a_18197_1051.t3 73.712
R3372 a_18197_1051.n0 a_18197_1051.t4 14.282
R3373 a_18197_1051.n0 a_18197_1051.t5 14.282
R3374 a_18197_1051.n1 a_18197_1051.t7 14.282
R3375 a_18197_1051.n1 a_18197_1051.t2 14.282
R3376 a_18197_1051.n5 a_18197_1051.t0 14.282
R3377 a_18197_1051.t1 a_18197_1051.n5 14.282
R3378 a_5863_103.n5 a_5863_103.n4 66.708
R3379 a_5863_103.n2 a_5863_103.n0 32.662
R3380 a_5863_103.n5 a_5863_103.n3 19.496
R3381 a_5863_103.t0 a_5863_103.n5 13.756
R3382 a_5863_103.t0 a_5863_103.n2 3.034
R3383 a_5863_103.n2 a_5863_103.n1 0.443
R3384 a_6144_210.n8 a_6144_210.n6 185.173
R3385 a_6144_210.t0 a_6144_210.n8 75.765
R3386 a_6144_210.n3 a_6144_210.n1 74.827
R3387 a_6144_210.n3 a_6144_210.n2 27.476
R3388 a_6144_210.n6 a_6144_210.n5 22.349
R3389 a_6144_210.t0 a_6144_210.n10 20.241
R3390 a_6144_210.t0 a_6144_210.n3 13.984
R3391 a_6144_210.n10 a_6144_210.n9 13.494
R3392 a_6144_210.n6 a_6144_210.n4 8.443
R3393 a_6144_210.t0 a_6144_210.n0 8.137
R3394 a_6144_210.n8 a_6144_210.n7 1.505
R3395 D.n5 D.t7 512.525
R3396 D.n2 D.t6 512.525
R3397 D.n0 D.t8 512.525
R3398 D.n6 D.t4 417.109
R3399 D.n3 D.t1 417.109
R3400 D.n1 D.t0 417.109
R3401 D.n5 D.t3 371.139
R3402 D.n2 D.t2 371.139
R3403 D.n0 D.t5 371.139
R3404 D.n6 D.n5 179.837
R3405 D.n3 D.n2 179.837
R3406 D.n1 D.n0 179.837
R3407 D.n4 D.n1 25.825
R3408 D.n7 D.n4 21.175
R3409 D.n4 D.n3 4.65
R3410 D.n7 D.n6 4.65
R3411 D.n7 D 0.046
R3412 a_11635_103.n5 a_11635_103.n4 66.708
R3413 a_11635_103.n2 a_11635_103.n0 32.662
R3414 a_11635_103.n5 a_11635_103.n3 19.496
R3415 a_11635_103.t0 a_11635_103.n5 13.756
R3416 a_11635_103.t0 a_11635_103.n2 3.034
R3417 a_11635_103.n2 a_11635_103.n1 0.443
R3418 a_16726_210.n10 a_16726_210.n8 171.558
R3419 a_16726_210.n8 a_16726_210.t1 75.764
R3420 a_16726_210.n3 a_16726_210.n2 27.476
R3421 a_16726_210.n10 a_16726_210.n9 27.2
R3422 a_16726_210.n11 a_16726_210.n0 23.498
R3423 a_16726_210.n11 a_16726_210.n10 22.4
R3424 a_16726_210.t1 a_16726_210.n5 20.241
R3425 a_16726_210.n7 a_16726_210.n6 19.952
R3426 a_16726_210.t1 a_16726_210.n3 13.984
R3427 a_16726_210.n5 a_16726_210.n4 13.494
R3428 a_16726_210.t1 a_16726_210.n1 7.04
R3429 a_16726_210.n8 a_16726_210.n7 1.505
R3430 a_7787_103.n5 a_7787_103.n4 66.708
R3431 a_7787_103.n2 a_7787_103.n0 32.662
R3432 a_7787_103.n5 a_7787_103.n3 19.496
R3433 a_7787_103.t0 a_7787_103.n5 13.756
R3434 a_7787_103.t0 a_7787_103.n2 3.034
R3435 a_7787_103.n2 a_7787_103.n1 0.443
R3436 a_8068_210.n10 a_8068_210.n8 171.558
R3437 a_8068_210.n8 a_8068_210.t1 75.764
R3438 a_8068_210.n11 a_8068_210.n0 49.6
R3439 a_8068_210.n3 a_8068_210.n2 27.476
R3440 a_8068_210.n10 a_8068_210.n9 27.2
R3441 a_8068_210.n11 a_8068_210.n10 22.4
R3442 a_8068_210.t1 a_8068_210.n5 20.241
R3443 a_8068_210.n7 a_8068_210.n6 19.952
R3444 a_8068_210.t1 a_8068_210.n3 13.984
R3445 a_8068_210.n5 a_8068_210.n4 13.494
R3446 a_8068_210.t1 a_8068_210.n1 7.04
R3447 a_8068_210.n8 a_8068_210.n7 1.505
R3448 a_9711_103.n5 a_9711_103.n4 66.708
R3449 a_9711_103.n2 a_9711_103.n0 32.662
R3450 a_9711_103.n5 a_9711_103.n3 19.496
R3451 a_9711_103.t0 a_9711_103.n5 13.756
R3452 a_9711_103.t0 a_9711_103.n2 3.034
R3453 a_9711_103.n2 a_9711_103.n1 0.443
R3454 QN.n13 QN.n12 227.387
R3455 QN.n2 QN.n1 165.613
R3456 QN.n13 QN.n2 132.893
R3457 QN.n12 QN.n11 127.909
R3458 QN.n10 QN.n5 126.225
R3459 QN.n10 QN.n9 112.771
R3460 QN.n2 QN.n0 99.355
R3461 QN.n9 QN.n8 30
R3462 QN.n7 QN.n6 24.383
R3463 QN.n9 QN.n7 23.684
R3464 QN.n5 QN.n4 22.578
R3465 QN.n0 QN.t3 14.282
R3466 QN.n0 QN.t4 14.282
R3467 QN.n1 QN.t1 14.282
R3468 QN.n1 QN.t0 14.282
R3469 QN.n5 QN.n3 8.58
R3470 QN.n12 QN.n10 7.053
R3471 QN.n14 QN.n13 4.65
R3472 QN.n14 QN 0.046
R3473 a_372_210.n9 a_372_210.n7 171.558
R3474 a_372_210.t0 a_372_210.n9 75.765
R3475 a_372_210.n3 a_372_210.n1 74.827
R3476 a_372_210.n3 a_372_210.n2 27.476
R3477 a_372_210.n7 a_372_210.n6 27.2
R3478 a_372_210.n5 a_372_210.n4 23.498
R3479 a_372_210.n7 a_372_210.n5 22.4
R3480 a_372_210.t0 a_372_210.n11 20.241
R3481 a_372_210.t0 a_372_210.n3 13.984
R3482 a_372_210.n11 a_372_210.n10 13.494
R3483 a_372_210.t0 a_372_210.n0 8.137
R3484 a_372_210.n9 a_372_210.n8 1.505
R3485 a_8749_103.n5 a_8749_103.n4 66.708
R3486 a_8749_103.n2 a_8749_103.n0 25.439
R3487 a_8749_103.n5 a_8749_103.n3 19.496
R3488 a_8749_103.t0 a_8749_103.n5 13.756
R3489 a_8749_103.n2 a_8749_103.n1 2.455
R3490 a_8749_103.t0 a_8749_103.n2 0.246
R3491 a_12597_103.n5 a_12597_103.n4 66.708
R3492 a_12597_103.n2 a_12597_103.n0 32.662
R3493 a_12597_103.n5 a_12597_103.n3 19.496
R3494 a_12597_103.t0 a_12597_103.n5 13.756
R3495 a_12597_103.t0 a_12597_103.n2 3.034
R3496 a_12597_103.n2 a_12597_103.n1 0.443
R3497 a_14521_103.n5 a_14521_103.n4 66.708
R3498 a_14521_103.n2 a_14521_103.n0 25.439
R3499 a_14521_103.n5 a_14521_103.n3 19.496
R3500 a_14521_103.t0 a_14521_103.n5 13.756
R3501 a_14521_103.n2 a_14521_103.n1 2.455
R3502 a_14521_103.t0 a_14521_103.n2 0.246
R3503 a_10673_103.t0 a_10673_103.n7 59.616
R3504 a_10673_103.n4 a_10673_103.n2 54.496
R3505 a_10673_103.n4 a_10673_103.n3 54.496
R3506 a_10673_103.n1 a_10673_103.n0 24.679
R3507 a_10673_103.n6 a_10673_103.n4 7.859
R3508 a_10673_103.t0 a_10673_103.n1 7.505
R3509 a_10673_103.t0 a_10673_103.n6 3.034
R3510 a_10673_103.n6 a_10673_103.n5 0.443
R3511 a_91_103.n5 a_91_103.n4 66.708
R3512 a_91_103.n2 a_91_103.n0 25.439
R3513 a_91_103.n5 a_91_103.n3 19.496
R3514 a_91_103.t0 a_91_103.n5 13.756
R3515 a_91_103.n2 a_91_103.n1 2.455
R3516 a_91_103.t0 a_91_103.n2 0.246
R3517 a_11916_210.n8 a_11916_210.n6 185.173
R3518 a_11916_210.t0 a_11916_210.n8 75.765
R3519 a_11916_210.n3 a_11916_210.n1 74.827
R3520 a_11916_210.n3 a_11916_210.n2 27.476
R3521 a_11916_210.n6 a_11916_210.n5 22.349
R3522 a_11916_210.t0 a_11916_210.n10 20.241
R3523 a_11916_210.t0 a_11916_210.n3 13.984
R3524 a_11916_210.n10 a_11916_210.n9 13.494
R3525 a_11916_210.n6 a_11916_210.n4 8.443
R3526 a_11916_210.t0 a_11916_210.n0 8.137
R3527 a_11916_210.n8 a_11916_210.n7 1.505
R3528 a_9992_210.n8 a_9992_210.n6 185.173
R3529 a_9992_210.t0 a_9992_210.n8 75.765
R3530 a_9992_210.n3 a_9992_210.n1 74.827
R3531 a_9992_210.n3 a_9992_210.n2 27.476
R3532 a_9992_210.n6 a_9992_210.n5 22.349
R3533 a_9992_210.t0 a_9992_210.n10 20.241
R3534 a_9992_210.t0 a_9992_210.n3 13.984
R3535 a_9992_210.n10 a_9992_210.n9 13.494
R3536 a_9992_210.n6 a_9992_210.n4 8.443
R3537 a_9992_210.t0 a_9992_210.n0 8.137
R3538 a_9992_210.n8 a_9992_210.n7 1.505
R3539 a_17428_101.n3 a_17428_101.n2 62.817
R3540 a_17428_101.n11 a_17428_101.n10 46.054
R3541 a_17428_101.n7 a_17428_101.n6 38.626
R3542 a_17428_101.n6 a_17428_101.n5 35.955
R3543 a_17428_101.n12 a_17428_101.n11 27.923
R3544 a_17428_101.n3 a_17428_101.n1 26.202
R3545 a_17428_101.t0 a_17428_101.n3 19.737
R3546 a_17428_101.t0 a_17428_101.n4 7.273
R3547 a_17428_101.n9 a_17428_101.n8 6.883
R3548 a_17428_101.t0 a_17428_101.n0 6.109
R3549 a_17428_101.t1 a_17428_101.n7 4.864
R3550 a_17428_101.t0 a_17428_101.n13 2.074
R3551 a_17428_101.t1 a_17428_101.n9 1.179
R3552 a_17428_101.t1 a_17428_101.n12 0.958
R3553 a_17428_101.n13 a_17428_101.t1 0.937
R3554 a_13559_103.t0 a_13559_103.n7 59.616
R3555 a_13559_103.n4 a_13559_103.n2 54.496
R3556 a_13559_103.n4 a_13559_103.n3 54.496
R3557 a_13559_103.n1 a_13559_103.n0 24.679
R3558 a_13559_103.t0 a_13559_103.n1 7.505
R3559 a_13559_103.n6 a_13559_103.n5 2.455
R3560 a_13559_103.n6 a_13559_103.n4 0.636
R3561 a_13559_103.t0 a_13559_103.n6 0.246
R3562 a_15483_103.n5 a_15483_103.n4 66.708
R3563 a_15483_103.n2 a_15483_103.n0 25.439
R3564 a_15483_103.n5 a_15483_103.n3 19.496
R3565 a_15483_103.t0 a_15483_103.n5 13.756
R3566 a_15483_103.n2 a_15483_103.n1 2.455
R3567 a_15483_103.t0 a_15483_103.n2 0.246
R3568 a_10954_210.n10 a_10954_210.n8 171.558
R3569 a_10954_210.n8 a_10954_210.t1 75.764
R3570 a_10954_210.n11 a_10954_210.n0 49.6
R3571 a_10954_210.n3 a_10954_210.n2 27.476
R3572 a_10954_210.n10 a_10954_210.n9 27.2
R3573 a_10954_210.n11 a_10954_210.n10 22.4
R3574 a_10954_210.t1 a_10954_210.n5 20.241
R3575 a_10954_210.n7 a_10954_210.n6 19.952
R3576 a_10954_210.t1 a_10954_210.n3 13.984
R3577 a_10954_210.n5 a_10954_210.n4 13.494
R3578 a_10954_210.t1 a_10954_210.n1 7.04
R3579 a_10954_210.n8 a_10954_210.n7 1.505
R3580 a_16445_103.t0 a_16445_103.n7 59.616
R3581 a_16445_103.n4 a_16445_103.n2 54.496
R3582 a_16445_103.n4 a_16445_103.n3 54.496
R3583 a_16445_103.n1 a_16445_103.n0 24.679
R3584 a_16445_103.t0 a_16445_103.n1 7.505
R3585 a_16445_103.n6 a_16445_103.n5 2.455
R3586 a_16445_103.n6 a_16445_103.n4 0.636
R3587 a_16445_103.t0 a_16445_103.n6 0.246
R3588 a_12878_210.n10 a_12878_210.n8 171.558
R3589 a_12878_210.n8 a_12878_210.t1 75.764
R3590 a_12878_210.n11 a_12878_210.n0 49.6
R3591 a_12878_210.n3 a_12878_210.n2 27.476
R3592 a_12878_210.n10 a_12878_210.n9 27.2
R3593 a_12878_210.n11 a_12878_210.n10 22.4
R3594 a_12878_210.t1 a_12878_210.n5 20.241
R3595 a_12878_210.n7 a_12878_210.n6 19.952
R3596 a_12878_210.t1 a_12878_210.n3 13.984
R3597 a_12878_210.n5 a_12878_210.n4 13.494
R3598 a_12878_210.t1 a_12878_210.n1 7.04
R3599 a_12878_210.n8 a_12878_210.n7 1.505
R3600 a_2296_210.n10 a_2296_210.n8 171.558
R3601 a_2296_210.n8 a_2296_210.t1 75.764
R3602 a_2296_210.n3 a_2296_210.n2 27.476
R3603 a_2296_210.n10 a_2296_210.n9 27.2
R3604 a_2296_210.n11 a_2296_210.n0 23.498
R3605 a_2296_210.n11 a_2296_210.n10 22.4
R3606 a_2296_210.t1 a_2296_210.n5 20.241
R3607 a_2296_210.n7 a_2296_210.n6 19.952
R3608 a_2296_210.t1 a_2296_210.n3 13.984
R3609 a_2296_210.n5 a_2296_210.n4 13.494
R3610 a_2296_210.t1 a_2296_210.n1 7.04
R3611 a_2296_210.n8 a_2296_210.n7 1.505
R3612 a_4220_210.n8 a_4220_210.n6 185.173
R3613 a_4220_210.t0 a_4220_210.n8 75.765
R3614 a_4220_210.n3 a_4220_210.n1 74.827
R3615 a_4220_210.n3 a_4220_210.n2 27.476
R3616 a_4220_210.n6 a_4220_210.n5 22.349
R3617 a_4220_210.t0 a_4220_210.n10 20.241
R3618 a_4220_210.t0 a_4220_210.n3 13.984
R3619 a_4220_210.n10 a_4220_210.n9 13.494
R3620 a_4220_210.n6 a_4220_210.n4 8.443
R3621 a_4220_210.t0 a_4220_210.n0 8.137
R3622 a_4220_210.n8 a_4220_210.n7 1.505
R3623 a_2015_103.t0 a_2015_103.n7 59.616
R3624 a_2015_103.n4 a_2015_103.n2 54.496
R3625 a_2015_103.n4 a_2015_103.n3 54.496
R3626 a_2015_103.n1 a_2015_103.n0 24.679
R3627 a_2015_103.t0 a_2015_103.n1 7.505
R3628 a_2015_103.n6 a_2015_103.n5 2.455
R3629 a_2015_103.n6 a_2015_103.n4 0.636
R3630 a_2015_103.t0 a_2015_103.n6 0.246
C11 SN GND 7.80fF
C12 RN GND 8.38fF
C13 VDD GND 31.90fF
C14 a_2015_103.n0 GND 0.08fF
C15 a_2015_103.n1 GND 0.07fF
C16 a_2015_103.n2 GND 0.04fF
C17 a_2015_103.n3 GND 0.06fF
C18 a_2015_103.n4 GND 0.03fF
C19 a_2015_103.n5 GND 0.04fF
C20 a_2015_103.n7 GND 0.08fF
C21 a_4220_210.n0 GND 0.07fF
C22 a_4220_210.n1 GND 0.09fF
C23 a_4220_210.n2 GND 0.12fF
C24 a_4220_210.n3 GND 0.08fF
C25 a_4220_210.n4 GND 0.02fF
C26 a_4220_210.n5 GND 0.03fF
C27 a_4220_210.n6 GND 0.05fF
C28 a_4220_210.n7 GND 0.02fF
C29 a_4220_210.n8 GND 0.14fF
C30 a_4220_210.n9 GND 0.08fF
C31 a_4220_210.n10 GND 0.02fF
C32 a_4220_210.t0 GND 0.31fF
C33 a_2296_210.n0 GND 0.02fF
C34 a_2296_210.n1 GND 0.09fF
C35 a_2296_210.n2 GND 0.12fF
C36 a_2296_210.n3 GND 0.08fF
C37 a_2296_210.n4 GND 0.08fF
C38 a_2296_210.n5 GND 0.02fF
C39 a_2296_210.t1 GND 0.29fF
C40 a_2296_210.n6 GND 0.09fF
C41 a_2296_210.n7 GND 0.02fF
C42 a_2296_210.n8 GND 0.13fF
C43 a_2296_210.n9 GND 0.02fF
C44 a_2296_210.n10 GND 0.03fF
C45 a_2296_210.n11 GND 0.03fF
C46 a_12878_210.n0 GND 0.02fF
C47 a_12878_210.n1 GND 0.09fF
C48 a_12878_210.n2 GND 0.12fF
C49 a_12878_210.n3 GND 0.08fF
C50 a_12878_210.n4 GND 0.08fF
C51 a_12878_210.n5 GND 0.02fF
C52 a_12878_210.t1 GND 0.29fF
C53 a_12878_210.n6 GND 0.09fF
C54 a_12878_210.n7 GND 0.02fF
C55 a_12878_210.n8 GND 0.13fF
C56 a_12878_210.n9 GND 0.02fF
C57 a_12878_210.n10 GND 0.03fF
C58 a_12878_210.n11 GND 0.02fF
C59 a_16445_103.n0 GND 0.08fF
C60 a_16445_103.n1 GND 0.07fF
C61 a_16445_103.n2 GND 0.04fF
C62 a_16445_103.n3 GND 0.06fF
C63 a_16445_103.n4 GND 0.03fF
C64 a_16445_103.n5 GND 0.04fF
C65 a_16445_103.n7 GND 0.08fF
C66 a_10954_210.n0 GND 0.02fF
C67 a_10954_210.n1 GND 0.09fF
C68 a_10954_210.n2 GND 0.12fF
C69 a_10954_210.n3 GND 0.08fF
C70 a_10954_210.n4 GND 0.08fF
C71 a_10954_210.n5 GND 0.02fF
C72 a_10954_210.t1 GND 0.29fF
C73 a_10954_210.n6 GND 0.09fF
C74 a_10954_210.n7 GND 0.02fF
C75 a_10954_210.n8 GND 0.13fF
C76 a_10954_210.n9 GND 0.02fF
C77 a_10954_210.n10 GND 0.03fF
C78 a_10954_210.n11 GND 0.02fF
C79 a_15483_103.n0 GND 0.11fF
C80 a_15483_103.n1 GND 0.04fF
C81 a_15483_103.n2 GND 0.03fF
C82 a_15483_103.n3 GND 0.07fF
C83 a_15483_103.n4 GND 0.08fF
C84 a_15483_103.n5 GND 0.03fF
C85 a_13559_103.n0 GND 0.08fF
C86 a_13559_103.n1 GND 0.07fF
C87 a_13559_103.n2 GND 0.04fF
C88 a_13559_103.n3 GND 0.06fF
C89 a_13559_103.n4 GND 0.03fF
C90 a_13559_103.n5 GND 0.04fF
C91 a_13559_103.n7 GND 0.08fF
C92 a_17428_101.n0 GND 0.02fF
C93 a_17428_101.n1 GND 0.09fF
C94 a_17428_101.n2 GND 0.07fF
C95 a_17428_101.n3 GND 0.03fF
C96 a_17428_101.n4 GND 0.01fF
C97 a_17428_101.n5 GND 0.03fF
C98 a_17428_101.n6 GND 0.04fF
C99 a_17428_101.n7 GND 0.02fF
C100 a_17428_101.n8 GND 0.04fF
C101 a_17428_101.n9 GND 0.08fF
C102 a_17428_101.n10 GND 0.04fF
C103 a_17428_101.n11 GND 0.12fF
C104 a_17428_101.n12 GND 0.14fF
C105 a_17428_101.n13 GND 0.01fF
C106 a_9992_210.n0 GND 0.07fF
C107 a_9992_210.n1 GND 0.09fF
C108 a_9992_210.n2 GND 0.12fF
C109 a_9992_210.n3 GND 0.08fF
C110 a_9992_210.n4 GND 0.02fF
C111 a_9992_210.n5 GND 0.03fF
C112 a_9992_210.n6 GND 0.05fF
C113 a_9992_210.n7 GND 0.02fF
C114 a_9992_210.n8 GND 0.14fF
C115 a_9992_210.n9 GND 0.08fF
C116 a_9992_210.n10 GND 0.02fF
C117 a_9992_210.t0 GND 0.31fF
C118 a_11916_210.n0 GND 0.07fF
C119 a_11916_210.n1 GND 0.09fF
C120 a_11916_210.n2 GND 0.12fF
C121 a_11916_210.n3 GND 0.08fF
C122 a_11916_210.n4 GND 0.02fF
C123 a_11916_210.n5 GND 0.03fF
C124 a_11916_210.n6 GND 0.05fF
C125 a_11916_210.n7 GND 0.02fF
C126 a_11916_210.n8 GND 0.14fF
C127 a_11916_210.n9 GND 0.08fF
C128 a_11916_210.n10 GND 0.02fF
C129 a_11916_210.t0 GND 0.31fF
C130 a_91_103.n0 GND 0.10fF
C131 a_91_103.n1 GND 0.03fF
C132 a_91_103.n2 GND 0.03fF
C133 a_91_103.n3 GND 0.07fF
C134 a_91_103.n4 GND 0.08fF
C135 a_91_103.n5 GND 0.03fF
C136 a_10673_103.n0 GND 0.08fF
C137 a_10673_103.n1 GND 0.07fF
C138 a_10673_103.n2 GND 0.04fF
C139 a_10673_103.n3 GND 0.06fF
C140 a_10673_103.n4 GND 0.11fF
C141 a_10673_103.n5 GND 0.04fF
C142 a_10673_103.n7 GND 0.08fF
C143 a_14521_103.n0 GND 0.11fF
C144 a_14521_103.n1 GND 0.04fF
C145 a_14521_103.n2 GND 0.03fF
C146 a_14521_103.n3 GND 0.07fF
C147 a_14521_103.n4 GND 0.08fF
C148 a_14521_103.n5 GND 0.03fF
C149 a_12597_103.n0 GND 0.13fF
C150 a_12597_103.n1 GND 0.04fF
C151 a_12597_103.n2 GND 0.09fF
C152 a_12597_103.n3 GND 0.07fF
C153 a_12597_103.n4 GND 0.08fF
C154 a_12597_103.n5 GND 0.03fF
C155 a_8749_103.n0 GND 0.11fF
C156 a_8749_103.n1 GND 0.04fF
C157 a_8749_103.n2 GND 0.03fF
C158 a_8749_103.n3 GND 0.07fF
C159 a_8749_103.n4 GND 0.08fF
C160 a_8749_103.n5 GND 0.03fF
C161 a_372_210.n0 GND 0.07fF
C162 a_372_210.n1 GND 0.09fF
C163 a_372_210.n2 GND 0.12fF
C164 a_372_210.n3 GND 0.08fF
C165 a_372_210.n4 GND 0.02fF
C166 a_372_210.n5 GND 0.03fF
C167 a_372_210.n6 GND 0.02fF
C168 a_372_210.n7 GND 0.03fF
C169 a_372_210.n8 GND 0.02fF
C170 a_372_210.n9 GND 0.13fF
C171 a_372_210.n10 GND 0.08fF
C172 a_372_210.n11 GND 0.02fF
C173 a_372_210.t0 GND 0.31fF
C174 QN.n0 GND 0.30fF
C175 QN.n1 GND 0.38fF
C176 QN.n2 GND 0.46fF
C177 QN.n3 GND 0.04fF
C178 QN.n4 GND 0.05fF
C179 QN.n5 GND 0.06fF
C180 QN.n6 GND 0.04fF
C181 QN.n7 GND 0.05fF
C182 QN.n8 GND 0.03fF
C183 QN.n9 GND 0.04fF
C184 QN.n10 GND 1.06fF
C185 QN.n11 GND 0.14fF
C186 QN.n12 GND 0.38fF
C187 QN.n13 GND 0.35fF
C188 QN.n14 GND 0.01fF
C189 a_9711_103.n0 GND 0.13fF
C190 a_9711_103.n1 GND 0.04fF
C191 a_9711_103.n2 GND 0.09fF
C192 a_9711_103.n3 GND 0.07fF
C193 a_9711_103.n4 GND 0.08fF
C194 a_9711_103.n5 GND 0.03fF
C195 a_8068_210.n0 GND 0.02fF
C196 a_8068_210.n1 GND 0.09fF
C197 a_8068_210.n2 GND 0.12fF
C198 a_8068_210.n3 GND 0.08fF
C199 a_8068_210.n4 GND 0.08fF
C200 a_8068_210.n5 GND 0.02fF
C201 a_8068_210.t1 GND 0.29fF
C202 a_8068_210.n6 GND 0.09fF
C203 a_8068_210.n7 GND 0.02fF
C204 a_8068_210.n8 GND 0.13fF
C205 a_8068_210.n9 GND 0.02fF
C206 a_8068_210.n10 GND 0.03fF
C207 a_8068_210.n11 GND 0.02fF
C208 a_7787_103.n0 GND 0.13fF
C209 a_7787_103.n1 GND 0.04fF
C210 a_7787_103.n2 GND 0.09fF
C211 a_7787_103.n3 GND 0.07fF
C212 a_7787_103.n4 GND 0.08fF
C213 a_7787_103.n5 GND 0.03fF
C214 a_16726_210.n0 GND 0.02fF
C215 a_16726_210.n1 GND 0.09fF
C216 a_16726_210.n2 GND 0.12fF
C217 a_16726_210.n3 GND 0.08fF
C218 a_16726_210.n4 GND 0.08fF
C219 a_16726_210.n5 GND 0.02fF
C220 a_16726_210.t1 GND 0.29fF
C221 a_16726_210.n6 GND 0.09fF
C222 a_16726_210.n7 GND 0.02fF
C223 a_16726_210.n8 GND 0.13fF
C224 a_16726_210.n9 GND 0.02fF
C225 a_16726_210.n10 GND 0.03fF
C226 a_16726_210.n11 GND 0.03fF
C227 a_11635_103.n0 GND 0.13fF
C228 a_11635_103.n1 GND 0.04fF
C229 a_11635_103.n2 GND 0.09fF
C230 a_11635_103.n3 GND 0.07fF
C231 a_11635_103.n4 GND 0.08fF
C232 a_11635_103.n5 GND 0.03fF
C233 a_6144_210.n0 GND 0.07fF
C234 a_6144_210.n1 GND 0.09fF
C235 a_6144_210.n2 GND 0.12fF
C236 a_6144_210.n3 GND 0.08fF
C237 a_6144_210.n4 GND 0.02fF
C238 a_6144_210.n5 GND 0.03fF
C239 a_6144_210.n6 GND 0.05fF
C240 a_6144_210.n7 GND 0.02fF
C241 a_6144_210.n8 GND 0.14fF
C242 a_6144_210.n9 GND 0.08fF
C243 a_6144_210.n10 GND 0.02fF
C244 a_6144_210.t0 GND 0.31fF
C245 a_5863_103.n0 GND 0.13fF
C246 a_5863_103.n1 GND 0.04fF
C247 a_5863_103.n2 GND 0.09fF
C248 a_5863_103.n3 GND 0.07fF
C249 a_5863_103.n4 GND 0.08fF
C250 a_5863_103.n5 GND 0.03fF
C251 a_18197_1051.n0 GND 0.28fF
C252 a_18197_1051.n1 GND 0.28fF
C253 a_18197_1051.n2 GND 0.45fF
C254 a_18197_1051.n3 GND 0.27fF
C255 a_18197_1051.n4 GND 0.70fF
C256 a_18197_1051.n5 GND 0.36fF
C257 a_18094_101.n0 GND 0.13fF
C258 a_18094_101.n1 GND 0.16fF
C259 a_18094_101.n2 GND 0.15fF
C260 a_18760_101.n0 GND 0.05fF
C261 a_18760_101.n1 GND 0.13fF
C262 a_18760_101.n2 GND 0.04fF
C263 a_18760_101.n3 GND 0.18fF
C264 a_4447_989.n0 GND 0.88fF
C265 a_4447_989.n1 GND 0.88fF
C266 a_4447_989.n2 GND 0.81fF
C267 a_4447_989.n3 GND 0.99fF
C268 a_4447_989.n4 GND 1.37fF
C269 a_4447_989.n5 GND 0.82fF
C270 a_4447_989.n6 GND 11.47fF
C271 a_4447_989.n7 GND 0.80fF
C272 a_4447_989.t12 GND 1.15fF
C273 a_4447_989.n8 GND 1.40fF
C274 a_4447_989.n9 GND 14.41fF
C275 a_4447_989.n10 GND 0.10fF
C276 a_4447_989.n11 GND 0.12fF
C277 a_4447_989.n12 GND 0.49fF
C278 a_4447_989.n13 GND 1.20fF
C279 a_4447_989.n14 GND 1.08fF
C280 a_4447_989.n15 GND 1.06fF
C281 a_4447_989.n16 GND 1.12fF
C282 a_4125_1050.n0 GND 0.38fF
C283 a_4125_1050.n1 GND 0.38fF
C284 a_4125_1050.n2 GND 0.32fF
C285 a_4125_1050.n3 GND 0.64fF
C286 a_4125_1050.n4 GND 0.33fF
C287 a_4125_1050.n5 GND 0.70fF
C288 a_4125_1050.n6 GND 0.44fF
C289 a_4125_1050.n7 GND 0.46fF
C290 a_4125_1050.n8 GND 0.49fF
C291 a_17533_1051.n0 GND 0.36fF
C292 a_17533_1051.n1 GND 0.32fF
C293 a_17533_1051.n2 GND 0.52fF
C294 a_17533_1051.n3 GND 0.30fF
C295 a_17533_1051.n4 GND 0.80fF
C296 a_17533_1051.n5 GND 0.43fF
C297 a_7973_1050.n0 GND 0.40fF
C298 a_7973_1050.n1 GND 0.40fF
C299 a_7973_1050.n2 GND 0.38fF
C300 a_7973_1050.n3 GND 0.65fF
C301 a_7973_1050.n4 GND 0.04fF
C302 a_7973_1050.n5 GND 0.05fF
C303 a_7973_1050.n6 GND 0.03fF
C304 a_7973_1050.n7 GND 0.17fF
C305 a_7973_1050.n8 GND 0.70fF
C306 a_7973_1050.n9 GND 0.52fF
C307 a_7973_1050.n10 GND 0.48fF
C308 a_7973_1050.n11 GND 0.50fF
C309 a_13840_210.n0 GND 0.02fF
C310 a_13840_210.n1 GND 0.09fF
C311 a_13840_210.n2 GND 0.12fF
C312 a_13840_210.n3 GND 0.08fF
C313 a_13840_210.n4 GND 0.08fF
C314 a_13840_210.n5 GND 0.02fF
C315 a_13840_210.t1 GND 0.29fF
C316 a_13840_210.n6 GND 0.09fF
C317 a_13840_210.n7 GND 0.02fF
C318 a_13840_210.n8 GND 0.13fF
C319 a_13840_210.n9 GND 0.02fF
C320 a_13840_210.n10 GND 0.03fF
C321 a_13840_210.n11 GND 0.03fF
C322 a_6049_1050.n0 GND 0.48fF
C323 a_6049_1050.n1 GND 0.83fF
C324 a_6049_1050.n2 GND 0.48fF
C325 a_6049_1050.n3 GND 0.60fF
C326 a_6049_1050.n4 GND 1.20fF
C327 a_6049_1050.n5 GND 0.05fF
C328 a_6049_1050.n6 GND 0.07fF
C329 a_6049_1050.n7 GND 0.04fF
C330 a_6049_1050.n8 GND 0.22fF
C331 a_6049_1050.n9 GND 0.72fF
C332 a_6049_1050.n10 GND 0.50fF
C333 a_6049_1050.n11 GND 0.64fF
C334 a_6049_1050.n12 GND 0.61fF
C335 a_6049_1050.n13 GND 0.66fF
C336 a_6049_1050.n14 GND 0.50fF
C337 a_3258_210.n0 GND 0.02fF
C338 a_3258_210.n1 GND 0.09fF
C339 a_3258_210.n2 GND 0.12fF
C340 a_3258_210.n3 GND 0.08fF
C341 a_3258_210.n4 GND 0.08fF
C342 a_3258_210.n5 GND 0.02fF
C343 a_3258_210.t1 GND 0.29fF
C344 a_3258_210.n6 GND 0.09fF
C345 a_3258_210.n7 GND 0.02fF
C346 a_3258_210.n8 GND 0.13fF
C347 a_3258_210.n9 GND 0.02fF
C348 a_3258_210.n10 GND 0.03fF
C349 a_3258_210.n11 GND 0.02fF
C350 a_2977_103.n0 GND 0.13fF
C351 a_2977_103.n1 GND 0.04fF
C352 a_2977_103.n2 GND 0.09fF
C353 a_2977_103.n3 GND 0.07fF
C354 a_2977_103.n4 GND 0.08fF
C355 a_2977_103.n5 GND 0.03fF
C356 a_15764_210.n0 GND 0.07fF
C357 a_15764_210.n1 GND 0.09fF
C358 a_15764_210.n2 GND 0.12fF
C359 a_15764_210.n3 GND 0.08fF
C360 a_15764_210.n4 GND 0.02fF
C361 a_15764_210.n5 GND 0.03fF
C362 a_15764_210.n6 GND 0.02fF
C363 a_15764_210.n7 GND 0.03fF
C364 a_15764_210.n8 GND 0.02fF
C365 a_15764_210.n9 GND 0.13fF
C366 a_15764_210.n10 GND 0.08fF
C367 a_15764_210.n11 GND 0.02fF
C368 a_15764_210.t0 GND 0.31fF
C369 a_15991_989.n0 GND 0.40fF
C370 a_15991_989.n1 GND 0.26fF
C371 a_15991_989.n2 GND 0.80fF
C372 a_15991_989.n3 GND 0.25fF
C373 a_15991_989.n4 GND 0.52fF
C374 a_15991_989.n5 GND 0.53fF
C375 a_15991_989.n6 GND 0.40fF
C376 a_15991_989.t7 GND 0.50fF
C377 a_15991_989.n7 GND 0.91fF
C378 a_15991_989.n8 GND 0.04fF
C379 a_15991_989.n9 GND 0.06fF
C380 a_15991_989.n10 GND 0.04fF
C381 a_15991_989.n11 GND 0.17fF
C382 a_15991_989.n12 GND 0.86fF
C383 a_15991_989.n13 GND 0.42fF
C384 a_15991_989.n14 GND 0.43fF
C385 a_15991_989.n15 GND 0.51fF
C386 a_15991_989.n16 GND 0.49fF
C387 a_15991_989.n17 GND 0.40fF
C388 a_1334_210.n0 GND 0.07fF
C389 a_1334_210.n1 GND 0.09fF
C390 a_1334_210.n2 GND 0.12fF
C391 a_1334_210.n3 GND 0.08fF
C392 a_1334_210.n4 GND 0.02fF
C393 a_1334_210.n5 GND 0.03fF
C394 a_1334_210.n6 GND 0.05fF
C395 a_1334_210.n7 GND 0.02fF
C396 a_1334_210.n8 GND 0.14fF
C397 a_1334_210.n9 GND 0.08fF
C398 a_1334_210.n10 GND 0.02fF
C399 a_1334_210.t0 GND 0.31fF
C400 a_1053_103.n0 GND 0.13fF
C401 a_1053_103.n1 GND 0.04fF
C402 a_1053_103.n2 GND 0.09fF
C403 a_1053_103.n3 GND 0.07fF
C404 a_1053_103.n4 GND 0.08fF
C405 a_1053_103.n5 GND 0.03fF
C406 a_7106_210.n0 GND 0.07fF
C407 a_7106_210.n1 GND 0.09fF
C408 a_7106_210.n2 GND 0.12fF
C409 a_7106_210.n3 GND 0.08fF
C410 a_7106_210.n4 GND 0.02fF
C411 a_7106_210.n5 GND 0.03fF
C412 a_7106_210.n6 GND 0.05fF
C413 a_7106_210.n7 GND 0.02fF
C414 a_7106_210.n8 GND 0.14fF
C415 a_7106_210.n9 GND 0.08fF
C416 a_7106_210.n10 GND 0.02fF
C417 a_7106_210.t0 GND 0.31fF
C418 a_6825_103.n0 GND 0.13fF
C419 a_6825_103.n1 GND 0.04fF
C420 a_6825_103.n2 GND 0.09fF
C421 a_6825_103.n3 GND 0.07fF
C422 a_6825_103.n4 GND 0.08fF
C423 a_6825_103.n5 GND 0.03fF
C424 a_5182_210.n0 GND 0.02fF
C425 a_5182_210.n1 GND 0.09fF
C426 a_5182_210.t1 GND 0.23fF
C427 a_5182_210.n2 GND 0.10fF
C428 a_5182_210.n3 GND 0.07fF
C429 a_5182_210.n4 GND 0.04fF
C430 a_5182_210.n5 GND 0.08fF
C431 a_5182_210.n6 GND 0.09fF
C432 a_5182_210.n7 GND 0.04fF
C433 a_5182_210.n8 GND 0.02fF
C434 a_5182_210.n9 GND 0.01fF
C435 a_5182_210.n10 GND 0.13fF
C436 a_5182_210.n11 GND 0.02fF
C437 a_5182_210.n12 GND 0.03fF
C438 a_5182_210.n13 GND 0.02fF
C439 a_4901_103.n0 GND 0.13fF
C440 a_4901_103.n1 GND 0.04fF
C441 a_4901_103.n2 GND 0.09fF
C442 a_4901_103.n3 GND 0.07fF
C443 a_4901_103.n4 GND 0.08fF
C444 a_4901_103.n5 GND 0.03fF
C445 a_6371_989.n0 GND 0.59fF
C446 a_6371_989.n1 GND 1.98fF
C447 a_6371_989.n2 GND 0.60fF
C448 a_6371_989.t11 GND 0.96fF
C449 a_6371_989.n3 GND 1.15fF
C450 a_6371_989.n4 GND 3.61fF
C451 a_6371_989.n5 GND 0.07fF
C452 a_6371_989.n6 GND 0.10fF
C453 a_6371_989.n7 GND 0.06fF
C454 a_6371_989.n8 GND 0.41fF
C455 a_6371_989.n9 GND 0.94fF
C456 a_6371_989.n10 GND 0.71fF
C457 a_6371_989.n11 GND 0.90fF
C458 a_6371_989.n12 GND 0.85fF
C459 a_6371_989.n13 GND 0.81fF
C460 a_6371_989.n14 GND 0.71fF
C461 a_10219_989.n0 GND 0.77fF
C462 a_10219_989.n1 GND 0.58fF
C463 a_10219_989.n2 GND 1.41fF
C464 a_10219_989.n3 GND 0.55fF
C465 a_10219_989.n4 GND 0.77fF
C466 a_10219_989.n5 GND 7.58fF
C467 a_10219_989.n6 GND 0.76fF
C468 a_10219_989.t13 GND 0.96fF
C469 a_10219_989.n7 GND 1.73fF
C470 a_10219_989.n8 GND 0.08fF
C471 a_10219_989.n9 GND 0.11fF
C472 a_10219_989.n10 GND 0.07fF
C473 a_10219_989.n11 GND 0.33fF
C474 a_10219_989.n12 GND 1.64fF
C475 a_10219_989.n13 GND 4.82fF
C476 a_10219_989.n14 GND 0.82fF
C477 a_10219_989.n15 GND 0.98fF
C478 a_10219_989.n16 GND 0.93fF
C479 a_10219_989.n17 GND 0.77fF
C480 SN.n0 GND 0.85fF
C481 SN.t10 GND 0.78fF
C482 SN.n1 GND 2.33fF
C483 SN.n2 GND 0.84fF
C484 SN.t12 GND 0.78fF
C485 SN.n3 GND 0.78fF
C486 SN.n4 GND 5.12fF
C487 SN.n5 GND 0.85fF
C488 SN.t9 GND 0.78fF
C489 SN.n6 GND 0.77fF
C490 SN.n7 GND 4.43fF
C491 SN.n8 GND 0.84fF
C492 SN.t3 GND 0.78fF
C493 SN.n9 GND 0.78fF
C494 SN.n10 GND 4.43fF
C495 SN.n11 GND 0.85fF
C496 SN.t1 GND 0.78fF
C497 SN.n12 GND 0.77fF
C498 SN.n13 GND 4.43fF
C499 SN.t17 GND 0.78fF
C500 SN.n14 GND 0.84fF
C501 SN.n15 GND 0.78fF
C502 SN.n16 GND 2.23fF
C503 a_2201_1050.n0 GND 0.36fF
C504 a_2201_1050.n1 GND 0.36fF
C505 a_2201_1050.n2 GND 0.35fF
C506 a_2201_1050.n3 GND 0.59fF
C507 a_2201_1050.n4 GND 0.04fF
C508 a_2201_1050.n5 GND 0.05fF
C509 a_2201_1050.n6 GND 0.03fF
C510 a_2201_1050.n7 GND 0.15fF
C511 a_2201_1050.n8 GND 0.64fF
C512 a_2201_1050.n9 GND 0.47fF
C513 a_2201_1050.n10 GND 0.43fF
C514 a_2201_1050.n11 GND 0.46fF
C515 a_277_1050.n0 GND 0.37fF
C516 a_277_1050.n1 GND 0.63fF
C517 a_277_1050.n2 GND 0.37fF
C518 a_277_1050.n3 GND 0.46fF
C519 a_277_1050.n4 GND 0.91fF
C520 a_277_1050.n5 GND 0.04fF
C521 a_277_1050.n6 GND 0.05fF
C522 a_277_1050.n7 GND 0.03fF
C523 a_277_1050.n8 GND 0.16fF
C524 a_277_1050.n9 GND 0.55fF
C525 a_277_1050.n10 GND 0.38fF
C526 a_277_1050.n11 GND 0.49fF
C527 a_277_1050.n12 GND 0.46fF
C528 a_277_1050.n13 GND 0.50fF
C529 a_277_1050.n14 GND 0.38fF
C530 a_13745_1050.n0 GND 0.40fF
C531 a_13745_1050.n1 GND 0.40fF
C532 a_13745_1050.n2 GND 0.38fF
C533 a_13745_1050.n3 GND 0.65fF
C534 a_13745_1050.n4 GND 0.04fF
C535 a_13745_1050.n5 GND 0.05fF
C536 a_13745_1050.n6 GND 0.03fF
C537 a_13745_1050.n7 GND 0.17fF
C538 a_13745_1050.n8 GND 0.70fF
C539 a_13745_1050.n9 GND 0.52fF
C540 a_13745_1050.n10 GND 0.48fF
C541 a_13745_1050.n11 GND 0.50fF
C542 a_7333_989.n0 GND 0.69fF
C543 a_7333_989.n1 GND 0.53fF
C544 a_7333_989.t15 GND 0.97fF
C545 a_7333_989.n2 GND 1.49fF
C546 a_7333_989.n3 GND 0.53fF
C547 a_7333_989.t13 GND 0.97fF
C548 a_7333_989.n4 GND 0.73fF
C549 a_7333_989.n5 GND 0.53fF
C550 a_7333_989.t12 GND 0.97fF
C551 a_7333_989.n6 GND 1.04fF
C552 a_7333_989.n7 GND 1.92fF
C553 a_7333_989.n8 GND 2.63fF
C554 a_7333_989.n9 GND 0.64fF
C555 a_7333_989.n10 GND 0.95fF
C556 a_7333_989.n11 GND 0.73fF
C557 a_7333_989.n12 GND 0.87fF
C558 a_7333_989.n13 GND 0.83fF
C559 a_7333_989.n14 GND 0.69fF
C560 a_9030_210.n0 GND 0.02fF
C561 a_9030_210.n1 GND 0.09fF
C562 a_9030_210.t1 GND 0.23fF
C563 a_9030_210.n2 GND 0.10fF
C564 a_9030_210.n3 GND 0.07fF
C565 a_9030_210.n4 GND 0.04fF
C566 a_9030_210.n5 GND 0.08fF
C567 a_9030_210.n6 GND 0.09fF
C568 a_9030_210.n7 GND 0.04fF
C569 a_9030_210.n8 GND 0.02fF
C570 a_9030_210.n9 GND 0.01fF
C571 a_9030_210.n10 GND 0.13fF
C572 a_9030_210.n11 GND 0.02fF
C573 a_9030_210.n12 GND 0.03fF
C574 a_9030_210.n13 GND 0.03fF
C575 a_11821_1050.n0 GND 0.48fF
C576 a_11821_1050.n1 GND 0.83fF
C577 a_11821_1050.n2 GND 0.48fF
C578 a_11821_1050.n3 GND 0.60fF
C579 a_11821_1050.n4 GND 1.20fF
C580 a_11821_1050.n5 GND 0.05fF
C581 a_11821_1050.n6 GND 0.07fF
C582 a_11821_1050.n7 GND 0.04fF
C583 a_11821_1050.n8 GND 0.22fF
C584 a_11821_1050.n9 GND 0.72fF
C585 a_11821_1050.n10 GND 0.50fF
C586 a_11821_1050.n11 GND 0.64fF
C587 a_11821_1050.n12 GND 0.61fF
C588 a_11821_1050.n13 GND 0.66fF
C589 a_11821_1050.n14 GND 0.50fF
C590 a_12143_989.n0 GND 0.70fF
C591 a_12143_989.n1 GND 0.58fF
C592 a_12143_989.n2 GND 1.96fF
C593 a_12143_989.n3 GND 0.59fF
C594 a_12143_989.t11 GND 0.95fF
C595 a_12143_989.n4 GND 1.13fF
C596 a_12143_989.n5 GND 3.56fF
C597 a_12143_989.n6 GND 0.07fF
C598 a_12143_989.n7 GND 0.10fF
C599 a_12143_989.n8 GND 0.06fF
C600 a_12143_989.n9 GND 0.40fF
C601 a_12143_989.n10 GND 0.93fF
C602 a_12143_989.n11 GND 0.80fF
C603 a_12143_989.n12 GND 0.89fF
C604 a_12143_989.n13 GND 0.84fF
C605 a_12143_989.n14 GND 0.70fF
C606 a_1561_989.n0 GND 0.63fF
C607 a_1561_989.n1 GND 0.49fF
C608 a_1561_989.t14 GND 0.89fF
C609 a_1561_989.n2 GND 1.37fF
C610 a_1561_989.n3 GND 0.49fF
C611 a_1561_989.t11 GND 0.89fF
C612 a_1561_989.n4 GND 0.67fF
C613 a_1561_989.n5 GND 0.49fF
C614 a_1561_989.t13 GND 0.89fF
C615 a_1561_989.n6 GND 0.96fF
C616 a_1561_989.n7 GND 1.76fF
C617 a_1561_989.n8 GND 2.42fF
C618 a_1561_989.n9 GND 0.06fF
C619 a_1561_989.n10 GND 0.09fF
C620 a_1561_989.n11 GND 0.05fF
C621 a_1561_989.n12 GND 0.41fF
C622 a_1561_989.n13 GND 0.84fF
C623 a_1561_989.n14 GND 0.67fF
C624 a_1561_989.n15 GND 0.80fF
C625 a_1561_989.n16 GND 0.76fF
C626 a_1561_989.n17 GND 0.63fF
C627 a_3939_103.n0 GND 0.13fF
C628 a_3939_103.n1 GND 0.04fF
C629 a_3939_103.n2 GND 0.09fF
C630 a_3939_103.n3 GND 0.07fF
C631 a_3939_103.n4 GND 0.08fF
C632 a_3939_103.n5 GND 0.03fF
C633 a_9897_1050.n0 GND 0.40fF
C634 a_9897_1050.n1 GND 0.33fF
C635 a_9897_1050.n2 GND 0.67fF
C636 a_9897_1050.n3 GND 0.35fF
C637 a_9897_1050.n4 GND 0.73fF
C638 a_9897_1050.n5 GND 0.46fF
C639 a_9897_1050.n6 GND 0.51fF
C640 a_9897_1050.n7 GND 0.48fF
C641 a_9897_1050.n8 GND 0.40fF
C642 a_599_989.n0 GND 0.53fF
C643 a_599_989.n1 GND 0.44fF
C644 a_599_989.n2 GND 1.48fF
C645 a_599_989.n3 GND 0.45fF
C646 a_599_989.t10 GND 0.72fF
C647 a_599_989.n4 GND 0.86fF
C648 a_599_989.n5 GND 2.70fF
C649 a_599_989.n6 GND 0.46fF
C650 a_599_989.n7 GND 0.73fF
C651 a_599_989.n8 GND 0.61fF
C652 a_599_989.n9 GND 0.68fF
C653 a_599_989.n10 GND 0.64fF
C654 a_599_989.n11 GND 0.53fF
C655 VDD.n1 GND 0.04fF
C656 VDD.n2 GND 0.14fF
C657 VDD.n3 GND 0.03fF
C658 VDD.n4 GND 0.02fF
C659 VDD.n5 GND 0.06fF
C660 VDD.n6 GND 0.02fF
C661 VDD.n7 GND 0.02fF
C662 VDD.n8 GND 0.02fF
C663 VDD.n9 GND 0.02fF
C664 VDD.n10 GND 0.02fF
C665 VDD.n11 GND 0.02fF
C666 VDD.n12 GND 0.02fF
C667 VDD.n13 GND 0.02fF
C668 VDD.n14 GND 0.04fF
C669 VDD.n15 GND 0.01fF
C670 VDD.n20 GND 0.49fF
C671 VDD.n21 GND 0.29fF
C672 VDD.n22 GND 0.02fF
C673 VDD.n23 GND 0.04fF
C674 VDD.n24 GND 0.26fF
C675 VDD.n25 GND 0.01fF
C676 VDD.n26 GND 0.02fF
C677 VDD.n27 GND 0.01fF
C678 VDD.n28 GND 0.18fF
C679 VDD.n29 GND 0.01fF
C680 VDD.n30 GND 0.02fF
C681 VDD.n31 GND 0.09fF
C682 VDD.n32 GND 0.02fF
C683 VDD.n33 GND 0.03fF
C684 VDD.n34 GND 0.03fF
C685 VDD.n35 GND 0.15fF
C686 VDD.n36 GND 0.02fF
C687 VDD.n37 GND 0.03fF
C688 VDD.n38 GND 0.03fF
C689 VDD.n39 GND 0.18fF
C690 VDD.n40 GND 0.01fF
C691 VDD.n41 GND 0.02fF
C692 VDD.n42 GND 0.02fF
C693 VDD.n43 GND 0.26fF
C694 VDD.n44 GND 0.01fF
C695 VDD.n45 GND 0.02fF
C696 VDD.n46 GND 0.02fF
C697 VDD.n47 GND 0.29fF
C698 VDD.n48 GND 0.01fF
C699 VDD.n49 GND 0.02fF
C700 VDD.n50 GND 0.04fF
C701 VDD.n51 GND 0.06fF
C702 VDD.n52 GND 0.02fF
C703 VDD.n53 GND 0.02fF
C704 VDD.n54 GND 0.02fF
C705 VDD.n55 GND 0.02fF
C706 VDD.n56 GND 0.02fF
C707 VDD.n57 GND 0.02fF
C708 VDD.n58 GND 0.02fF
C709 VDD.n59 GND 0.02fF
C710 VDD.n60 GND 0.02fF
C711 VDD.n61 GND 0.02fF
C712 VDD.n62 GND 0.02fF
C713 VDD.n63 GND 0.03fF
C714 VDD.n64 GND 0.03fF
C715 VDD.n65 GND 0.23fF
C716 VDD.n66 GND 0.02fF
C717 VDD.n67 GND 0.02fF
C718 VDD.n69 GND 0.02fF
C719 VDD.n73 GND 0.29fF
C720 VDD.n74 GND 0.29fF
C721 VDD.n75 GND 0.01fF
C722 VDD.n76 GND 0.02fF
C723 VDD.n77 GND 0.04fF
C724 VDD.n78 GND 0.26fF
C725 VDD.n79 GND 0.01fF
C726 VDD.n80 GND 0.02fF
C727 VDD.n81 GND 0.02fF
C728 VDD.n82 GND 0.18fF
C729 VDD.n83 GND 0.01fF
C730 VDD.n84 GND 0.02fF
C731 VDD.n85 GND 0.02fF
C732 VDD.n86 GND 0.15fF
C733 VDD.n87 GND 0.02fF
C734 VDD.n88 GND 0.03fF
C735 VDD.n89 GND 0.03fF
C736 VDD.n90 GND 0.02fF
C737 VDD.n91 GND 0.03fF
C738 VDD.n92 GND 0.03fF
C739 VDD.n93 GND 0.18fF
C740 VDD.n94 GND 0.01fF
C741 VDD.n95 GND 0.02fF
C742 VDD.n96 GND 0.02fF
C743 VDD.n97 GND 0.26fF
C744 VDD.n98 GND 0.01fF
C745 VDD.n99 GND 0.02fF
C746 VDD.n100 GND 0.02fF
C747 VDD.n101 GND 0.29fF
C748 VDD.n102 GND 0.01fF
C749 VDD.n103 GND 0.02fF
C750 VDD.n104 GND 0.04fF
C751 VDD.n105 GND 0.23fF
C752 VDD.n106 GND 0.02fF
C753 VDD.n107 GND 0.02fF
C754 VDD.n108 GND 0.02fF
C755 VDD.n109 GND 0.06fF
C756 VDD.n110 GND 0.02fF
C757 VDD.n111 GND 0.02fF
C758 VDD.n112 GND 0.02fF
C759 VDD.n113 GND 0.02fF
C760 VDD.n114 GND 0.02fF
C761 VDD.n115 GND 0.02fF
C762 VDD.n116 GND 0.02fF
C763 VDD.n117 GND 0.02fF
C764 VDD.n118 GND 0.02fF
C765 VDD.n119 GND 0.02fF
C766 VDD.n120 GND 0.03fF
C767 VDD.n121 GND 0.03fF
C768 VDD.n122 GND 0.02fF
C769 VDD.n126 GND 0.29fF
C770 VDD.n127 GND 0.29fF
C771 VDD.n128 GND 0.01fF
C772 VDD.n129 GND 0.02fF
C773 VDD.n130 GND 0.04fF
C774 VDD.n131 GND 0.07fF
C775 VDD.n132 GND 0.26fF
C776 VDD.n133 GND 0.01fF
C777 VDD.n134 GND 0.01fF
C778 VDD.n135 GND 0.02fF
C779 VDD.n136 GND 0.18fF
C780 VDD.n137 GND 0.01fF
C781 VDD.n138 GND 0.02fF
C782 VDD.n139 GND 0.02fF
C783 VDD.n140 GND 0.09fF
C784 VDD.n141 GND 0.05fF
C785 VDD.n142 GND 0.02fF
C786 VDD.n143 GND 0.02fF
C787 VDD.n144 GND 0.03fF
C788 VDD.n145 GND 0.15fF
C789 VDD.n146 GND 0.02fF
C790 VDD.n147 GND 0.02fF
C791 VDD.n148 GND 0.03fF
C792 VDD.n149 GND 0.18fF
C793 VDD.n150 GND 0.01fF
C794 VDD.n151 GND 0.02fF
C795 VDD.n152 GND 0.02fF
C796 VDD.n153 GND 0.07fF
C797 VDD.n154 GND 0.26fF
C798 VDD.n155 GND 0.01fF
C799 VDD.n156 GND 0.01fF
C800 VDD.n157 GND 0.02fF
C801 VDD.n158 GND 0.29fF
C802 VDD.n159 GND 0.01fF
C803 VDD.n160 GND 0.02fF
C804 VDD.n161 GND 0.04fF
C805 VDD.n162 GND 0.28fF
C806 VDD.n163 GND 0.02fF
C807 VDD.n164 GND 0.02fF
C808 VDD.n165 GND 0.02fF
C809 VDD.n166 GND 0.06fF
C810 VDD.n167 GND 0.02fF
C811 VDD.n168 GND 0.02fF
C812 VDD.n169 GND 0.02fF
C813 VDD.n170 GND 0.02fF
C814 VDD.n171 GND 0.02fF
C815 VDD.n172 GND 0.02fF
C816 VDD.n173 GND 0.02fF
C817 VDD.n174 GND 0.02fF
C818 VDD.n175 GND 0.02fF
C819 VDD.n176 GND 0.02fF
C820 VDD.n177 GND 0.03fF
C821 VDD.n178 GND 0.03fF
C822 VDD.n179 GND 0.02fF
C823 VDD.n183 GND 0.29fF
C824 VDD.n184 GND 0.29fF
C825 VDD.n185 GND 0.01fF
C826 VDD.n186 GND 0.02fF
C827 VDD.n187 GND 0.04fF
C828 VDD.n188 GND 0.29fF
C829 VDD.n189 GND 0.01fF
C830 VDD.n190 GND 0.02fF
C831 VDD.n191 GND 0.02fF
C832 VDD.n192 GND 0.24fF
C833 VDD.n193 GND 0.01fF
C834 VDD.n194 GND 0.07fF
C835 VDD.n195 GND 0.02fF
C836 VDD.n196 GND 0.18fF
C837 VDD.n197 GND 0.01fF
C838 VDD.n198 GND 0.02fF
C839 VDD.n199 GND 0.02fF
C840 VDD.n200 GND 0.17fF
C841 VDD.n201 GND 0.01fF
C842 VDD.n202 GND 0.09fF
C843 VDD.n203 GND 0.05fF
C844 VDD.n204 GND 0.02fF
C845 VDD.n205 GND 0.02fF
C846 VDD.n206 GND 0.15fF
C847 VDD.n207 GND 0.02fF
C848 VDD.n208 GND 0.02fF
C849 VDD.n209 GND 0.03fF
C850 VDD.n210 GND 0.16fF
C851 VDD.n211 GND 0.02fF
C852 VDD.n212 GND 0.02fF
C853 VDD.n213 GND 0.03fF
C854 VDD.n214 GND 0.09fF
C855 VDD.n215 GND 0.05fF
C856 VDD.n216 GND 0.17fF
C857 VDD.n217 GND 0.01fF
C858 VDD.n218 GND 0.02fF
C859 VDD.n219 GND 0.02fF
C860 VDD.n220 GND 0.18fF
C861 VDD.n221 GND 0.01fF
C862 VDD.n222 GND 0.02fF
C863 VDD.n223 GND 0.02fF
C864 VDD.n224 GND 0.07fF
C865 VDD.n225 GND 0.24fF
C866 VDD.n226 GND 0.01fF
C867 VDD.n227 GND 0.01fF
C868 VDD.n228 GND 0.02fF
C869 VDD.n229 GND 0.29fF
C870 VDD.n230 GND 0.01fF
C871 VDD.n231 GND 0.02fF
C872 VDD.n232 GND 0.02fF
C873 VDD.n233 GND 0.29fF
C874 VDD.n234 GND 0.01fF
C875 VDD.n235 GND 0.02fF
C876 VDD.n236 GND 0.04fF
C877 VDD.n237 GND 0.33fF
C878 VDD.n238 GND 0.02fF
C879 VDD.n239 GND 0.02fF
C880 VDD.n240 GND 0.02fF
C881 VDD.n241 GND 0.06fF
C882 VDD.n242 GND 0.02fF
C883 VDD.n243 GND 0.02fF
C884 VDD.n244 GND 0.02fF
C885 VDD.n245 GND 0.02fF
C886 VDD.n246 GND 0.02fF
C887 VDD.n247 GND 0.02fF
C888 VDD.n248 GND 0.02fF
C889 VDD.n249 GND 0.02fF
C890 VDD.n250 GND 0.02fF
C891 VDD.n251 GND 0.02fF
C892 VDD.n252 GND 0.03fF
C893 VDD.n253 GND 0.03fF
C894 VDD.n254 GND 0.02fF
C895 VDD.n258 GND 0.29fF
C896 VDD.n259 GND 0.29fF
C897 VDD.n260 GND 0.01fF
C898 VDD.n261 GND 0.02fF
C899 VDD.n262 GND 0.04fF
C900 VDD.n263 GND 0.29fF
C901 VDD.n264 GND 0.01fF
C902 VDD.n265 GND 0.02fF
C903 VDD.n266 GND 0.02fF
C904 VDD.n267 GND 0.24fF
C905 VDD.n268 GND 0.01fF
C906 VDD.n269 GND 0.07fF
C907 VDD.n270 GND 0.02fF
C908 VDD.n271 GND 0.18fF
C909 VDD.n272 GND 0.01fF
C910 VDD.n273 GND 0.02fF
C911 VDD.n274 GND 0.02fF
C912 VDD.n275 GND 0.17fF
C913 VDD.n276 GND 0.01fF
C914 VDD.n277 GND 0.09fF
C915 VDD.n278 GND 0.05fF
C916 VDD.n279 GND 0.02fF
C917 VDD.n280 GND 0.02fF
C918 VDD.n281 GND 0.15fF
C919 VDD.n282 GND 0.02fF
C920 VDD.n283 GND 0.02fF
C921 VDD.n284 GND 0.03fF
C922 VDD.n285 GND 0.16fF
C923 VDD.n286 GND 0.02fF
C924 VDD.n287 GND 0.02fF
C925 VDD.n288 GND 0.03fF
C926 VDD.n289 GND 0.09fF
C927 VDD.n290 GND 0.05fF
C928 VDD.n291 GND 0.17fF
C929 VDD.n292 GND 0.01fF
C930 VDD.n293 GND 0.02fF
C931 VDD.n294 GND 0.02fF
C932 VDD.n295 GND 0.18fF
C933 VDD.n296 GND 0.01fF
C934 VDD.n297 GND 0.02fF
C935 VDD.n298 GND 0.02fF
C936 VDD.n299 GND 0.07fF
C937 VDD.n300 GND 0.24fF
C938 VDD.n301 GND 0.01fF
C939 VDD.n302 GND 0.01fF
C940 VDD.n303 GND 0.02fF
C941 VDD.n304 GND 0.29fF
C942 VDD.n305 GND 0.01fF
C943 VDD.n306 GND 0.02fF
C944 VDD.n307 GND 0.02fF
C945 VDD.n308 GND 0.29fF
C946 VDD.n309 GND 0.01fF
C947 VDD.n310 GND 0.02fF
C948 VDD.n311 GND 0.04fF
C949 VDD.n312 GND 0.33fF
C950 VDD.n313 GND 0.02fF
C951 VDD.n314 GND 0.02fF
C952 VDD.n315 GND 0.02fF
C953 VDD.n316 GND 0.06fF
C954 VDD.n317 GND 0.02fF
C955 VDD.n318 GND 0.02fF
C956 VDD.n319 GND 0.02fF
C957 VDD.n320 GND 0.02fF
C958 VDD.n321 GND 0.02fF
C959 VDD.n322 GND 0.02fF
C960 VDD.n323 GND 0.02fF
C961 VDD.n324 GND 0.02fF
C962 VDD.n325 GND 0.02fF
C963 VDD.n326 GND 0.02fF
C964 VDD.n327 GND 0.03fF
C965 VDD.n328 GND 0.03fF
C966 VDD.n329 GND 0.02fF
C967 VDD.n333 GND 0.29fF
C968 VDD.n334 GND 0.29fF
C969 VDD.n335 GND 0.01fF
C970 VDD.n336 GND 0.02fF
C971 VDD.n337 GND 0.04fF
C972 VDD.n338 GND 0.29fF
C973 VDD.n339 GND 0.01fF
C974 VDD.n340 GND 0.02fF
C975 VDD.n341 GND 0.02fF
C976 VDD.n342 GND 0.24fF
C977 VDD.n343 GND 0.01fF
C978 VDD.n344 GND 0.07fF
C979 VDD.n345 GND 0.02fF
C980 VDD.n346 GND 0.18fF
C981 VDD.n347 GND 0.01fF
C982 VDD.n348 GND 0.02fF
C983 VDD.n349 GND 0.02fF
C984 VDD.n350 GND 0.17fF
C985 VDD.n351 GND 0.01fF
C986 VDD.n352 GND 0.09fF
C987 VDD.n353 GND 0.05fF
C988 VDD.n354 GND 0.02fF
C989 VDD.n355 GND 0.02fF
C990 VDD.n356 GND 0.15fF
C991 VDD.n357 GND 0.02fF
C992 VDD.n358 GND 0.02fF
C993 VDD.n359 GND 0.03fF
C994 VDD.n360 GND 0.16fF
C995 VDD.n361 GND 0.02fF
C996 VDD.n362 GND 0.02fF
C997 VDD.n363 GND 0.03fF
C998 VDD.n364 GND 0.09fF
C999 VDD.n365 GND 0.05fF
C1000 VDD.n366 GND 0.17fF
C1001 VDD.n367 GND 0.01fF
C1002 VDD.n368 GND 0.02fF
C1003 VDD.n369 GND 0.02fF
C1004 VDD.n370 GND 0.18fF
C1005 VDD.n371 GND 0.01fF
C1006 VDD.n372 GND 0.02fF
C1007 VDD.n373 GND 0.02fF
C1008 VDD.n374 GND 0.07fF
C1009 VDD.n375 GND 0.24fF
C1010 VDD.n376 GND 0.01fF
C1011 VDD.n377 GND 0.01fF
C1012 VDD.n378 GND 0.02fF
C1013 VDD.n379 GND 0.29fF
C1014 VDD.n380 GND 0.01fF
C1015 VDD.n381 GND 0.02fF
C1016 VDD.n382 GND 0.02fF
C1017 VDD.n383 GND 0.29fF
C1018 VDD.n384 GND 0.01fF
C1019 VDD.n385 GND 0.02fF
C1020 VDD.n386 GND 0.04fF
C1021 VDD.n387 GND 0.33fF
C1022 VDD.n388 GND 0.02fF
C1023 VDD.n389 GND 0.02fF
C1024 VDD.n390 GND 0.02fF
C1025 VDD.n391 GND 0.06fF
C1026 VDD.n392 GND 0.02fF
C1027 VDD.n393 GND 0.02fF
C1028 VDD.n394 GND 0.02fF
C1029 VDD.n395 GND 0.02fF
C1030 VDD.n396 GND 0.02fF
C1031 VDD.n397 GND 0.02fF
C1032 VDD.n398 GND 0.02fF
C1033 VDD.n399 GND 0.02fF
C1034 VDD.n400 GND 0.02fF
C1035 VDD.n401 GND 0.02fF
C1036 VDD.n402 GND 0.03fF
C1037 VDD.n403 GND 0.03fF
C1038 VDD.n404 GND 0.02fF
C1039 VDD.n408 GND 0.29fF
C1040 VDD.n409 GND 0.29fF
C1041 VDD.n410 GND 0.01fF
C1042 VDD.n411 GND 0.02fF
C1043 VDD.n412 GND 0.04fF
C1044 VDD.n413 GND 0.29fF
C1045 VDD.n414 GND 0.01fF
C1046 VDD.n415 GND 0.02fF
C1047 VDD.n416 GND 0.02fF
C1048 VDD.n417 GND 0.24fF
C1049 VDD.n418 GND 0.01fF
C1050 VDD.n419 GND 0.07fF
C1051 VDD.n420 GND 0.02fF
C1052 VDD.n421 GND 0.18fF
C1053 VDD.n422 GND 0.01fF
C1054 VDD.n423 GND 0.02fF
C1055 VDD.n424 GND 0.02fF
C1056 VDD.n425 GND 0.17fF
C1057 VDD.n426 GND 0.01fF
C1058 VDD.n427 GND 0.09fF
C1059 VDD.n428 GND 0.05fF
C1060 VDD.n429 GND 0.02fF
C1061 VDD.n430 GND 0.02fF
C1062 VDD.n431 GND 0.15fF
C1063 VDD.n432 GND 0.02fF
C1064 VDD.n433 GND 0.02fF
C1065 VDD.n434 GND 0.03fF
C1066 VDD.n435 GND 0.16fF
C1067 VDD.n436 GND 0.02fF
C1068 VDD.n437 GND 0.02fF
C1069 VDD.n438 GND 0.03fF
C1070 VDD.n439 GND 0.09fF
C1071 VDD.n440 GND 0.05fF
C1072 VDD.n441 GND 0.17fF
C1073 VDD.n442 GND 0.01fF
C1074 VDD.n443 GND 0.02fF
C1075 VDD.n444 GND 0.02fF
C1076 VDD.n445 GND 0.18fF
C1077 VDD.n446 GND 0.01fF
C1078 VDD.n447 GND 0.02fF
C1079 VDD.n448 GND 0.02fF
C1080 VDD.n449 GND 0.07fF
C1081 VDD.n450 GND 0.24fF
C1082 VDD.n451 GND 0.01fF
C1083 VDD.n452 GND 0.01fF
C1084 VDD.n453 GND 0.02fF
C1085 VDD.n454 GND 0.29fF
C1086 VDD.n455 GND 0.01fF
C1087 VDD.n456 GND 0.02fF
C1088 VDD.n457 GND 0.02fF
C1089 VDD.n458 GND 0.29fF
C1090 VDD.n459 GND 0.01fF
C1091 VDD.n460 GND 0.02fF
C1092 VDD.n461 GND 0.04fF
C1093 VDD.n462 GND 0.33fF
C1094 VDD.n463 GND 0.02fF
C1095 VDD.n464 GND 0.02fF
C1096 VDD.n465 GND 0.02fF
C1097 VDD.n466 GND 0.06fF
C1098 VDD.n467 GND 0.02fF
C1099 VDD.n468 GND 0.02fF
C1100 VDD.n469 GND 0.02fF
C1101 VDD.n470 GND 0.02fF
C1102 VDD.n471 GND 0.02fF
C1103 VDD.n472 GND 0.02fF
C1104 VDD.n473 GND 0.02fF
C1105 VDD.n474 GND 0.02fF
C1106 VDD.n475 GND 0.02fF
C1107 VDD.n476 GND 0.02fF
C1108 VDD.n477 GND 0.03fF
C1109 VDD.n478 GND 0.03fF
C1110 VDD.n479 GND 0.02fF
C1111 VDD.n483 GND 0.29fF
C1112 VDD.n484 GND 0.29fF
C1113 VDD.n485 GND 0.01fF
C1114 VDD.n486 GND 0.02fF
C1115 VDD.n487 GND 0.04fF
C1116 VDD.n488 GND 0.29fF
C1117 VDD.n489 GND 0.01fF
C1118 VDD.n490 GND 0.02fF
C1119 VDD.n491 GND 0.02fF
C1120 VDD.n492 GND 0.24fF
C1121 VDD.n493 GND 0.01fF
C1122 VDD.n494 GND 0.07fF
C1123 VDD.n495 GND 0.02fF
C1124 VDD.n496 GND 0.18fF
C1125 VDD.n497 GND 0.01fF
C1126 VDD.n498 GND 0.02fF
C1127 VDD.n499 GND 0.02fF
C1128 VDD.n500 GND 0.17fF
C1129 VDD.n501 GND 0.01fF
C1130 VDD.n502 GND 0.09fF
C1131 VDD.n503 GND 0.05fF
C1132 VDD.n504 GND 0.02fF
C1133 VDD.n505 GND 0.02fF
C1134 VDD.n506 GND 0.15fF
C1135 VDD.n507 GND 0.02fF
C1136 VDD.n508 GND 0.02fF
C1137 VDD.n509 GND 0.03fF
C1138 VDD.n510 GND 0.16fF
C1139 VDD.n511 GND 0.02fF
C1140 VDD.n512 GND 0.02fF
C1141 VDD.n513 GND 0.03fF
C1142 VDD.n514 GND 0.09fF
C1143 VDD.n515 GND 0.05fF
C1144 VDD.n516 GND 0.17fF
C1145 VDD.n517 GND 0.01fF
C1146 VDD.n518 GND 0.02fF
C1147 VDD.n519 GND 0.02fF
C1148 VDD.n520 GND 0.18fF
C1149 VDD.n521 GND 0.01fF
C1150 VDD.n522 GND 0.02fF
C1151 VDD.n523 GND 0.02fF
C1152 VDD.n524 GND 0.07fF
C1153 VDD.n525 GND 0.24fF
C1154 VDD.n526 GND 0.01fF
C1155 VDD.n527 GND 0.01fF
C1156 VDD.n528 GND 0.02fF
C1157 VDD.n529 GND 0.29fF
C1158 VDD.n530 GND 0.01fF
C1159 VDD.n531 GND 0.02fF
C1160 VDD.n532 GND 0.02fF
C1161 VDD.n533 GND 0.29fF
C1162 VDD.n534 GND 0.01fF
C1163 VDD.n535 GND 0.02fF
C1164 VDD.n536 GND 0.04fF
C1165 VDD.n537 GND 0.33fF
C1166 VDD.n538 GND 0.02fF
C1167 VDD.n539 GND 0.02fF
C1168 VDD.n540 GND 0.02fF
C1169 VDD.n541 GND 0.06fF
C1170 VDD.n542 GND 0.02fF
C1171 VDD.n543 GND 0.02fF
C1172 VDD.n544 GND 0.02fF
C1173 VDD.n545 GND 0.02fF
C1174 VDD.n546 GND 0.02fF
C1175 VDD.n547 GND 0.02fF
C1176 VDD.n548 GND 0.02fF
C1177 VDD.n549 GND 0.02fF
C1178 VDD.n550 GND 0.02fF
C1179 VDD.n551 GND 0.02fF
C1180 VDD.n552 GND 0.03fF
C1181 VDD.n553 GND 0.03fF
C1182 VDD.n554 GND 0.02fF
C1183 VDD.n558 GND 0.29fF
C1184 VDD.n559 GND 0.29fF
C1185 VDD.n560 GND 0.01fF
C1186 VDD.n561 GND 0.02fF
C1187 VDD.n562 GND 0.04fF
C1188 VDD.n563 GND 0.29fF
C1189 VDD.n564 GND 0.01fF
C1190 VDD.n565 GND 0.02fF
C1191 VDD.n566 GND 0.02fF
C1192 VDD.n567 GND 0.24fF
C1193 VDD.n568 GND 0.01fF
C1194 VDD.n569 GND 0.07fF
C1195 VDD.n570 GND 0.02fF
C1196 VDD.n571 GND 0.18fF
C1197 VDD.n572 GND 0.01fF
C1198 VDD.n573 GND 0.02fF
C1199 VDD.n574 GND 0.02fF
C1200 VDD.n575 GND 0.17fF
C1201 VDD.n576 GND 0.01fF
C1202 VDD.n577 GND 0.09fF
C1203 VDD.n578 GND 0.05fF
C1204 VDD.n579 GND 0.02fF
C1205 VDD.n580 GND 0.02fF
C1206 VDD.n581 GND 0.15fF
C1207 VDD.n582 GND 0.02fF
C1208 VDD.n583 GND 0.02fF
C1209 VDD.n584 GND 0.03fF
C1210 VDD.n585 GND 0.16fF
C1211 VDD.n586 GND 0.02fF
C1212 VDD.n587 GND 0.02fF
C1213 VDD.n588 GND 0.03fF
C1214 VDD.n589 GND 0.09fF
C1215 VDD.n590 GND 0.05fF
C1216 VDD.n591 GND 0.17fF
C1217 VDD.n592 GND 0.01fF
C1218 VDD.n593 GND 0.02fF
C1219 VDD.n594 GND 0.02fF
C1220 VDD.n595 GND 0.18fF
C1221 VDD.n596 GND 0.01fF
C1222 VDD.n597 GND 0.02fF
C1223 VDD.n598 GND 0.02fF
C1224 VDD.n599 GND 0.07fF
C1225 VDD.n600 GND 0.24fF
C1226 VDD.n601 GND 0.01fF
C1227 VDD.n602 GND 0.01fF
C1228 VDD.n603 GND 0.02fF
C1229 VDD.n604 GND 0.29fF
C1230 VDD.n605 GND 0.01fF
C1231 VDD.n606 GND 0.02fF
C1232 VDD.n607 GND 0.02fF
C1233 VDD.n608 GND 0.29fF
C1234 VDD.n609 GND 0.01fF
C1235 VDD.n610 GND 0.02fF
C1236 VDD.n611 GND 0.04fF
C1237 VDD.n612 GND 0.33fF
C1238 VDD.n613 GND 0.02fF
C1239 VDD.n614 GND 0.02fF
C1240 VDD.n615 GND 0.02fF
C1241 VDD.n616 GND 0.06fF
C1242 VDD.n617 GND 0.02fF
C1243 VDD.n618 GND 0.02fF
C1244 VDD.n619 GND 0.02fF
C1245 VDD.n620 GND 0.02fF
C1246 VDD.n621 GND 0.02fF
C1247 VDD.n622 GND 0.02fF
C1248 VDD.n623 GND 0.02fF
C1249 VDD.n624 GND 0.02fF
C1250 VDD.n625 GND 0.02fF
C1251 VDD.n626 GND 0.02fF
C1252 VDD.n627 GND 0.03fF
C1253 VDD.n628 GND 0.03fF
C1254 VDD.n629 GND 0.02fF
C1255 VDD.n633 GND 0.29fF
C1256 VDD.n634 GND 0.29fF
C1257 VDD.n635 GND 0.01fF
C1258 VDD.n636 GND 0.02fF
C1259 VDD.n637 GND 0.04fF
C1260 VDD.n638 GND 0.29fF
C1261 VDD.n639 GND 0.01fF
C1262 VDD.n640 GND 0.02fF
C1263 VDD.n641 GND 0.02fF
C1264 VDD.n642 GND 0.24fF
C1265 VDD.n643 GND 0.01fF
C1266 VDD.n644 GND 0.07fF
C1267 VDD.n645 GND 0.02fF
C1268 VDD.n646 GND 0.18fF
C1269 VDD.n647 GND 0.01fF
C1270 VDD.n648 GND 0.02fF
C1271 VDD.n649 GND 0.02fF
C1272 VDD.n650 GND 0.17fF
C1273 VDD.n651 GND 0.01fF
C1274 VDD.n652 GND 0.09fF
C1275 VDD.n653 GND 0.05fF
C1276 VDD.n654 GND 0.02fF
C1277 VDD.n655 GND 0.02fF
C1278 VDD.n656 GND 0.15fF
C1279 VDD.n657 GND 0.02fF
C1280 VDD.n658 GND 0.02fF
C1281 VDD.n659 GND 0.03fF
C1282 VDD.n660 GND 0.16fF
C1283 VDD.n661 GND 0.02fF
C1284 VDD.n662 GND 0.02fF
C1285 VDD.n663 GND 0.03fF
C1286 VDD.n664 GND 0.09fF
C1287 VDD.n665 GND 0.05fF
C1288 VDD.n666 GND 0.17fF
C1289 VDD.n667 GND 0.01fF
C1290 VDD.n668 GND 0.02fF
C1291 VDD.n669 GND 0.02fF
C1292 VDD.n670 GND 0.18fF
C1293 VDD.n671 GND 0.01fF
C1294 VDD.n672 GND 0.02fF
C1295 VDD.n673 GND 0.02fF
C1296 VDD.n674 GND 0.07fF
C1297 VDD.n675 GND 0.24fF
C1298 VDD.n676 GND 0.01fF
C1299 VDD.n677 GND 0.01fF
C1300 VDD.n678 GND 0.02fF
C1301 VDD.n679 GND 0.29fF
C1302 VDD.n680 GND 0.01fF
C1303 VDD.n681 GND 0.02fF
C1304 VDD.n682 GND 0.02fF
C1305 VDD.n683 GND 0.29fF
C1306 VDD.n684 GND 0.01fF
C1307 VDD.n685 GND 0.02fF
C1308 VDD.n686 GND 0.04fF
C1309 VDD.n687 GND 0.33fF
C1310 VDD.n688 GND 0.02fF
C1311 VDD.n689 GND 0.02fF
C1312 VDD.n690 GND 0.02fF
C1313 VDD.n691 GND 0.06fF
C1314 VDD.n692 GND 0.02fF
C1315 VDD.n693 GND 0.02fF
C1316 VDD.n694 GND 0.02fF
C1317 VDD.n695 GND 0.02fF
C1318 VDD.n696 GND 0.02fF
C1319 VDD.n697 GND 0.02fF
C1320 VDD.n698 GND 0.02fF
C1321 VDD.n699 GND 0.02fF
C1322 VDD.n700 GND 0.02fF
C1323 VDD.n701 GND 0.02fF
C1324 VDD.n702 GND 0.03fF
C1325 VDD.n703 GND 0.03fF
C1326 VDD.n704 GND 0.02fF
C1327 VDD.n708 GND 0.29fF
C1328 VDD.n709 GND 0.29fF
C1329 VDD.n710 GND 0.01fF
C1330 VDD.n711 GND 0.02fF
C1331 VDD.n712 GND 0.04fF
C1332 VDD.n713 GND 0.29fF
C1333 VDD.n714 GND 0.01fF
C1334 VDD.n715 GND 0.02fF
C1335 VDD.n716 GND 0.02fF
C1336 VDD.n717 GND 0.24fF
C1337 VDD.n718 GND 0.01fF
C1338 VDD.n719 GND 0.07fF
C1339 VDD.n720 GND 0.02fF
C1340 VDD.n721 GND 0.18fF
C1341 VDD.n722 GND 0.01fF
C1342 VDD.n723 GND 0.02fF
C1343 VDD.n724 GND 0.02fF
C1344 VDD.n725 GND 0.17fF
C1345 VDD.n726 GND 0.01fF
C1346 VDD.n727 GND 0.09fF
C1347 VDD.n728 GND 0.05fF
C1348 VDD.n729 GND 0.02fF
C1349 VDD.n730 GND 0.02fF
C1350 VDD.n731 GND 0.15fF
C1351 VDD.n732 GND 0.02fF
C1352 VDD.n733 GND 0.02fF
C1353 VDD.n734 GND 0.03fF
C1354 VDD.n735 GND 0.16fF
C1355 VDD.n736 GND 0.02fF
C1356 VDD.n737 GND 0.02fF
C1357 VDD.n738 GND 0.03fF
C1358 VDD.n739 GND 0.09fF
C1359 VDD.n740 GND 0.05fF
C1360 VDD.n741 GND 0.17fF
C1361 VDD.n742 GND 0.01fF
C1362 VDD.n743 GND 0.02fF
C1363 VDD.n744 GND 0.02fF
C1364 VDD.n745 GND 0.18fF
C1365 VDD.n746 GND 0.01fF
C1366 VDD.n747 GND 0.02fF
C1367 VDD.n748 GND 0.02fF
C1368 VDD.n749 GND 0.07fF
C1369 VDD.n750 GND 0.24fF
C1370 VDD.n751 GND 0.01fF
C1371 VDD.n752 GND 0.01fF
C1372 VDD.n753 GND 0.02fF
C1373 VDD.n754 GND 0.29fF
C1374 VDD.n755 GND 0.01fF
C1375 VDD.n756 GND 0.02fF
C1376 VDD.n757 GND 0.02fF
C1377 VDD.n758 GND 0.33fF
C1378 VDD.n759 GND 0.02fF
C1379 VDD.n760 GND 0.02fF
C1380 VDD.n761 GND 0.02fF
C1381 VDD.n762 GND 0.06fF
C1382 VDD.n763 GND 0.02fF
C1383 VDD.n764 GND 0.02fF
C1384 VDD.n765 GND 0.02fF
C1385 VDD.n766 GND 0.02fF
C1386 VDD.n767 GND 0.02fF
C1387 VDD.n768 GND 0.02fF
C1388 VDD.n769 GND 0.02fF
C1389 VDD.n770 GND 0.02fF
C1390 VDD.n771 GND 0.02fF
C1391 VDD.n772 GND 0.02fF
C1392 VDD.n773 GND 0.03fF
C1393 VDD.n774 GND 0.03fF
C1394 VDD.n775 GND 0.02fF
C1395 VDD.n779 GND 0.29fF
C1396 VDD.n780 GND 0.29fF
C1397 VDD.n781 GND 0.01fF
C1398 VDD.n782 GND 0.02fF
C1399 VDD.n783 GND 0.02fF
C1400 VDD.n784 GND 0.19fF
C1401 VDD.n785 GND 0.02fF
C1402 VDD.n786 GND 0.02fF
C1403 VDD.n787 GND 0.06fF
C1404 VDD.n788 GND 0.02fF
C1405 VDD.n789 GND 0.02fF
C1406 VDD.n790 GND 0.02fF
C1407 VDD.n791 GND 0.02fF
C1408 VDD.n792 GND 0.02fF
C1409 VDD.n793 GND 0.02fF
C1410 VDD.n794 GND 0.02fF
C1411 VDD.n795 GND 0.02fF
C1412 VDD.n796 GND 0.04fF
C1413 VDD.n797 GND 0.04fF
C1414 VDD.n798 GND 0.02fF
C1415 VDD.n802 GND 0.49fF
C1416 VDD.n803 GND 0.29fF
C1417 VDD.n804 GND 0.02fF
C1418 VDD.n805 GND 0.03fF
C1419 VDD.n806 GND 0.03fF
C1420 VDD.n807 GND 0.29fF
C1421 VDD.n808 GND 0.01fF
C1422 VDD.n809 GND 0.02fF
C1423 VDD.n810 GND 0.02fF
C1424 VDD.n811 GND 0.07fF
C1425 VDD.n812 GND 0.24fF
C1426 VDD.n813 GND 0.01fF
C1427 VDD.n814 GND 0.01fF
C1428 VDD.n815 GND 0.02fF
C1429 VDD.n816 GND 0.18fF
C1430 VDD.n817 GND 0.01fF
C1431 VDD.n818 GND 0.02fF
C1432 VDD.n819 GND 0.02fF
C1433 VDD.n820 GND 0.09fF
C1434 VDD.n821 GND 0.05fF
C1435 VDD.n822 GND 0.17fF
C1436 VDD.n823 GND 0.01fF
C1437 VDD.n824 GND 0.02fF
C1438 VDD.n825 GND 0.02fF
C1439 VDD.n826 GND 0.16fF
C1440 VDD.n827 GND 0.02fF
C1441 VDD.n828 GND 0.02fF
C1442 VDD.n829 GND 0.03fF
C1443 VDD.n830 GND 0.15fF
C1444 VDD.n831 GND 0.02fF
C1445 VDD.n832 GND 0.02fF
C1446 VDD.n833 GND 0.03fF
C1447 VDD.n834 GND 0.17fF
C1448 VDD.n835 GND 0.01fF
C1449 VDD.n836 GND 0.09fF
C1450 VDD.n837 GND 0.05fF
C1451 VDD.n838 GND 0.02fF
C1452 VDD.n839 GND 0.02fF
C1453 VDD.n840 GND 0.18fF
C1454 VDD.n841 GND 0.01fF
C1455 VDD.n842 GND 0.02fF
C1456 VDD.n843 GND 0.02fF
C1457 VDD.n844 GND 0.24fF
C1458 VDD.n845 GND 0.01fF
C1459 VDD.n846 GND 0.07fF
C1460 VDD.n847 GND 0.02fF
C1461 VDD.n848 GND 0.29fF
C1462 VDD.n849 GND 0.01fF
C1463 VDD.n850 GND 0.02fF
C1464 VDD.n851 GND 0.02fF
C1465 VDD.n852 GND 0.29fF
C1466 VDD.n853 GND 0.01fF
C1467 VDD.n854 GND 0.02fF
C1468 VDD.n855 GND 0.04fF
C1469 VDD.n856 GND 0.06fF
C1470 VDD.n857 GND 0.02fF
C1471 VDD.n858 GND 0.02fF
C1472 VDD.n859 GND 0.02fF
C1473 VDD.n860 GND 0.02fF
C1474 VDD.n861 GND 0.02fF
C1475 VDD.n862 GND 0.02fF
C1476 VDD.n863 GND 0.02fF
C1477 VDD.n864 GND 0.02fF
C1478 VDD.n865 GND 0.02fF
C1479 VDD.n866 GND 0.02fF
C1480 VDD.n867 GND 0.02fF
C1481 VDD.n868 GND 0.03fF
C1482 VDD.n869 GND 0.03fF
C1483 VDD.n872 GND 0.02fF
C1484 VDD.n874 GND 0.02fF
C1485 VDD.n875 GND 0.33fF
C1486 VDD.n876 GND 0.02fF
C1487 VDD.n878 GND 0.29fF
C1488 VDD.n879 GND 0.29fF
C1489 VDD.n880 GND 0.01fF
C1490 VDD.n881 GND 0.02fF
C1491 VDD.n882 GND 0.04fF
C1492 VDD.n883 GND 0.29fF
C1493 VDD.n884 GND 0.01fF
C1494 VDD.n885 GND 0.02fF
C1495 VDD.n886 GND 0.02fF
C1496 VDD.n887 GND 0.07fF
C1497 VDD.n888 GND 0.24fF
C1498 VDD.n889 GND 0.01fF
C1499 VDD.n890 GND 0.01fF
C1500 VDD.n891 GND 0.02fF
C1501 VDD.n892 GND 0.18fF
C1502 VDD.n893 GND 0.01fF
C1503 VDD.n894 GND 0.02fF
C1504 VDD.n895 GND 0.02fF
C1505 VDD.n896 GND 0.09fF
C1506 VDD.n897 GND 0.05fF
C1507 VDD.n898 GND 0.17fF
C1508 VDD.n899 GND 0.01fF
C1509 VDD.n900 GND 0.02fF
C1510 VDD.n901 GND 0.02fF
C1511 VDD.n902 GND 0.16fF
C1512 VDD.n903 GND 0.02fF
C1513 VDD.n904 GND 0.02fF
C1514 VDD.n905 GND 0.03fF
C1515 VDD.n906 GND 0.15fF
C1516 VDD.n907 GND 0.02fF
C1517 VDD.n908 GND 0.02fF
C1518 VDD.n909 GND 0.03fF
C1519 VDD.n910 GND 0.17fF
C1520 VDD.n911 GND 0.01fF
C1521 VDD.n912 GND 0.09fF
C1522 VDD.n913 GND 0.05fF
C1523 VDD.n914 GND 0.02fF
C1524 VDD.n915 GND 0.02fF
C1525 VDD.n916 GND 0.18fF
C1526 VDD.n917 GND 0.01fF
C1527 VDD.n918 GND 0.02fF
C1528 VDD.n919 GND 0.02fF
C1529 VDD.n920 GND 0.24fF
C1530 VDD.n921 GND 0.01fF
C1531 VDD.n922 GND 0.07fF
C1532 VDD.n923 GND 0.02fF
C1533 VDD.n924 GND 0.29fF
C1534 VDD.n925 GND 0.01fF
C1535 VDD.n926 GND 0.02fF
C1536 VDD.n927 GND 0.02fF
C1537 VDD.n928 GND 0.29fF
C1538 VDD.n929 GND 0.01fF
C1539 VDD.n930 GND 0.02fF
C1540 VDD.n931 GND 0.04fF
C1541 VDD.n932 GND 0.33fF
C1542 VDD.n933 GND 0.02fF
C1543 VDD.n934 GND 0.02fF
C1544 VDD.n935 GND 0.02fF
C1545 VDD.n936 GND 0.06fF
C1546 VDD.n937 GND 0.02fF
C1547 VDD.n938 GND 0.02fF
C1548 VDD.n939 GND 0.02fF
C1549 VDD.n940 GND 0.02fF
C1550 VDD.n941 GND 0.02fF
C1551 VDD.n942 GND 0.02fF
C1552 VDD.n943 GND 0.02fF
C1553 VDD.n944 GND 0.02fF
C1554 VDD.n945 GND 0.02fF
C1555 VDD.n946 GND 0.02fF
C1556 VDD.n947 GND 0.03fF
C1557 VDD.n948 GND 0.03fF
C1558 VDD.n949 GND 0.02fF
C1559 VDD.n953 GND 0.29fF
C1560 VDD.n954 GND 0.29fF
C1561 VDD.n955 GND 0.01fF
C1562 VDD.n956 GND 0.02fF
C1563 VDD.n957 GND 0.04fF
C1564 VDD.n958 GND 0.29fF
C1565 VDD.n959 GND 0.01fF
C1566 VDD.n960 GND 0.02fF
C1567 VDD.n961 GND 0.02fF
C1568 VDD.n962 GND 0.07fF
C1569 VDD.n963 GND 0.24fF
C1570 VDD.n964 GND 0.01fF
C1571 VDD.n965 GND 0.01fF
C1572 VDD.n966 GND 0.02fF
C1573 VDD.n967 GND 0.18fF
C1574 VDD.n968 GND 0.01fF
C1575 VDD.n969 GND 0.02fF
C1576 VDD.n970 GND 0.02fF
C1577 VDD.n971 GND 0.09fF
C1578 VDD.n972 GND 0.05fF
C1579 VDD.n973 GND 0.17fF
C1580 VDD.n974 GND 0.01fF
C1581 VDD.n975 GND 0.02fF
C1582 VDD.n976 GND 0.02fF
C1583 VDD.n977 GND 0.16fF
C1584 VDD.n978 GND 0.02fF
C1585 VDD.n979 GND 0.02fF
C1586 VDD.n980 GND 0.03fF
C1587 VDD.n981 GND 0.15fF
C1588 VDD.n982 GND 0.02fF
C1589 VDD.n983 GND 0.02fF
C1590 VDD.n984 GND 0.03fF
C1591 VDD.n985 GND 0.17fF
C1592 VDD.n986 GND 0.01fF
C1593 VDD.n987 GND 0.09fF
C1594 VDD.n988 GND 0.05fF
C1595 VDD.n989 GND 0.02fF
C1596 VDD.n990 GND 0.02fF
C1597 VDD.n991 GND 0.18fF
C1598 VDD.n992 GND 0.01fF
C1599 VDD.n993 GND 0.02fF
C1600 VDD.n994 GND 0.02fF
C1601 VDD.n995 GND 0.24fF
C1602 VDD.n996 GND 0.01fF
C1603 VDD.n997 GND 0.07fF
C1604 VDD.n998 GND 0.02fF
C1605 VDD.n999 GND 0.29fF
C1606 VDD.n1000 GND 0.01fF
C1607 VDD.n1001 GND 0.02fF
C1608 VDD.n1002 GND 0.02fF
C1609 VDD.n1003 GND 0.29fF
C1610 VDD.n1004 GND 0.01fF
C1611 VDD.n1005 GND 0.02fF
C1612 VDD.n1006 GND 0.04fF
C1613 VDD.n1007 GND 0.33fF
C1614 VDD.n1008 GND 0.02fF
C1615 VDD.n1009 GND 0.02fF
C1616 VDD.n1010 GND 0.02fF
C1617 VDD.n1011 GND 0.06fF
C1618 VDD.n1012 GND 0.02fF
C1619 VDD.n1013 GND 0.02fF
C1620 VDD.n1014 GND 0.02fF
C1621 VDD.n1015 GND 0.02fF
C1622 VDD.n1016 GND 0.02fF
C1623 VDD.n1017 GND 0.02fF
C1624 VDD.n1018 GND 0.02fF
C1625 VDD.n1019 GND 0.02fF
C1626 VDD.n1020 GND 0.02fF
C1627 VDD.n1021 GND 0.02fF
C1628 VDD.n1022 GND 0.03fF
C1629 VDD.n1023 GND 0.03fF
C1630 VDD.n1024 GND 0.02fF
C1631 VDD.n1028 GND 0.29fF
C1632 VDD.n1029 GND 0.29fF
C1633 VDD.n1030 GND 0.01fF
C1634 VDD.n1031 GND 0.02fF
C1635 VDD.n1032 GND 0.04fF
C1636 VDD.n1033 GND 0.29fF
C1637 VDD.n1034 GND 0.01fF
C1638 VDD.n1035 GND 0.02fF
C1639 VDD.n1036 GND 0.02fF
C1640 VDD.n1037 GND 0.07fF
C1641 VDD.n1038 GND 0.24fF
C1642 VDD.n1039 GND 0.01fF
C1643 VDD.n1040 GND 0.01fF
C1644 VDD.n1041 GND 0.02fF
C1645 VDD.n1042 GND 0.18fF
C1646 VDD.n1043 GND 0.01fF
C1647 VDD.n1044 GND 0.02fF
C1648 VDD.n1045 GND 0.02fF
C1649 VDD.n1046 GND 0.09fF
C1650 VDD.n1047 GND 0.05fF
C1651 VDD.n1048 GND 0.17fF
C1652 VDD.n1049 GND 0.01fF
C1653 VDD.n1050 GND 0.02fF
C1654 VDD.n1051 GND 0.02fF
C1655 VDD.n1052 GND 0.16fF
C1656 VDD.n1053 GND 0.02fF
C1657 VDD.n1054 GND 0.02fF
C1658 VDD.n1055 GND 0.03fF
C1659 VDD.n1056 GND 0.15fF
C1660 VDD.n1057 GND 0.02fF
C1661 VDD.n1058 GND 0.02fF
C1662 VDD.n1059 GND 0.03fF
C1663 VDD.n1060 GND 0.17fF
C1664 VDD.n1061 GND 0.01fF
C1665 VDD.n1062 GND 0.09fF
C1666 VDD.n1063 GND 0.05fF
C1667 VDD.n1064 GND 0.02fF
C1668 VDD.n1065 GND 0.02fF
C1669 VDD.n1066 GND 0.18fF
C1670 VDD.n1067 GND 0.01fF
C1671 VDD.n1068 GND 0.02fF
C1672 VDD.n1069 GND 0.02fF
C1673 VDD.n1070 GND 0.24fF
C1674 VDD.n1071 GND 0.01fF
C1675 VDD.n1072 GND 0.07fF
C1676 VDD.n1073 GND 0.02fF
C1677 VDD.n1074 GND 0.29fF
C1678 VDD.n1075 GND 0.01fF
C1679 VDD.n1076 GND 0.02fF
C1680 VDD.n1077 GND 0.02fF
C1681 VDD.n1078 GND 0.29fF
C1682 VDD.n1079 GND 0.01fF
C1683 VDD.n1080 GND 0.02fF
C1684 VDD.n1081 GND 0.04fF
C1685 VDD.n1082 GND 0.33fF
C1686 VDD.n1083 GND 0.02fF
C1687 VDD.n1084 GND 0.02fF
C1688 VDD.n1085 GND 0.02fF
C1689 VDD.n1086 GND 0.06fF
C1690 VDD.n1087 GND 0.02fF
C1691 VDD.n1088 GND 0.02fF
C1692 VDD.n1089 GND 0.02fF
C1693 VDD.n1090 GND 0.02fF
C1694 VDD.n1091 GND 0.02fF
C1695 VDD.n1092 GND 0.02fF
C1696 VDD.n1093 GND 0.02fF
C1697 VDD.n1094 GND 0.02fF
C1698 VDD.n1095 GND 0.02fF
C1699 VDD.n1096 GND 0.02fF
C1700 VDD.n1097 GND 0.03fF
C1701 VDD.n1098 GND 0.03fF
C1702 VDD.n1099 GND 0.02fF
C1703 VDD.n1103 GND 0.29fF
C1704 VDD.n1104 GND 0.29fF
C1705 VDD.n1105 GND 0.01fF
C1706 VDD.n1106 GND 0.02fF
C1707 VDD.n1107 GND 0.04fF
C1708 VDD.n1108 GND 0.29fF
C1709 VDD.n1109 GND 0.01fF
C1710 VDD.n1110 GND 0.02fF
C1711 VDD.n1111 GND 0.02fF
C1712 VDD.n1112 GND 0.07fF
C1713 VDD.n1113 GND 0.24fF
C1714 VDD.n1114 GND 0.01fF
C1715 VDD.n1115 GND 0.01fF
C1716 VDD.n1116 GND 0.02fF
C1717 VDD.n1117 GND 0.18fF
C1718 VDD.n1118 GND 0.01fF
C1719 VDD.n1119 GND 0.02fF
C1720 VDD.n1120 GND 0.02fF
C1721 VDD.n1121 GND 0.09fF
C1722 VDD.n1122 GND 0.05fF
C1723 VDD.n1123 GND 0.17fF
C1724 VDD.n1124 GND 0.01fF
C1725 VDD.n1125 GND 0.02fF
C1726 VDD.n1126 GND 0.02fF
C1727 VDD.n1127 GND 0.16fF
C1728 VDD.n1128 GND 0.02fF
C1729 VDD.n1129 GND 0.02fF
C1730 VDD.n1130 GND 0.03fF
C1731 VDD.n1131 GND 0.15fF
C1732 VDD.n1132 GND 0.02fF
C1733 VDD.n1133 GND 0.02fF
C1734 VDD.n1134 GND 0.03fF
C1735 VDD.n1135 GND 0.17fF
C1736 VDD.n1136 GND 0.01fF
C1737 VDD.n1137 GND 0.09fF
C1738 VDD.n1138 GND 0.05fF
C1739 VDD.n1139 GND 0.02fF
C1740 VDD.n1140 GND 0.02fF
C1741 VDD.n1141 GND 0.18fF
C1742 VDD.n1142 GND 0.01fF
C1743 VDD.n1143 GND 0.02fF
C1744 VDD.n1144 GND 0.02fF
C1745 VDD.n1145 GND 0.24fF
C1746 VDD.n1146 GND 0.01fF
C1747 VDD.n1147 GND 0.07fF
C1748 VDD.n1148 GND 0.02fF
C1749 VDD.n1149 GND 0.29fF
C1750 VDD.n1150 GND 0.01fF
C1751 VDD.n1151 GND 0.02fF
C1752 VDD.n1152 GND 0.02fF
C1753 VDD.n1153 GND 0.29fF
C1754 VDD.n1154 GND 0.01fF
C1755 VDD.n1155 GND 0.02fF
C1756 VDD.n1156 GND 0.04fF
C1757 VDD.n1157 GND 0.33fF
C1758 VDD.n1158 GND 0.02fF
C1759 VDD.n1159 GND 0.02fF
C1760 VDD.n1160 GND 0.02fF
C1761 VDD.n1161 GND 0.06fF
C1762 VDD.n1162 GND 0.02fF
C1763 VDD.n1163 GND 0.02fF
C1764 VDD.n1164 GND 0.02fF
C1765 VDD.n1165 GND 0.02fF
C1766 VDD.n1166 GND 0.02fF
C1767 VDD.n1167 GND 0.02fF
C1768 VDD.n1168 GND 0.02fF
C1769 VDD.n1169 GND 0.02fF
C1770 VDD.n1170 GND 0.02fF
C1771 VDD.n1171 GND 0.02fF
C1772 VDD.n1172 GND 0.03fF
C1773 VDD.n1173 GND 0.03fF
C1774 VDD.n1174 GND 0.02fF
C1775 VDD.n1178 GND 0.29fF
C1776 VDD.n1179 GND 0.29fF
C1777 VDD.n1180 GND 0.01fF
C1778 VDD.n1181 GND 0.02fF
C1779 VDD.n1182 GND 0.04fF
C1780 VDD.n1183 GND 0.29fF
C1781 VDD.n1184 GND 0.01fF
C1782 VDD.n1185 GND 0.02fF
C1783 VDD.n1186 GND 0.02fF
C1784 VDD.n1187 GND 0.07fF
C1785 VDD.n1188 GND 0.24fF
C1786 VDD.n1189 GND 0.01fF
C1787 VDD.n1190 GND 0.01fF
C1788 VDD.n1191 GND 0.02fF
C1789 VDD.n1192 GND 0.18fF
C1790 VDD.n1193 GND 0.01fF
C1791 VDD.n1194 GND 0.02fF
C1792 VDD.n1195 GND 0.02fF
C1793 VDD.n1196 GND 0.09fF
C1794 VDD.n1197 GND 0.05fF
C1795 VDD.n1198 GND 0.17fF
C1796 VDD.n1199 GND 0.01fF
C1797 VDD.n1200 GND 0.02fF
C1798 VDD.n1201 GND 0.02fF
C1799 VDD.n1202 GND 0.16fF
C1800 VDD.n1203 GND 0.02fF
C1801 VDD.n1204 GND 0.02fF
C1802 VDD.n1205 GND 0.03fF
C1803 VDD.n1206 GND 0.15fF
C1804 VDD.n1207 GND 0.02fF
C1805 VDD.n1208 GND 0.02fF
C1806 VDD.n1209 GND 0.03fF
C1807 VDD.n1210 GND 0.17fF
C1808 VDD.n1211 GND 0.01fF
C1809 VDD.n1212 GND 0.09fF
C1810 VDD.n1213 GND 0.05fF
C1811 VDD.n1214 GND 0.02fF
C1812 VDD.n1215 GND 0.02fF
C1813 VDD.n1216 GND 0.18fF
C1814 VDD.n1217 GND 0.01fF
C1815 VDD.n1218 GND 0.02fF
C1816 VDD.n1219 GND 0.02fF
C1817 VDD.n1220 GND 0.24fF
C1818 VDD.n1221 GND 0.01fF
C1819 VDD.n1222 GND 0.07fF
C1820 VDD.n1223 GND 0.02fF
C1821 VDD.n1224 GND 0.29fF
C1822 VDD.n1225 GND 0.01fF
C1823 VDD.n1226 GND 0.02fF
C1824 VDD.n1227 GND 0.02fF
C1825 VDD.n1228 GND 0.29fF
C1826 VDD.n1229 GND 0.01fF
C1827 VDD.n1230 GND 0.02fF
C1828 VDD.n1231 GND 0.04fF
C1829 VDD.n1232 GND 0.33fF
C1830 VDD.n1233 GND 0.02fF
C1831 VDD.n1234 GND 0.02fF
C1832 VDD.n1235 GND 0.02fF
C1833 VDD.n1236 GND 0.06fF
C1834 VDD.n1237 GND 0.02fF
C1835 VDD.n1238 GND 0.02fF
C1836 VDD.n1239 GND 0.02fF
C1837 VDD.n1240 GND 0.02fF
C1838 VDD.n1241 GND 0.02fF
C1839 VDD.n1242 GND 0.02fF
C1840 VDD.n1243 GND 0.02fF
C1841 VDD.n1244 GND 0.02fF
C1842 VDD.n1245 GND 0.02fF
C1843 VDD.n1246 GND 0.02fF
C1844 VDD.n1247 GND 0.03fF
C1845 VDD.n1248 GND 0.03fF
C1846 VDD.n1249 GND 0.02fF
C1847 VDD.n1253 GND 0.29fF
C1848 VDD.n1254 GND 0.29fF
C1849 VDD.n1255 GND 0.01fF
C1850 VDD.n1256 GND 0.02fF
C1851 VDD.n1257 GND 0.04fF
C1852 VDD.n1258 GND 0.29fF
C1853 VDD.n1259 GND 0.01fF
C1854 VDD.n1260 GND 0.02fF
C1855 VDD.n1261 GND 0.02fF
C1856 VDD.n1262 GND 0.07fF
C1857 VDD.n1263 GND 0.24fF
C1858 VDD.n1264 GND 0.01fF
C1859 VDD.n1265 GND 0.01fF
C1860 VDD.n1266 GND 0.02fF
C1861 VDD.n1267 GND 0.18fF
C1862 VDD.n1268 GND 0.01fF
C1863 VDD.n1269 GND 0.02fF
C1864 VDD.n1270 GND 0.02fF
C1865 VDD.n1271 GND 0.09fF
C1866 VDD.n1272 GND 0.05fF
C1867 VDD.n1273 GND 0.17fF
C1868 VDD.n1274 GND 0.01fF
C1869 VDD.n1275 GND 0.02fF
C1870 VDD.n1276 GND 0.02fF
C1871 VDD.n1277 GND 0.16fF
C1872 VDD.n1278 GND 0.02fF
C1873 VDD.n1279 GND 0.02fF
C1874 VDD.n1280 GND 0.03fF
C1875 VDD.n1281 GND 0.15fF
C1876 VDD.n1282 GND 0.02fF
C1877 VDD.n1283 GND 0.02fF
C1878 VDD.n1284 GND 0.03fF
C1879 VDD.n1285 GND 0.17fF
C1880 VDD.n1286 GND 0.01fF
C1881 VDD.n1287 GND 0.09fF
C1882 VDD.n1288 GND 0.05fF
C1883 VDD.n1289 GND 0.02fF
C1884 VDD.n1290 GND 0.02fF
C1885 VDD.n1291 GND 0.18fF
C1886 VDD.n1292 GND 0.01fF
C1887 VDD.n1293 GND 0.02fF
C1888 VDD.n1294 GND 0.02fF
C1889 VDD.n1295 GND 0.24fF
C1890 VDD.n1296 GND 0.01fF
C1891 VDD.n1297 GND 0.07fF
C1892 VDD.n1298 GND 0.02fF
C1893 VDD.n1299 GND 0.29fF
C1894 VDD.n1300 GND 0.01fF
C1895 VDD.n1301 GND 0.02fF
C1896 VDD.n1302 GND 0.02fF
C1897 VDD.n1303 GND 0.29fF
C1898 VDD.n1304 GND 0.01fF
C1899 VDD.n1305 GND 0.02fF
C1900 VDD.n1306 GND 0.04fF
C1901 VDD.n1307 GND 0.33fF
C1902 VDD.n1308 GND 0.02fF
C1903 VDD.n1309 GND 0.02fF
C1904 VDD.n1310 GND 0.02fF
C1905 VDD.n1311 GND 0.06fF
C1906 VDD.n1312 GND 0.02fF
C1907 VDD.n1313 GND 0.02fF
C1908 VDD.n1314 GND 0.02fF
C1909 VDD.n1315 GND 0.02fF
C1910 VDD.n1316 GND 0.02fF
C1911 VDD.n1317 GND 0.02fF
C1912 VDD.n1318 GND 0.02fF
C1913 VDD.n1319 GND 0.02fF
C1914 VDD.n1320 GND 0.02fF
C1915 VDD.n1321 GND 0.02fF
C1916 VDD.n1322 GND 0.03fF
C1917 VDD.n1323 GND 0.03fF
C1918 VDD.n1324 GND 0.02fF
C1919 VDD.n1328 GND 0.29fF
C1920 VDD.n1329 GND 0.29fF
C1921 VDD.n1330 GND 0.01fF
C1922 VDD.n1331 GND 0.02fF
C1923 VDD.n1332 GND 0.04fF
C1924 VDD.n1333 GND 0.29fF
C1925 VDD.n1334 GND 0.01fF
C1926 VDD.n1335 GND 0.02fF
C1927 VDD.n1336 GND 0.02fF
C1928 VDD.n1337 GND 0.07fF
C1929 VDD.n1338 GND 0.24fF
C1930 VDD.n1339 GND 0.01fF
C1931 VDD.n1340 GND 0.01fF
C1932 VDD.n1341 GND 0.02fF
C1933 VDD.n1342 GND 0.18fF
C1934 VDD.n1343 GND 0.01fF
C1935 VDD.n1344 GND 0.02fF
C1936 VDD.n1345 GND 0.02fF
C1937 VDD.n1346 GND 0.09fF
C1938 VDD.n1347 GND 0.05fF
C1939 VDD.n1348 GND 0.17fF
C1940 VDD.n1349 GND 0.01fF
C1941 VDD.n1350 GND 0.02fF
C1942 VDD.n1351 GND 0.02fF
C1943 VDD.n1352 GND 0.16fF
C1944 VDD.n1353 GND 0.02fF
C1945 VDD.n1354 GND 0.02fF
C1946 VDD.n1355 GND 0.03fF
C1947 VDD.n1356 GND 0.15fF
C1948 VDD.n1357 GND 0.02fF
C1949 VDD.n1358 GND 0.02fF
C1950 VDD.n1359 GND 0.03fF
C1951 VDD.n1360 GND 0.17fF
C1952 VDD.n1361 GND 0.01fF
C1953 VDD.n1362 GND 0.09fF
C1954 VDD.n1363 GND 0.05fF
C1955 VDD.n1364 GND 0.02fF
C1956 VDD.n1365 GND 0.02fF
C1957 VDD.n1366 GND 0.18fF
C1958 VDD.n1367 GND 0.01fF
C1959 VDD.n1368 GND 0.02fF
C1960 VDD.n1369 GND 0.02fF
C1961 VDD.n1370 GND 0.24fF
C1962 VDD.n1371 GND 0.01fF
C1963 VDD.n1372 GND 0.07fF
C1964 VDD.n1373 GND 0.02fF
C1965 VDD.n1374 GND 0.29fF
C1966 VDD.n1375 GND 0.01fF
C1967 VDD.n1376 GND 0.02fF
C1968 VDD.n1377 GND 0.02fF
C1969 VDD.n1378 GND 0.29fF
C1970 VDD.n1379 GND 0.01fF
C1971 VDD.n1380 GND 0.02fF
C1972 VDD.n1381 GND 0.04fF
C1973 VDD.n1382 GND 0.33fF
C1974 VDD.n1383 GND 0.02fF
C1975 VDD.n1384 GND 0.02fF
C1976 VDD.n1385 GND 0.02fF
C1977 VDD.n1386 GND 0.06fF
C1978 VDD.n1387 GND 0.02fF
C1979 VDD.n1388 GND 0.02fF
C1980 VDD.n1389 GND 0.02fF
C1981 VDD.n1390 GND 0.02fF
C1982 VDD.n1391 GND 0.02fF
C1983 VDD.n1392 GND 0.02fF
C1984 VDD.n1393 GND 0.02fF
C1985 VDD.n1394 GND 0.02fF
C1986 VDD.n1395 GND 0.02fF
C1987 VDD.n1396 GND 0.02fF
C1988 VDD.n1397 GND 0.03fF
C1989 VDD.n1398 GND 0.03fF
C1990 VDD.n1399 GND 0.02fF
C1991 VDD.n1403 GND 0.29fF
C1992 VDD.n1404 GND 0.29fF
C1993 VDD.n1405 GND 0.01fF
C1994 VDD.n1406 GND 0.02fF
C1995 VDD.n1407 GND 0.04fF
C1996 VDD.n1408 GND 0.29fF
C1997 VDD.n1409 GND 0.01fF
C1998 VDD.n1410 GND 0.02fF
C1999 VDD.n1411 GND 0.02fF
C2000 VDD.n1412 GND 0.07fF
C2001 VDD.n1413 GND 0.24fF
C2002 VDD.n1414 GND 0.01fF
C2003 VDD.n1415 GND 0.01fF
C2004 VDD.n1416 GND 0.02fF
C2005 VDD.n1417 GND 0.18fF
C2006 VDD.n1418 GND 0.01fF
C2007 VDD.n1419 GND 0.02fF
C2008 VDD.n1420 GND 0.02fF
C2009 VDD.n1421 GND 0.09fF
C2010 VDD.n1422 GND 0.05fF
C2011 VDD.n1423 GND 0.17fF
C2012 VDD.n1424 GND 0.01fF
C2013 VDD.n1425 GND 0.02fF
C2014 VDD.n1426 GND 0.02fF
C2015 VDD.n1427 GND 0.16fF
C2016 VDD.n1428 GND 0.02fF
C2017 VDD.n1429 GND 0.02fF
C2018 VDD.n1430 GND 0.03fF
C2019 VDD.n1431 GND 0.15fF
C2020 VDD.n1432 GND 0.02fF
C2021 VDD.n1433 GND 0.02fF
C2022 VDD.n1434 GND 0.03fF
C2023 VDD.n1435 GND 0.17fF
C2024 VDD.n1436 GND 0.01fF
C2025 VDD.n1437 GND 0.09fF
C2026 VDD.n1438 GND 0.05fF
C2027 VDD.n1439 GND 0.02fF
C2028 VDD.n1440 GND 0.02fF
C2029 VDD.n1441 GND 0.18fF
C2030 VDD.n1442 GND 0.01fF
C2031 VDD.n1443 GND 0.02fF
C2032 VDD.n1444 GND 0.02fF
C2033 VDD.n1445 GND 0.24fF
C2034 VDD.n1446 GND 0.01fF
C2035 VDD.n1447 GND 0.07fF
C2036 VDD.n1448 GND 0.02fF
C2037 VDD.n1449 GND 0.29fF
C2038 VDD.n1450 GND 0.01fF
C2039 VDD.n1451 GND 0.02fF
C2040 VDD.n1452 GND 0.02fF
C2041 VDD.n1453 GND 0.29fF
C2042 VDD.n1454 GND 0.01fF
C2043 VDD.n1455 GND 0.02fF
C2044 VDD.n1456 GND 0.04fF
C2045 VDD.n1457 GND 0.33fF
C2046 VDD.n1458 GND 0.02fF
C2047 VDD.n1459 GND 0.02fF
C2048 VDD.n1460 GND 0.02fF
C2049 VDD.n1461 GND 0.06fF
C2050 VDD.n1462 GND 0.02fF
C2051 VDD.n1463 GND 0.02fF
C2052 VDD.n1464 GND 0.02fF
C2053 VDD.n1465 GND 0.02fF
C2054 VDD.n1466 GND 0.02fF
C2055 VDD.n1467 GND 0.02fF
C2056 VDD.n1468 GND 0.02fF
C2057 VDD.n1469 GND 0.02fF
C2058 VDD.n1470 GND 0.02fF
C2059 VDD.n1471 GND 0.02fF
C2060 VDD.n1472 GND 0.03fF
C2061 VDD.n1473 GND 0.03fF
C2062 VDD.n1474 GND 0.02fF
C2063 VDD.n1478 GND 0.29fF
C2064 VDD.n1479 GND 0.29fF
C2065 VDD.n1480 GND 0.01fF
C2066 VDD.n1481 GND 0.02fF
C2067 VDD.n1482 GND 0.04fF
C2068 VDD.n1483 GND 0.29fF
C2069 VDD.n1484 GND 0.01fF
C2070 VDD.n1485 GND 0.02fF
C2071 VDD.n1486 GND 0.02fF
C2072 VDD.n1487 GND 0.07fF
C2073 VDD.n1488 GND 0.24fF
C2074 VDD.n1489 GND 0.01fF
C2075 VDD.n1490 GND 0.01fF
C2076 VDD.n1491 GND 0.02fF
C2077 VDD.n1492 GND 0.18fF
C2078 VDD.n1493 GND 0.01fF
C2079 VDD.n1494 GND 0.02fF
C2080 VDD.n1495 GND 0.02fF
C2081 VDD.n1496 GND 0.09fF
C2082 VDD.n1497 GND 0.05fF
C2083 VDD.n1498 GND 0.17fF
C2084 VDD.n1499 GND 0.01fF
C2085 VDD.n1500 GND 0.02fF
C2086 VDD.n1501 GND 0.02fF
C2087 VDD.n1502 GND 0.16fF
C2088 VDD.n1503 GND 0.02fF
C2089 VDD.n1504 GND 0.02fF
C2090 VDD.n1505 GND 0.03fF
C2091 VDD.n1506 GND 0.15fF
C2092 VDD.n1507 GND 0.02fF
C2093 VDD.n1508 GND 0.02fF
C2094 VDD.n1509 GND 0.03fF
C2095 VDD.n1510 GND 0.17fF
C2096 VDD.n1511 GND 0.01fF
C2097 VDD.n1512 GND 0.09fF
C2098 VDD.n1513 GND 0.05fF
C2099 VDD.n1514 GND 0.02fF
C2100 VDD.n1515 GND 0.02fF
C2101 VDD.n1516 GND 0.18fF
C2102 VDD.n1517 GND 0.01fF
C2103 VDD.n1518 GND 0.02fF
C2104 VDD.n1519 GND 0.02fF
C2105 VDD.n1520 GND 0.24fF
C2106 VDD.n1521 GND 0.01fF
C2107 VDD.n1522 GND 0.07fF
C2108 VDD.n1523 GND 0.02fF
C2109 VDD.n1524 GND 0.29fF
C2110 VDD.n1525 GND 0.01fF
C2111 VDD.n1526 GND 0.02fF
C2112 VDD.n1527 GND 0.02fF
C2113 VDD.n1528 GND 0.29fF
C2114 VDD.n1529 GND 0.01fF
C2115 VDD.n1530 GND 0.02fF
C2116 VDD.n1531 GND 0.03fF
C2117 a_15669_1050.n0 GND 0.38fF
C2118 a_15669_1050.n1 GND 0.38fF
C2119 a_15669_1050.n2 GND 0.48fF
C2120 a_15669_1050.n3 GND 0.45fF
C2121 a_15669_1050.n4 GND 0.43fF
C2122 a_15669_1050.n5 GND 0.31fF
C2123 a_15669_1050.n6 GND 0.63fF
C2124 a_15669_1050.n7 GND 0.68fF
C2125 a_15669_1050.n8 GND 0.08fF
C2126 a_15669_1050.n9 GND 0.21fF
C2127 a_15669_1050.n10 GND 0.04fF
C2128 a_13105_989.n0 GND 0.65fF
C2129 a_13105_989.n1 GND 0.65fF
C2130 a_13105_989.n2 GND 0.82fF
C2131 a_13105_989.n3 GND 0.78fF
C2132 a_13105_989.n4 GND 0.69fF
C2133 a_13105_989.n5 GND 0.50fF
C2134 a_13105_989.t9 GND 0.91fF
C2135 a_13105_989.n6 GND 1.40fF
C2136 a_13105_989.n7 GND 0.50fF
C2137 a_13105_989.t8 GND 0.91fF
C2138 a_13105_989.n8 GND 0.68fF
C2139 a_13105_989.n9 GND 0.50fF
C2140 a_13105_989.t15 GND 0.91fF
C2141 a_13105_989.n10 GND 0.98fF
C2142 a_13105_989.n11 GND 1.80fF
C2143 a_13105_989.n12 GND 2.47fF
C2144 a_13105_989.n13 GND 0.87fF
C2145 a_13105_989.n14 GND 0.14fF
C2146 a_13105_989.n15 GND 0.41fF
C2147 a_13105_989.n16 GND 0.07fF
C2148 a_14802_210.n0 GND 0.02fF
C2149 a_14802_210.n1 GND 0.09fF
C2150 a_14802_210.t1 GND 0.23fF
C2151 a_14802_210.n2 GND 0.10fF
C2152 a_14802_210.n3 GND 0.07fF
C2153 a_14802_210.n4 GND 0.04fF
C2154 a_14802_210.n5 GND 0.08fF
C2155 a_14802_210.n6 GND 0.09fF
C2156 a_14802_210.n7 GND 0.04fF
C2157 a_14802_210.n8 GND 0.02fF
C2158 a_14802_210.n9 GND 0.01fF
C2159 a_14802_210.n10 GND 0.13fF
C2160 a_14802_