magic
tech sky130
magscale 1 2
timestamp 1645389040
<< nmos >>
rect 55 222 85 273
tri 85 222 101 238 sw
rect 55 192 161 222
tri 161 192 191 222 sw
rect 55 92 85 192
tri 85 176 101 192 nw
tri 145 176 161 192 ne
tri 85 92 101 108 sw
tri 145 92 161 108 se
rect 161 92 191 192
tri 55 62 85 92 ne
rect 85 62 161 92
tri 161 62 191 92 nw
<< ndiff >>
rect 5 62 55 273
rect 85 238 241 273
tri 85 222 101 238 ne
rect 101 222 241 238
tri 161 192 191 222 ne
tri 85 176 101 192 se
rect 101 176 145 192
tri 145 176 161 192 sw
rect 85 108 161 176
tri 85 92 101 108 ne
rect 101 92 145 108
tri 145 92 161 108 nw
tri 55 62 85 92 sw
tri 161 62 191 92 se
rect 191 62 241 222
rect 5 12 241 62
<< poly >>
rect 55 273 85 309
<< end >>
