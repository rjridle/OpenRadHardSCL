magic
tech sky130A
magscale 1 2
timestamp 1642388399
<< error_p >>
rect 609 322 610 323
rect 610 321 611 322
rect 127 318 128 319
rect 311 318 312 319
rect 128 317 129 318
rect 312 317 313 318
rect 625 291 626 292
rect 660 291 661 292
rect 143 287 144 288
rect 178 287 179 288
rect 327 287 328 288
rect 362 287 363 288
rect 625 188 626 189
rect 660 188 661 189
rect 143 184 144 185
rect 178 184 179 185
rect 327 184 328 185
rect 362 184 363 185
<< nwell >>
rect 0 591 796 1353
<< nmos >>
rect 98 318 128 368
rect 98 288 194 318
tri 194 288 224 318 sw
rect 282 318 312 368
rect 98 184 128 288
tri 128 272 144 288 nw
tri 178 272 194 288 ne
tri 128 184 144 200 sw
tri 178 184 194 200 se
rect 194 184 224 288
rect 282 288 378 318
tri 378 288 408 318 sw
tri 98 154 128 184 ne
rect 128 154 194 184
tri 194 154 224 184 nw
rect 282 184 312 288
tri 312 272 328 288 nw
tri 362 272 378 288 ne
tri 312 184 328 200 sw
tri 362 184 378 200 se
rect 378 184 408 288
tri 282 154 312 184 ne
rect 312 154 378 184
tri 378 154 408 184 nw
rect 580 322 610 372
rect 580 292 676 322
tri 676 292 706 322 sw
rect 580 188 610 292
tri 610 276 626 292 nw
tri 660 276 676 292 ne
tri 610 188 626 204 sw
tri 660 188 676 204 se
rect 676 188 706 292
tri 580 158 610 188 ne
rect 610 158 676 188
tri 676 158 706 188 nw
<< pmos >>
rect 98 629 128 1229
rect 186 629 216 1229
rect 282 629 312 1229
rect 370 629 400 1229
rect 580 629 610 1229
rect 668 629 698 1229
<< ndiff >>
rect 36 347 98 368
rect 36 313 52 347
rect 86 313 98 347
rect 128 347 282 368
rect 128 318 236 347
rect 36 279 98 313
tri 194 288 224 318 ne
rect 224 313 236 318
rect 270 313 282 347
rect 312 347 470 368
rect 312 318 420 347
rect 36 245 52 279
rect 86 245 98 279
rect 36 211 98 245
rect 36 177 52 211
rect 86 177 98 211
tri 128 272 144 288 se
rect 144 272 178 288
tri 178 272 194 288 sw
rect 128 240 194 272
rect 128 206 140 240
rect 174 206 194 240
rect 128 200 194 206
tri 128 184 144 200 ne
rect 144 184 178 200
tri 178 184 194 200 nw
rect 224 279 282 313
tri 378 288 408 318 ne
rect 408 313 420 318
rect 454 313 470 347
rect 224 245 236 279
rect 270 245 282 279
rect 224 211 282 245
rect 36 154 98 177
tri 98 154 128 184 sw
tri 194 154 224 184 se
rect 224 177 236 211
rect 270 177 282 211
tri 312 272 328 288 se
rect 328 272 362 288
tri 362 272 378 288 sw
rect 312 240 378 272
rect 312 206 324 240
rect 358 206 378 240
rect 312 200 378 206
tri 312 184 328 200 ne
rect 328 184 362 200
tri 362 184 378 200 nw
rect 408 279 470 313
rect 408 245 420 279
rect 454 245 470 279
rect 408 211 470 245
rect 224 154 282 177
tri 282 154 312 184 sw
tri 378 154 408 184 se
rect 408 177 420 211
rect 454 177 470 211
rect 408 154 470 177
rect 36 143 470 154
rect 36 109 52 143
rect 86 109 144 143
rect 178 109 236 143
rect 270 109 420 143
rect 454 109 470 143
rect 36 101 470 109
rect 524 298 580 372
rect 610 322 760 372
rect 524 264 534 298
rect 568 264 580 298
tri 676 292 706 322 ne
rect 706 298 760 322
rect 524 215 580 264
rect 524 181 534 215
rect 568 181 580 215
tri 610 276 626 292 se
rect 626 276 660 292
tri 660 276 676 292 sw
rect 610 244 676 276
rect 610 210 622 244
rect 656 210 676 244
rect 610 204 676 210
tri 610 188 626 204 ne
rect 626 188 660 204
tri 660 188 676 204 nw
rect 706 264 718 298
rect 752 264 760 298
rect 706 215 760 264
rect 524 158 580 181
tri 580 158 610 188 sw
tri 676 158 706 188 se
rect 706 181 718 215
rect 752 181 760 215
rect 706 158 760 181
rect 524 147 760 158
rect 524 113 534 147
rect 568 113 622 147
rect 656 113 718 147
rect 752 113 760 147
rect 524 101 760 113
<< pdiff >>
rect 42 1213 98 1229
rect 42 1179 52 1213
rect 86 1179 98 1213
rect 42 1145 98 1179
rect 42 1111 52 1145
rect 86 1111 98 1145
rect 42 1077 98 1111
rect 42 1043 52 1077
rect 86 1043 98 1077
rect 42 1009 98 1043
rect 42 975 52 1009
rect 86 975 98 1009
rect 42 941 98 975
rect 42 907 52 941
rect 86 907 98 941
rect 42 873 98 907
rect 42 839 52 873
rect 86 839 98 873
rect 42 805 98 839
rect 42 771 52 805
rect 86 771 98 805
rect 42 737 98 771
rect 42 703 52 737
rect 86 703 98 737
rect 42 629 98 703
rect 128 1213 186 1229
rect 128 1179 140 1213
rect 174 1179 186 1213
rect 128 1145 186 1179
rect 128 1111 140 1145
rect 174 1111 186 1145
rect 128 1077 186 1111
rect 128 1043 140 1077
rect 174 1043 186 1077
rect 128 1009 186 1043
rect 128 975 140 1009
rect 174 975 186 1009
rect 128 941 186 975
rect 128 907 140 941
rect 174 907 186 941
rect 128 873 186 907
rect 128 839 140 873
rect 174 839 186 873
rect 128 805 186 839
rect 128 771 140 805
rect 174 771 186 805
rect 128 737 186 771
rect 128 703 140 737
rect 174 703 186 737
rect 128 629 186 703
rect 216 1213 282 1229
rect 216 1179 236 1213
rect 270 1179 282 1213
rect 216 1145 282 1179
rect 216 1111 236 1145
rect 270 1111 282 1145
rect 216 1077 282 1111
rect 216 1043 236 1077
rect 270 1043 282 1077
rect 216 1009 282 1043
rect 216 975 236 1009
rect 270 975 282 1009
rect 216 941 282 975
rect 216 907 236 941
rect 270 907 282 941
rect 216 873 282 907
rect 216 839 236 873
rect 270 839 282 873
rect 216 805 282 839
rect 216 771 236 805
rect 270 771 282 805
rect 216 737 282 771
rect 216 703 236 737
rect 270 703 282 737
rect 216 629 282 703
rect 312 1213 370 1229
rect 312 1179 324 1213
rect 358 1179 370 1213
rect 312 1145 370 1179
rect 312 1111 324 1145
rect 358 1111 370 1145
rect 312 1077 370 1111
rect 312 1043 324 1077
rect 358 1043 370 1077
rect 312 1009 370 1043
rect 312 975 324 1009
rect 358 975 370 1009
rect 312 941 370 975
rect 312 907 324 941
rect 358 907 370 941
rect 312 873 370 907
rect 312 839 324 873
rect 358 839 370 873
rect 312 805 370 839
rect 312 771 324 805
rect 358 771 370 805
rect 312 737 370 771
rect 312 703 324 737
rect 358 703 370 737
rect 312 629 370 703
rect 400 1213 454 1229
rect 400 1179 412 1213
rect 446 1179 454 1213
rect 400 1145 454 1179
rect 400 1111 412 1145
rect 446 1111 454 1145
rect 400 1077 454 1111
rect 400 1043 412 1077
rect 446 1043 454 1077
rect 400 1009 454 1043
rect 400 975 412 1009
rect 446 975 454 1009
rect 400 941 454 975
rect 400 907 412 941
rect 446 907 454 941
rect 400 873 454 907
rect 400 839 412 873
rect 446 839 454 873
rect 400 805 454 839
rect 400 771 412 805
rect 446 771 454 805
rect 400 737 454 771
rect 400 703 412 737
rect 446 703 454 737
rect 400 629 454 703
rect 524 1213 580 1229
rect 524 1179 534 1213
rect 568 1179 580 1213
rect 524 1145 580 1179
rect 524 1111 534 1145
rect 568 1111 580 1145
rect 524 1077 580 1111
rect 524 1043 534 1077
rect 568 1043 580 1077
rect 524 1009 580 1043
rect 524 975 534 1009
rect 568 975 580 1009
rect 524 941 580 975
rect 524 907 534 941
rect 568 907 580 941
rect 524 873 580 907
rect 524 839 534 873
rect 568 839 580 873
rect 524 805 580 839
rect 524 771 534 805
rect 568 771 580 805
rect 524 737 580 771
rect 524 703 534 737
rect 568 703 580 737
rect 524 629 580 703
rect 610 1213 668 1229
rect 610 1179 622 1213
rect 656 1179 668 1213
rect 610 1145 668 1179
rect 610 1111 622 1145
rect 656 1111 668 1145
rect 610 1077 668 1111
rect 610 1043 622 1077
rect 656 1043 668 1077
rect 610 1009 668 1043
rect 610 975 622 1009
rect 656 975 668 1009
rect 610 941 668 975
rect 610 907 622 941
rect 656 907 668 941
rect 610 873 668 907
rect 610 839 622 873
rect 656 839 668 873
rect 610 805 668 839
rect 610 771 622 805
rect 656 771 668 805
rect 610 737 668 771
rect 610 703 622 737
rect 656 703 668 737
rect 610 629 668 703
rect 698 1213 752 1229
rect 698 1179 710 1213
rect 744 1179 752 1213
rect 698 1145 752 1179
rect 698 1111 710 1145
rect 744 1111 752 1145
rect 698 1077 752 1111
rect 698 1043 710 1077
rect 744 1043 752 1077
rect 698 1009 752 1043
rect 698 975 710 1009
rect 744 975 752 1009
rect 698 941 752 975
rect 698 907 710 941
rect 744 907 752 941
rect 698 873 752 907
rect 698 839 710 873
rect 744 839 752 873
rect 698 805 752 839
rect 698 771 710 805
rect 744 771 752 805
rect 698 737 752 771
rect 698 703 710 737
rect 744 703 752 737
rect 698 629 752 703
<< ndiffc >>
rect 52 313 86 347
rect 236 313 270 347
rect 52 245 86 279
rect 52 177 86 211
rect 140 206 174 240
rect 420 313 454 347
rect 236 245 270 279
rect 236 177 270 211
rect 324 206 358 240
rect 420 245 454 279
rect 420 177 454 211
rect 52 109 86 143
rect 144 109 178 143
rect 236 109 270 143
rect 420 109 454 143
rect 534 264 568 298
rect 534 181 568 215
rect 622 210 656 244
rect 718 264 752 298
rect 718 181 752 215
rect 534 113 568 147
rect 622 113 656 147
rect 718 113 752 147
<< pdiffc >>
rect 52 1179 86 1213
rect 52 1111 86 1145
rect 52 1043 86 1077
rect 52 975 86 1009
rect 52 907 86 941
rect 52 839 86 873
rect 52 771 86 805
rect 52 703 86 737
rect 140 1179 174 1213
rect 140 1111 174 1145
rect 140 1043 174 1077
rect 140 975 174 1009
rect 140 907 174 941
rect 140 839 174 873
rect 140 771 174 805
rect 140 703 174 737
rect 236 1179 270 1213
rect 236 1111 270 1145
rect 236 1043 270 1077
rect 236 975 270 1009
rect 236 907 270 941
rect 236 839 270 873
rect 236 771 270 805
rect 236 703 270 737
rect 324 1179 358 1213
rect 324 1111 358 1145
rect 324 1043 358 1077
rect 324 975 358 1009
rect 324 907 358 941
rect 324 839 358 873
rect 324 771 358 805
rect 324 703 358 737
rect 412 1179 446 1213
rect 412 1111 446 1145
rect 412 1043 446 1077
rect 412 975 446 1009
rect 412 907 446 941
rect 412 839 446 873
rect 412 771 446 805
rect 412 703 446 737
rect 534 1179 568 1213
rect 534 1111 568 1145
rect 534 1043 568 1077
rect 534 975 568 1009
rect 534 907 568 941
rect 534 839 568 873
rect 534 771 568 805
rect 534 703 568 737
rect 622 1179 656 1213
rect 622 1111 656 1145
rect 622 1043 656 1077
rect 622 975 656 1009
rect 622 907 656 941
rect 622 839 656 873
rect 622 771 656 805
rect 622 703 656 737
rect 710 1179 744 1213
rect 710 1111 744 1145
rect 710 1043 744 1077
rect 710 975 744 1009
rect 710 907 744 941
rect 710 839 744 873
rect 710 771 744 805
rect 710 703 744 737
<< psubdiff >>
rect 36 13 60 47
rect 94 13 129 47
rect 163 13 205 47
rect 239 13 273 47
rect 307 13 342 47
rect 376 13 410 47
rect 444 13 548 47
rect 582 13 617 47
rect 651 13 693 47
rect 727 13 760 47
<< nsubdiff >>
rect 36 1283 60 1317
rect 94 1283 128 1317
rect 162 1283 196 1317
rect 231 1283 265 1317
rect 299 1283 333 1317
rect 367 1283 401 1317
rect 435 1283 469 1317
rect 503 1283 537 1317
rect 572 1283 606 1317
rect 640 1283 674 1317
rect 708 1283 760 1317
<< psubdiffcont >>
rect 60 13 94 47
rect 129 13 163 47
rect 205 13 239 47
rect 273 13 307 47
rect 342 13 376 47
rect 410 13 444 47
rect 548 13 582 47
rect 617 13 651 47
rect 693 13 727 47
<< nsubdiffcont >>
rect 60 1283 94 1317
rect 128 1283 162 1317
rect 196 1283 231 1317
rect 265 1283 299 1317
rect 333 1283 367 1317
rect 401 1283 435 1317
rect 469 1283 503 1317
rect 537 1283 572 1317
rect 606 1283 640 1317
rect 674 1283 708 1317
<< poly >>
rect 98 1229 128 1255
rect 186 1229 216 1255
rect 282 1229 312 1255
rect 370 1229 400 1255
rect 580 1229 610 1255
rect 668 1229 698 1255
rect 98 612 128 629
rect 186 612 216 629
rect 98 582 216 612
rect 282 612 312 629
rect 370 612 400 629
rect 282 582 400 612
rect 580 612 610 629
rect 668 612 698 629
rect 580 582 698 612
rect 98 568 128 582
rect 62 552 128 568
rect 62 518 72 552
rect 106 518 128 552
rect 62 502 128 518
rect 98 368 128 502
rect 282 494 312 582
rect 580 578 610 582
rect 544 562 610 578
rect 544 528 554 562
rect 588 528 610 562
rect 544 512 610 528
rect 249 478 312 494
rect 249 444 259 478
rect 293 444 312 478
rect 249 428 312 444
rect 282 368 312 428
rect 580 372 610 512
<< polycont >>
rect 72 518 106 552
rect 554 528 588 562
rect 259 444 293 478
<< locali >>
rect 36 1317 760 1332
rect 36 1283 60 1317
rect 94 1283 128 1317
rect 162 1283 196 1317
rect 231 1283 265 1317
rect 299 1283 333 1317
rect 367 1283 401 1317
rect 435 1283 469 1317
rect 503 1283 537 1317
rect 572 1283 606 1317
rect 640 1283 674 1317
rect 708 1283 760 1317
rect 36 1270 760 1283
rect 52 1213 86 1270
rect 52 1145 86 1179
rect 52 1077 86 1111
rect 52 1009 86 1043
rect 52 941 86 975
rect 52 873 86 907
rect 52 805 86 839
rect 52 737 86 771
rect 52 687 86 703
rect 140 1213 174 1229
rect 140 1145 174 1179
rect 140 1077 174 1111
rect 140 1009 174 1043
rect 140 941 174 975
rect 140 873 174 907
rect 140 805 174 839
rect 140 737 174 771
rect 140 684 174 703
rect 236 1213 270 1270
rect 236 1145 270 1179
rect 236 1077 270 1111
rect 236 1009 270 1043
rect 236 941 270 975
rect 236 873 270 907
rect 236 805 270 839
rect 236 737 270 771
rect 236 687 270 703
rect 324 1213 358 1229
rect 324 1145 358 1179
rect 324 1077 358 1111
rect 324 1009 358 1043
rect 324 941 358 975
rect 324 873 358 907
rect 324 805 358 839
rect 324 737 358 771
rect 324 684 358 703
rect 412 1213 446 1270
rect 412 1145 446 1179
rect 412 1077 446 1111
rect 412 1009 446 1043
rect 412 941 446 975
rect 412 873 446 907
rect 412 805 446 839
rect 412 737 446 771
rect 72 552 106 568
rect 72 502 106 518
rect 140 562 174 650
rect 412 627 446 703
rect 534 1213 568 1270
rect 534 1145 568 1179
rect 534 1077 568 1111
rect 534 1009 568 1043
rect 534 941 568 975
rect 534 873 568 907
rect 534 805 568 839
rect 534 737 568 771
rect 534 627 568 703
rect 622 1213 656 1229
rect 622 1145 656 1179
rect 622 1077 656 1111
rect 622 1009 656 1043
rect 622 941 656 975
rect 622 873 656 907
rect 622 805 656 839
rect 622 737 656 771
rect 622 684 656 703
rect 554 562 588 578
rect 140 528 554 562
rect 52 347 86 363
rect 52 279 86 313
rect 52 211 86 245
rect 140 240 174 528
rect 554 512 588 528
rect 259 478 293 494
rect 259 428 293 444
rect 140 190 174 206
rect 236 347 454 363
rect 270 329 420 347
rect 236 279 270 313
rect 236 211 270 245
rect 52 143 86 177
rect 236 143 270 177
rect 324 240 358 280
rect 36 109 52 143
rect 86 109 144 143
rect 178 109 236 143
rect 270 109 286 143
rect 324 62 358 206
rect 420 279 454 313
rect 420 211 454 245
rect 420 143 454 177
rect 534 298 568 343
rect 534 215 568 264
rect 622 244 656 650
rect 710 1213 744 1270
rect 710 1145 744 1179
rect 710 1077 744 1111
rect 710 1009 744 1043
rect 710 941 744 975
rect 710 873 744 907
rect 710 805 744 839
rect 710 737 744 771
rect 710 627 744 703
rect 622 194 656 210
rect 718 298 752 343
rect 718 215 752 264
rect 534 147 568 181
rect 718 147 752 181
rect 404 109 420 143
rect 454 109 470 143
rect 568 113 622 147
rect 656 113 718 147
rect 534 62 568 113
rect 718 62 752 113
rect 36 47 760 62
rect 36 13 60 47
rect 94 13 129 47
rect 163 13 205 47
rect 239 13 273 47
rect 307 13 342 47
rect 376 13 410 47
rect 444 13 548 47
rect 582 13 617 47
rect 651 13 693 47
rect 727 13 760 47
rect 36 0 760 13
<< viali >>
rect 60 1283 94 1317
rect 128 1283 162 1317
rect 196 1283 231 1317
rect 265 1283 299 1317
rect 333 1283 367 1317
rect 401 1283 435 1317
rect 469 1283 503 1317
rect 537 1283 572 1317
rect 606 1283 640 1317
rect 674 1283 708 1317
rect 140 650 174 684
rect 324 650 358 684
rect 72 518 106 552
rect 622 650 656 684
rect 259 444 293 478
rect 60 13 94 47
rect 129 13 163 47
rect 205 13 239 47
rect 273 13 307 47
rect 342 13 376 47
rect 410 13 444 47
rect 548 13 582 47
rect 617 13 651 47
rect 693 13 727 47
<< metal1 >>
rect 36 1317 760 1332
rect 36 1283 60 1317
rect 94 1283 128 1317
rect 162 1283 196 1317
rect 231 1283 265 1317
rect 299 1283 333 1317
rect 367 1283 401 1317
rect 435 1283 469 1317
rect 503 1283 537 1317
rect 572 1283 606 1317
rect 640 1283 674 1317
rect 708 1283 760 1317
rect 36 1270 760 1283
rect 622 690 656 696
rect 134 684 180 690
rect 318 684 364 690
rect 616 684 662 690
rect 128 650 140 684
rect 174 650 324 684
rect 358 650 370 684
rect 616 650 622 684
rect 656 650 662 684
rect 134 649 364 650
rect 134 644 180 649
rect 318 644 364 649
rect 616 644 662 650
rect 622 614 656 644
rect 72 559 106 573
rect 62 552 112 559
rect 62 518 72 552
rect 106 518 112 552
rect 62 511 112 518
rect 72 497 106 511
rect 259 485 293 499
rect 249 478 299 485
rect 249 444 259 478
rect 293 444 299 478
rect 249 437 299 444
rect 259 423 293 437
rect 36 47 760 62
rect 36 13 60 47
rect 94 13 129 47
rect 163 13 205 47
rect 239 13 273 47
rect 307 13 342 47
rect 376 13 410 47
rect 444 13 548 47
rect 582 13 617 47
rect 651 13 693 47
rect 727 13 760 47
rect 36 0 760 13
<< labels >>
rlabel metal1 72 518 106 552 1 A
rlabel metal1 259 444 293 478 1 B
rlabel metal1 622 650 656 684 1 Y
rlabel metal1 42 29 42 29 1 VSS
rlabel metal1 39 1298 39 1298 1 VDD
<< end >>
