magic
tech sky130A
magscale 1 2
timestamp 1649546427
<< nwell >>
rect 84 1554 363 1575
rect 31 1492 413 1554
rect 84 832 363 1492
<< pdiffc >>
rect 117 1106 151 1140
rect 205 1106 239 1140
rect 293 1106 327 1140
<< psubdiff >>
rect 17 510 427 572
rect 31 13 55 47
rect 89 13 127 47
rect 161 13 205 47
rect 239 13 283 47
rect 317 13 355 47
rect 389 13 413 47
<< nsubdiff >>
rect 31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 205 1539
rect 239 1505 283 1539
rect 317 1505 355 1539
rect 389 1505 413 1539
rect -31 868 475 930
<< psubdiffcont >>
rect 55 13 89 47
rect 127 13 161 47
rect 205 13 239 47
rect 283 13 317 47
rect 355 13 389 47
<< nsubdiffcont >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 205 1505 239 1539
rect 283 1505 317 1539
rect 355 1505 389 1539
<< poly >>
rect 155 409 185 441
<< locali >>
rect 31 1539 413 1554
rect 31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 205 1539
rect 239 1505 283 1539
rect 317 1505 355 1539
rect 389 1505 413 1539
rect 31 1492 413 1505
rect 205 1450 239 1492
rect 117 1140 151 1157
rect 117 1046 151 1106
rect 205 1140 239 1157
rect 205 1062 239 1106
rect 293 1140 327 1157
rect 293 1062 327 1106
rect 117 1012 165 1046
rect 131 477 165 1012
rect 205 262 239 561
rect 279 395 313 953
rect 279 377 337 395
rect 279 361 313 377
rect 109 62 143 101
rect 205 62 239 117
rect 303 62 337 101
rect 31 47 413 62
rect 31 13 55 47
rect 89 13 127 47
rect 161 13 205 47
rect 239 13 283 47
rect 317 13 355 47
rect 389 13 413 47
rect 31 0 413 13
<< viali >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 205 1505 239 1539
rect 283 1505 317 1539
rect 355 1505 389 1539
rect 55 13 89 47
rect 127 13 161 47
rect 205 13 239 47
rect 283 13 317 47
rect 355 13 389 47
<< metal1 >>
rect 31 1539 413 1554
rect 31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 205 1539
rect 239 1505 283 1539
rect 317 1505 355 1539
rect 389 1505 413 1539
rect 31 1492 413 1505
rect 205 575 239 609
rect 31 47 413 62
rect 31 13 55 47
rect 89 13 127 47
rect 161 13 205 47
rect 239 13 283 47
rect 317 13 355 47
rect 389 13 413 47
rect 31 0 413 13
use li1_M1_contact  li1_M1_contact_0 pcells
timestamp 1648061256
transform -1 0 222 0 -1 592
box -53 -33 29 33
use nmos_top  nmos_top_0 pcells
timestamp 1648061425
transform -1 0 345 0 1 101
box 0 0 246 308
use pmos2  pmos2_0 pcells
timestamp 1648061063
transform 1 0 19 0 1 1450
box 52 -461 352 42
use diff_ring_side  diff_ring_side_1 pcells
timestamp 1648063806
transform 1 0 0 0 1 0
box -84 0 84 1575
use diff_ring_side  diff_ring_side_0
timestamp 1648063806
transform 1 0 444 0 1 0
box -84 0 84 1575
use poly_li1_contact  poly_li1_contact_0 pcells
timestamp 1648060378
transform 0 1 297 -1 0 987
box -32 -28 34 26
use poly_li1_contact  poly_li1_contact_1
timestamp 1648060378
transform 0 1 149 -1 0 445
box -32 -28 34 26
<< labels >>
rlabel metal1 205 575 239 609 1 YN
port 1 n
rlabel nwell 55 1505 89 1539 1 VDD
port 2 n
rlabel metal1 55 13 89 47 1 VSS
port 3 n
<< end >>
