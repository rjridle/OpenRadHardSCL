* SPICE3 file created from NAND3X1.ext - technology: sky130A

.subckt NAND3X1 Y A B VDD VSS
X0 VDD B Y VDD sky130_fd_pr__pfet_01v8 ad=2.26p pd=1.826u as=1.74p ps=1.374u w=2u l=0.15u M=2
X1 VDD a_599_989# Y VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X2 Y a_599_989# a_372_210# VSS sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=0p ps=0u w=3u l=0.15u
X3 Y A VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X4 VSS A a_91_103# VSS sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=0p ps=0u w=3u l=0.15u
X5 a_372_210# B a_91_103# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
C0 VDD Y 2.50fF
.ends
