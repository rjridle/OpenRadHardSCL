magic
tech sky130A
magscale 1 2
timestamp 1647328323
<< metal1 >>
rect 55 1505 89 1539
rect 131 649 165 683
rect 279 649 313 683
rect 55 13 89 47
use li1_M1_contact  li1_M1_contact_0 pcells
timestamp 1646004885
transform 1 0 148 0 1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_1
timestamp 1646004885
transform -1 0 296 0 -1 666
box -53 -33 29 33
use invx1_pcell  invx1_pcell_0 pcells
timestamp 1647328248
transform 1 0 0 0 1 0
box -84 0 528 1575
<< labels >>
rlabel metal1 148 666 148 666 1 A
port 1 n
rlabel metal1 296 666 296 666 1 Y
port 2 n
rlabel metal1 72 30 72 30 1 VSS
port 3 n
rlabel metal1 72 1522 72 1522 1 VDD
port 4 n
<< end >>
