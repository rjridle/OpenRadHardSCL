magic
tech sky130A
magscale 1 2
timestamp 1648048163
<< nwell >>
rect 55 1505 89 1539
<< psubdiffcont >>
rect 55 13 89 47
<< nsubdiffcont >>
rect 55 1505 89 1539
<< viali >>
rect 55 1505 89 1539
rect 55 13 89 47
<< metal1 >>
rect 833 871 1131 905
rect 1161 871 3979 905
rect 717 797 3058 831
rect 4349 797 4383 831
rect 4385 797 4831 831
rect 479 723 4683 757
rect 1389 649 1423 683
rect 1611 649 1645 683
rect 1681 649 3765 683
rect 4237 649 5012 683
rect 5015 649 5049 683
rect 268 575 2103 609
rect 2461 575 2762 609
use nand3x1_pcell  nand3x1_pcell_0 pcells
timestamp 1647328266
transform 1 0 962 0 1 0
box -84 0 1046 1575
use nand3x1_pcell  nand3x1_pcell_3
timestamp 1647328266
transform 1 0 0 0 1 0
box -84 0 1046 1575
use li1_M1_contact  li1_M1_contact_21 pcells
timestamp 1646004885
transform -1 0 222 0 -1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_12
timestamp 1646004885
transform -1 0 444 0 -1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_10
timestamp 1646004885
transform -1 0 666 0 -1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_4
timestamp 1646004885
transform -1 0 814 0 -1 888
box -53 -33 29 33
use nand2x1_pcell  nand2x1_pcell_0 pcells
timestamp 1647328257
transform 1 0 1924 0 1 0
box -84 0 750 1575
use li1_M1_contact  li1_M1_contact_20
timestamp 1646004885
transform 1 0 1406 0 1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_2
timestamp 1646004885
transform -1 0 1628 0 -1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_7
timestamp 1646004885
transform 1 0 2146 0 1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_6
timestamp 1646004885
transform -1 0 1776 0 -1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_3
timestamp 1646004885
transform 1 0 1184 0 1 888
box -53 -33 29 33
use nand3x1_pcell  nand3x1_pcell_2
timestamp 1647328266
transform 1 0 2590 0 1 0
box -84 0 1046 1575
use li1_M1_contact  li1_M1_contact_19
timestamp 1646004885
transform 1 0 2812 0 1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_18
timestamp 1646004885
transform -1 0 2442 0 -1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_1
timestamp 1646004885
transform 1 0 3256 0 1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_8
timestamp 1646004885
transform 1 0 3034 0 1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_11
timestamp 1646004885
transform -1 0 2294 0 -1 740
box -53 -33 29 33
use nand3x1_pcell  nand3x1_pcell_1
timestamp 1647328266
transform 1 0 3552 0 1 0
box -84 0 1046 1575
use nand2x1_pcell  nand2x1_pcell_1
timestamp 1647328257
transform 1 0 4514 0 1 0
box -84 0 750 1575
use li1_M1_contact  li1_M1_contact_16
timestamp 1646004885
transform -1 0 4218 0 -1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_14
timestamp 1646004885
transform -1 0 4366 0 -1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_9
timestamp 1646004885
transform -1 0 3404 0 -1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1646004885
transform 1 0 3774 0 1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_5
timestamp 1646004885
transform 1 0 3996 0 1 888
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_15
timestamp 1646004885
transform 1 0 4884 0 1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_13
timestamp 1646004885
transform 1 0 4736 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_17
timestamp 1646004885
transform 1 0 5032 0 1 666
box -53 -33 29 33
<< labels >>
rlabel metal1 649 797 683 831 1 CLK
port 1 n
rlabel metal1 1611 649 1645 683 1 RN
port 2 n
rlabel metal1 55 13 89 47 1 VSS
port 3 n
rlabel metal1 55 1505 89 1539 1 VDD
port 4 n
rlabel metal1 1389 649 1423 683 1 D
port 5 n
rlabel metal1 5015 649 5049 683 1 Q
port 6 n
rlabel metal1 4349 797 4383 831 1 QN
port 7 n
<< end >>
