* SPICE3 file created from TMRDFFSNQNX1.ext - technology: sky130A

.subckt TMRDFFSNQNX1 QN D CLK SN VDD GND
X0 VDD.t9 a_8357_1050.t5 a_8483_411.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X1 VDD.t112 D.t0 a_5101_1050.t4 VDD.t111 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X2 a_5227_411.t6 CLK.t0 VDD.t36 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X3 a_14869_1051.t7 a_3599_411.t7 a_15533_1051.t5  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X4 VDD.t80 D.t1 a_217_1050.t2 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X5 VDD.t130 a_1265_989.t5 a_1905_1050.t5  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X6 a_9985_1050.t1 a_10111_411.t7 VDD.t1 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X7 GND a_9985_1050.t6 a_11487_103.t0 GND sky130_fd_pr__nfet_01v8 ad=3.7611p pd=3.297u as=0p ps=0u w=0u l=0u
X8 VDD.t44 a_5101_1050.t5 a_6789_1050.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X9 a_15533_1051.t3 a_13367_411.t7 QN.t5 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X10 a_6789_1050.t2 a_6149_989.t5 VDD.t66  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X11 VDD.t177 a_11033_989.t5 a_11673_1050.t6 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X12 a_3599_411.t1 a_1265_989.t6 VDD.t128  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X13 a_13241_1050.t1 a_10111_411.t8 VDD.t191 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X14 a_1905_1050.t1 a_217_1050.t5 VDD.t84  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X15 VDD.t48 a_11673_1050.t7 a_11033_989.t0 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X16 a_14869_1051.t3 a_8483_411.t8 a_15533_1051.t2  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X17 VDD.t5 a_343_411.t7 a_217_1050.t0 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X18 VDD.t54 a_5227_411.t7 a_5101_1050.t2  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X19 GND a_11673_1050.t8 a_12470_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X20 a_11673_1050.t5 a_11033_989.t6 VDD.t56 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X21 VDD.t132 a_217_1050.t6 a_343_411.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X22 a_3473_1050.t1 a_3599_411.t9 VDD.t110 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X23 VDD.t70 a_13241_1050.t5 a_13367_411.t2  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X24 a_10111_411.t6 CLK.t2 VDD.t159 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X25 GND a_8483_411.t11 a_15430_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X26 a_5227_411.t2 a_6149_989.t7 VDD.t90  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X27 VDD.t76 a_11033_989.t7 a_10111_411.t1 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X28 VDD.t104 a_5227_411.t8 a_8357_1050.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X29 a_13241_1050.t4 a_13367_411.t9 VDD.t116 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X30 a_6149_989.t3 CLK.t3 VDD.t11  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X31 a_14869_1051.t1 a_8483_411.t9 VDD.t23 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X32 a_13367_411.t1 a_13241_1050.t6 VDD.t68  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X33 VDD.t74 a_6149_989.t8 a_8483_411.t4 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X34 GND a_217_1050.t7 a_757_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X35 QN a_13367_411.t11 a_16096_101.t0 GND sky130_fd_pr__nfet_01v8 ad=5.373p pd=4.72u as=0p ps=0u w=0u l=0u
X36 VDD.t58 a_13367_411.t10 a_14869_1051.t5  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X37 GND D.t3 a_112_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X38 VDD.t34 CLK.t5 a_343_411.t3 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X39 a_3473_1050.t4 a_343_411.t8 VDD.t14  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X40 VDD.t60 a_1905_1050.t7 a_1265_989.t0 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X41 a_8483_411.t6 SN.t2 VDD.t167  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X42 VDD.t165 SN.t3 a_13367_411.t4 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X43 a_10111_411.t2 a_9985_1050.t7 VDD.t94  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X44 GND a_343_411.t9 a_3368_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X45 a_15533_1051.t1 a_8483_411.t10 a_14869_1051.t2 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X46 VDD.t62 a_10111_411.t9 a_9985_1050.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X47 GND a_8357_1050.t7 a_8897_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X48 VDD.t163 SN.t4 a_11673_1050.t1 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X49 a_6149_989.t1 a_6789_1050.t8 VDD.t46  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X50 VDD.t169 a_3473_1050.t5 a_3599_411.t4 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X51 VDD.t64 a_1265_989.t9 a_3599_411.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X52 VDD.t40 a_1265_989.t10 a_343_411.t6 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X53 a_8483_411.t0 a_8357_1050.t6 VDD.t7  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X54 VDD.t179 a_11033_989.t9 a_13367_411.t6 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X55 VDD.t134 a_5101_1050.t6 a_5227_411.t4  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X56 a_15533_1051.t4 a_3599_411.t10 a_14869_1051.t6 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X57 a_8483_411.t2 a_6149_989.t10 VDD.t32  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X58 a_217_1050.t1 D.t4 VDD.t82 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X59 VDD.t137 D.t5 a_9985_1050.t4  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X60 a_1905_1050.t4 a_1265_989.t11 VDD.t114 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X61 GND D.t6 a_9880_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X62 a_6789_1050.t0 a_5101_1050.t7 VDD.t3  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X63 VDD.t96 a_9985_1050.t8 a_11673_1050.t3 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X64 GND a_217_1050.t8 a_1719_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X65 QN.t4 a_13367_411.t12 a_15533_1051.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X66 QN a_3599_411.t12 a_15430_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X67 VDD.t161 SN.t7 a_3599_411.t3 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X68 VDD.t122 SN.t8 a_6789_1050.t5  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X69 a_11033_989.t1 a_11673_1050.t9 VDD.t72 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X70 a_1905_1050.t3 SN.t9 VDD.t157  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X71 a_5101_1050.t1 a_5227_411.t10 VDD.t52 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X72 a_217_1050.t4 a_343_411.t10 VDD.t173  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X73 GND a_10111_411.t12 a_13136_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X74 GND a_1905_1050.t8 a_2702_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X75 a_6789_1050.t6 SN.t10 VDD.t155 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X76 QN.t2 a_3599_411.t11 a_15533_1051.t6  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X77 VDD.t108 a_9985_1050.t9 a_10111_411.t3 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X78 GND a_13241_1050.t7 a_13781_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X79 a_343_411.t0 a_217_1050.t9 VDD.t139  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X80 VDD.t20 a_8483_411.t12 a_8357_1050.t4 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X81 GND a_5227_411.t12 a_8252_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X82 VDD.t88 a_6149_989.t12 a_6789_1050.t3  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X83 GND a_5101_1050.t8 a_5641_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X84 VDD.t184 a_10111_411.t11 a_13241_1050.t0 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X85 a_10111_411.t4 a_11033_989.t11 VDD.t141  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X86 VDD.t118 a_217_1050.t10 a_1905_1050.t0 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X87 a_8357_1050.t3 a_5227_411.t11 VDD.t188  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X88 VDD.t195 a_6789_1050.t9 a_6149_989.t0 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X89 a_11033_989.t3 CLK.t8 VDD.t50  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X90 GND a_8483_411.t15 a_14764_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X91 a_5101_1050.t3 D.t7 VDD.t27 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X92 a_343_411.t2 CLK.t10 VDD.t102  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X93 a_14869_1051.t4 a_13367_411.t13 VDD.t29 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X94 a_9985_1050.t3 D.t8 VDD.t38  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X95 a_13367_411.t3 SN.t12 VDD.t153 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X96 a_1265_989.t1 a_1905_1050.t9 VDD.t120  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X97 VDD.t106 a_3599_411.t13 a_3473_1050.t0 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X98 VDD.t181 CLK.t11 a_10111_411.t5  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X99 a_11673_1050.t0 SN.t13 VDD.t151 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X100 VDD.t126 CLK.t12 a_1265_989.t3  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X101 GND a_5101_1050.t10 a_6603_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X102 VDD.t86 a_6149_989.t13 a_5227_411.t1 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X103 VDD.t143 a_13367_411.t14 a_13241_1050.t3  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X104 a_8357_1050.t0 a_8483_411.t13 VDD.t18 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X105 a_3599_411.t6 a_3473_1050.t6 VDD.t193  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X106 VDD.t78 CLK.t13 a_6149_989.t2 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X107 GND a_3473_1050.t7 a_4013_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X108 VDD.t16 a_8483_411.t14 a_14869_1051.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X109 QN a_13367_411.t15 a_14764_101.t1 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X110 a_343_411.t5 a_1265_989.t13 VDD.t92 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X111 VDD.t171 a_343_411.t12 a_3473_1050.t3  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X112 a_5227_411.t3 a_5101_1050.t9 VDD.t124 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X113 a_13367_411.t0 a_11033_989.t13 VDD.t42  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X114 VDD.t149 SN.t15 a_8483_411.t5 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X115 GND a_6789_1050.t7 a_7586_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X116 a_1265_989.t2 CLK.t14 VDD.t100  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X117 VDD.t147 SN.t16 a_1905_1050.t2 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X118 GND a_9985_1050.t5 a_10525_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X119 GND a_3599_411.t8 a_16096_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X120 GND D.t2 a_4996_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X121 a_11673_1050.t2 a_9985_1050.t10 VDD.t175  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X122 VDD.t186 CLK.t15 a_5227_411.t5 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X123 a_15533_1051.t7 a_3599_411.t15 QN.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X124 a_3599_411.t2 SN.t17 VDD.t145 0<��� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X125 VDD.t98 CLK.t17 a_11033_989.t2  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
C0 CLK SN 0.46fF
C1 QN VDD 0.73fF
C2 VDD D 0.95fF
C3 VDD CLK 7.98fF
C4 D CLK 0.39fF
C5 VDD SN 1.76fF
C6 D SN 9.38fF
R0 a_8357_1050.n3 a_8357_1050.t5 512.525
R1 a_8357_1050.n4 a_8357_1050.t7 417.109
R2 a_8357_1050.n3 a_8357_1050.t6 371.139
R3 a_8357_1050.n7 a_8357_1050.n5 367.82
R4 a_8357_1050.n4 a_8357_1050.n3 179.837
R5 a_8357_1050.n2 a_8357_1050.n1 157.964
R6 a_8357_1050.n5 a_8357_1050.n2 104.282
R7 a_8357_1050.n2 a_8357_1050.n0 91.706
R8 a_8357_1050.n7 a_8357_1050.n6 15.218
R9 a_8357_1050.n0 a_8357_1050.t4 14.282
R10 a_8357_1050.n0 a_8357_1050.t0 14.282
R11 a_8357_1050.n1 a_8357_1050.t1 14.282
R12 a_8357_1050.n1 a_8357_1050.t3 14.282
R13 a_8357_1050.n8 a_8357_1050.n7 12.014
R14 a_8357_1050.n5 a_8357_1050.n4 10.615
R15 a_8483_411.n8 a_8483_411.t14 512.525
R16 a_8483_411.n6 a_8483_411.t8 477.179
R17 a_8483_411.n11 a_8483_411.t12 472.359
R18 a_8483_411.n7 a_8483_411.t11 440.954
R19 a_8483_411.n6 a_8483_411.t10 406.485
R20 a_8483_411.n11 a_8483_411.t13 384.527
R21 a_8483_411.n8 a_8483_411.t9 371.139
R22 a_8483_411.n10 a_8483_411.t15 350.777
R23 a_8483_411.n12 a_8483_411.t7 314.896
R24 a_8483_411.n16 a_8483_411.n14 308.216
R25 a_8483_411.n12 a_8483_411.n11 182.814
R26 a_8483_411.n14 a_8483_411.n5 179.199
R27 a_8483_411.n4 a_8483_411.n3 161.352
R28 a_8483_411.n5 a_8483_411.n1 95.095
R29 a_8483_411.n4 a_8483_411.n2 95.095
R30 a_8483_411.n10 a_8483_411.n9 83.75
R31 a_8483_411.n9 a_8483_411.n8 77.972
R32 a_8483_411.n5 a_8483_411.n4 66.258
R33 a_8483_411.n17 a_8483_411.n0 55.263
R34 a_8483_411.n16 a_8483_411.n15 30
R35 a_8483_411.n17 a_8483_411.n16 23.684
R36 a_8483_411.n13 a_8483_411.n10 23.649
R37 a_8483_411.n7 a_8483_411.n6 21.4
R38 a_8483_411.n1 a_8483_411.t4 14.282
R39 a_8483_411.n1 a_8483_411.t2 14.282
R40 a_8483_411.n2 a_8483_411.t5 14.282
R41 a_8483_411.n2 a_8483_411.t6 14.282
R42 a_8483_411.n3 a_8483_411.t1 14.282
R43 a_8483_411.n3 a_8483_411.t0 14.282
R44 a_8483_411.n13 a_8483_411.n12 8.685
R45 a_8483_411.n9 a_8483_411.n7 6.833
R46 a_8483_411.n14 a_8483_411.n13 4.65
R47 VDD.n759 VDD.n748 144.705
R48 VDD.n834 VDD.n827 144.705
R49 VDD.n909 VDD.n902 144.705
R50 VDD.n966 VDD.n959 144.705
R51 VDD.n1023 VDD.n1016 144.705
R52 VDD.n1098 VDD.n1091 144.705
R53 VDD.n1155 VDD.n1148 144.705
R54 VDD.n1230 VDD.n1223 144.705
R55 VDD.n1305 VDD.n1298 144.705
R56 VDD.n656 VDD.n649 144.705
R57 VDD.n1362 VDD.n1355 144.705
R58 VDD.n581 VDD.n574 144.705
R59 VDD.n524 VDD.n517 144.705
R60 VDD.n449 VDD.n442 144.705
R61 VDD.n374 VDD.n367 144.705
R62 VDD.n317 VDD.n310 144.705
R63 VDD.n260 VDD.n253 144.705
R64 VDD.n185 VDD.n178 144.705
R65 VDD.n128 VDD.n121 144.705
R66 VDD.n75 VDD.n64 144.705
R67 VDD.n801 VDD.t40 143.754
R68 VDD.n876 VDD.t130 143.754
R69 VDD.n1065 VDD.t64 143.754
R70 VDD.n1197 VDD.t86 143.754
R71 VDD.n1272 VDD.t88 143.754
R72 VDD.n590 VDD.t74 143.754
R73 VDD.n458 VDD.t76 143.754
R74 VDD.n383 VDD.t177 143.754
R75 VDD.n194 VDD.t179 143.754
R76 VDD.n726 VDD.t5 143.754
R77 VDD.n934 VDD.t126 143.754
R78 VDD.n991 VDD.t106 143.754
R79 VDD.n1123 VDD.t54 143.754
R80 VDD.n1330 VDD.t78 143.754
R81 VDD.n659 VDD.t20 143.754
R82 VDD.n527 VDD.t62 143.754
R83 VDD.n320 VDD.t98 143.754
R84 VDD.n263 VDD.t143 143.754
R85 VDD.n153 VDD.t23 135.539
R86 VDD.n131 VDD.t58 135.539
R87 VDD.n704 VDD.t82 135.17
R88 VDD.n766 VDD.t139 135.17
R89 VDD.n841 VDD.t84 135.17
R90 VDD.n912 VDD.t120 135.17
R91 VDD.n969 VDD.t14 135.17
R92 VDD.n1030 VDD.t193 135.17
R93 VDD.n1101 VDD.t27 135.17
R94 VDD.n1162 VDD.t124 135.17
R95 VDD.n1237 VDD.t3 135.17
R96 VDD.n1308 VDD.t46 135.17
R97 VDD.n1365 VDD.t188 135.17
R98 VDD.n620 VDD.t7 135.17
R99 VDD.n549 VDD.t38 135.17
R100 VDD.n488 VDD.t94 135.17
R101 VDD.n413 VDD.t175 135.17
R102 VDD.n342 VDD.t72 135.17
R103 VDD.n285 VDD.t191 135.17
R104 VDD.n224 VDD.t68 135.17
R105 VDD.n141 VDD.n140 129.849
R106 VDD.n718 VDD.n717 129.472
R107 VDD.n776 VDD.n775 129.472
R108 VDD.n792 VDD.n791 129.472
R109 VDD.n851 VDD.n850 129.472
R110 VDD.n867 VDD.n866 129.472
R111 VDD.n926 VDD.n925 129.472
R112 VDD.n983 VDD.n982 129.472
R113 VDD.n1040 VDD.n1039 129.472
R114 VDD.n1056 VDD.n1055 129.472
R115 VDD.n1115 VDD.n1114 129.472
R116 VDD.n1172 VDD.n1171 129.472
R117 VDD.n1188 VDD.n1187 129.472
R118 VDD.n1247 VDD.n1246 129.472
R119 VDD.n1263 VDD.n1262 129.472
R120 VDD.n1322 VDD.n1321 129.472
R121 VDD.n669 VDD.n668 129.472
R122 VDD.n611 VDD.n610 129.472
R123 VDD.n599 VDD.n598 129.472
R124 VDD.n537 VDD.n536 129.472
R125 VDD.n479 VDD.n478 129.472
R126 VDD.n467 VDD.n466 129.472
R127 VDD.n404 VDD.n403 129.472
R128 VDD.n392 VDD.n391 129.472
R129 VDD.n330 VDD.n329 129.472
R130 VDD.n273 VDD.n272 129.472
R131 VDD.n215 VDD.n214 129.472
R132 VDD.n203 VDD.n202 129.472
R133 VDD.n60 VDD.n59 92.5
R134 VDD.n58 VDD.n57 92.5
R135 VDD.n56 VDD.n55 92.5
R136 VDD.n54 VDD.n53 92.5
R137 VDD.n62 VDD.n61 92.5
R138 VDD.n117 VDD.n116 92.5
R139 VDD.n115 VDD.n114 92.5
R140 VDD.n113 VDD.n112 92.5
R141 VDD.n111 VDD.n110 92.5
R142 VDD.n119 VDD.n118 92.5
R143 VDD.n174 VDD.n173 92.5
R144 VDD.n172 VDD.n171 92.5
R145 VDD.n170 VDD.n169 92.5
R146 VDD.n168 VDD.n167 92.5
R147 VDD.n176 VDD.n175 92.5
R148 VDD.n249 VDD.n248 92.5
R149 VDD.n247 VDD.n246 92.5
R150 VDD.n245 VDD.n244 92.5
R151 VDD.n243 VDD.n242 92.5
R152 VDD.n251 VDD.n250 92.5
R153 VDD.n306 VDD.n305 92.5
R154 VDD.n304 VDD.n303 92.5
R155 VDD.n302 VDD.n301 92.5
R156 VDD.n300 VDD.n299 92.5
R157 VDD.n308 VDD.n307 92.5
R158 VDD.n363 VDD.n362 92.5
R159 VDD.n361 VDD.n360 92.5
R160 VDD.n359 VDD.n358 92.5
R161 VDD.n357 VDD.n356 92.5
R162 VDD.n365 VDD.n364 92.5
R163 VDD.n438 VDD.n437 92.5
R164 VDD.n436 VDD.n435 92.5
R165 VDD.n434 VDD.n433 92.5
R166 VDD.n432 VDD.n431 92.5
R167 VDD.n440 VDD.n439 92.5
R168 VDD.n513 VDD.n512 92.5
R169 VDD.n511 VDD.n510 92.5
R170 VDD.n509 VDD.n508 92.5
R171 VDD.n507 VDD.n506 92.5
R172 VDD.n515 VDD.n514 92.5
R173 VDD.n570 VDD.n569 92.5
R174 VDD.n568 VDD.n567 92.5
R175 VDD.n566 VDD.n565 92.5
R176 VDD.n564 VDD.n563 92.5
R177 VDD.n572 VDD.n571 92.5
R178 VDD.n645 VDD.n644 92.5
R179 VDD.n643 VDD.n642 92.5
R180 VDD.n641 VDD.n640 92.5
R181 VDD.n639 VDD.n638 92.5
R182 VDD.n647 VDD.n646 92.5
R183 VDD.n1351 VDD.n1350 92.5
R184 VDD.n1349 VDD.n1348 92.5
R185 VDD.n1347 VDD.n1346 92.5
R186 VDD.n1345 VDD.n1344 92.5
R187 VDD.n1353 VDD.n1352 92.5
R188 VDD.n1294 VDD.n1293 92.5
R189 VDD.n1292 VDD.n1291 92.5
R190 VDD.n1290 VDD.n1289 92.5
R191 VDD.n1288 VDD.n1287 92.5
R192 VDD.n1296 VDD.n1295 92.5
R193 VDD.n1219 VDD.n1218 92.5
R194 VDD.n1217 VDD.n1216 92.5
R195 VDD.n1215 VDD.n1214 92.5
R196 VDD.n1213 VDD.n1212 92.5
R197 VDD.n1221 VDD.n1220 92.5
R198 VDD.n1144 VDD.n1143 92.5
R199 VDD.n1142 VDD.n1141 92.5
R200 VDD.n1140 VDD.n1139 92.5
R201 VDD.n1138 VDD.n1137 92.5
R202 VDD.n1146 VDD.n1145 92.5
R203 VDD.n1087 VDD.n1086 92.5
R204 VDD.n1085 VDD.n1084 92.5
R205 VDD.n1083 VDD.n1082 92.5
R206 VDD.n1081 VDD.n1080 92.5
R207 VDD.n1089 VDD.n1088 92.5
R208 VDD.n1012 VDD.n1011 92.5
R209 VDD.n1010 VDD.n1009 92.5
R210 VDD.n1008 VDD.n1007 92.5
R211 VDD.n1006 VDD.n1005 92.5
R212 VDD.n1014 VDD.n1013 92.5
R213 VDD.n955 VDD.n954 92.5
R214 VDD.n953 VDD.n952 92.5
R215 VDD.n951 VDD.n950 92.5
R216 VDD.n949 VDD.n948 92.5
R217 VDD.n957 VDD.n956 92.5
R218 VDD.n898 VDD.n897 92.5
R219 VDD.n896 VDD.n895 92.5
R220 VDD.n894 VDD.n893 92.5
R221 VDD.n892 VDD.n891 92.5
R222 VDD.n900 VDD.n899 92.5
R223 VDD.n823 VDD.n822 92.5
R224 VDD.n821 VDD.n820 92.5
R225 VDD.n819 VDD.n818 92.5
R226 VDD.n817 VDD.n816 92.5
R227 VDD.n825 VDD.n824 92.5
R228 VDD.n744 VDD.n743 92.5
R229 VDD.n742 VDD.n741 92.5
R230 VDD.n740 VDD.n739 92.5
R231 VDD.n738 VDD.n737 92.5
R232 VDD.n746 VDD.n745 92.5
R233 VDD.n692 VDD.n691 92.5
R234 VDD.n690 VDD.n689 92.5
R235 VDD.n688 VDD.n687 92.5
R236 VDD.n686 VDD.n685 92.5
R237 VDD.n694 VDD.n693 92.5
R238 VDD.n14 VDD.n1 92.5
R239 VDD.n5 VDD.n4 92.5
R240 VDD.n7 VDD.n6 92.5
R241 VDD.n9 VDD.n8 92.5
R242 VDD.n11 VDD.n10 92.5
R243 VDD.n13 VDD.n12 92.5
R244 VDD.n21 VDD.n20 92.059
R245 VDD.n74 VDD.n73 92.059
R246 VDD.n127 VDD.n126 92.059
R247 VDD.n184 VDD.n183 92.059
R248 VDD.n259 VDD.n258 92.059
R249 VDD.n316 VDD.n315 92.059
R250 VDD.n373 VDD.n372 92.059
R251 VDD.n448 VDD.n447 92.059
R252 VDD.n523 VDD.n522 92.059
R253 VDD.n580 VDD.n579 92.059
R254 VDD.n655 VDD.n654 92.059
R255 VDD.n1361 VDD.n1360 92.059
R256 VDD.n1304 VDD.n1303 92.059
R257 VDD.n1229 VDD.n1228 92.059
R258 VDD.n1154 VDD.n1153 92.059
R259 VDD.n1097 VDD.n1096 92.059
R260 VDD.n1022 VDD.n1021 92.059
R261 VDD.n965 VDD.n964 92.059
R262 VDD.n908 VDD.n907 92.059
R263 VDD.n833 VDD.n832 92.059
R264 VDD.n758 VDD.n757 92.059
R265 VDD.n700 VDD.n699 92.059
R266 VDD.n20 VDD.n16 67.194
R267 VDD.n20 VDD.n17 67.194
R268 VDD.n20 VDD.n18 67.194
R269 VDD.n20 VDD.n19 67.194
R270 VDD.n684 VDD.n683 44.141
R271 VDD.n815 VDD.n814 44.141
R272 VDD.n890 VDD.n889 44.141
R273 VDD.n947 VDD.n946 44.141
R274 VDD.n1004 VDD.n1003 44.141
R275 VDD.n1079 VDD.n1078 44.141
R276 VDD.n1136 VDD.n1135 44.141
R277 VDD.n1211 VDD.n1210 44.141
R278 VDD.n1286 VDD.n1285 44.141
R279 VDD.n1343 VDD.n1342 44.141
R280 VDD.n637 VDD.n636 44.141
R281 VDD.n562 VDD.n561 44.141
R282 VDD.n505 VDD.n504 44.141
R283 VDD.n430 VDD.n429 44.141
R284 VDD.n355 VDD.n354 44.141
R285 VDD.n298 VDD.n297 44.141
R286 VDD.n241 VDD.n240 44.141
R287 VDD.n166 VDD.n165 44.141
R288 VDD.n109 VDD.n108 44.141
R289 VDD.n5 VDD.n3 44.141
R290 VDD.n814 VDD.n812 44.107
R291 VDD.n889 VDD.n887 44.107
R292 VDD.n946 VDD.n944 44.107
R293 VDD.n1003 VDD.n1001 44.107
R294 VDD.n1078 VDD.n1076 44.107
R295 VDD.n1135 VDD.n1133 44.107
R296 VDD.n1210 VDD.n1208 44.107
R297 VDD.n1285 VDD.n1283 44.107
R298 VDD.n1342 VDD.n1340 44.107
R299 VDD.n636 VDD.n634 44.107
R300 VDD.n561 VDD.n559 44.107
R301 VDD.n504 VDD.n502 44.107
R302 VDD.n429 VDD.n427 44.107
R303 VDD.n354 VDD.n352 44.107
R304 VDD.n297 VDD.n295 44.107
R305 VDD.n240 VDD.n238 44.107
R306 VDD.n165 VDD.n163 44.107
R307 VDD.n108 VDD.n106 44.107
R308 VDD.n683 VDD.n681 44.107
R309 VDD.n3 VDD.n2 44.107
R310 VDD.n20 VDD.n15 41.052
R311 VDD.n68 VDD.n66 39.742
R312 VDD.n68 VDD.n67 39.742
R313 VDD.n70 VDD.n69 39.742
R314 VDD.n123 VDD.n122 39.742
R315 VDD.n180 VDD.n179 39.742
R316 VDD.n255 VDD.n254 39.742
R317 VDD.n312 VDD.n311 39.742
R318 VDD.n369 VDD.n368 39.742
R319 VDD.n444 VDD.n443 39.742
R320 VDD.n519 VDD.n518 39.742
R321 VDD.n576 VDD.n575 39.742
R322 VDD.n651 VDD.n650 39.742
R323 VDD.n1357 VDD.n1356 39.742
R324 VDD.n1300 VDD.n1299 39.742
R325 VDD.n1225 VDD.n1224 39.742
R326 VDD.n1150 VDD.n1149 39.742
R327 VDD.n1093 VDD.n1092 39.742
R328 VDD.n1018 VDD.n1017 39.742
R329 VDD.n961 VDD.n960 39.742
R330 VDD.n904 VDD.n903 39.742
R331 VDD.n829 VDD.n828 39.742
R332 VDD.n696 VDD.n695 39.742
R333 VDD.n756 VDD.n753 39.742
R334 VDD.n756 VDD.n755 39.742
R335 VDD.n752 VDD.n751 39.742
R336 VDD.n108 VDD.n107 38
R337 VDD.n165 VDD.n164 38
R338 VDD.n240 VDD.n239 38
R339 VDD.n297 VDD.n296 38
R340 VDD.n354 VDD.n353 38
R341 VDD.n429 VDD.n428 38
R342 VDD.n504 VDD.n503 38
R343 VDD.n561 VDD.n560 38
R344 VDD.n636 VDD.n635 38
R345 VDD.n1342 VDD.n1341 38
R346 VDD.n1285 VDD.n1284 38
R347 VDD.n1210 VDD.n1209 38
R348 VDD.n1135 VDD.n1134 38
R349 VDD.n1078 VDD.n1077 38
R350 VDD.n1003 VDD.n1002 38
R351 VDD.n946 VDD.n945 38
R352 VDD.n889 VDD.n888 38
R353 VDD.n814 VDD.n813 38
R354 VDD.n683 VDD.n682 38
R355 VDD.n812 VDD.n811 36.774
R356 VDD.n887 VDD.n886 36.774
R357 VDD.n944 VDD.n943 36.774
R358 VDD.n1001 VDD.n1000 36.774
R359 VDD.n1076 VDD.n1075 36.774
R360 VDD.n1133 VDD.n1132 36.774
R361 VDD.n1208 VDD.n1207 36.774
R362 VDD.n1283 VDD.n1282 36.774
R363 VDD.n1340 VDD.n1339 36.774
R364 VDD.n634 VDD.n633 36.774
R365 VDD.n559 VDD.n558 36.774
R366 VDD.n502 VDD.n501 36.774
R367 VDD.n427 VDD.n426 36.774
R368 VDD.n352 VDD.n351 36.774
R369 VDD.n295 VDD.n294 36.774
R370 VDD.n238 VDD.n237 36.774
R371 VDD.n163 VDD.n162 36.774
R372 VDD.n106 VDD.n105 36.774
R373 VDD.n66 VDD.n65 36.774
R374 VDD.n755 VDD.n754 36.774
R375 VDD.n196 0<��� 35.8
R376 VDD.n385 0<��� 35.8
R377 VDD.n460 0<��� 35.8
R378 VDD.n592 0<��� 35.8
R379 VDD.n1266  35.8
R380 VDD.n1191 0<��� 35.8
R381 VDD.n1059  35.8
R382 VDD.n870  35.8
R383 VDD.n795 0<��� 35.8
R384 VDD.n220  33.243
R385 VDD.n409  33.243
R386 VDD.n484  33.243
R387 VDD.n616  33.243
R388 VDD.n1242  33.243
R389 VDD.n1167 0<��� 33.243
R390 VDD.n1035  33.243
R391 VDD.n846  33.243
R392 VDD.n771  33.243
R393 VDD.n1 VDD.n0 30.923
R394 VDD.n73 VDD.n71 26.38
R395 VDD.n73 VDD.n70 26.38
R396 VDD.n73 VDD.n68 26.38
R397 VDD.n73 VDD.n72 26.38
R398 VDD.n126 VDD.n124 26.38
R399 VDD.n126 VDD.n123 26.38
R400 VDD.n126 VDD.n125 26.38
R401 VDD.n183 VDD.n181 26.38
R402 VDD.n183 VDD.n180 26.38
R403 VDD.n183 VDD.n182 26.38
R404 VDD.n258 VDD.n256 26.38
R405 VDD.n258 VDD.n255 26.38
R406 VDD.n258 VDD.n257 26.38
R407 VDD.n315 VDD.n313 26.38
R408 VDD.n315 VDD.n312 26.38
R409 VDD.n315 VDD.n314 26.38
R410 VDD.n372 VDD.n370 26.38
R411 VDD.n372 VDD.n369 26.38
R412 VDD.n372 VDD.n371 26.38
R413 VDD.n447 VDD.n445 26.38
R414 VDD.n447 VDD.n444 26.38
R415 VDD.n447 VDD.n446 26.38
R416 VDD.n522 VDD.n520 26.38
R417 VDD.n522 VDD.n519 26.38
R418 VDD.n522 VDD.n521 26.38
R419 VDD.n579 VDD.n577 26.38
R420 VDD.n579 VDD.n576 26.38
R421 VDD.n579 VDD.n578 26.38
R422 VDD.n654 VDD.n652 26.38
R423 VDD.n654 VDD.n651 26.38
R424 VDD.n654 VDD.n653 26.38
R425 VDD.n1360 VDD.n1358 26.38
R426 VDD.n1360 VDD.n1357 26.38
R427 VDD.n1360 VDD.n1359 26.38
R428 VDD.n1303 VDD.n1301 26.38
R429 VDD.n1303 VDD.n1300 26.38
R430 VDD.n1303 VDD.n1302 26.38
R431 VDD.n1228 VDD.n1226 26.38
R432 VDD.n1228 VDD.n1225 26.38
R433 VDD.n1228 VDD.n1227 26.38
R434 VDD.n1153 VDD.n1151 26.38
R435 VDD.n1153 VDD.n1150 26.38
R436 VDD.n1153 VDD.n1152 26.38
R437 VDD.n1096 VDD.n1094 26.38
R438 VDD.n1096 VDD.n1093 26.38
R439 VDD.n1096 VDD.n1095 26.38
R440 VDD.n1021 VDD.n1019 26.38
R441 VDD.n1021 VDD.n1018 26.38
R442 VDD.n1021 VDD.n1020 26.38
R443 VDD.n964 VDD.n962 26.38
R444 VDD.n964 VDD.n961 26.38
R445 VDD.n964 VDD.n963 26.38
R446 VDD.n907 VDD.n905 26.38
R447 VDD.n907 VDD.n904 26.38
R448 VDD.n907 VDD.n906 26.38
R449 VDD.n832 VDD.n830 26.38
R450 VDD.n832 VDD.n829 26.38
R451 VDD.n832 VDD.n831 26.38
R452 VDD.n699 VDD.n697 26.38
R453 VDD.n699 VDD.n696 26.38
R454 VDD.n699 VDD.n698 26.38
R455 VDD.n757 VDD.n756 26.38
R456 VDD.n757 VDD.n752 26.38
R457 VDD.n757 VDD.n750 26.38
R458 VDD.n757 VDD.n749 26.38
R459 VDD.n702 VDD.n694 22.915
R460 VDD.n23 VDD.n14 22.915
R461 VDD.n28 0<��� 20.457
R462 VDD.n93 0<��� 20.457
R463 VDD.n136  20.457
R464 VDD.n268  20.457
R465 VDD.n325  20.457
R466 VDD.n532  20.457
R467 VDD.n664 0<��� 20.457
R468 VDD.n1326 0<��� 20.457
R469 VDD.n1119  20.457
R470 VDD.n987 0<��� 20.457
R471 VDD.n930  20.457
R472 VDD.n722 0<��� 20.457
R473 VDD.n39  17.9
R474 VDD.n82  17.9
R475 VDD.n149 0<��� 17.9
R476 VDD.n281 0<��� 17.9
R477 VDD.n338 0<��� 17.9
R478 VDD.n545  17.9
R479 VDD.n677  17.9
R480 VDD.n1313  17.9
R481 VDD.n1106 0<��� 17.9
R482 VDD.n974  17.9
R483 VDD.n917  17.9
R484 VDD.n709 0<��� 17.9
R485 VDD.n200  15.343
R486 VDD.n389 0<��� 15.343
R487 VDD.n464  15.343
R488 VDD.n596  15.343
R489 VDD.n1260  15.343
R490 VDD.n1185  15.343
R491 VDD.n1053  15.343
R492 VDD.n864 0<��� 15.343
R493 VDD.n789 0<��� 15.343
R494 VDD.n694 VDD.n692 14.864
R495 VDD.n692 VDD.n690 14.864
R496 VDD.n690 VDD.n688 14.864
R497 VDD.n688 VDD.n686 14.864
R498 VDD.n686 VDD.n684 14.864
R499 VDD.n825 VDD.n823 14.864
R500 VDD.n823 VDD.n821 14.864
R501 VDD.n821 VDD.n819 14.864
R502 VDD.n819 VDD.n817 14.864
R503 VDD.n817 VDD.n815 14.864
R504 VDD.n900 VDD.n898 14.864
R505 VDD.n898 VDD.n896 14.864
R506 VDD.n896 VDD.n894 14.864
R507 VDD.n894 VDD.n892 14.864
R508 VDD.n892 VDD.n890 14.864
R509 VDD.n957 VDD.n955 14.864
R510 VDD.n955 VDD.n953 14.864
R511 VDD.n953 VDD.n951 14.864
R512 VDD.n951 VDD.n949 14.864
R513 VDD.n949 VDD.n947 14.864
R514 VDD.n1014 VDD.n1012 14.864
R515 VDD.n1012 VDD.n1010 14.864
R516 VDD.n1010 VDD.n1008 14.864
R517 VDD.n1008 VDD.n1006 14.864
R518 VDD.n1006 VDD.n1004 14.864
R519 VDD.n1089 VDD.n1087 14.864
R520 VDD.n1087 VDD.n1085 14.864
R521 VDD.n1085 VDD.n1083 14.864
R522 VDD.n1083 VDD.n1081 14.864
R523 VDD.n1081 VDD.n1079 14.864
R524 VDD.n1146 VDD.n1144 14.864
R525 VDD.n1144 VDD.n1142 14.864
R526 VDD.n1142 VDD.n1140 14.864
R527 VDD.n1140 VDD.n1138 14.864
R528 VDD.n1138 VDD.n1136 14.864
R529 VDD.n1221 VDD.n1219 14.864
R530 VDD.n1219 VDD.n1217 14.864
R531 VDD.n1217 VDD.n1215 14.864
R532 VDD.n1215 VDD.n1213 14.864
R533 VDD.n1213 VDD.n1211 14.864
R534 VDD.n1296 VDD.n1294 14.864
R535 VDD.n1294 VDD.n1292 14.864
R536 VDD.n1292 VDD.n1290 14.864
R537 VDD.n1290 VDD.n1288 14.864
R538 VDD.n1288 VDD.n1286 14.864
R539 VDD.n1353 VDD.n1351 14.864
R540 VDD.n1351 VDD.n1349 14.864
R541 VDD.n1349 VDD.n1347 14.864
R542 VDD.n1347 VDD.n1345 14.864
R543 VDD.n1345 VDD.n1343 14.864
R544 VDD.n647 VDD.n645 14.864
R545 VDD.n645 VDD.n643 14.864
R546 VDD.n643 VDD.n641 14.864
R547 VDD.n641 VDD.n639 14.864
R548 VDD.n639 VDD.n637 14.864
R549 VDD.n572 VDD.n570 14.864
R550 VDD.n570 VDD.n568 14.864
R551 VDD.n568 VDD.n566 14.864
R552 VDD.n566 VDD.n564 14.864
R553 VDD.n564 VDD.n562 14.864
R554 VDD.n515 VDD.n513 14.864
R555 VDD.n513 VDD.n511 14.864
R556 VDD.n511 VDD.n509 14.864
R557 VDD.n509 VDD.n507 14.864
R558 VDD.n507 VDD.n505 14.864
R559 VDD.n440 VDD.n438 14.864
R560 VDD.n438 VDD.n436 14.864
R561 VDD.n436 VDD.n434 14.864
R562 VDD.n434 VDD.n432 14.864
R563 VDD.n432 VDD.n430 14.864
R564 VDD.n365 VDD.n363 14.864
R565 VDD.n363 VDD.n361 14.864
R566 VDD.n361 VDD.n359 14.864
R567 VDD.n359 VDD.n357 14.864
R568 VDD.n357 VDD.n355 14.864
R569 VDD.n308 VDD.n306 14.864
R570 VDD.n306 VDD.n304 14.864
R571 VDD.n304 VDD.n302 14.864
R572 VDD.n302 VDD.n300 14.864
R573 VDD.n300 VDD.n298 14.864
R574 VDD.n251 VDD.n249 14.864
R575 VDD.n249 VDD.n247 14.864
R576 VDD.n247 VDD.n245 14.864
R577 VDD.n245 VDD.n243 14.864
R578 VDD.n243 VDD.n241 14.864
R579 VDD.n176 VDD.n174 14.864
R580 VDD.n174 VDD.n172 14.864
R581 VDD.n172 VDD.n170 14.864
R582 VDD.n170 VDD.n168 14.864
R583 VDD.n168 VDD.n166 14.864
R584 VDD.n119 VDD.n117 14.864
R585 VDD.n117 VDD.n115 14.864
R586 VDD.n115 VDD.n113 14.864
R587 VDD.n113 VDD.n111 14.864
R588 VDD.n111 VDD.n109 14.864
R589 VDD.n62 VDD.n60 14.864
R590 VDD.n60 VDD.n58 14.864
R591 VDD.n58 VDD.n56 14.864
R592 VDD.n56 VDD.n54 14.864
R593 VDD.n54 VDD.n52 14.864
R594 VDD.n52 VDD.n51 14.864
R595 VDD.n746 VDD.n744 14.864
R596 VDD.n744 VDD.n742 14.864
R597 VDD.n742 VDD.n740 14.864
R598 VDD.n740 VDD.n738 14.864
R599 VDD.n738 VDD.n736 14.864
R600 VDD.n736 VDD.n735 14.864
R601 VDD.n14 VDD.n13 14.864
R602 VDD.n13 VDD.n11 14.864
R603 VDD.n11 VDD.n9 14.864
R604 VDD.n9 VDD.n7 14.864
R605 VDD.n7 VDD.n5 14.864
R606 VDD.n76 VDD.n63 14.864
R607 VDD.n129 VDD.n120 14.864
R608 VDD.n186 VDD.n177 14.864
R609 VDD.n261 VDD.n252 14.864
R610 VDD.n318 VDD.n309 14.864
R611 VDD.n375 VDD.n366 14.864
R612 VDD.n450 VDD.n441 14.864
R613 VDD.n525 VDD.n516 14.864
R614 VDD.n582 VDD.n573 14.864
R615 VDD.n657 VDD.n648 14.864
R616 VDD.n1363 VDD.n1354 14.864
R617 VDD.n1306 VDD.n1297 14.864
R618 VDD.n1231 VDD.n1222 14.864
R619 VDD.n1156 VDD.n1147 14.864
R620 VDD.n1099 VDD.n1090 14.864
R621 VDD.n1024 VDD.n1015 14.864
R622 VDD.n967 VDD.n958 14.864
R623 VDD.n910 VDD.n901 14.864
R624 VDD.n835 VDD.n826 14.864
R625 VDD.n760 VDD.n747 14.864
R626 VDD.n717 VDD.t173 14.282
R627 VDD.n717 VDD.t80 14.282
R628 VDD.n775 VDD.t102 14.282
R629 VDD.n775 VDD.t132 14.282
R630 VDD.n791 VDD.t92 14.282
R631 VDD.n791 VDD.t34 14.282
R632 VDD.n850 VDD.t157 14.282
R633 VDD.n850 VDD.t118 14.282
R634 VDD.n866 VDD.t114 14.282
R635 VDD.n866 VDD.t147 14.282
R636 VDD.n925 VDD.t100 14.282
R637 VDD.n925 VDD.t60 14.282
R638 VDD.n982 VDD.t110 14.282
R639 VDD.n982 VDD.t171 14.282
R640 VDD.n1039 VDD.t145 14.282
R641 VDD.n1039 VDD.t169 14.282
R642 VDD.n1055 VDD.t128 14.282
R643 VDD.n1055 VDD.t161 14.282
R644 VDD.n1114 VDD.t52 14.282
R645 VDD.n1114 VDD.t112 14.282
R646 VDD.n1171 VDD.t36 14.282
R647 VDD.n1171 VDD.t134 14.282
R648 VDD.n1187 VDD.t90 14.282
R649 VDD.n1187 VDD.t186 14.282
R650 VDD.n1246 VDD.t155 14.282
R651 VDD.n1246 VDD.t44 14.282
R652 VDD.n1262 VDD.t66 14.282
R653 VDD.n1262 VDD.t122 14.282
R654 VDD.n1321 VDD.t11 14.282
R655 VDD.n1321 VDD.t195 14.282
R656 VDD.n668 VDD.t18 14.282
R657 VDD.n668 VDD.t104 14.282
R658 VDD.n610 VDD.t167 14.282
R659 VDD.n610 VDD.t9 14.282
R660 VDD.n598 VDD.t32 14.282
R661 VDD.n598 VDD.t149 14.282
R662 VDD.n536 VDD.t1 14.282
R663 VDD.n536 VDD.t137 14.282
R664 VDD.n478 VDD.t159 14.282
R665 VDD.n478 VDD.t108 14.282
R666 VDD.n466 VDD.t141 14.282
R667 VDD.n466 VDD.t181 14.282
R668 VDD.n403 VDD.t151 14.282
R669 VDD.n403 VDD.t96 14.282
R670 VDD.n391 VDD.t56 14.282
R671 VDD.n391 VDD.t163 14.282
R672 VDD.n329 VDD.t50 14.282
R673 VDD.n329 VDD.t48 14.282
R674 VDD.n272 VDD.t116 14.282
R675 VDD.n272 VDD.t184 14.282
R676 VDD.n214 VDD.t153 14.282
R677 VDD.n214 VDD.t70 14.282
R678 VDD.n202 VDD.t42 14.282
R679 VDD.n202 VDD.t165 14.282
R680 VDD.n140 VDD.t29 14.282
R681 VDD.n140 VDD.t16 14.282
R682 VDD.n216  12.786
R683 VDD.n405 0<��� 12.786
R684 VDD.n480 0<��� 12.786
R685 VDD.n612 ���V 12.786
R686 VDD.n1248  12.786
R687 VDD.n1173  12.786
R688 VDD.n1041 0<��� 12.786
R689 VDD.n852 0<��� 12.786
R690 VDD.n777  12.786
R691 VDD.n143 VDD.n141 9.083
R692 VDD.n275 VDD.n273 9.083
R693 VDD.n332 VDD.n330 9.083
R694 VDD.n539 VDD.n537 9.083
R695 VDD.n671 VDD.n669 9.083
R696 VDD.n1324 VDD.n1322 9.083
R697 VDD.n1117 VDD.n1115 9.083
R698 VDD.n985 VDD.n983 9.083
R699 VDD.n928 VDD.n926 9.083
R700 VDD.n720 VDD.n718 9.083
R701 VDD.n23 VDD.n22 8.855
R702 VDD.n22 VDD.n21 8.855
R703 VDD.n26 VDD.n25 8.855
R704 VDD.n25 VDD.n24 8.855
R705 VDD.n30 VDD.n29 8.855
R706 VDD.n29 VDD.n28 8.855
R707 VDD.n33 VDD.n32 8.855
R708 VDD.n32  8.855
R709 VDD.n37 VDD.n36 8.855
R710 VDD.n36 VDD.n35 8.855
R711 VDD.n41 VDD.n40 8.855
R712 VDD.n40 VDD.n39 8.855
R713 VDD.n45 VDD.n44 8.855
R714 VDD.n44 VDD.n43 8.855
R715 VDD.n49 VDD.n48 8.855
R716 VDD.n48 VDD.n47 8.855
R717 VDD.n76 VDD.n75 8.855
R718 VDD.n75 VDD.n74 8.855
R719 VDD.n80 VDD.n79 8.855
R720 VDD.n79 VDD.n78 8.855
R721 VDD.n84 VDD.n83 8.855
R722 VDD.n83 VDD.n82 8.855
R723 VDD.n88 VDD.n87 8.855
R724 VDD.n87 VDD.n86 8.855
R725 VDD.n91 VDD.n90 8.855
R726 VDD.n90  8.855
R727 VDD.n95 VDD.n94 8.855
R728 VDD.n94 VDD.n93 8.855
R729 VDD.n99 VDD.n98 8.855
R730 VDD.n98 VDD.n97 8.855
R731 VDD.n103 VDD.n102 8.855
R732 VDD.n102 VDD.n101 8.855
R733 VDD.n129 VDD.n128 8.855
R734 VDD.n128 VDD.n127 8.855
R735 VDD.n134 VDD.n133 8.855
R736 VDD.n133 VDD.n132 8.855
R737 VDD.n138 VDD.n137 8.855
R738 VDD.n137 VDD.n136 8.855
R739 VDD.n143 VDD.n142 8.855
R740 VDD.n142 0<��� 8.855
R741 VDD.n147 VDD.n146 8.855
R742 VDD.n146 VDD.n145 8.855
R743 VDD.n151 VDD.n150 8.855
R744 VDD.n150 VDD.n149 8.855
R745 VDD.n156 VDD.n155 8.855
R746 VDD.n155 VDD.n154 8.855
R747 VDD.n160 VDD.n159 8.855
R748 VDD.n159 VDD.n158 8.855
R749 VDD.n186 VDD.n185 8.855
R750 VDD.n185 VDD.n184 8.855
R751 VDD.n190 VDD.n189 8.855
R752 VDD.n189 VDD.n188 8.855
R753 VDD.n194 VDD.n193 8.855
R754 VDD.n193 VDD.n192 8.855
R755 VDD.n198 VDD.n197 8.855
R756 VDD.n197 VDD.n196 8.855
R757 VDD.n204 VDD.n201 8.855
R758 VDD.n201 VDD.n200 8.855
R759 VDD.n208 VDD.n207 8.855
R760 VDD.n207 VDD.n206 8.855
R761 VDD.n212 VDD.n211 8.855
R762 VDD.n211 VDD.n210 8.855
R763 VDD.n218 VDD.n217 8.855
R764 VDD.n217 VDD.n216 8.855
R765 VDD.n222 VDD.n221 8.855
R766 VDD.n221 VDD.n220 8.855
R767 VDD.n227 VDD.n226 8.855
R768 VDD.n226 VDD.n225 8.855
R769 VDD.n231 VDD.n230 8.855
R770 VDD.n230 VDD.n229 8.855
R771 VDD.n235 VDD.n234 8.855
R772 VDD.n234 VDD.n233 8.855
R773 VDD.n261 VDD.n260 8.855
R774 VDD.n260 VDD.n259 8.855
R775 VDD.n266 VDD.n265 8.855
R776 VDD.n265 VDD.n264 8.855
R777 VDD.n270 VDD.n269 8.855
R778 VDD.n269 VDD.n268 8.855
R779 VDD.n275 VDD.n274 8.855
R780 VDD.n274 0<��� 8.855
R781 VDD.n279 VDD.n278 8.855
R782 VDD.n278 VDD.n277 8.855
R783 VDD.n283 VDD.n282 8.855
R784 VDD.n282 VDD.n281 8.855
R785 VDD.n288 VDD.n287 8.855
R786 VDD.n287 VDD.n286 8.855
R787 VDD.n292 VDD.n291 8.855
R788 VDD.n291 VDD.n290 8.855
R789 VDD.n318 VDD.n317 8.855
R790 VDD.n317 VDD.n316 8.855
R791 VDD.n323 VDD.n322 8.855
R792 VDD.n322 VDD.n321 8.855
R793 VDD.n327 VDD.n326 8.855
R794 VDD.n326 VDD.n325 8.855
R795 VDD.n332 VDD.n331 8.855
R796 VDD.n331  8.855
R797 VDD.n336 VDD.n335 8.855
R798 VDD.n335 VDD.n334 8.855
R799 VDD.n340 VDD.n339 8.855
R800 VDD.n339 VDD.n338 8.855
R801 VDD.n345 VDD.n344 8.855
R802 VDD.n344 VDD.n343 8.855
R803 VDD.n349 VDD.n348 8.855
R804 VDD.n348 VDD.n347 8.855
R805 VDD.n375 VDD.n374 8.855
R806 VDD.n374 VDD.n373 8.855
R807 VDD.n379 VDD.n378 8.855
R808 VDD.n378 VDD.n377 8.855
R809 VDD.n383 VDD.n382 8.855
R810 VDD.n382 VDD.n381 8.855
R811 VDD.n387 VDD.n386 8.855
R812 VDD.n386 VDD.n385 8.855
R813 VDD.n393 VDD.n390 8.855
R814 VDD.n390 VDD.n389 8.855
R815 VDD.n397 VDD.n396 8.855
R816 VDD.n396 VDD.n395 8.855
R817 VDD.n401 VDD.n400 8.855
R818 VDD.n400 VDD.n399 8.855
R819 VDD.n407 VDD.n406 8.855
R820 VDD.n406 VDD.n405 8.855
R821 VDD.n411 VDD.n410 8.855
R822 VDD.n410 VDD.n409 8.855
R823 VDD.n416 VDD.n415 8.855
R824 VDD.n415 VDD.n414 8.855
R825 VDD.n420 VDD.n419 8.855
R826 VDD.n419 VDD.n418 8.855
R827 VDD.n424 VDD.n423 8.855
R828 VDD.n423 VDD.n422 8.855
R829 VDD.n450 VDD.n449 8.855
R830 VDD.n449 VDD.n448 8.855
R831 VDD.n454 VDD.n453 8.855
R832 VDD.n453 VDD.n452 8.855
R833 VDD.n458 VDD.n457 8.855
R834 VDD.n457 VDD.n456 8.855
R835 VDD.n462 VDD.n461 8.855
R836 VDD.n461 VDD.n460 8.855
R837 VDD.n468 VDD.n465 8.855
R838 VDD.n465 VDD.n464 8.855
R839 VDD.n472 VDD.n471 8.855
R840 VDD.n471 VDD.n470 8.855
R841 VDD.n476 VDD.n475 8.855
R842 VDD.n475 VDD.n474 8.855
R843 VDD.n482 VDD.n481 8.855
R844 VDD.n481 VDD.n480 8.855
R845 VDD.n486 VDD.n485 8.855
R846 VDD.n485 VDD.n484 8.855
R847 VDD.n491 VDD.n490 8.855
R848 VDD.n490 VDD.n489 8.855
R849 VDD.n495 VDD.n494 8.855
R850 VDD.n494 VDD.n493 8.855
R851 VDD.n499 VDD.n498 8.855
R852 VDD.n498 VDD.n497 8.855
R853 VDD.n525 VDD.n524 8.855
R854 VDD.n524 VDD.n523 8.855
R855 VDD.n530 VDD.n529 8.855
R856 VDD.n529 VDD.n528 8.855
R857 VDD.n534 VDD.n533 8.855
R858 VDD.n533 VDD.n532 8.855
R859 VDD.n539 VDD.n538 8.855
R860 VDD.n538 0<��� 8.855
R861 VDD.n543 VDD.n542 8.855
R862 VDD.n542 VDD.n541 8.855
R863 VDD.n547 VDD.n546 8.855
R864 VDD.n546 VDD.n545 8.855
R865 VDD.n552 VDD.n551 8.855
R866 VDD.n551 VDD.n550 8.855
R867 VDD.n556 VDD.n555 8.855
R868 VDD.n555 VDD.n554 8.855
R869 VDD.n582 VDD.n581 8.855
R870 VDD.n581 VDD.n580 8.855
R871 VDD.n586 VDD.n585 8.855
R872 VDD.n585 VDD.n584 8.855
R873 VDD.n590 VDD.n589 8.855
R874 VDD.n589 VDD.n588 8.855
R875 VDD.n594 VDD.n593 8.855
R876 VDD.n593 VDD.n592 8.855
R877 VDD.n600 VDD.n597 8.855
R878 VDD.n597 VDD.n596 8.855
R879 VDD.n604 VDD.n603 8.855
R880 VDD.n603 VDD.n602 8.855
R881 VDD.n608 VDD.n607 8.855
R882 VDD.n607 VDD.n606 8.855
R883 VDD.n614 VDD.n613 8.855
R884 VDD.n613 VDD.n612 8.855
R885 VDD.n618 VDD.n617 8.855
R886 VDD.n617 VDD.n616 8.855
R887 VDD.n623 VDD.n622 8.855
R888 VDD.n622 VDD.n621 8.855
R889 VDD.n627 VDD.n626 8.855
R890 VDD.n626 VDD.n625 8.855
R891 VDD.n631 VDD.n630 8.855
R892 VDD.n630 VDD.n629 8.855
R893 VDD.n657 VDD.n656 8.855
R894 VDD.n656 VDD.n655 8.855
R895 VDD.n662 VDD.n661 8.855
R896 VDD.n661 VDD.n660 8.855
R897 VDD.n666 VDD.n665 8.855
R898 VDD.n665 VDD.n664 8.855
R899 VDD.n671 VDD.n670 8.855
R900 VDD.n670 0<��� 8.855
R901 VDD.n675 VDD.n674 8.855
R902 VDD.n674 VDD.n673 8.855
R903 VDD.n679 VDD.n678 8.855
R904 VDD.n678 VDD.n677 8.855
R905 VDD.n1368 VDD.n1367 8.855
R906 VDD.n1367 VDD.n1366 8.855
R907 VDD.n1363 VDD.n1362 8.855
R908 VDD.n1362 VDD.n1361 8.855
R909 VDD.n1337 VDD.n1336 8.855
R910 VDD.n1336 VDD.n1335 8.855
R911 VDD.n1333 VDD.n1332 8.855
R912 VDD.n1332 VDD.n1331 8.855
R913 VDD.n1328 VDD.n1327 8.855
R914 VDD.n1327 VDD.n1326 8.855
R915 VDD.n1324 VDD.n1323 8.855
R916 VDD.n1323  8.855
R917 VDD.n1319 VDD.n1318 8.855
R918 VDD.n1318 VDD.n1317 8.855
R919 VDD.n1315 VDD.n1314 8.855
R920 VDD.n1314 VDD.n1313 8.855
R921 VDD.n1311 VDD.n1310 8.855
R922 VDD.n1310 VDD.n1309 8.855
R923 VDD.n1306 VDD.n1305 8.855
R924 VDD.n1305 VDD.n1304 8.855
R925 VDD.n1280 VDD.n1279 8.855
R926 VDD.n1279 VDD.n1278 8.855
R927 VDD.n1276 VDD.n1275 8.855
R928 VDD.n1275 VDD.n1274 8.855
R929 VDD.n1272 VDD.n1271 8.855
R930 VDD.n1271 VDD.n1270 8.855
R931 VDD.n1268 VDD.n1267 8.855
R932 VDD.n1267 VDD.n1266 8.855
R933 VDD.n1264 VDD.n1261 8.855
R934 VDD.n1261 VDD.n1260 8.855
R935 VDD.n1258 VDD.n1257 8.855
R936 VDD.n1257 VDD.n1256 8.855
R937 VDD.n1254 VDD.n1253 8.855
R938 VDD.n1253 VDD.n1252 8.855
R939 VDD.n1250 VDD.n1249 8.855
R940 VDD.n1249 VDD.n1248 8.855
R941 VDD.n1244 VDD.n1243 8.855
R942 VDD.n1243 VDD.n1242 8.855
R943 VDD.n1240 VDD.n1239 8.855
R944 VDD.n1239 VDD.n1238 8.855
R945 VDD.n1235 VDD.n1234 8.855
R946 VDD.n1234 VDD.n1233 8.855
R947 VDD.n1231 VDD.n1230 8.855
R948 VDD.n1230 VDD.n1229 8.855
R949 VDD.n1205 VDD.n1204 8.855
R950 VDD.n1204 VDD.n1203 8.855
R951 VDD.n1201 VDD.n1200 8.855
R952 VDD.n1200 VDD.n1199 8.855
R953 VDD.n1197 VDD.n1196 8.855
R954 VDD.n1196 VDD.n1195 8.855
R955 VDD.n1193 VDD.n1192 8.855
R956 VDD.n1192 VDD.n1191 8.855
R957 VDD.n1189 VDD.n1186 8.855
R958 VDD.n1186 VDD.n1185 8.855
R959 VDD.n1183 VDD.n1182 8.855
R960 VDD.n1182 VDD.n1181 8.855
R961 VDD.n1179 VDD.n1178 8.855
R962 VDD.n1178 VDD.n1177 8.855
R963 VDD.n1175 VDD.n1174 8.855
R964 VDD.n1174 VDD.n1173 8.855
R965 VDD.n1169 VDD.n1168 8.855
R966 VDD.n1168 VDD.n1167 8.855
R967 VDD.n1165 VDD.n1164 8.855
R968 VDD.n1164 VDD.n1163 8.855
R969 VDD.n1160 VDD.n1159 8.855
R970 VDD.n1159 VDD.n1158 8.855
R971 VDD.n1156 VDD.n1155 8.855
R972 VDD.n1155 VDD.n1154 8.855
R973 VDD.n1130 VDD.n1129 8.855
R974 VDD.n1129 VDD.n1128 8.855
R975 VDD.n1126 VDD.n1125 8.855
R976 VDD.n1125 VDD.n1124 8.855
R977 VDD.n1121 VDD.n1120 8.855
R978 VDD.n1120 VDD.n1119 8.855
R979 VDD.n1117 VDD.n1116 8.855
R980 VDD.n1116 0<��� 8.855
R981 VDD.n1112 VDD.n1111 8.855
R982 VDD.n1111 VDD.n1110 8.855
R983 VDD.n1108 VDD.n1107 8.855
R984 VDD.n1107 VDD.n1106 8.855
R985 VDD.n1104 VDD.n1103 8.855
R986 VDD.n1103 VDD.n1102 8.855
R987 VDD.n1099 VDD.n1098 8.855
R988 VDD.n1098 VDD.n1097 8.855
R989 VDD.n1073 VDD.n1072 8.855
R990 VDD.n1072 VDD.n1071 8.855
R991 VDD.n1069 VDD.n1068 8.855
R992 VDD.n1068 VDD.n1067 8.855
R993 VDD.n1065 VDD.n1064 8.855
R994 VDD.n1064 VDD.n1063 8.855
R995 VDD.n1061 VDD.n1060 8.855
R996 VDD.n1060 VDD.n1059 8.855
R997 VDD.n1057 VDD.n1054 8.855
R998 VDD.n1054 VDD.n1053 8.855
R999 VDD.n1051 VDD.n1050 8.855
R1000 VDD.n1050 VDD.n1049 8.855
R1001 VDD.n1047 VDD.n1046 8.855
R1002 VDD.n1046 VDD.n1045 8.855
R1003 VDD.n1043 VDD.n1042 8.855
R1004 VDD.n1042 VDD.n1041 8.855
R1005 VDD.n1037 VDD.n1036 8.855
R1006 VDD.n1036 VDD.n1035 8.855
R1007 VDD.n1033 VDD.n1032 8.855
R1008 VDD.n1032 VDD.n1031 8.855
R1009 VDD.n1028 VDD.n1027 8.855
R1010 VDD.n1027 VDD.n1026 8.855
R1011 VDD.n1024 VDD.n1023 8.855
R1012 VDD.n1023 VDD.n1022 8.855
R1013 VDD.n998 VDD.n997 8.855
R1014 VDD.n997 VDD.n996 8.855
R1015 VDD.n994 VDD.n993 8.855
R1016 VDD.n993 VDD.n992 8.855
R1017 VDD.n989 VDD.n988 8.855
R1018 VDD.n988 VDD.n987 8.855
R1019 VDD.n985 VDD.n984 8.855
R1020 VDD.n984 0<��� 8.855
R1021 VDD.n980 VDD.n979 8.855
R1022 VDD.n979 VDD.n978 8.855
R1023 VDD.n976 VDD.n975 8.855
R1024 VDD.n975 VDD.n974 8.855
R1025 VDD.n972 VDD.n971 8.855
R1026 VDD.n971 VDD.n970 8.855
R1027 VDD.n967 VDD.n966 8.855
R1028 VDD.n966 VDD.n965 8.855
R1029 VDD.n941 VDD.n940 8.855
R1030 VDD.n940 VDD.n939 8.855
R1031 VDD.n937 VDD.n936 8.855
R1032 VDD.n936 VDD.n935 8.855
R1033 VDD.n932 VDD.n931 8.855
R1034 VDD.n931 VDD.n930 8.855
R1035 VDD.n928 VDD.n927 8.855
R1036 VDD.n927  8.855
R1037 VDD.n923 VDD.n922 8.855
R1038 VDD.n922 VDD.n921 8.855
R1039 VDD.n919 VDD.n918 8.855
R1040 VDD.n918 VDD.n917 8.855
R1041 VDD.n915 VDD.n914 8.855
R1042 VDD.n914 VDD.n913 8.855
R1043 VDD.n910 VDD.n909 8.855
R1044 VDD.n909 VDD.n908 8.855
R1045 VDD.n884 VDD.n883 8.855
R1046 VDD.n883 VDD.n882 8.855
R1047 VDD.n880 VDD.n879 8.855
R1048 VDD.n879 VDD.n878 8.855
R1049 VDD.n876 VDD.n875 8.855
R1050 VDD.n875 VDD.n874 8.855
R1051 VDD.n872 VDD.n871 8.855
R1052 VDD.n871 VDD.n870 8.855
R1053 VDD.n868 VDD.n865 8.855
R1054 VDD.n865 VDD.n864 8.855
R1055 VDD.n862 VDD.n861 8.855
R1056 VDD.n861 VDD.n860 8.855
R1057 VDD.n858 VDD.n857 8.855
R1058 VDD.n857 VDD.n856 8.855
R1059 VDD.n854 VDD.n853 8.855
R1060 VDD.n853 VDD.n852 8.855
R1061 VDD.n848 VDD.n847 8.855
R1062 VDD.n847 VDD.n846 8.855
R1063 VDD.n844 VDD.n843 8.855
R1064 VDD.n843 VDD.n842 8.855
R1065 VDD.n839 VDD.n838 8.855
R1066 VDD.n838 VDD.n837 8.855
R1067 VDD.n835 VDD.n834 8.855
R1068 VDD.n834 VDD.n833 8.855
R1069 VDD.n809 VDD.n808 8.855
R1070 VDD.n808 VDD.n807 8.855
R1071 VDD.n805 VDD.n804 8.855
R1072 VDD.n804 VDD.n803 8.855
R1073 VDD.n801 VDD.n800 8.855
R1074 VDD.n800 VDD.n799 8.855
R1075 VDD.n797 VDD.n796 8.855
R1076 VDD.n796 VDD.n795 8.855
R1077 VDD.n793 VDD.n790 8.855
R1078 VDD.n790 VDD.n789 8.855
R1079 VDD.n787 VDD.n786 8.855
R1080 VDD.n786 VDD.n785 8.855
R1081 VDD.n783 VDD.n782 8.855
R1082 VDD.n782 VDD.n781 8.855
R1083 VDD.n779 VDD.n778 8.855
R1084 VDD.n778 VDD.n777 8.855
R1085 VDD.n773 VDD.n772 8.855
R1086 VDD.n772 VDD.n771 8.855
R1087 VDD.n769 VDD.n768 8.855
R1088 VDD.n768 VDD.n767 8.855
R1089 VDD.n764 VDD.n763 8.855
R1090 VDD.n763 VDD.n762 8.855
R1091 VDD.n760 VDD.n759 8.855
R1092 VDD.n759 VDD.n758 8.855
R1093 VDD.n733 VDD.n732 8.855
R1094 VDD.n732 VDD.n731 8.855
R1095 VDD.n729 VDD.n728 8.855
R1096 VDD.n728 VDD.n727 8.855
R1097 VDD.n724 VDD.n723 8.855
R1098 VDD.n723 VDD.n722 8.855
R1099 VDD.n720 VDD.n719 8.855
R1100 VDD.n719  8.855
R1101 VDD.n715 VDD.n714 8.855
R1102 VDD.n714 VDD.n713 8.855
R1103 VDD.n711 VDD.n710 8.855
R1104 VDD.n710 VDD.n709 8.855
R1105 VDD.n707 VDD.n706 8.855
R1106 VDD.n706 VDD.n705 8.855
R1107 VDD.n702 VDD.n701 8.855
R1108 VDD.n701 VDD.n700 8.855
R1109 VDD.n826 VDD.n825 8.051
R1110 VDD.n901 VDD.n900 8.051
R1111 VDD.n958 VDD.n957 8.051
R1112 VDD.n1015 VDD.n1014 8.051
R1113 VDD.n1090 VDD.n1089 8.051
R1114 VDD.n1147 VDD.n1146 8.051
R1115 VDD.n1222 VDD.n1221 8.051
R1116 VDD.n1297 VDD.n1296 8.051
R1117 VDD.n1354 VDD.n1353 8.051
R1118 VDD.n648 VDD.n647 8.051
R1119 VDD.n573 VDD.n572 8.051
R1120 VDD.n516 VDD.n515 8.051
R1121 VDD.n441 VDD.n440 8.051
R1122 VDD.n366 VDD.n365 8.051
R1123 VDD.n309 VDD.n308 8.051
R1124 VDD.n252 VDD.n251 8.051
R1125 VDD.n177 VDD.n176 8.051
R1126 VDD.n120 VDD.n119 8.051
R1127 VDD.n63 VDD.n62 8.051
R1128 VDD.n747 VDD.n746 8.051
R1129 VDD.n210 0<��� 7.671
R1130 VDD.n399 0<��� 7.671
R1131 VDD.n474 0<��� 7.671
R1132 VDD.n606  7.671
R1133 VDD.n1252 0<��� 7.671
R1134 VDD.n1177 0<��� 7.671
R1135 VDD.n1045 0<��� 7.671
R1136 VDD.n856  7.671
R1137 VDD.n781  7.671
R1138 VDD.n218 VDD.n215 7.019
R1139 VDD.n407 VDD.n404 7.019
R1140 VDD.n482 VDD.n479 7.019
R1141 VDD.n614 VDD.n611 7.019
R1142 VDD.n1250 VDD.n1247 7.019
R1143 VDD.n1175 VDD.n1172 7.019
R1144 VDD.n1043 VDD.n1040 7.019
R1145 VDD.n854 VDD.n851 7.019
R1146 VDD.n779 VDD.n776 7.019
R1147 VDD.n204 VDD.n203 6.606
R1148 VDD.n393 VDD.n392 6.606
R1149 VDD.n468 VDD.n467 6.606
R1150 VDD.n600 VDD.n599 6.606
R1151 VDD.n1264 VDD.n1263 6.606
R1152 VDD.n1189 VDD.n1188 6.606
R1153 VDD.n1057 VDD.n1056 6.606
R1154 VDD.n868 VDD.n867 6.606
R1155 VDD.n793 VDD.n792 6.606
R1156 VDD.n206 0<��� 5.114
R1157 VDD.n395 0<��� 5.114
R1158 VDD.n470  5.114
R1159 VDD.n602 0<��� 5.114
R1160 VDD.n1256  5.114
R1161 VDD.n1181 0<��� 5.114
R1162 VDD.n1049 0<��� 5.114
R1163 VDD.n860 0<��� 5.114
R1164 VDD.n785 0<��� 5.114
R1165 VDD.n31 VDD.n30 4.65
R1166 VDD.n34 VDD.n33 4.65
R1167 VDD.n38 VDD.n37 4.65
R1168 VDD.n42 VDD.n41 4.65
R1169 VDD.n46 VDD.n45 4.65
R1170 VDD.n50 VDD.n49 4.65
R1171 VDD.n77 VDD.n76 4.65
R1172 VDD.n81 VDD.n80 4.65
R1173 VDD.n85 VDD.n84 4.65
R1174 VDD.n89 VDD.n88 4.65
R1175 VDD.n92 VDD.n91 4.65
R1176 VDD.n96 VDD.n95 4.65
R1177 VDD.n100 VDD.n99 4.65
R1178 VDD.n104 VDD.n103 4.65
R1179 VDD.n130 VDD.n129 4.65
R1180 VDD.n135 VDD.n134 4.65
R1181 VDD.n139 VDD.n138 4.65
R1182 VDD.n144 VDD.n143 4.65
R1183 VDD.n148 VDD.n147 4.65
R1184 VDD.n152 VDD.n151 4.65
R1185 VDD.n157 VDD.n156 4.65
R1186 VDD.n161 VDD.n160 4.65
R1187 VDD.n187 VDD.n186 4.65
R1188 VDD.n191 VDD.n190 4.65
R1189 VDD.n195 VDD.n194 4.65
R1190 VDD.n199 VDD.n198 4.65
R1191 VDD.n205 VDD.n204 4.65
R1192 VDD.n209 VDD.n208 4.65
R1193 VDD.n213 VDD.n212 4.65
R1194 VDD.n219 VDD.n218 4.65
R1195 VDD.n223 VDD.n222 4.65
R1196 VDD.n228 VDD.n227 4.65
R1197 VDD.n232 VDD.n231 4.65
R1198 VDD.n236 VDD.n235 4.65
R1199 VDD.n262 VDD.n261 4.65
R1200 VDD.n267 VDD.n266 4.65
R1201 VDD.n271 VDD.n270 4.65
R1202 VDD.n276 VDD.n275 4.65
R1203 VDD.n280 VDD.n279 4.65
R1204 VDD.n284 VDD.n283 4.65
R1205 VDD.n289 VDD.n288 4.65
R1206 VDD.n293 VDD.n292 4.65
R1207 VDD.n319 VDD.n318 4.65
R1208 VDD.n324 VDD.n323 4.65
R1209 VDD.n328 VDD.n327 4.65
R1210 VDD.n333 VDD.n332 4.65
R1211 VDD.n337 VDD.n336 4.65
R1212 VDD.n341 VDD.n340 4.65
R1213 VDD.n346 VDD.n345 4.65
R1214 VDD.n350 VDD.n349 4.65
R1215 VDD.n376 VDD.n375 4.65
R1216 VDD.n380 VDD.n379 4.65
R1217 VDD.n384 VDD.n383 4.65
R1218 VDD.n388 VDD.n387 4.65
R1219 VDD.n394 VDD.n393 4.65
R1220 VDD.n398 VDD.n397 4.65
R1221 VDD.n402 VDD.n401 4.65
R1222 VDD.n408 VDD.n407 4.65
R1223 VDD.n412 VDD.n411 4.65
R1224 VDD.n417 VDD.n416 4.65
R1225 VDD.n421 VDD.n420 4.65
R1226 VDD.n425 VDD.n424 4.65
R1227 VDD.n451 VDD.n450 4.65
R1228 VDD.n455 VDD.n454 4.65
R1229 VDD.n459 VDD.n458 4.65
R1230 VDD.n463 VDD.n462 4.65
R1231 VDD.n469 VDD.n468 4.65
R1232 VDD.n473 VDD.n472 4.65
R1233 VDD.n477 VDD.n476 4.65
R1234 VDD.n483 VDD.n482 4.65
R1235 VDD.n487 VDD.n486 4.65
R1236 VDD.n492 VDD.n491 4.65
R1237 VDD.n496 VDD.n495 4.65
R1238 VDD.n500 VDD.n499 4.65
R1239 VDD.n526 VDD.n525 4.65
R1240 VDD.n531 VDD.n530 4.65
R1241 VDD.n535 VDD.n534 4.65
R1242 VDD.n540 VDD.n539 4.65
R1243 VDD.n544 VDD.n543 4.65
R1244 VDD.n548 VDD.n547 4.65
R1245 VDD.n553 VDD.n552 4.65
R1246 VDD.n557 VDD.n556 4.65
R1247 VDD.n583 VDD.n582 4.65
R1248 VDD.n587 VDD.n586 4.65
R1249 VDD.n591 VDD.n590 4.65
R1250 VDD.n595 VDD.n594 4.65
R1251 VDD.n601 VDD.n600 4.65
R1252 VDD.n605 VDD.n604 4.65
R1253 VDD.n609 VDD.n608 4.65
R1254 VDD.n615 VDD.n614 4.65
R1255 VDD.n619 VDD.n618 4.65
R1256 VDD.n624 VDD.n623 4.65
R1257 VDD.n628 VDD.n627 4.65
R1258 VDD.n632 VDD.n631 4.65
R1259 VDD.n658 VDD.n657 4.65
R1260 VDD.n663 VDD.n662 4.65
R1261 VDD.n667 VDD.n666 4.65
R1262 VDD.n672 VDD.n671 4.65
R1263 VDD.n676 VDD.n675 4.65
R1264 VDD.n680 VDD.n679 4.65
R1265 VDD.n1369 VDD.n1368 4.65
R1266 VDD.n1364 VDD.n1363 4.65
R1267 VDD.n1338 VDD.n1337 4.65
R1268 VDD.n1334 VDD.n1333 4.65
R1269 VDD.n1329 VDD.n1328 4.65
R1270 VDD.n1325 VDD.n1324 4.65
R1271 VDD.n1320 VDD.n1319 4.65
R1272 VDD.n1316 VDD.n1315 4.65
R1273 VDD.n1312 VDD.n1311 4.65
R1274 VDD.n1307 VDD.n1306 4.65
R1275 VDD.n1281 VDD.n1280 4.65
R1276 VDD.n1277 VDD.n1276 4.65
R1277 VDD.n1273 VDD.n1272 4.65
R1278 VDD.n1269 VDD.n1268 4.65
R1279 VDD.n1265 VDD.n1264 4.65
R1280 VDD.n1259 VDD.n1258 4.65
R1281 VDD.n1255 VDD.n1254 4.65
R1282 VDD.n1251 VDD.n1250 4.65
R1283 VDD.n1245 VDD.n1244 4.65
R1284 VDD.n1241 VDD.n1240 4.65
R1285 VDD.n1236 VDD.n1235 4.65
R1286 VDD.n1232 VDD.n1231 4.65
R1287 VDD.n1206 VDD.n1205 4.65
R1288 VDD.n1202 VDD.n1201 4.65
R1289 VDD.n1198 VDD.n1197 4.65
R1290 VDD.n1194 VDD.n1193 4.65
R1291 VDD.n1190 VDD.n1189 4.65
R1292 VDD.n1184 VDD.n1183 4.65
R1293 VDD.n1180 VDD.n1179 4.65
R1294 VDD.n1176 VDD.n1175 4.65
R1295 VDD.n1170 VDD.n1169 4.65
R1296 VDD.n1166 VDD.n1165 4.65
R1297 VDD.n1161 VDD.n1160 4.65
R1298 VDD.n1157 VDD.n1156 4.65
R1299 VDD.n1131 VDD.n1130 4.65
R1300 VDD.n1127 VDD.n1126 4.65
R1301 VDD.n1122 VDD.n1121 4.65
R1302 VDD.n1118 VDD.n1117 4.65
R1303 VDD.n1113 VDD.n1112 4.65
R1304 VDD.n1109 VDD.n1108 4.65
R1305 VDD.n1105 VDD.n1104 4.65
R1306 VDD.n1100 VDD.n1099 4.65
R1307 VDD.n1074 VDD.n1073 4.65
R1308 VDD.n1070 VDD.n1069 4.65
R1309 VDD.n1066 VDD.n1065 4.65
R1310 VDD.n1062 VDD.n1061 4.65
R1311 VDD.n1058 VDD.n1057 4.65
R1312 VDD.n1052 VDD.n1051 4.65
R1313 VDD.n1048 VDD.n1047 4.65
R1314 VDD.n1044 VDD.n1043 4.65
R1315 VDD.n1038 VDD.n1037 4.65
R1316 VDD.n1034 VDD.n1033 4.65
R1317 VDD.n1029 VDD.n1028 4.65
R1318 VDD.n1025 VDD.n1024 4.65
R1319 VDD.n999 VDD.n998 4.65
R1320 VDD.n995 VDD.n994 4.65
R1321 VDD.n990 VDD.n989 4.65
R1322 VDD.n986 VDD.n985 4.65
R1323 VDD.n981 VDD.n980 4.65
R1324 VDD.n977 VDD.n976 4.65
R1325 VDD.n973 VDD.n972 4.65
R1326 VDD.n968 VDD.n967 4.65
R1327 VDD.n942 VDD.n941 4.65
R1328 VDD.n938 VDD.n937 4.65
R1329 VDD.n933 VDD.n932 4.65
R1330 VDD.n929 VDD.n928 4.65
R1331 VDD.n924 VDD.n923 4.65
R1332 VDD.n920 VDD.n919 4.65
R1333 VDD.n916 VDD.n915 4.65
R1334 VDD.n911 VDD.n910 4.65
R1335 VDD.n885 VDD.n884 4.65
R1336 VDD.n881 VDD.n880 4.65
R1337 VDD.n877 VDD.n876 4.65
R1338 VDD.n873 VDD.n872 4.65
R1339 VDD.n869 VDD.n868 4.65
R1340 VDD.n863 VDD.n862 4.65
R1341 VDD.n859 VDD.n858 4.65
R1342 VDD.n855 VDD.n854 4.65
R1343 VDD.n849 VDD.n848 4.65
R1344 VDD.n845 VDD.n844 4.65
R1345 VDD.n840 VDD.n839 4.65
R1346 VDD.n836 VDD.n835 4.65
R1347 VDD.n810 VDD.n809 4.65
R1348 VDD.n806 VDD.n805 4.65
R1349 VDD.n802 VDD.n801 4.65
R1350 VDD.n798 VDD.n797 4.65
R1351 VDD.n794 VDD.n793 4.65
R1352 VDD.n788 VDD.n787 4.65
R1353 VDD.n784 VDD.n783 4.65
R1354 VDD.n780 VDD.n779 4.65
R1355 VDD.n774 VDD.n773 4.65
R1356 VDD.n770 VDD.n769 4.65
R1357 VDD.n765 VDD.n764 4.65
R1358 VDD.n761 VDD.n760 4.65
R1359 VDD.n734 VDD.n733 4.65
R1360 VDD.n730 VDD.n729 4.65
R1361 VDD.n725 VDD.n724 4.65
R1362 VDD.n721 VDD.n720 4.65
R1363 VDD.n716 VDD.n715 4.65
R1364 VDD.n712 VDD.n711 4.65
R1365 VDD.n708 VDD.n707 4.65
R1366 VDD.n703 VDD.n702 4.65
R1367 VDD.n27 VDD.n23 2.933
R1368 VDD.n156 VDD.n153 2.89
R1369 VDD.n288 VDD.n285 2.89
R1370 VDD.n345 VDD.n342 2.89
R1371 VDD.n552 VDD.n549 2.89
R1372 VDD.n1368 VDD.n1365 2.89
R1373 VDD.n1311 VDD.n1308 2.89
R1374 VDD.n1104 VDD.n1101 2.89
R1375 VDD.n972 VDD.n969 2.89
R1376 VDD.n915 VDD.n912 2.89
R1377 VDD.n707 VDD.n704 2.89
R1378 VDD.n27 VDD.n26 2.844
R1379 VDD.n35  2.557
R1380 VDD.n86 0<��� 2.557
R1381 VDD.n145  2.557
R1382 VDD.n277 0<��� 2.557
R1383 VDD.n334 0<��� 2.557
R1384 VDD.n541  2.557
R1385 VDD.n673  2.557
R1386 VDD.n1317 0<��� 2.557
R1387 VDD.n1110 VDD.t111 2.557
R1388 VDD.n978  2.557
R1389 VDD.n921 0<��� 2.557
R1390 VDD.n713 0<��� 2.557
R1391 VDD.n134 VDD.n131 2.477
R1392 VDD.n266 VDD.n263 2.477
R1393 VDD.n323 VDD.n320 2.477
R1394 VDD.n530 VDD.n527 2.477
R1395 VDD.n662 VDD.n659 2.477
R1396 VDD.n1333 VDD.n1330 2.477
R1397 VDD.n1126 VDD.n1123 2.477
R1398 VDD.n994 VDD.n991 2.477
R1399 VDD.n937 VDD.n934 2.477
R1400 VDD.n729 VDD.n726 2.477
R1401 VDD.n31 VDD.n27 1.063
R1402 VDD.n227 VDD.n224 0.412
R1403 VDD.n416 VDD.n413 0.412
R1404 VDD.n491 VDD.n488 0.412
R1405 VDD.n623 VDD.n620 0.412
R1406 VDD.n1240 VDD.n1237 0.412
R1407 VDD.n1165 VDD.n1162 0.412
R1408 VDD.n1033 VDD.n1030 0.412
R1409 VDD.n844 VDD.n841 0.412
R1410 VDD.n769 VDD.n766 0.412
R1411 VDD.n77 VDD.n50 0.29
R1412 VDD.n130 VDD.n104 0.29
R1413 VDD.n187 VDD.n161 0.29
R1414 VDD.n262 VDD.n236 0.29
R1415 VDD.n319 VDD.n293 0.29
R1416 VDD.n376 VDD.n350 0.29
R1417 VDD.n451 VDD.n425 0.29
R1418 VDD.n526 VDD.n500 0.29
R1419 VDD.n583 VDD.n557 0.29
R1420 VDD.n658 VDD.n632 0.29
R1421 VDD.n1364 VDD.n1338 0.29
R1422 VDD.n1307 VDD.n1281 0.29
R1423 VDD.n1232 VDD.n1206 0.29
R1424 VDD.n1157 VDD.n1131 0.29
R1425 VDD.n1100 VDD.n1074 0.29
R1426 VDD.n1025 VDD.n999 0.29
R1427 VDD.n968 VDD.n942 0.29
R1428 VDD.n911 VDD.n885 0.29
R1429 VDD.n836 VDD.n810 0.29
R1430 VDD.n761 VDD.n734 0.29
R1431 VDD.n703 VDD 0.207
R1432 VDD.n213 VDD.n209 0.197
R1433 VDD.n402 VDD.n398 0.197
R1434 VDD.n477 VDD.n473 0.197
R1435 VDD.n609 VDD.n605 0.197
R1436 VDD.n1259 VDD.n1255 0.197
R1437 VDD.n1184 VDD.n1180 0.197
R1438 VDD.n1052 VDD.n1048 0.197
R1439 VDD.n863 VDD.n859 0.197
R1440 VDD.n788 VDD.n784 0.197
R1441 VDD.n38 VDD.n34 0.181
R1442 VDD.n92 VDD.n89 0.181
R1443 VDD.n148 VDD.n144 0.181
R1444 VDD.n280 VDD.n276 0.181
R1445 VDD.n337 VDD.n333 0.181
R1446 VDD.n544 VDD.n540 0.181
R1447 VDD.n676 VDD.n672 0.181
R1448 VDD.n1325 VDD.n1320 0.181
R1449 VDD.n1118 VDD.n1113 0.181
R1450 VDD.n986 VDD.n981 0.181
R1451 VDD.n929 VDD.n924 0.181
R1452 VDD.n721 VDD.n716 0.181
R1453 VDD.n34 VDD.n31 0.145
R1454 VDD.n42 VDD.n38 0.145
R1455 VDD.n46 VDD.n42 0.145
R1456 VDD.n50 VDD.n46 0.145
R1457 VDD.n81 VDD.n77 0.145
R1458 VDD.n85 VDD.n81 0.145
R1459 VDD.n89 VDD.n85 0.145
R1460 VDD.n96 VDD.n92 0.145
R1461 VDD.n100 VDD.n96 0.145
R1462 VDD.n104 VDD.n100 0.145
R1463 VDD.n135 VDD.n130 0.145
R1464 VDD.n139 VDD.n135 0.145
R1465 VDD.n144 VDD.n139 0.145
R1466 VDD.n152 VDD.n148 0.145
R1467 VDD.n157 VDD.n152 0.145
R1468 VDD.n161 VDD.n157 0.145
R1469 VDD.n191 VDD.n187 0.145
R1470 VDD.n195 VDD.n191 0.145
R1471 VDD.n199 VDD.n195 0.145
R1472 VDD.n205 VDD.n199 0.145
R1473 VDD.n209 VDD.n205 0.145
R1474 VDD.n219 VDD.n213 0.145
R1475 VDD.n223 VDD.n219 0.145
R1476 VDD.n228 VDD.n223 0.145
R1477 VDD.n232 VDD.n228 0.145
R1478 VDD.n236 VDD.n232 0.145
R1479 VDD.n267 VDD.n262 0.145
R1480 VDD.n271 VDD.n267 0.145
R1481 VDD.n276 VDD.n271 0.145
R1482 VDD.n284 VDD.n280 0.145
R1483 VDD.n289 VDD.n284 0.145
R1484 VDD.n293 VDD.n289 0.145
R1485 VDD.n324 VDD.n319 0.145
R1486 VDD.n328 VDD.n324 0.145
R1487 VDD.n333 VDD.n328 0.145
R1488 VDD.n341 VDD.n337 0.145
R1489 VDD.n346 VDD.n341 0.145
R1490 VDD.n350 VDD.n346 0.145
R1491 VDD.n380 VDD.n376 0.145
R1492 VDD.n384 VDD.n380 0.145
R1493 VDD.n388 VDD.n384 0.145
R1494 VDD.n394 VDD.n388 0.145
R1495 VDD.n398 VDD.n394 0.145
R1496 VDD.n408 VDD.n402 0.145
R1497 VDD.n412 VDD.n408 0.145
R1498 VDD.n417 VDD.n412 0.145
R1499 VDD.n421 VDD.n417 0.145
R1500 VDD.n425 VDD.n421 0.145
R1501 VDD.n455 VDD.n451 0.145
R1502 VDD.n459 VDD.n455 0.145
R1503 VDD.n463 VDD.n459 0.145
R1504 VDD.n469 VDD.n463 0.145
R1505 VDD.n473 VDD.n469 0.145
R1506 VDD.n483 VDD.n477 0.145
R1507 VDD.n487 VDD.n483 0.145
R1508 VDD.n492 VDD.n487 0.145
R1509 VDD.n496 VDD.n492 0.145
R1510 VDD.n500 VDD.n496 0.145
R1511 VDD.n531 VDD.n526 0.145
R1512 VDD.n535 VDD.n531 0.145
R1513 VDD.n540 VDD.n535 0.145
R1514 VDD.n548 VDD.n544 0.145
R1515 VDD.n553 VDD.n548 0.145
R1516 VDD.n557 VDD.n553 0.145
R1517 VDD.n587 VDD.n583 0.145
R1518 VDD.n591 VDD.n587 0.145
R1519 VDD.n595 VDD.n591 0.145
R1520 VDD.n601 VDD.n595 0.145
R1521 VDD.n605 VDD.n601 0.145
R1522 VDD.n615 VDD.n609 0.145
R1523 VDD.n619 VDD.n615 0.145
R1524 VDD.n624 VDD.n619 0.145
R1525 VDD.n628 VDD.n624 0.145
R1526 VDD.n632 VDD.n628 0.145
R1527 VDD.n663 VDD.n658 0.145
R1528 VDD.n667 VDD.n663 0.145
R1529 VDD.n672 VDD.n667 0.145
R1530 VDD.n680 VDD.n676 0.145
R1531 VDD.n1369 VDD.n1364 0.145
R1532 VDD.n1338 VDD.n1334 0.145
R1533 VDD.n1334 VDD.n1329 0.145
R1534 VDD.n1329 VDD.n1325 0.145
R1535 VDD.n1320 VDD.n1316 0.145
R1536 VDD.n1316 VDD.n1312 0.145
R1537 VDD.n1312 VDD.n1307 0.145
R1538 VDD.n1281 VDD.n1277 0.145
R1539 VDD.n1277 VDD.n1273 0.145
R1540 VDD.n1273 VDD.n1269 0.145
R1541 VDD.n1269 VDD.n1265 0.145
R1542 VDD.n1265 VDD.n1259 0.145
R1543 VDD.n1255 VDD.n1251 0.145
R1544 VDD.n1251 VDD.n1245 0.145
R1545 VDD.n1245 VDD.n1241 0.145
R1546 VDD.n1241 VDD.n1236 0.145
R1547 VDD.n1236 VDD.n1232 0.145
R1548 VDD.n1206 VDD.n1202 0.145
R1549 VDD.n1202 VDD.n1198 0.145
R1550 VDD.n1198 VDD.n1194 0.145
R1551 VDD.n1194 VDD.n1190 0.145
R1552 VDD.n1190 VDD.n1184 0.145
R1553 VDD.n1180 VDD.n1176 0.145
R1554 VDD.n1176 VDD.n1170 0.145
R1555 VDD.n1170 VDD.n1166 0.145
R1556 VDD.n1166 VDD.n1161 0.145
R1557 VDD.n1161 VDD.n1157 0.145
R1558 VDD.n1131 VDD.n1127 0.145
R1559 VDD.n1127 VDD.n1122 0.145
R1560 VDD.n1122 VDD.n1118 0.145
R1561 VDD.n1113 VDD.n1109 0.145
R1562 VDD.n1109 VDD.n1105 0.145
R1563 VDD.n1105 VDD.n1100 0.145
R1564 VDD.n1074 VDD.n1070 0.145
R1565 VDD.n1070 VDD.n1066 0.145
R1566 VDD.n1066 VDD.n1062 0.145
R1567 VDD.n1062 VDD.n1058 0.145
R1568 VDD.n1058 VDD.n1052 0.145
R1569 VDD.n1048 VDD.n1044 0.145
R1570 VDD.n1044 VDD.n1038 0.145
R1571 VDD.n1038 VDD.n1034 0.145
R1572 VDD.n1034 VDD.n1029 0.145
R1573 VDD.n1029 VDD.n1025 0.145
R1574 VDD.n999 VDD.n995 0.145
R1575 VDD.n995 VDD.n990 0.145
R1576 VDD.n990 VDD.n986 0.145
R1577 VDD.n981 VDD.n977 0.145
R1578 VDD.n977 VDD.n973 0.145
R1579 VDD.n973 VDD.n968 0.145
R1580 VDD.n942 VDD.n938 0.145
R1581 VDD.n938 VDD.n933 0.145
R1582 VDD.n933 VDD.n929 0.145
R1583 VDD.n924 VDD.n920 0.145
R1584 VDD.n920 VDD.n916 0.145
R1585 VDD.n916 VDD.n911 0.145
R1586 VDD.n885 VDD.n881 0.145
R1587 VDD.n881 VDD.n877 0.145
R1588 VDD.n877 VDD.n873 0.145
R1589 VDD.n873 VDD.n869 0.145
R1590 VDD.n869 VDD.n863 0.145
R1591 VDD.n859 VDD.n855 0.145
R1592 VDD.n855 VDD.n849 0.145
R1593 VDD.n849 VDD.n845 0.145
R1594 VDD.n845 VDD.n840 0.145
R1595 VDD.n840 VDD.n836 0.145
R1596 VDD.n810 VDD.n806 0.145
R1597 VDD.n806 VDD.n802 0.145
R1598 VDD.n802 VDD.n798 0.145
R1599 VDD.n798 VDD.n794 0.145
R1600 VDD.n794 VDD.n788 0.145
R1601 VDD.n784 VDD.n780 0.145
R1602 VDD.n780 VDD.n774 0.145
R1603 VDD.n774 VDD.n770 0.145
R1604 VDD.n770 VDD.n765 0.145
R1605 VDD.n765 VDD.n761 0.145
R1606 VDD.n734 VDD.n730 0.145
R1607 VDD.n730 VDD.n725 0.145
R1608 VDD.n725 VDD.n721 0.145
R1609 VDD.n716 VDD.n712 0.145
R1610 VDD.n712 VDD.n708 0.145
R1611 VDD.n708 VDD.n703 0.145
R1612 VDD VDD.n1369 0.082
R1613 VDD VDD.n680 0.062
R1614 a_6789_1050.n5 a_6789_1050.t9 480.392
R1615 a_6789_1050.n5 a_6789_1050.t8 403.272
R1616 a_6789_1050.n6 a_6789_1050.t7 301.486
R1617 a_6789_1050.n9 a_6789_1050.n7 259.02
R1618 a_6789_1050.n7 a_6789_1050.n4 234.917
R1619 a_6789_1050.n6 a_6789_1050.n5 227.006
R1620 a_6789_1050.n3 a_6789_1050.n2 161.352
R1621 a_6789_1050.n4 a_6789_1050.n0 95.095
R1622 a_6789_1050.n3 a_6789_1050.n1 95.095
R1623 a_6789_1050.n4 a_6789_1050.n3 66.258
R1624 a_6789_1050.n9 a_6789_1050.n8 15.218
R1625 a_6789_1050.n0 a_6789_1050.t3 14.282
R1626 a_6789_1050.n0 a_6789_1050.t2 14.282
R1627 a_6789_1050.n1 a_6789_1050.t5 14.282
R1628 a_6789_1050.n1 a_6789_1050.t6 14.282
R1629 a_6789_1050.n2 a_6789_1050.t1 14.282
R1630 a_6789_1050.n2 a_6789_1050.t0 14.282
R1631 a_6789_1050.n10 a_6789_1050.n9 12.014
R1632 a_6789_1050.n7 a_6789_1050.n6 10.615
R1633 a_7586_101.t0 a_7586_101.n1 93.333
R1634 a_7586_101.n4 a_7586_101.n2 79.092
R1635 a_7586_101.t0 a_7586_101.n0 8.137
R1636 a_7586_101.n4 a_7586_101.n3 4.614
R1637 a_7586_101.t0 a_7586_101.n4 0.111
R1638 GND.n28 GND.n27 237.558
R1639 GND.n414 GND.n413 237.558
R1640 GND.n458 GND.n457 237.558
R1641 GND.n500 GND.n499 237.558
R1642 GND.n532 GND.n531 237.558
R1643 GND.n562 GND.n561 237.558
R1644 GND.n607 GND.n606 237.558
R1645 GND.n639 GND.n638 237.558
R1646 GND.n683 GND.n682 237.558
R1647 GND.n727 GND.n726 237.558
R1648 GND.n363 GND.n362 237.558
R1649 GND.n759 GND.n758 237.558
R1650 GND.n318 GND.n317 237.558
R1651 GND.n286 GND.n285 237.558
R1652 GND.n242 GND.n241 237.558
R1653 GND.n198 GND.n197 237.558
R1654 GND.n168 GND.n167 237.558
R1655 GND.n136 GND.n135 237.558
R1656 GND.n94 GND.n93 237.558
R1657 GND.n61 GND.n60 237.558
R1658 GND.n25 GND.n24 210.82
R1659 GND.n58 GND.n57 210.82
R1660 GND.n416 GND.n415 210.82
R1661 GND.n460 GND.n459 210.82
R1662 GND.n502 GND.n501 210.82
R1663 GND.n534 GND.n533 210.82
R1664 GND.n564 GND.n563 210.82
R1665 GND.n609 GND.n608 210.82
R1666 GND.n641 GND.n640 210.82
R1667 GND.n685 GND.n684 210.82
R1668 GND.n729 GND.n728 210.82
R1669 GND.n761 GND.n760 210.82
R1670 GND.n360 GND.n359 210.82
R1671 GND.n315 GND.n314 210.82
R1672 GND.n283 GND.n282 210.82
R1673 GND.n239 GND.n238 210.82
R1674 GND.n195 GND.n194 210.82
R1675 GND.n165 GND.n164 210.82
R1676 GND.n133 GND.n132 210.82
R1677 GND.n91 GND.n90 210.82
R1678 GND.n123 GND.n122 173.365
R1679 GND.n469 GND.n468 173.365
R1680 GND.n184 GND.n183 172.612
R1681 GND.n542 GND.n541 172.612
R1682 GND.n14 GND.n13 172.612
R1683 GND.n229 GND.n228 167.358
R1684 GND.n273 GND.n272 167.358
R1685 GND.n696 GND.n695 167.358
R1686 GND.n652 GND.n651 167.358
R1687 GND.n427 GND.n426 167.358
R1688 GND.n154 GND.n153 166.605
R1689 GND.n304 GND.n303 166.605
R1690 GND.n381 GND.n380 166.605
R1691 GND.n739 GND.n738 166.605
R1692 GND.n619 GND.n618 166.605
R1693 GND.n512 GND.n511 166.605
R1694 GND.n394 GND.n393 166.605
R1695 GND.n350 GND.n349 152.358
R1696 GND.n576 GND.n575 152.358
R1697 GND.n47 GND.n46 151.605
R1698 GND.n80 GND.n79 151.605
R1699 GND.n46 GND.n45 28.421
R1700 GND.n79 GND.n78 28.421
R1701 GND.n349 GND.n348 28.421
R1702 GND.n575 GND.n574 28.421
R1703 GND.n46 GND.n44 25.263
R1704 GND.n79 GND.n77 25.263
R1705 GND.n349 GND.n347 25.263
R1706 GND.n575 GND.n573 25.263
R1707 GND.n44 GND.n43 24.383
R1708 GND.n77 GND.n76 24.383
R1709 GND.n347 GND.n346 24.383
R1710 GND.n573 GND.n572 24.383
R1711 GND.n153 GND.n151 23.03
R1712 GND.n228 GND.n226 23.03
R1713 GND.n272 GND.n270 23.03
R1714 GND.n303 GND.n301 23.03
R1715 GND.n380 GND.n378 23.03
R1716 GND.n738 GND.n736 23.03
R1717 GND.n695 GND.n693 23.03
R1718 GND.n651 GND.n649 23.03
R1719 GND.n618 GND.n616 23.03
R1720 GND.n511 GND.n509 23.03
R1721 GND.n426 GND.n424 23.03
R1722 GND.n393 GND.n391 23.03
R1723 GND.n26 GND.n25 18.953
R1724 GND.n59 GND.n58 18.953
R1725 GND.n417 GND.n416 18.953
R1726 GND.n461 GND.n460 18.953
R1727 GND.n503 GND.n502 18.953
R1728 GND.n535 GND.n534 18.953
R1729 GND.n565 GND.n564 18.953
R1730 GND.n610 GND.n609 18.953
R1731 GND.n642 GND.n641 18.953
R1732 GND.n686 GND.n685 18.953
R1733 GND.n730 GND.n729 18.953
R1734 GND.n762 GND.n761 18.953
R1735 GND.n361 GND.n360 18.953
R1736 GND.n316 GND.n315 18.953
R1737 GND.n284 GND.n283 18.953
R1738 GND.n240 GND.n239 18.953
R1739 GND.n196 GND.n195 18.953
R1740 GND.n166 GND.n165 18.953
R1741 GND.n134 GND.n133 18.953
R1742 GND.n92 GND.n91 18.953
R1743 GND.n29 GND.n26 14.864
R1744 GND.n62 GND.n59 14.864
R1745 GND.n95 GND.n92 14.864
R1746 GND.n137 GND.n134 14.864
R1747 GND.n169 GND.n166 14.864
R1748 GND.n199 GND.n196 14.864
R1749 GND.n243 GND.n240 14.864
R1750 GND.n287 GND.n284 14.864
R1751 GND.n319 GND.n316 14.864
R1752 GND.n364 GND.n361 14.864
R1753 GND.n763 GND.n762 14.864
R1754 GND.n731 GND.n730 14.864
R1755 GND.n687 GND.n686 14.864
R1756 GND.n643 GND.n642 14.864
R1757 GND.n611 GND.n610 14.864
R1758 GND.n566 GND.n565 14.864
R1759 GND.n536 GND.n535 14.864
R1760 GND.n504 GND.n503 14.864
R1761 GND.n462 GND.n461 14.864
R1762 GND.n418 GND.n417 14.864
R1763 GND.n389 GND.n388 9.154
R1764 GND.n396 GND.n395 9.154
R1765 GND.n399 GND.n398 9.154
R1766 GND.n402 GND.n401 9.154
R1767 GND.n405 GND.n404 9.154
R1768 GND.n408 GND.n407 9.154
R1769 GND.n411 GND.n410 9.154
R1770 GND.n418 GND.n414 9.154
R1771 GND.n421 GND.n420 9.154
R1772 GND.n428 GND.n423 9.154
R1773 GND.n431 GND.n430 9.154
R1774 GND.n434 GND.n433 9.154
R1775 GND.n437 GND.n436 9.154
R1776 GND.n440 GND.n439 9.154
R1777 GND.n443 GND.n442 9.154
R1778 GND.n446 GND.n445 9.154
R1779 GND.n449 GND.n448 9.154
R1780 GND.n452 GND.n451 9.154
R1781 GND.n455 GND.n454 9.154
R1782 GND.n462 GND.n458 9.154
R1783 GND.n465 GND.n464 9.154
R1784 GND.n470 GND.n467 9.154
R1785 GND.n473 GND.n472 9.154
R1786 GND.n476 GND.n475 9.154
R1787 GND.n479 GND.n478 9.154
R1788 GND.n482 GND.n481 9.154
R1789 GND.n485 GND.n484 9.154
R1790 GND.n488 GND.n487 9.154
R1791 GND.n491 GND.n490 9.154
R1792 GND.n494 GND.n493 9.154
R1793 GND.n497 GND.n496 9.154
R1794 GND.n504 GND.n500 9.154
R1795 GND.n507 GND.n506 9.154
R1796 GND.n514 GND.n513 9.154
R1797 GND.n517 GND.n516 9.154
R1798 GND.n520 GND.n519 9.154
R1799 GND.n523 GND.n522 9.154
R1800 GND.n526 GND.n525 9.154
R1801 GND.n529 GND.n528 9.154
R1802 GND.n536 GND.n532 9.154
R1803 GND.n539 GND.n538 9.154
R1804 GND.n544 GND.n543 9.154
R1805 GND.n547 GND.n546 9.154
R1806 GND.n550 GND.n549 9.154
R1807 GND.n553 GND.n552 9.154
R1808 GND.n556 GND.n555 9.154
R1809 GND.n559 GND.n558 9.154
R1810 GND.n566 GND.n562 9.154
R1811 GND.n569 GND.n568 9.154
R1812 GND.n577 GND.n571 9.154
R1813 GND.n580 GND.n579 9.154
R1814 GND.n583 GND.n582 9.154
R1815 GND.n586 GND.n585 9.154
R1816 GND.n589 GND.n588 9.154
R1817 GND.n592 GND.n591 9.154
R1818 GND.n595 GND.n594 9.154
R1819 GND.n598 GND.n597 9.154
R1820 GND.n601 GND.n600 9.154
R1821 GND.n604 GND.n603 9.154
R1822 GND.n611 GND.n607 9.154
R1823 GND.n614 GND.n613 9.154
R1824 GND.n621 GND.n620 9.154
R1825 GND.n624 GND.n623 9.154
R1826 GND.n627 GND.n626 9.154
R1827 GND.n630 GND.n629 9.154
R1828 GND.n633 GND.n632 9.154
R1829 GND.n636 GND.n635 9.154
R1830 GND.n643 GND.n639 9.154
R1831 GND.n646 GND.n645 9.154
R1832 GND.n653 GND.n648 9.154
R1833 GND.n656 GND.n655 9.154
R1834 GND.n659 GND.n658 9.154
R1835 GND.n662 GND.n661 9.154
R1836 GND.n665 GND.n664 9.154
R1837 GND.n668 GND.n667 9.154
R1838 GND.n671 GND.n670 9.154
R1839 GND.n674 GND.n673 9.154
R1840 GND.n677 GND.n676 9.154
R1841 GND.n680 GND.n679 9.154
R1842 GND.n687 GND.n683 9.154
R1843 GND.n690 GND.n689 9.154
R1844 GND.n697 GND.n692 9.154
R1845 GND.n700 GND.n699 9.154
R1846 GND.n703 GND.n702 9.154
R1847 GND.n706 GND.n705 9.154
R1848 GND.n709 GND.n708 9.154
R1849 GND.n712 GND.n711 9.154
R1850 GND.n715 GND.n714 9.154
R1851 GND.n718 GND.n717 9.154
R1852 GND.n721 GND.n720 9.154
R1853 GND.n724 GND.n723 9.154
R1854 GND.n731 GND.n727 9.154
R1855 GND.n734 GND.n733 9.154
R1856 GND.n741 GND.n740 9.154
R1857 GND.n744 GND.n743 9.154
R1858 GND.n747 GND.n746 9.154
R1859 GND.n750 GND.n749 9.154
R1860 GND.n753 GND.n752 9.154
R1861 GND.n756 GND.n755 9.154
R1862 GND.n763 GND.n759 9.154
R1863 GND.n766 GND.n765 9.154
R1864 GND.n383 GND.n382 9.154
R1865 GND.n376 GND.n375 9.154
R1866 GND.n373 GND.n372 9.154
R1867 GND.n370 GND.n369 9.154
R1868 GND.n367 GND.n366 9.154
R1869 GND.n364 GND.n363 9.154
R1870 GND.n357 GND.n356 9.154
R1871 GND.n354 GND.n353 9.154
R1872 GND.n351 GND.n345 9.154
R1873 GND.n343 GND.n342 9.154
R1874 GND.n340 GND.n339 9.154
R1875 GND.n337 GND.n336 9.154
R1876 GND.n334 GND.n333 9.154
R1877 GND.n331 GND.n330 9.154
R1878 GND.n328 GND.n327 9.154
R1879 GND.n325 GND.n324 9.154
R1880 GND.n322 GND.n321 9.154
R1881 GND.n319 GND.n318 9.154
R1882 GND.n312 GND.n311 9.154
R1883 GND.n309 GND.n308 9.154
R1884 GND.n306 GND.n305 9.154
R1885 GND.n299 GND.n298 9.154
R1886 GND.n296 GND.n295 9.154
R1887 GND.n293 GND.n292 9.154
R1888 GND.n290 GND.n289 9.154
R1889 GND.n287 GND.n286 9.154
R1890 GND.n280 GND.n279 9.154
R1891 GND.n277 GND.n276 9.154
R1892 GND.n274 GND.n269 9.154
R1893 GND.n267 GND.n266 9.154
R1894 GND.n264 GND.n263 9.154
R1895 GND.n261 GND.n260 9.154
R1896 GND.n258 GND.n257 9.154
R1897 GND.n255 GND.n254 9.154
R1898 GND.n252 GND.n251 9.154
R1899 GND.n249 GND.n248 9.154
R1900 GND.n246 GND.n245 9.154
R1901 GND.n243 GND.n242 9.154
R1902 GND.n236 GND.n235 9.154
R1903 GND.n233 GND.n232 9.154
R1904 GND.n230 GND.n225 9.154
R1905 GND.n223 GND.n222 9.154
R1906 GND.n220 GND.n219 9.154
R1907 GND.n217 GND.n216 9.154
R1908 GND.n214 GND.n213 9.154
R1909 GND.n211 GND.n210 9.154
R1910 GND.n208 GND.n207 9.154
R1911 GND.n205 GND.n204 9.154
R1912 GND.n202 GND.n201 9.154
R1913 GND.n199 GND.n198 9.154
R1914 GND.n192 GND.n191 9.154
R1915 GND.n189 GND.n188 9.154
R1916 GND.n186 GND.n185 9.154
R1917 GND.n181 GND.n180 9.154
R1918 GND.n178 GND.n177 9.154
R1919 GND.n175 GND.n174 9.154
R1920 GND.n172 GND.n171 9.154
R1921 GND.n169 GND.n168 9.154
R1922 GND.n162 GND.n161 9.154
R1923 GND.n159 GND.n158 9.154
R1924 GND.n156 GND.n155 9.154
R1925 GND.n149 GND.n148 9.154
R1926 GND.n146 GND.n145 9.154
R1927 GND.n143 GND.n142 9.154
R1928 GND.n140 GND.n139 9.154
R1929 GND.n137 GND.n136 9.154
R1930 GND.n130 GND.n129 9.154
R1931 GND.n127 GND.n126 9.154
R1932 GND.n124 GND.n121 9.154
R1933 GND.n119 GND.n118 9.154
R1934 GND.n116 GND.n115 9.154
R1935 GND.n113 GND.n112 9.154
R1936 GND.n110 GND.n109 9.154
R1937 GND.n107 GND.n106 9.154
R1938 GND.n104 GND.n103 9.154
R1939 GND.n101 GND.n100 9.154
R1940 GND.n98 GND.n97 9.154
R1941 GND.n95 GND.n94 9.154
R1942 GND.n88 GND.n87 9.154
R1943 GND.n85 GND.n84 9.154
R1944 GND.n82 GND.n81 9.154
R1945 GND.n74 GND.n73 9.154
R1946 GND.n71 GND.n70 9.154
R1947 GND.n68 GND.n67 9.154
R1948 GND.n65 GND.n64 9.154
R1949 GND.n62 GND.n61 9.154
R1950 GND.n55 GND.n54 9.154
R1951 GND.n52 GND.n51 9.154
R1952 GND.n49 GND.n48 9.154
R1953 GND.n41 GND.n40 9.154
R1954 GND.n38 GND.n37 9.154
R1955 GND.n1 GND.n0 9.154
R1956 GND.n5 GND.n4 9.154
R1957 GND.n8 GND.n7 9.154
R1958 GND.n11 GND.n10 9.154
R1959 GND.n16 GND.n15 9.154
R1960 GND.n19 GND.n18 9.154
R1961 GND.n22 GND.n21 9.154
R1962 GND.n29 GND.n28 9.154
R1963 GND.n32 GND.n31 9.154
R1964 GND.n35 GND.n34 9.154
R1965 GND.n153 GND.n152 8.128
R1966 GND.n228 GND.n227 8.128
R1967 GND.n272 GND.n271 8.128
R1968 GND.n303 GND.n302 8.128
R1969 GND.n380 GND.n379 8.128
R1970 GND.n738 GND.n737 8.128
R1971 GND.n695 GND.n694 8.128
R1972 GND.n651 GND.n650 8.128
R1973 GND.n618 GND.n617 8.128
R1974 GND.n511 GND.n510 8.128
R1975 GND.n426 GND.n425 8.128
R1976 GND.n393 GND.n392 8.128
R1977 GND.n387 GND.n386 4.65
R1978 GND.n39 GND.n38 4.65
R1979 GND.n42 GND.n41 4.65
R1980 GND.n50 GND.n49 4.65
R1981 GND.n53 GND.n52 4.65
R1982 GND.n56 GND.n55 4.65
R1983 GND.n63 GND.n62 4.65
R1984 GND.n66 GND.n65 4.65
R1985 GND.n69 GND.n68 4.65
R1986 GND.n72 GND.n71 4.65
R1987 GND.n75 GND.n74 4.65
R1988 GND.n83 GND.n82 4.65
R1989 GND.n86 GND.n85 4.65
R1990 GND.n89 GND.n88 4.65
R1991 GND.n96 GND.n95 4.65
R1992 GND.n99 GND.n98 4.65
R1993 GND.n102 GND.n101 4.65
R1994 GND.n105 GND.n104 4.65
R1995 GND.n108 GND.n107 4.65
R1996 GND.n111 GND.n110 4.65
R1997 GND.n114 GND.n113 4.65
R1998 GND.n117 GND.n116 4.65
R1999 GND.n120 GND.n119 4.65
R2000 GND.n125 GND.n124 4.65
R2001 GND.n128 GND.n127 4.65
R2002 GND.n131 GND.n130 4.65
R2003 GND.n138 GND.n137 4.65
R2004 GND.n141 GND.n140 4.65
R2005 GND.n144 GND.n143 4.65
R2006 GND.n147 GND.n146 4.65
R2007 GND.n150 GND.n149 4.65
R2008 GND.n157 GND.n156 4.65
R2009 GND.n160 GND.n159 4.65
R2010 GND.n163 GND.n162 4.65
R2011 GND.n170 GND.n169 4.65
R2012 GND.n173 GND.n172 4.65
R2013 GND.n176 GND.n175 4.65
R2014 GND.n179 GND.n178 4.65
R2015 GND.n182 GND.n181 4.65
R2016 GND.n187 GND.n186 4.65
R2017 GND.n190 GND.n189 4.65
R2018 GND.n193 GND.n192 4.65
R2019 GND.n200 GND.n199 4.65
R2020 GND.n203 GND.n202 4.65
R2021 GND.n206 GND.n205 4.65
R2022 GND.n209 GND.n208 4.65
R2023 GND.n212 GND.n211 4.65
R2024 GND.n215 GND.n214 4.65
R2025 GND.n218 GND.n217 4.65
R2026 GND.n221 GND.n220 4.65
R2027 GND.n224 GND.n223 4.65
R2028 GND.n231 GND.n230 4.65
R2029 GND.n234 GND.n233 4.65
R2030 GND.n237 GND.n236 4.65
R2031 GND.n244 GND.n243 4.65
R2032 GND.n247 GND.n246 4.65
R2033 GND.n250 GND.n249 4.65
R2034 GND.n253 GND.n252 4.65
R2035 GND.n256 GND.n255 4.65
R2036 GND.n259 GND.n258 4.65
R2037 GND.n262 GND.n261 4.65
R2038 GND.n265 GND.n264 4.65
R2039 GND.n268 GND.n267 4.65
R2040 GND.n275 GND.n274 4.65
R2041 GND.n278 GND.n277 4.65
R2042 GND.n281 GND.n280 4.65
R2043 GND.n288 GND.n287 4.65
R2044 GND.n291 GND.n290 4.65
R2045 GND.n294 GND.n293 4.65
R2046 GND.n297 GND.n296 4.65
R2047 GND.n300 GND.n299 4.65
R2048 GND.n307 GND.n306 4.65
R2049 GND.n310 GND.n309 4.65
R2050 GND.n313 GND.n312 4.65
R2051 GND.n320 GND.n319 4.65
R2052 GND.n323 GND.n322 4.65
R2053 GND.n326 GND.n325 4.65
R2054 GND.n329 GND.n328 4.65
R2055 GND.n332 GND.n331 4.65
R2056 GND.n335 GND.n334 4.65
R2057 GND.n338 GND.n337 4.65
R2058 GND.n341 GND.n340 4.65
R2059 GND.n344 GND.n343 4.65
R2060 GND.n352 GND.n351 4.65
R2061 GND.n355 GND.n354 4.65
R2062 GND.n358 GND.n357 4.65
R2063 GND.n365 GND.n364 4.65
R2064 GND.n368 GND.n367 4.65
R2065 GND.n371 GND.n370 4.65
R2066 GND.n374 GND.n373 4.65
R2067 GND.n377 GND.n376 4.65
R2068 GND.n384 GND.n383 4.65
R2069 GND.n767 GND.n766 4.65
R2070 GND.n764 GND.n763 4.65
R2071 GND.n757 GND.n756 4.65
R2072 GND.n754 GND.n753 4.65
R2073 GND.n751 GND.n750 4.65
R2074 GND.n748 GND.n747 4.65
R2075 GND.n745 GND.n744 4.65
R2076 GND.n742 GND.n741 4.65
R2077 GND.n735 GND.n734 4.65
R2078 GND.n732 GND.n731 4.65
R2079 GND.n725 GND.n724 4.65
R2080 GND.n722 GND.n721 4.65
R2081 GND.n719 GND.n718 4.65
R2082 GND.n716 GND.n715 4.65
R2083 GND.n713 GND.n712 4.65
R2084 GND.n710 GND.n709 4.65
R2085 GND.n707 GND.n706 4.65
R2086 GND.n704 GND.n703 4.65
R2087 GND.n701 GND.n700 4.65
R2088 GND.n698 GND.n697 4.65
R2089 GND.n691 GND.n690 4.65
R2090 GND.n688 GND.n687 4.65
R2091 GND.n681 GND.n680 4.65
R2092 GND.n678 GND.n677 4.65
R2093 GND.n675 GND.n674 4.65
R2094 GND.n672 GND.n671 4.65
R2095 GND.n669 GND.n668 4.65
R2096 GND.n666 GND.n665 4.65
R2097 GND.n663 GND.n662 4.65
R2098 GND.n660 GND.n659 4.65
R2099 GND.n657 GND.n656 4.65
R2100 GND.n654 GND.n653 4.65
R2101 GND.n647 GND.n646 4.65
R2102 GND.n644 GND.n643 4.65
R2103 GND.n637 GND.n636 4.65
R2104 GND.n634 GND.n633 4.65
R2105 GND.n631 GND.n630 4.65
R2106 GND.n628 GND.n627 4.65
R2107 GND.n625 GND.n624 4.65
R2108 GND.n622 GND.n621 4.65
R2109 GND.n615 GND.n614 4.65
R2110 GND.n612 GND.n611 4.65
R2111 GND.n605 GND.n604 4.65
R2112 GND.n602 GND.n601 4.65
R2113 GND.n599 GND.n598 4.65
R2114 GND.n596 GND.n595 4.65
R2115 GND.n593 GND.n592 4.65
R2116 GND.n590 GND.n589 4.65
R2117 GND.n587 GND.n586 4.65
R2118 GND.n584 GND.n583 4.65
R2119 GND.n581 GND.n580 4.65
R2120 GND.n578 GND.n577 4.65
R2121 GND.n570 GND.n569 4.65
R2122 GND.n567 GND.n566 4.65
R2123 GND.n560 GND.n559 4.65
R2124 GND.n557 GND.n556 4.65
R2125 GND.n554 GND.n553 4.65
R2126 GND.n551 GND.n550 4.65
R2127 GND.n548 GND.n547 4.65
R2128 GND.n545 GND.n544 4.65
R2129 GND.n540 GND.n539 4.65
R2130 GND.n537 GND.n536 4.65
R2131 GND.n530 GND.n529 4.65
R2132 GND.n527 GND.n526 4.65
R2133 GND.n524 GND.n523 4.65
R2134 GND.n521 GND.n520 4.65
R2135 GND.n518 GND.n517 4.65
R2136 GND.n515 GND.n514 4.65
R2137 GND.n508 GND.n507 4.65
R2138 GND.n505 GND.n504 4.65
R2139 GND.n498 GND.n497 4.65
R2140 GND.n495 GND.n494 4.65
R2141 GND.n492 GND.n491 4.65
R2142 GND.n489 GND.n488 4.65
R2143 GND.n486 GND.n485 4.65
R2144 GND.n483 GND.n482 4.65
R2145 GND.n480 GND.n479 4.65
R2146 GND.n477 GND.n476 4.65
R2147 GND.n474 GND.n473 4.65
R2148 GND.n471 GND.n470 4.65
R2149 GND.n466 GND.n465 4.65
R2150 GND.n463 GND.n462 4.65
R2151 GND.n456 GND.n455 4.65
R2152 GND.n453 GND.n452 4.65
R2153 GND.n450 GND.n449 4.65
R2154 GND.n447 GND.n446 4.65
R2155 GND.n444 GND.n443 4.65
R2156 GND.n441 GND.n440 4.65
R2157 GND.n438 GND.n437 4.65
R2158 GND.n435 GND.n434 4.65
R2159 GND.n432 GND.n431 4.65
R2160 GND.n429 GND.n428 4.65
R2161 GND.n422 GND.n421 4.65
R2162 GND.n419 GND.n418 4.65
R2163 GND.n412 GND.n411 4.65
R2164 GND.n409 GND.n408 4.65
R2165 GND.n406 GND.n405 4.65
R2166 GND.n403 GND.n402 4.65
R2167 GND.n400 GND.n399 4.65
R2168 GND.n397 GND.n396 4.65
R2169 GND.n390 GND.n389 4.65
R2170 GND.n6 GND.n5 4.65
R2171 GND.n9 GND.n8 4.65
R2172 GND.n12 GND.n11 4.65
R2173 GND.n17 GND.n16 4.65
R2174 GND.n20 GND.n19 4.65
R2175 GND.n23 GND.n22 4.65
R2176 GND.n30 GND.n29 4.65
R2177 GND.n33 GND.n32 4.65
R2178 GND.n36 GND.n35 4.65
R2179 GND.n16 GND.n14 4.129
R2180 GND.n49 GND.n47 4.129
R2181 GND.n82 GND.n80 4.129
R2182 GND.n156 GND.n154 4.129
R2183 GND.n186 GND.n184 4.129
R2184 GND.n306 GND.n304 4.129
R2185 GND.n383 GND.n381 4.129
R2186 GND.n741 GND.n739 4.129
R2187 GND.n621 GND.n619 4.129
R2188 GND.n544 GND.n542 4.129
R2189 GND.n514 GND.n512 4.129
R2190 GND.n396 GND.n394 4.129
R2191 GND.n3 GND.n2 3.408
R2192 GND.n3 GND.n1 2.844
R2193 GND.n6 GND.n3 1.063
R2194 GND.n386 GND.n385 0.474
R2195 GND.n30 GND.n23 0.29
R2196 GND.n63 GND.n56 0.29
R2197 GND.n96 GND.n89 0.29
R2198 GND.n138 GND.n131 0.29
R2199 GND.n170 GND.n163 0.29
R2200 GND.n200 GND.n193 0.29
R2201 GND.n244 GND.n237 0.29
R2202 GND.n288 GND.n281 0.29
R2203 GND.n320 GND.n313 0.29
R2204 GND.n365 GND.n358 0.29
R2205 GND.n764 GND.n757 0.29
R2206 GND.n732 GND.n725 0.29
R2207 GND.n688 GND.n681 0.29
R2208 GND.n644 GND.n637 0.29
R2209 GND.n612 GND.n605 0.29
R2210 GND.n567 GND.n560 0.29
R2211 GND.n537 GND.n530 0.29
R2212 GND.n505 GND.n498 0.29
R2213 GND.n463 GND.n456 0.29
R2214 GND.n419 GND.n412 0.29
R2215 GND.n387 GND 0.207
R2216 GND.n124 GND.n123 0.206
R2217 GND.n230 GND.n229 0.206
R2218 GND.n274 GND.n273 0.206
R2219 GND.n351 GND.n350 0.206
R2220 GND.n697 GND.n696 0.206
R2221 GND.n653 GND.n652 0.206
R2222 GND.n577 GND.n576 0.206
R2223 GND.n470 GND.n469 0.206
R2224 GND.n428 GND.n427 0.206
R2225 GND.n114 GND.n111 0.197
R2226 GND.n218 GND.n215 0.197
R2227 GND.n262 GND.n259 0.197
R2228 GND.n338 GND.n335 0.197
R2229 GND.n710 GND.n707 0.197
R2230 GND.n666 GND.n663 0.197
R2231 GND.n590 GND.n587 0.197
R2232 GND.n483 GND.n480 0.197
R2233 GND.n441 GND.n438 0.197
R2234 GND.n12 GND.n9 0.181
R2235 GND.n42 GND.n39 0.181
R2236 GND.n75 GND.n72 0.181
R2237 GND.n150 GND.n147 0.181
R2238 GND.n182 GND.n179 0.181
R2239 GND.n300 GND.n297 0.181
R2240 GND.n377 GND.n374 0.181
R2241 GND.n748 GND.n745 0.181
R2242 GND.n628 GND.n625 0.181
R2243 GND.n551 GND.n548 0.181
R2244 GND.n521 GND.n518 0.181
R2245 GND.n403 GND.n400 0.181
R2246 GND.n9 GND.n6 0.145
R2247 GND.n17 GND.n12 0.145
R2248 GND.n20 GND.n17 0.145
R2249 GND.n23 GND.n20 0.145
R2250 GND.n33 GND.n30 0.145
R2251 GND.n36 GND.n33 0.145
R2252 GND.n39 GND.n36 0.145
R2253 GND.n50 GND.n42 0.145
R2254 GND.n53 GND.n50 0.145
R2255 GND.n56 GND.n53 0.145
R2256 GND.n66 GND.n63 0.145
R2257 GND.n69 GND.n66 0.145
R2258 GND.n72 GND.n69 0.145
R2259 GND.n83 GND.n75 0.145
R2260 GND.n86 GND.n83 0.145
R2261 GND.n89 GND.n86 0.145
R2262 GND.n99 GND.n96 0.145
R2263 GND.n102 GND.n99 0.145
R2264 GND.n105 GND.n102 0.145
R2265 GND.n108 GND.n105 0.145
R2266 GND.n111 GND.n108 0.145
R2267 GND.n117 GND.n114 0.145
R2268 GND.n120 GND.n117 0.145
R2269 GND.n125 GND.n120 0.145
R2270 GND.n128 GND.n125 0.145
R2271 GND.n131 GND.n128 0.145
R2272 GND.n141 GND.n138 0.145
R2273 GND.n144 GND.n141 0.145
R2274 GND.n147 GND.n144 0.145
R2275 GND.n157 GND.n150 0.145
R2276 GND.n160 GND.n157 0.145
R2277 GND.n163 GND.n160 0.145
R2278 GND.n173 GND.n170 0.145
R2279 GND.n176 GND.n173 0.145
R2280 GND.n179 GND.n176 0.145
R2281 GND.n187 GND.n182 0.145
R2282 GND.n190 GND.n187 0.145
R2283 GND.n193 GND.n190 0.145
R2284 GND.n203 GND.n200 0.145
R2285 GND.n206 GND.n203 0.145
R2286 GND.n209 GND.n206 0.145
R2287 GND.n212 GND.n209 0.145
R2288 GND.n215 GND.n212 0.145
R2289 GND.n221 GND.n218 0.145
R2290 GND.n224 GND.n221 0.145
R2291 GND.n231 GND.n224 0.145
R2292 GND.n234 GND.n231 0.145
R2293 GND.n237 GND.n234 0.145
R2294 GND.n247 GND.n244 0.145
R2295 GND.n250 GND.n247 0.145
R2296 GND.n253 GND.n250 0.145
R2297 GND.n256 GND.n253 0.145
R2298 GND.n259 GND.n256 0.145
R2299 GND.n265 GND.n262 0.145
R2300 GND.n268 GND.n265 0.145
R2301 GND.n275 GND.n268 0.145
R2302 GND.n278 GND.n275 0.145
R2303 GND.n281 GND.n278 0.145
R2304 GND.n291 GND.n288 0.145
R2305 GND.n294 GND.n291 0.145
R2306 GND.n297 GND.n294 0.145
R2307 GND.n307 GND.n300 0.145
R2308 GND.n310 GND.n307 0.145
R2309 GND.n313 GND.n310 0.145
R2310 GND.n323 GND.n320 0.145
R2311 GND.n326 GND.n323 0.145
R2312 GND.n329 GND.n326 0.145
R2313 GND.n332 GND.n329 0.145
R2314 GND.n335 GND.n332 0.145
R2315 GND.n341 GND.n338 0.145
R2316 GND.n344 GND.n341 0.145
R2317 GND.n352 GND.n344 0.145
R2318 GND.n355 GND.n352 0.145
R2319 GND.n358 GND.n355 0.145
R2320 GND.n368 GND.n365 0.145
R2321 GND.n371 GND.n368 0.145
R2322 GND.n374 GND.n371 0.145
R2323 GND.n384 GND.n377 0.145
R2324 GND.n767 GND.n764 0.145
R2325 GND.n757 GND.n754 0.145
R2326 GND.n754 GND.n751 0.145
R2327 GND.n751 GND.n748 0.145
R2328 GND.n745 GND.n742 0.145
R2329 GND.n742 GND.n735 0.145
R2330 GND.n735 GND.n732 0.145
R2331 GND.n725 GND.n722 0.145
R2332 GND.n722 GND.n719 0.145
R2333 GND.n719 GND.n716 0.145
R2334 GND.n716 GND.n713 0.145
R2335 GND.n713 GND.n710 0.145
R2336 GND.n707 GND.n704 0.145
R2337 GND.n704 GND.n701 0.145
R2338 GND.n701 GND.n698 0.145
R2339 GND.n698 GND.n691 0.145
R2340 GND.n691 GND.n688 0.145
R2341 GND.n681 GND.n678 0.145
R2342 GND.n678 GND.n675 0.145
R2343 GND.n675 GND.n672 0.145
R2344 GND.n672 GND.n669 0.145
R2345 GND.n669 GND.n666 0.145
R2346 GND.n663 GND.n660 0.145
R2347 GND.n660 GND.n657 0.145
R2348 GND.n657 GND.n654 0.145
R2349 GND.n654 GND.n647 0.145
R2350 GND.n647 GND.n644 0.145
R2351 GND.n637 GND.n634 0.145
R2352 GND.n634 GND.n631 0.145
R2353 GND.n631 GND.n628 0.145
R2354 GND.n625 GND.n622 0.145
R2355 GND.n622 GND.n615 0.145
R2356 GND.n615 GND.n612 0.145
R2357 GND.n605 GND.n602 0.145
R2358 GND.n602 GND.n599 0.145
R2359 GND.n599 GND.n596 0.145
R2360 GND.n596 GND.n593 0.145
R2361 GND.n593 GND.n590 0.145
R2362 GND.n587 GND.n584 0.145
R2363 GND.n584 GND.n581 0.145
R2364 GND.n581 GND.n578 0.145
R2365 GND.n578 GND.n570 0.145
R2366 GND.n570 GND.n567 0.145
R2367 GND.n560 GND.n557 0.145
R2368 GND.n557 GND.n554 0.145
R2369 GND.n554 GND.n551 0.145
R2370 GND.n548 GND.n545 0.145
R2371 GND.n545 GND.n540 0.145
R2372 GND.n540 GND.n537 0.145
R2373 GND.n530 GND.n527 0.145
R2374 GND.n527 GND.n524 0.145
R2375 GND.n524 GND.n521 0.145
R2376 GND.n518 GND.n515 0.145
R2377 GND.n515 GND.n508 0.145
R2378 GND.n508 GND.n505 0.145
R2379 GND.n498 GND.n495 0.145
R2380 GND.n495 GND.n492 0.145
R2381 GND.n492 GND.n489 0.145
R2382 GND.n489 GND.n486 0.145
R2383 GND.n486 GND.n483 0.145
R2384 GND.n480 GND.n477 0.145
R2385 GND.n477 GND.n474 0.145
R2386 GND.n474 GND.n471 0.145
R2387 GND.n471 GND.n466 0.145
R2388 GND.n466 GND.n463 0.145
R2389 GND.n456 GND.n453 0.145
R2390 GND.n453 GND.n450 0.145
R2391 GND.n450 GND.n447 0.145
R2392 GND.n447 GND.n444 0.145
R2393 GND.n444 GND.n441 0.145
R2394 GND.n438 GND.n435 0.145
R2395 GND.n435 GND.n432 0.145
R2396 GND.n432 GND.n429 0.145
R2397 GND.n429 GND.n422 0.145
R2398 GND.n422 GND.n419 0.145
R2399 GND.n412 GND.n409 0.145
R2400 GND.n409 GND.n406 0.145
R2401 GND.n406 GND.n403 0.145
R2402 GND.n400 GND.n397 0.145
R2403 GND.n397 GND.n390 0.145
R2404 GND.n390 GND.n387 0.145
R2405 GND GND.n767 0.082
R2406 GND GND.n384 0.062
R2407 D.n5 D.t1 480.392
R2408 D.n2 D.t0 480.392
R2409 D.n0 D.t5 480.392
R2410 D.n5 D.t4 403.272
R2411 D.n2 D.t7 403.272
R2412 D.n0 D.t8 403.272
R2413 D.n6 D.n5 282.724
R2414 D.n3 D.n2 282.724
R2415 D.n1 D.n0 282.724
R2416 D.n6 D.t3 178.533
R2417 D.n3 D.t2 178.533
R2418 D.n1 D.t6 178.533
R2419 D.n4 D.n1 22.56
R2420 D.n7 D.n4 17.91
R2421 D.n4 D.n3 4.65
R2422 D.n7 D.n6 4.65
R2423 D.n7 D 0.046
R2424 a_5101_1050.n3 a_5101_1050.t6 512.525
R2425 a_5101_1050.n1 a_5101_1050.t5 512.525
R2426 a_5101_1050.n3 a_5101_1050.t9 371.139
R2427 a_5101_1050.n1 a_5101_1050.t7 371.139
R2428 a_5101_1050.n2 a_5101_1050.t10 305.674
R2429 a_5101_1050.n4 a_5101_1050.t8 305.298
R2430 a_5101_1050.n4 a_5101_1050.n3 291.648
R2431 a_5101_1050.n2 a_5101_1050.n1 291.272
R2432 a_5101_1050.n7 a_5101_1050.n6 271.602
R2433 a_5101_1050.n8 a_5101_1050.n7 215.717
R2434 a_5101_1050.n9 a_5101_1050.n8 157.963
R2435 a_5101_1050.n8 a_5101_1050.n0 91.706
R2436 a_5101_1050.n0 a_5101_1050.t2 14.282
R2437 a_5101_1050.n0 a_5101_1050.t1 14.282
R2438 a_5101_1050.t4 a_5101_1050.n9 14.282
R2439 a_5101_1050.n9 a_5101_1050.t3 14.282
R2440 a_5101_1050.n5 a_5101_1050.n2 8.138
R2441 a_5101_1050.n7 a_5101_1050.n5 5.964
R2442 a_5101_1050.n5 a_5101_1050.n4 4.65
R2443 CLK.n15 CLK.t12 472.359
R2444 CLK.n6 CLK.t13 472.359
R2445 CLK.n0 CLK.t17 472.359
R2446 CLK.n20 CLK.t5 459.505
R2447 CLK.n11 CLK.t15 459.505
R2448 CLK.n2 CLK.t11 459.505
R2449 CLK.n21 CLK.t9 399.181
R2450 CLK.n12 CLK.t16 399.181
R2451 CLK.n3 CLK.t4 399.181
R2452 CLK.n1 CLK.t7 398.558
R2453 CLK.n17 CLK.t1 397.101
R2454 CLK.n8 CLK.t6 397.101
R2455 CLK.n20 CLK.t10 384.527
R2456 CLK.n15 CLK.t14 384.527
R2457 CLK.n11 CLK.t0 384.527
R2458 CLK.n6 CLK.t3 384.527
R2459 CLK.n2 CLK.t2 384.527
R2460 CLK.n0 CLK.t8 384.527
R2461 CLK.n21 CLK.n20 33.832
R2462 CLK.n3 CLK.n2 33.832
R2463 CLK.n12 CLK.n11 33.832
R2464 CLK.n1 CLK.n0 32.394
R2465 CLK.n16 CLK.n15 30.822
R2466 CLK.n7 CLK.n6 30.822
R2467 CLK.n5 CLK.n4 11.101
R2468 CLK.n14 CLK.n13 11.101
R2469 CLK.n4 CLK.n1 8.215
R2470 CLK.n13 CLK.n10 6.718
R2471 CLK.n22 CLK.n19 6.718
R2472 CLK.n17 CLK.n16 4.577
R2473 CLK.n8 CLK.n7 4.577
R2474 CLK.n9 CLK.n8 4.282
R2475 CLK.n18 CLK.n17 4.282
R2476 CLK.n4 CLK.n3 2.079
R2477 CLK.n13 CLK.n12 2.079
R2478 CLK.n22 CLK.n21 2.079
R2479 CLK.n22 CLK 0.046
R2480 CLK.n10 CLK.n9 0.038
R2481 CLK.n19 CLK.n18 0.038
R2482 CLK.n9 CLK.n5 0.008
R2483 CLK.n18 CLK.n14 0.008
R2484 a_5227_411.n2 a_5227_411.t8 480.392
R2485 a_5227_411.n4 a_5227_411.t7 472.359
R2486 a_5227_411.n3 a_5227_411.t12 412.921
R2487 a_5227_411.n2 a_5227_411.t11 403.272
R2488 a_5227_411.n4 a_5227_411.t10 384.527
R2489 a_5227_411.n10 a_5227_411.n9 379.101
R2490 a_5227_411.n5 a_5227_411.t9 370.613
R2491 a_5227_411.n13 a_5227_411.n12 161.352
R2492 a_5227_411.n5 a_5227_411.n4 127.096
R2493 a_5227_411.n11 a_5227_411.n10 123.126
R2494 a_5227_411.n3 a_5227_411.n2 115.571
R2495 a_5227_411.n11 a_5227_411.n1 95.095
R2496 a_5227_411.n12 a_5227_411.n0 95.095
R2497 a_5227_411.n12 a_5227_411.n11 66.258
R2498 a_5227_411.n9 a_5227_411.n8 22.578
R2499 a_5227_411.n1 a_5227_411.t1 14.282
R2500 a_5227_411.n1 a_5227_411.t2 14.282
R2501 a_5227_411.n0 a_5227_411.t5 14.282
R2502 a_5227_411.n0 a_5227_411.t6 14.282
R2503 a_5227_411.t4 a_5227_411.n13 14.282
R2504 a_5227_411.n13 a_5227_411.t3 14.282
R2505 a_5227_411.n6 a_5227_411.n3 11.954
R2506 a_5227_411.n6 a_5227_411.n5 8.682
R2507 a_5227_411.n9 a_5227_411.n7 8.58
R2508 a_5227_411.n10 a_5227_411.n6 4.65
R2509 a_3599_411.n7 a_3599_411.t15 512.525
R2510 a_3599_411.n6 a_3599_411.t10 512.525
R2511 a_3599_411.n11 a_3599_411.t13 472.359
R2512 a_3599_411.n11 a_3599_411.t9 384.527
R2513 a_3599_411.n7 a_3599_411.t11 371.139
R2514 a_3599_411.n6 a_3599_411.t7 371.139
R2515 a_3599_411.n8 a_3599_411.n7 343.521
R2516 a_3599_411.n12 a_3599_411.t14 287.037
R2517 a_3599_411.n16 a_3599_411.n14 280.357
R2518 a_3599_411.n10 a_3599_411.n6 259.945
R2519 a_3599_411.n12 a_3599_411.n11 210.673
R2520 a_3599_411.n14 a_3599_411.n5 207.058
R2521 a_3599_411.n8 a_3599_411.t8 172.106
R2522 a_3599_411.n9 a_3599_411.t12 165.68
R2523 a_3599_411.n4 a_3599_411.n3 161.352
R2524 a_3599_411.n5 a_3599_411.n1 95.095
R2525 a_3599_411.n4 a_3599_411.n2 95.095
R2526 a_3599_411.n10 a_3599_411.n9 83.576
R2527 a_3599_411.n5 a_3599_411.n4 66.258
R2528 a_3599_411.n17 a_3599_411.n0 55.263
R2529 a_3599_411.n13 a_3599_411.n10 45.413
R2530 a_3599_411.n16 a_3599_411.n15 30
R2531 a_3599_411.n17 a_3599_411.n16 23.684
R2532 a_3599_411.n1 a_3599_411.t0 14.282
R2533 a_3599_411.n1 a_3599_411.t1 14.282
R2534 a_3599_411.n2 a_3599_411.t3 14.282
R2535 a_3599_411.n2 a_3599_411.t2 14.282
R2536 a_3599_411.n3 a_3599_411.t4 14.282
R2537 a_3599_411.n3 a_3599_411.t6 14.282
R2538 a_3599_411.n9 a_3599_411.n8 10.343
R2539 a_3599_411.n13 a_3599_411.n12 8.685
R2540 a_3599_411.n14 a_3599_411.n13 4.65
R2541 a_15533_1051.n4 a_15533_1051.t3 179.895
R2542 a_15533_1051.n2 a_15533_1051.n1 165.613
R2543 a_15533_1051.n2 a_15533_1051.n0 142.653
R2544 a_15533_1051.n4 a_15533_1051.n3 106.183
R2545 a_15533_1051.n5 a_15533_1051.n4 99.358
R2546 a_15533_1051.n3 a_15533_1051.n2 82.665
R2547 a_15533_1051.n3 a_15533_1051.t6 73.712
R2548 a_15533_1051.n0 a_15533_1051.t5 14.282
R2549 a_15533_1051.n0 a_15533_1051.t4 14.282
R2550 a_15533_1051.n1 a_15533_1051.t2 14.282
R2551 a_15533_1051.n1 a_15533_1051.t1 14.282
R2552 a_15533_1051.t0 a_15533_1051.n5 14.282
R2553 a_15533_1051.n5 a_15533_1051.t7 14.282
R2554 a_14869_1051.n2 a_14869_1051.t7 179.895
R2555 a_14869_1051.n5 a_14869_1051.n4 157.021
R2556 a_14869_1051.n4 a_14869_1051.n0 124.955
R2557 a_14869_1051.n3 a_14869_1051.n2 106.183
R2558 a_14869_1051.n2 a_14869_1051.n1 99.355
R2559 a_14869_1051.n4 a_14869_1051.n3 82.65
R2560 a_14869_1051.n3 a_14869_1051.t2 73.712
R2561 a_14869_1051.n0 a_14869_1051.t5 14.282
R2562 a_14869_1051.n0 a_14869_1051.t4 14.282
R2563 a_14869_1051.n1 a_14869_1051.t6 14.282
R2564 a_14869_1051.n1 a_14869_1051.t3 14.282
R2565 a_14869_1051.n5 a_14869_1051.t0 14.282
R2566 a_14869_1051.t1 a_14869_1051.n5 14.282
R2567 a_217_1050.n3 a_217_1050.t6 512.525
R2568 a_217_1050.n1 a_217_1050.t10 512.525
R2569 a_217_1050.n3 a_217_1050.t9 371.139
R2570 a_217_1050.n1 a_217_1050.t5 371.139
R2571 a_217_1050.n2 a_217_1050.t8 305.674
R2572 a_217_1050.n4 a_217_1050.t7 305.298
R2573 a_217_1050.n4 a_217_1050.n3 291.648
R2574 a_217_1050.n2 a_217_1050.n1 291.272
R2575 a_217_1050.n7 a_217_1050.n6 271.602
R2576 a_217_1050.n8 a_217_1050.n7 215.717
R2577 a_217_1050.n9 a_217_1050.n8 157.963
R2578 a_217_1050.n8 a_217_1050.n0 91.706
R2579 a_217_1050.n0 a_217_1050.t0 14.282
R2580 a_217_1050.n0 a_217_1050.t4 14.282
R2581 a_217_1050.t2 a_217_1050.n9 14.282
R2582 a_217_1050.n9 a_217_1050.t1 14.282
R2583 a_217_1050.n5 a_217_1050.n2 8.138
R2584 a_217_1050.n7 a_217_1050.n5 5.964
R2585 a_217_1050.n5 a_217_1050.n4 4.65
R2586 a_1265_989.n2 a_1265_989.t11 454.685
R2587 a_1265_989.n4 a_1265_989.t13 454.685
R2588 a_1265_989.n0 a_1265_989.t6 454.685
R2589 a_1265_989.n2 a_1265_989.t5 428.979
R2590 a_1265_989.n4 a_1265_989.t10 428.979
R2591 a_1265_989.n0 a_1265_989.t9 428.979
R2592 a_1265_989.n3 a_1265_989.t7 339.542
R2593 a_1265_989.n5 a_1265_989.t8 339.542
R2594 a_1265_989.n1 a_1265_989.t12 339.542
R2595 a_1265_989.n12 a_1265_989.n11 333.44
R2596 a_1265_989.n14 a_1265_989.n13 157.964
R2597 a_1265_989.n3 a_1265_989.n2 143.429
R2598 a_1265_989.n5 a_1265_989.n4 143.429
R2599 a_1265_989.n1 a_1265_989.n0 143.429
R2600 a_1265_989.n14 a_1265_989.n12 132.141
R2601 a_1265_989.n15 a_1265_989.n14 91.705
R2602 a_1265_989.n11 a_1265_989.n10 30
R2603 a_1265_989.n9 a_1265_989.n8 24.383
R2604 a_1265_989.n11 a_1265_989.n9 23.684
R2605 a_1265_989.n13 a_1265_989.t0 14.282
R2606 a_1265_989.n13 a_1265_989.t1 14.282
R2607 a_1265_989.t3 a_1265_989.n15 14.282
R2608 a_1265_989.n15 a_1265_989.t2 14.282
R2609 a_1265_989.n7 a_1265_989.n1 10.046
R2610 a_1265_989.n6 a_1265_989.n5 8.141
R2611 a_1265_989.n6 a_1265_989.n3 4.65
R2612 a_1265_989.n12 a_1265_989.n7 4.65
R2613 a_1265_989.n7 a_1265_989.n6 2.947
R2614 a_1905_1050.n2 a_1905_1050.t7 480.392
R2615 a_1905_1050.n2 a_1905_1050.t9 403.272
R2616 a_1905_1050.n3 a_1905_1050.t8 301.486
R2617 a_1905_1050.n8 a_1905_1050.n7 252.498
R2618 a_1905_1050.n9 a_1905_1050.n8 234.917
R2619 a_1905_1050.n3 a_1905_1050.n2 227.006
R2620 a_1905_1050.n11 a_1905_1050.n10 161.352
R2621 a_1905_1050.n9 a_1905_1050.n1 95.095
R2622 a_1905_1050.n10 a_1905_1050.n0 95.095
R2623 a_1905_1050.n10 a_1905_1050.n9 66.258
R2624 a_1905_1050.n7 a_1905_1050.n6 30
R2625 a_1905_1050.n5 a_1905_1050.n4 24.383
R2626 a_1905_1050.n7 a_1905_1050.n5 23.684
R2627 a_1905_1050.n1 a_1905_1050.t5 14.282
R2628 a_1905_1050.n1 a_1905_1050.t4 14.282
R2629 a_1905_1050.n0 a_1905_1050.t2 14.282
R2630 a_1905_1050.n0 a_1905_1050.t3 14.282
R2631 a_1905_1050.n11 a_1905_1050.t0 14.282
R2632 a_1905_1050.t1 a_1905_1050.n11 14.282
R2633 a_1905_1050.n8 a_1905_1050.n3 10.615
R2634 a_10111_411.n1 a_10111_411.t11 480.392
R2635 a_10111_411.n3 a_10111_411.t9 472.359
R2636 a_10111_411.n2 a_10111_411.t12 412.921
R2637 a_10111_411.n1 a_10111_411.t8 403.272
R2638 a_10111_411.n3 a_10111_411.t7 384.527
R2639 a_10111_411.n9 a_10111_411.n8 379.101
R2640 a_10111_411.n4 a_10111_411.t10 370.613
R2641 a_10111_411.n12 a_10111_411.n11 161.352
R2642 a_10111_411.n4 a_10111_411.n3 127.096
R2643 a_10111_411.n10 a_10111_411.n9 123.126
R2644 a_10111_411.n2 a_10111_411.n1 115.571
R2645 a_10111_411.n10 a_10111_411.n0 95.095
R2646 a_10111_411.n13 a_10111_411.n12 95.094
R2647 a_10111_411.n12 a_10111_411.n10 66.258
R2648 a_10111_411.n8 a_10111_411.n7 22.578
R2649 a_10111_411.n0 a_10111_411.t1 14.282
R2650 a_10111_411.n0 a_10111_411.t4 14.282
R2651 a_10111_411.n11 a_10111_411.t3 14.282
R2652 a_10111_411.n11 a_10111_411.t2 14.282
R2653 a_10111_411.n13 a_10111_411.t5 14.282
R2654 a_10111_411.t6 a_10111_411.n13 14.282
R2655 a_10111_411.n5 a_10111_411.n2 11.954
R2656 a_10111_411.n5 a_10111_411.n4 8.682
R2657 a_10111_411.n8 a_10111_411.n6 8.58
R2658 a_10111_411.n9 a_10111_411.n5 4.65
R2659 a_9985_1050.n2 a_9985_1050.t9 512.525
R2660 a_9985_1050.n0 a_9985_1050.t8 512.525
R2661 a_9985_1050.n2 a_9985_1050.t7 371.139
R2662 a_9985_1050.n0 a_9985_1050.t10 371.139
R2663 a_9985_1050.n1 a_9985_1050.t6 305.674
R2664 a_9985_1050.n3 a_9985_1050.t5 305.298
R2665 a_9985_1050.n3 a_9985_1050.n2 291.648
R2666 a_9985_1050.n1 a_9985_1050.n0 291.272
R2667 a_9985_1050.n9 a_9985_1050.n8 249.863
R2668 a_9985_1050.n11 a_9985_1050.n9 215.717
R2669 a_9985_1050.n11 a_9985_1050.n10 157.964
R2670 a_9985_1050.n12 a_9985_1050.n11 91.705
R2671 a_9985_1050.n8 a_9985_1050.n7 30
R2672 a_9985_1050.n6 a_9985_1050.n5 24.383
R2673 a_9985_1050.n8 a_9985_1050.n6 23.684
R2674 a_9985_1050.n10 a_9985_1050.t4 14.282
R2675 a_9985_1050.n10 a_9985_1050.t3 14.282
R2676 a_9985_1050.n12 a_9985_1050.t0 14.282
R2677 a_9985_1050.t1 a_9985_1050.n12 14.282
R2678 a_9985_1050.n4 a_9985_1050.n1 8.138
R2679 a_9985_1050.n9 a_9985_1050.n4 5.964
R2680 a_9985_1050.n4 a_9985_1050.n3 4.65
R2681 a_10525_103.t0 a_10525_103.n7 59.616
R2682 a_10525_103.n4 a_10525_103.n2 54.496
R2683 a_10525_103.n4 a_10525_103.n3 54.496
R2684 a_10525_103.n1 a_10525_103.n0 24.679
R2685 a_10525_103.n6 a_10525_103.n4 7.859
R2686 a_10525_103.t0 a_10525_103.n1 7.505
R2687 a_10525_103.t0 a_10525_103.n6 3.034
R2688 a_10525_103.n6 a_10525_103.n5 0.443
R2689 a_16096_101.n3 a_16096_101.n1 42.788
R2690 a_16096_101.t0 a_16096_101.n0 8.137
R2691 a_16096_101.n3 a_16096_101.n2 4.665
R2692 a_16096_101.t0 a_16096_101.n3 0.06
R2693 a_4996_101.n11 a_4996_101.n10 68.43
R2694 a_4996_101.n3 a_4996_101.n2 62.817
R2695 a_4996_101.n7 a_4996_101.n6 38.626
R2696 a_4996_101.n6 a_4996_101.n5 35.955
R2697 a_4996_101.n3 a_4996_101.n1 26.202
R2698 a_4996_101.t0 a_4996_101.n3 19.737
R2699 a_4996_101.t1 a_4996_101.n8 8.137
R2700 a_4996_101.t0 a_4996_101.n4 7.273
R2701 a_4996_101.t0 a_4996_101.n0 6.109
R2702 a_4996_101.t1 a_4996_101.n7 4.864
R2703 a_4996_101.t0 a_4996_101.n12 2.074
R2704 a_4996_101.n12 a_4996_101.t1 0.937
R2705 a_4996_101.t1 a_4996_101.n11 0.763
R2706 a_4996_101.n11 a_4996_101.n9 0.185
R2707 a_13367_411.n6 a_13367_411.t7 475.572
R2708 a_13367_411.n11 a_13367_411.t14 472.359
R2709 a_13367_411.n8 a_13367_411.t10 469.145
R2710 a_13367_411.n11 a_13367_411.t9 384.527
R2711 a_13367_411.n8 a_13367_411.t13 384.527
R2712 a_13367_411.n6 a_13367_411.t12 384.527
R2713 a_13367_411.n12 a_13367_411.t8 370.613
R2714 a_13367_411.n9 a_13367_411.t15 370.613
R2715 a_13367_411.n7 a_13367_411.t11 370.613
R2716 a_13367_411.n16 a_13367_411.n14 363.934
R2717 a_13367_411.n4 a_13367_411.n3 161.352
R2718 a_13367_411.n7 a_13367_411.n6 128.028
R2719 a_13367_411.n12 a_13367_411.n11 127.096
R2720 a_13367_411.n9 a_13367_411.n8 126.97
R2721 a_13367_411.n14 a_13367_411.n5 123.481
R2722 a_13367_411.n5 a_13367_411.n1 95.095
R2723 a_13367_411.n4 a_13367_411.n2 95.095
R2724 a_13367_411.n5 a_13367_411.n4 66.258
R2725 a_13367_411.n17 a_13367_411.n0 55.263
R2726 a_13367_411.n16 a_13367_411.n15 30
R2727 a_13367_411.n17 a_13367_411.n16 23.684
R2728 a_13367_411.n1 a_13367_411.t6 14.282
R2729 a_13367_411.n1 a_13367_411.t0 14.282
R2730 a_13367_411.n2 a_13367_411.t4 14.282
R2731 a_13367_411.n2 a_13367_411.t3 14.282
R2732 a_13367_411.n3 a_13367_411.t2 14.282
R2733 a_13367_411.n3 a_13367_411.t1 14.282
R2734 a_13367_411.n10 a_13367_411.n7 9.501
R2735 a_13367_411.n13 a_13367_411.n12 8.685
R2736 a_13367_411.n10 a_13367_411.n9 4.65
R2737 a_13367_411.n14 a_13367_411.n13 4.65
R2738 a_13367_411.n13 a_13367_411.n10 1.859
R2739 QN.n14 QN.n13 227.387
R2740 QN.n2 QN.n1 165.613
R2741 QN.n14 QN.n2 132.893
R2742 QN.n13 QN.n12 127.909
R2743 QN.n11 QN.n10 112.771
R2744 QN.n11 QN.n6 110.702
R2745 QN.n2 QN.n0 99.355
R2746 QN.n6 QN.n5 30
R2747 QN.n10 QN.n9 30
R2748 QN.n4 QN.n3 24.383
R2749 QN.n8 QN.n7 24.383
R2750 QN.n6 QN.n4 23.684
R2751 QN.n10 QN.n8 23.684
R2752 QN.n0 QN.t5 14.282
R2753 QN.n0 QN.t4 14.282
R2754 QN.n1 QN.t1 14.282
R2755 QN.n1 QN.t2 14.282
R2756 QN.n13 QN.n11 7.053
R2757 QN.n15 QN.n14 4.65
R2758 QN.n15 QN 0.046
R2759 a_6149_989.n3 a_6149_989.t5 454.685
R2760 a_6149_989.n5 a_6149_989.t7 454.685
R2761 a_6149_989.n1 a_6149_989.t10 454.685
R2762 a_6149_989.n3 a_6149_989.t12 428.979
R2763 a_6149_989.n5 a_6149_989.t13 428.979
R2764 a_6149_989.n1 a_6149_989.t8 428.979
R2765 a_6149_989.n12 a_6149_989.n11 348.963
R2766 a_6149_989.n4 a_6149_989.t11 339.542
R2767 a_6149_989.n6 a_6149_989.t9 339.542
R2768 a_6149_989.n2 a_6149_989.t6 339.542
R2769 a_6149_989.n14 a_6149_989.n13 157.963
R2770 a_6149_989.n4 a_6149_989.n3 143.429
R2771 a_6149_989.n6 a_6149_989.n5 143.429
R2772 a_6149_989.n2 a_6149_989.n1 143.429
R2773 a_6149_989.n13 a_6149_989.n12 132.141
R2774 a_6149_989.n13 a_6149_989.n0 91.706
R2775 a_6149_989.n11 a_6149_989.n9 22.578
R2776 a_6149_989.n0 a_6149_989.t2 14.282
R2777 a_6149_989.n0 a_6149_989.t3 14.282
R2778 a_6149_989.n14 a_6149_989.t0 14.282
R2779 a_6149_989.t1 a_6149_989.n14 14.282
R2780 a_6149_989.n8 a_6149_989.n2 10.046
R2781 a_6149_989.n11 a_6149_989.n10 8.58
R2782 a_6149_989.n7 a_6149_989.n6 8.141
R2783 a_6149_989.n7 a_6149_989.n4 4.65
R2784 a_6149_989.n12 a_6149_989.n8 4.65
R2785 a_6149_989.n8 a_6149_989.n7 2.947
R2786 a_11033_989.n2 a_11033_989.t6 454.685
R2787 a_11033_989.n4 a_11033_989.t11 454.685
R2788 a_11033_989.n0 a_11033_989.t13 454.685
R2789 a_11033_989.n2 a_11033_989.t5 428.979
R2790 a_11033_989.n4 a_11033_989.t7 428.979
R2791 a_11033_989.n0 a_11033_989.t9 428.979
R2792 a_11033_989.n3 a_11033_989.t12 339.542
R2793 a_11033_989.n5 a_11033_989.t10 339.542
R2794 a_11033_989.n1 a_11033_989.t8 339.542
R2795 a_11033_989.n12 a_11033_989.n11 333.44
R2796 a_11033_989.n14 a_11033_989.n13 157.964
R2797 a_11033_989.n3 a_11033_989.n2 143.429
R2798 a_11033_989.n5 a_11033_989.n4 143.429
R2799 a_11033_989.n1 a_11033_989.n0 143.429
R2800 a_11033_989.n14 a_11033_989.n12 132.141
R2801 a_11033_989.n15 a_11033_989.n14 91.705
R2802 a_11033_989.n11 a_11033_989.n10 30
R2803 a_11033_989.n9 a_11033_989.n8 24.383
R2804 a_11033_989.n11 a_11033_989.n9 23.684
R2805 a_11033_989.n13 a_11033_989.t0 14.282
R2806 a_11033_989.n13 a_11033_989.t1 14.282
R2807 a_11033_989.n15 a_11033_989.t2 14.282
R2808 a_11033_989.t3 a_11033_989.n15 14.282
R2809 a_11033_989.n7 a_11033_989.n1 10.046
R2810 a_11033_989.n6 a_11033_989.n5 8.141
R2811 a_11033_989.n6 a_11033_989.n3 4.65
R2812 a_11033_989.n12 a_11033_989.n7 4.65
R2813 a_11033_989.n7 a_11033_989.n6 2.947
R2814 a_11673_1050.n2 a_11673_1050.t7 480.392
R2815 a_11673_1050.n2 a_11673_1050.t9 403.272
R2816 a_11673_1050.n3 a_11673_1050.t8 301.486
R2817 a_11673_1050.n8 a_11673_1050.n7 252.498
R2818 a_11673_1050.n9 a_11673_1050.n8 234.917
R2819 a_11673_1050.n3 a_11673_1050.n2 227.006
R2820 a_11673_1050.n11 a_11673_1050.n10 161.352
R2821 a_11673_1050.n9 a_11673_1050.n1 95.095
R2822 a_11673_1050.n10 a_11673_1050.n0 95.095
R2823 a_11673_1050.n10 a_11673_1050.n9 66.258
R2824 a_11673_1050.n7 a_11673_1050.n6 30
R2825 a_11673_1050.n5 a_11673_1050.n4 24.383
R2826 a_11673_1050.n7 a_11673_1050.n5 23.684
R2827 a_11673_1050.n1 a_11673_1050.t6 14.282
R2828 a_11673_1050.n1 a_11673_1050.t5 14.282
R2829 a_11673_1050.n0 a_11673_1050.t1 14.282
R2830 a_11673_1050.n0 a_11673_1050.t0 14.282
R2831 a_11673_1050.t3 a_11673_1050.n11 14.282
R2832 a_11673_1050.n11 a_11673_1050.t2 14.282
R2833 a_11673_1050.n8 a_11673_1050.n3 10.615
R2834 a_2702_101.n11 a_2702_101.n10 68.43
R2835 a_2702_101.n3 a_2702_101.n2 62.817
R2836 a_2702_101.n7 a_2702_101.n6 38.626
R2837 a_2702_101.n6 a_2702_101.n5 35.955
R2838 a_2702_101.n3 a_2702_101.n1 26.202
R2839 a_2702_101.t0 a_2702_101.n3 19.737
R2840 a_2702_101.t1 a_2702_101.n8 8.137
R2841 a_2702_101.t0 a_2702_101.n4 7.273
R2842 a_2702_101.t0 a_2702_101.n0 6.109
R2843 a_2702_101.t1 a_2702_101.n7 4.864
R2844 a_2702_101.t0 a_2702_101.n12 2.074
R2845 a_2702_101.n12 a_2702_101.t1 0.937
R2846 a_2702_101.t1 a_2702_101.n11 0.763
R2847 a_2702_101.n11 a_2702_101.n9 0.185
R2848 a_9178_210.n10 a_9178_210.n8 171.558
R2849 a_9178_210.n8 a_9178_210.t1 75.764
R2850 a_9178_210.n11 a_9178_210.n0 49.6
R2851 a_9178_210.n3 a_9178_210.n2 27.476
R2852 a_9178_210.n10 a_9178_210.n9 27.2
R2853 a_9178_210.n11 a_9178_210.n10 22.4
R2854 a_9178_210.t1 a_9178_210.n5 20.241
R2855 a_9178_210.n7 a_9178_210.n6 19.952
R2856 a_9178_210.t1 a_9178_210.n3 13.984
R2857 a_9178_210.n5 a_9178_210.n4 13.494
R2858 a_9178_210.t1 a_9178_210.n1 7.04
R2859 a_9178_210.n8 a_9178_210.n7 1.505
R2860 a_8252_101.n3 a_8252_101.n1 42.788
R2861 a_8252_101.t0 a_8252_101.n0 8.137
R2862 a_8252_101.n3 a_8252_101.n2 4.665
R2863 a_8252_101.t0 a_8252_101.n3 0.06
R2864 a_13241_1050.n1 a_13241_1050.t5 512.525
R2865 a_13241_1050.n2 a_13241_1050.t7 445.142
R2866 a_13241_1050.n7 a_13241_1050.n6 389.157
R2867 a_13241_1050.n1 a_13241_1050.t6 371.139
R2868 a_13241_1050.n9 a_13241_1050.n8 157.963
R2869 a_13241_1050.n8 a_13241_1050.n0 91.706
R2870 a_13241_1050.n2 a_13241_1050.n1 85.101
R2871 a_13241_1050.n8 a_13241_1050.n7 76.423
R2872 a_13241_1050.n6 a_13241_1050.n5 30
R2873 a_13241_1050.n4 a_13241_1050.n3 24.383
R2874 a_13241_1050.n6 a_13241_1050.n4 23.684
R2875 a_13241_1050.n0 a_13241_1050.t3 14.282
R2876 a_13241_1050.n0 a_13241_1050.t4 14.282
R2877 a_13241_1050.n9 a_13241_1050.t0 14.282
R2878 a_13241_1050.t1 a_13241_1050.n9 14.282
R2879 a_13241_1050.n7 a_13241_1050.n2 8.044
R2880 SN.n14 SN.t16 479.223
R2881 SN.n11 SN.t7 479.223
R2882 SN.n8 SN.t8 479.223
R2883 SN.n5 SN.t15 479.223
R2884 SN.n2 SN.t4 479.223
R2885 SN.n0 SN.t3 479.223
R2886 SN.n14 SN.t9 375.52
R2887 SN.n11 SN.t17 375.52
R2888 SN.n8 SN.t10 375.52
R2889 SN.n5 SN.t2 375.52
R2890 SN.n2 SN.t13 375.52
R2891 SN.n0 SN.t12 375.52
R2892 SN.n15 SN.n14 252.188
R2893 SN.n12 SN.n11 252.188
R2894 SN.n9 SN.n8 252.188
R2895 SN.n6 SN.n5 252.188
R2896 SN.n3 SN.n2 252.188
R2897 SN.n1 SN.n0 252.188
R2898 SN.n15 SN.t14 231.854
R2899 SN.n12 SN.t1 231.854
R2900 SN.n9 SN.t0 231.854
R2901 SN.n6 SN.t6 231.854
R2902 SN.n3 SN.t5 231.854
R2903 SN.n1 SN.t11 231.854
R2904 SN.n4 SN.n1 13.038
R2905 SN.n7 SN.n4 9.476
R2906 SN.n13 SN.n10 9.476
R2907 SN.n10 SN.n7 8.388
R2908 SN.n16 SN.n13 8.388
R2909 SN.n4 SN.n3 4.65
R2910 SN.n7 SN.n6 4.65
R2911 SN.n10 SN.n9 4.65
R2912 SN.n13 SN.n12 4.65
R2913 SN.n16 SN.n15 4.65
R2914 SN.n16 SN 0.046
R2915 a_6603_103.t0 a_6603_103.n7 59.616
R2916 a_6603_103.n4 a_6603_103.n2 54.496
R2917 a_6603_103.n4 a_6603_103.n3 54.496
R2918 a_6603_103.n1 a_6603_103.n0 24.679
R2919 a_6603_103.n6 a_6603_103.n4 7.859
R2920 a_6603_103.t0 a_6603_103.n1 7.505
R2921 a_6603_103.t0 a_6603_103.n6 3.034
R2922 a_6603_103.n6 a_6603_103.n5 0.443
R2923 a_6884_210.n10 a_6884_210.n8 171.558
R2924 a_6884_210.n8 a_6884_210.t1 75.764
R2925 a_6884_210.n11 a_6884_210.n0 49.6
R2926 a_6884_210.n3 a_6884_210.n2 27.476
R2927 a_6884_210.n10 a_6884_210.n9 27.2
R2928 a_6884_210.n11 a_6884_210.n10 22.4
R2929 a_6884_210.t1 a_6884_210.n5 20.241
R2930 a_6884_210.n7 a_6884_210.n6 19.952
R2931 a_6884_210.t1 a_6884_210.n3 13.984
R2932 a_6884_210.n5 a_6884_210.n4 13.494
R2933 a_6884_210.t1 a_6884_210.n1 7.04
R2934 a_6884_210.n8 a_6884_210.n7 1.505
R2935 a_13136_101.n11 a_13136_101.n10 68.43
R2936 a_13136_101.n3 a_13136_101.n2 62.817
R2937 a_13136_101.n7 a_13136_101.n6 38.626
R2938 a_13136_101.n6 a_13136_101.n5 35.955
R2939 a_13136_101.n3 a_13136_101.n1 26.202
R2940 a_13136_101.t0 a_13136_101.n3 19.737
R2941 a_13136_101.t1 a_13136_101.n8 8.137
R2942 a_13136_101.t0 a_13136_101.n4 7.273
R2943 a_13136_101.t0 a_13136_101.n0 6.109
R2944 a_13136_101.t1 a_13136_101.n7 4.864
R2945 a_13136_101.t0 a_13136_101.n12 2.074
R2946 a_13136_101.n12 a_13136_101.t1 0.937
R2947 a_13136_101.t1 a_13136_101.n11 0.763
R2948 a_13136_101.n11 a_13136_101.n9 0.185
R2949 a_4013_103.n5 a_4013_103.n4 66.708
R2950 a_4013_103.n2 a_4013_103.n0 32.662
R2951 a_4013_103.n5 a_4013_103.n3 19.496
R2952 a_4013_103.t0 a_4013_103.n5 13.756
R2953 a_4013_103.t0 a_4013_103.n2 3.034
R2954 a_4013_103.n2 a_4013_103.n1 0.443
R2955 a_4294_210.n10 a_4294_210.n8 171.558
R2956 a_4294_210.n8 a_4294_210.t1 75.764
R2957 a_4294_210.n11 a_4294_210.n0 49.6
R2958 a_4294_210.n3 a_4294_210.n2 27.476
R2959 a_4294_210.n10 a_4294_210.n9 27.2
R2960 a_4294_210.n11 a_4294_210.n10 22.4
R2961 a_4294_210.t1 a_4294_210.n5 20.241
R2962 a_4294_210.n7 a_4294_210.n6 19.952
R2963 a_4294_210.t1 a_4294_210.n3 13.984
R2964 a_4294_210.n5 a_4294_210.n4 13.494
R2965 a_4294_210.t1 a_4294_210.n1 7.04
R2966 a_4294_210.n8 a_4294_210.n7 1.505
R2967 a_343_411.n2 a_343_411.t12 480.392
R2968 a_343_411.n4 a_343_411.t7 472.359
R2969 a_343_411.n3 a_343_411.t9 412.921
R2970 a_343_411.n2 a_343_411.t8 403.272
R2971 a_343_411.n4 a_343_411.t10 384.527
R2972 a_343_411.n5 a_343_411.t11 370.613
R2973 a_343_411.n11 a_343_411.n10 363.578
R2974 a_343_411.n14 a_343_411.n13 161.352
R2975 a_343_411.n5 a_343_411.n4 127.096
R2976 a_343_411.n12 a_343_411.n11 123.126
R2977 a_343_411.n3 a_343_411.n2 115.571
R2978 a_343_411.n12 a_343_411.n1 95.095
R2979 a_343_411.n13 a_343_411.n0 95.095
R2980 a_343_411.n13 a_343_411.n12 66.258
R2981 a_343_411.n10 a_343_411.n9 30
R2982 a_343_411.n8 a_343_411.n7 24.383
R2983 a_343_411.n10 a_343_411.n8 23.684
R2984 a_343_411.n1 a_343_411.t6 14.282
R2985 a_343_411.n1 a_343_411.t5 14.282
R2986 a_343_411.n0 a_343_411.t3 14.282
R2987 a_343_411.n0 a_343_411.t2 14.282
R2988 a_343_411.t1 a_343_411.n14 14.282
R2989 a_343_411.n14 a_343_411.t0 14.282
R2990 a_343_411.n6 a_343_411.n3 11.954
R2991 a_343_411.n6 a_343_411.n5 8.682
R2992 a_343_411.n11 a_343_411.n6 4.65
R2993 a_11487_103.t0 a_11487_103.n7 59.616
R2994 a_11487_103.n4 a_11487_103.n2 54.496
R2995 a_11487_103.n4 a_11487_103.n3 54.496
R2996 a_11487_103.n1 a_11487_103.n0 24.679
R2997 a_11487_103.n6 a_11487_103.n4 7.859
R2998 a_11487_103.t0 a_11487_103.n1 7.505
R2999 a_11487_103.t0 a_11487_103.n6 3.034
R3000 a_11487_103.n6 a_11487_103.n5 0.443
R3001 a_3473_1050.n0 a_3473_1050.t5 512.525
R3002 a_3473_1050.n1 a_3473_1050.t7 417.109
R3003 a_3473_1050.n0 a_3473_1050.t6 371.139
R3004 a_3473_1050.n6 a_3473_1050.n5 361.298
R3005 a_3473_1050.n1 a_3473_1050.n0 179.837
R3006 a_3473_1050.n8 a_3473_1050.n7 157.964
R3007 a_3473_1050.n8 a_3473_1050.n6 104.282
R3008 a_3473_1050.n9 a_3473_1050.n8 91.705
R3009 a_3473_1050.n5 a_3473_1050.n4 30
R3010 a_3473_1050.n3 a_3473_1050.n2 24.383
R3011 a_3473_1050.n5 a_3473_1050.n3 23.684
R3012 a_3473_1050.n7 a_3473_1050.t3 14.282
R3013 a_3473_1050.n7 a_3473_1050.t4 14.282
R3014 a_3473_1050.n9 a_3473_1050.t0 14.282
R3015 a_3473_1050.t1 a_3473_1050.n9 14.282
R3016 a_3473_1050.n6 a_3473_1050.n1 10.615
R3017 a_2000_210.n10 a_2000_210.n8 171.558
R3018 a_2000_210.n8 a_2000_210.t1 75.764
R3019 a_2000_210.n3 a_2000_210.n2 27.476
R3020 a_2000_210.n10 a_2000_210.n9 27.2
R3021 a_2000_210.n11 a_2000_210.n0 23.498
R3022 a_2000_210.n11 a_2000_210.n10 22.4
R3023 a_2000_210.t1 a_2000_210.n5 20.241
R3024 a_2000_210.n7 a_2000_210.n6 19.952
R3025 a_2000_210.t1 a_2000_210.n3 13.984
R3026 a_2000_210.n5 a_2000_210.n4 13.494
R3027 a_2000_210.t1 a_2000_210.n1 7.04
R3028 a_2000_210.n8 a_2000_210.n7 1.505
R3029 a_10806_210.n10 a_10806_210.n8 171.558
R3030 a_10806_210.n8 a_10806_210.t1 75.764
R3031 a_10806_210.n11 a_10806_210.n0 49.6
R3032 a_10806_210.n3 a_10806_210.n2 27.476
R3033 a_10806_210.n10 a_10806_210.n9 27.2
R3034 a_10806_210.n11 a_10806_210.n10 22.4
R3035 a_10806_210.t1 a_10806_210.n5 20.241
R3036 a_10806_210.n7 a_10806_210.n6 19.952
R3037 a_10806_210.t1 a_10806_210.n3 13.984
R3038 a_10806_210.n5 a_10806_210.n4 13.494
R3039 a_10806_210.t1 a_10806_210.n1 7.04
R3040 a_10806_210.n8 a_10806_210.n7 1.505
R3041 a_12470_101.n3 a_12470_101.n1 42.788
R3042 a_12470_101.t0 a_12470_101.n0 8.137
R3043 a_12470_101.n3 a_12470_101.n2 4.665
R3044 a_12470_101.t0 a_12470_101.n3 0.06
R3045 a_15430_101.n2 a_15430_101.n0 42.755
R3046 a_15430_101.n2 a_15430_101.n1 2.198
R3047 a_15430_101.t0 a_15430_101.n2 0.106
R3048 a_1038_210.n10 a_1038_210.n8 171.558
R3049 a_1038_210.n8 a_1038_210.t1 75.764
R3050 a_1038_210.n3 a_1038_210.n2 27.476
R3051 a_1038_210.n10 a_1038_210.n9 27.2
R3052 a_1038_210.n11 a_1038_210.n0 23.498
R3053 a_1038_210.n11 a_1038_210.n10 22.4
R3054 a_1038_210.t1 a_1038_210.n5 20.241
R3055 a_1038_210.n7 a_1038_210.n6 19.952
R3056 a_1038_210.t1 a_1038_210.n3 13.984
R3057 a_1038_210.n5 a_1038_210.n4 13.494
R3058 a_1038_210.t1 a_1038_210.n1 7.04
R3059 a_1038_210.n8 a_1038_210.n7 1.505
R3060 a_14062_210.n10 a_14062_210.n8 171.558
R3061 a_14062_210.n8 a_14062_210.t1 75.764
R3062 a_14062_210.n3 a_14062_210.n2 27.476
R3063 a_14062_210.n10 a_14062_210.n9 27.2
R3064 a_14062_210.n11 a_14062_210.n0 23.498
R3065 a_14062_210.n11 a_14062_210.n10 22.4
R3066 a_14062_210.t1 a_14062_210.n5 20.241
R3067 a_14062_210.n7 a_14062_210.n6 19.952
R3068 a_14062_210.t1 a_14062_210.n3 13.984
R3069 a_14062_210.n5 a_14062_210.n4 13.494
R3070 a_14062_210.t1 a_14062_210.n1 7.04
R3071 a_14062_210.n8 a_14062_210.n7 1.505
R3072 a_11768_210.n10 a_11768_210.n8 171.558
R3073 a_11768_210.n8 a_11768_210.t1 75.764
R3074 a_11768_210.n11 a_11768_210.n0 49.6
R3075 a_11768_210.n3 a_11768_210.n2 27.476
R3076 a_11768_210.n10 a_11768_210.n9 27.2
R3077 a_11768_210.n11 a_11768_210.n10 22.4
R3078 a_11768_210.t1 a_11768_210.n5 20.241
R3079 a_11768_210.n7 a_11768_210.n6 19.952
R3080 a_11768_210.t1 a_11768_210.n3 13.984
R3081 a_11768_210.n5 a_11768_210.n4 13.494
R3082 a_11768_210.t1 a_11768_210.n1 7.04
R3083 a_11768_210.n8 a_11768_210.n7 1.505
R3084 a_757_103.n5 a_757_103.n4 66.708
R3085 a_757_103.n2 a_757_103.n0 25.439
R3086 a_757_103.n5 a_757_103.n3 19.496
R3087 a_757_103.t0 a_757_103.n5 13.756
R3088 a_757_103.n2 a_757_103.n1 2.455
R3089 a_757_103.t0 a_757_103.n2 0.246
R3090 a_5922_210.n10 a_5922_210.n8 171.558
R3091 a_5922_210.n8 a_5922_210.t1 75.764
R3092 a_5922_210.n3 a_5922_210.n2 27.476
R3093 a_5922_210.n10 a_5922_210.n9 27.2
R3094 a_5922_210.n11 a_5922_210.n0 23.498
R3095 a_5922_210.n11 a_5922_210.n10 22.4
R3096 a_5922_210.t1 a_5922_210.n5 20.241
R3097 a_5922_210.n7 a_5922_210.n6 19.952
R3098 a_5922_210.t1 a_5922_210.n3 13.984
R3099 a_5922_210.n5 a_5922_210.n4 13.494
R3100 a_5922_210.t1 a_5922_210.n1 7.04
R3101 a_5922_210.n8 a_5922_210.n7 1.505
R3102 a_112_101.n11 a_112_101.n10 68.43
R3103 a_112_101.n3 a_112_101.n2 62.817
R3104 a_112_101.n7 a_112_101.n6 38.626
R3105 a_112_101.n6 a_112_101.n5 35.955
R3106 a_112_101.n3 a_112_101.n1 26.202
R3107 a_112_101.t0 a_112_101.n3 19.737
R3108 a_112_101.t1 a_112_101.n8 8.137
R3109 a_112_101.t0 a_112_101.n4 7.273
R3110 a_112_101.t0 a_112_101.n0 6.109
R3111 a_112_101.t1 a_112_101.n7 4.864
R3112 a_112_101.t0 a_112_101.n12 2.074
R3113 a_112_101.n12 a_112_101.t1 0.937
R3114 a_112_101.t1 a_112_101.n11 0.763
R3115 a_112_101.n11 a_112_101.n9 0.185
R3116 a_8897_103.n5 a_8897_103.n4 66.708
R3117 a_8897_103.n2 a_8897_103.n0 25.439
R3118 a_8897_103.n5 a_8897_103.n3 19.496
R3119 a_8897_103.t0 a_8897_103.n5 13.756
R3120 a_8897_103.n2 a_8897_103.n1 2.455
R3121 a_8897_103.t0 a_8897_103.n2 0.246
R3122 a_3368_101.n3 a_3368_101.n1 42.788
R3123 a_3368_101.t0 a_3368_101.n0 8.137
R3124 a_3368_101.n3 a_3368_101.n2 4.665
R3125 a_3368_101.t0 a_3368_101.n3 0.06
R3126 a_9880_101.n3 a_9880_101.n1 42.788
R3127 a_9880_101.t0 a_9880_101.n0 8.137
R3128 a_9880_101.n3 a_9880_101.n2 4.665
R3129 a_9880_101.t0 a_9880_101.n3 0.06
R3130 a_1719_103.t0 a_1719_103.n7 59.616
R3131 a_1719_103.n4 a_1719_103.n2 54.496
R3132 a_1719_103.n4 a_1719_103.n3 54.496
R3133 a_1719_103.n1 a_1719_103.n0 24.679
R3134 a_1719_103.t0 a_1719_103.n1 7.505
R3135 a_1719_103.n6 a_1719_103.n5 2.455
R3136 a_1719_103.n6 a_1719_103.n4 0.636
R3137 a_1719_103.t0 a_1719_103.n6 0.246
R3138 a_13781_103.t0 a_13781_103.n7 59.616
R3139 a_13781_103.n4 a_13781_103.n2 54.496
R3140 a_13781_103.n4 a_13781_103.n3 54.496
R3141 a_13781_103.n1 a_13781_103.n0 24.679
R3142 a_13781_103.t0 a_13781_103.n1 7.505
R3143 a_13781_103.n6 a_13781_103.n5 2.455
R3144 a_13781_103.n6 a_13781_103.n4 0.636
R3145 a_13781_103.t0 a_13781_103.n6 0.246
R3146 a_5641_103.n5 a_5641_103.n4 66.708
R3147 a_5641_103.n2 a_5641_103.n0 25.439
R3148 a_5641_103.n5 a_5641_103.n3 19.496
R3149 a_5641_103.t0 a_5641_103.n5 13.756
R3150 a_5641_103.n2 a_5641_103.n1 2.455
R3151 a_5641_103.t0 a_5641_103.n2 0.246
R3152 a_14764_101.n3 a_14764_101.n2 62.817
R3153 a_14764_101.n11 a_14764_101.n10 46.054
R3154 a_14764_101.n7 a_14764_101.n6 38.626
R3155 a_14764_101.n6 a_14764_101.n5 35.955
R3156 a_14764_101.n12 a_14764_101.n11 27.923
R3157 a_14764_101.n3 a_14764_101.n1 26.202
R3158 a_14764_101.t0 a_14764_101.n3 19.737
R3159 a_14764_101.t0 a_14764_101.n4 7.273
R3160 a_14764_101.n9 a_14764_101.n8 6.883
R3161 a_14764_101.t0 a_14764_101.n0 6.109
R3162 a_14764_101.t1 a_14764_101.n7 4.864
R3163 a_14764_101.t0 a_14764_101.n13 2.074
R3164 a_14764_101.t1 a_14764_101.n9 1.179
R3165 a_14764_101.t1 a_14764_101.n12 0.958
R3166 a_14764_101.n13 a_14764_101.t1 0.937
C7 SN GND 6.35fF
C8 VDD GND 27.09fF
C9 a_14764_101.n0 GND 0.02fF
C10 a_14764_101.n1 GND 0.09fF
C11 a_14764_101.n2 GND 0.07fF
C12 a_14764_101.n3 GND 0.03fF
C13 a_14764_101.n4 GND 0.01fF
C14 a_14764_101.n5 GND 0.03fF
C15 a_14764_101.n6 GND 0.04fF
C16 a_14764_101.n7 GND 0.02fF
C17 a_14764_101.n8 GND 0.04fF
C18 a_14764_101.n9 GND 0.08fF
C19 a_14764_101.n10 GND 0.04fF
C20 a_14764_101.n11 GND 0.12fF
C21 a_14764_101.n12 GND 0.14fF
C22 a_14764_101.n13 GND 0.01fF
C23 a_5641_103.n0 GND 0.11fF
C24 a_5641_103.n1 GND 0.04fF
C25 a_5641_103.n2 GND 0.03fF
C26 a_5641_103.n3 GND 0.07fF
C27 a_5641_103.n4 GND 0.08fF
C28 a_5641_103.n5 GND 0.03fF
C29 a_13781_103.n0 GND 0.08fF
C30 a_13781_103.n1 GND 0.07fF
C31 a_13781_103.n2 GND 0.04fF
C32 a_13781_103.n3 GND 0.06fF
C33 a_13781_103.n4 GND 0.03fF
C34 a_13781_103.n5 GND 0.04fF
C35 a_13781_103.n7 GND 0.08fF
C36 a_1719_103.n0 GND 0.08fF
C37 a_1719_103.n1 GND 0.07fF
C38 a_1719_103.n2 GND 0.04fF
C39 a_1719_103.n3 GND 0.06fF
C40 a_1719_103.n4 GND 0.03fF
C41 a_1719_103.n5 GND 0.04fF
C42 a_1719_103.n7 GND 0.08fF
C43 a_9880_101.n0 GND 0.05fF
C44 a_9880_101.n1 GND 0.12fF
C45 a_9880_101.n2 GND 0.04fF
C46 a_9880_101.n3 GND 0.17fF
C47 a_3368_101.n0 GND 0.05fF
C48 a_3368_101.n1 GND 0.12fF
C49 a_3368_101.n2 GND 0.04fF
C50 a_3368_101.n3 GND 0.17fF
C51 a_8897_103.n0 GND 0.11fF
C52 a_8897_103.n1 GND 0.04fF
C53 a_8897_103.n2 GND 0.03fF
C54 a_8897_103.n3 GND 0.07fF
C55 a_8897_103.n4 GND 0.08fF
C56 a_8897_103.n5 GND 0.03fF
C57 a_112_101.n0 GND 0.02fF
C58 a_112_101.n1 GND 0.09fF
C59 a_112_101.n2 GND 0.08fF
C60 a_112_101.n3 GND 0.03fF
C61 a_112_101.n4 GND 0.01fF
C62 a_112_101.n5 GND 0.04fF
C63 a_112_101.n6 GND 0.04fF
C64 a_112_101.n7 GND 0.02fF
C65 a_112_101.n8 GND 0.05fF
C66 a_112_101.n9 GND 0.14fF
C67 a_112_101.n10 GND 0.08fF
C68 a_112_101.n11 GND 0.08fF
C69 a_112_101.t1 GND 0.22fF
C70 a_112_101.n12 GND 0.01fF
C71 a_5922_210.n0 GND 0.02fF
C72 a_5922_210.n1 GND 0.09fF
C73 a_5922_210.n2 GND 0.12fF
C74 a_5922_210.n3 GND 0.08fF
C75 a_5922_210.n4 GND 0.08fF
C76 a_5922_210.n5 GND 0.02fF
C77 a_5922_210.t1 GND 0.29fF
C78 a_5922_210.n6 GND 0.09fF
C79 a_5922_210.n7 GND 0.02fF
C80 a_5922_210.n8 GND 0.13fF
C81 a_5922_210.n9 GND 0.02fF
C82 a_5922_210.n10 GND 0.03fF
C83 a_5922_210.n11 GND 0.03fF
C84 a_757_103.n0 GND 0.11fF
C85 a_757_103.n1 GND 0.04fF
C86 a_757_103.n2 GND 0.03fF
C87 a_757_103.n3 GND 0.07fF
C88 a_757_103.n4 GND 0.08fF
C89 a_757_103.n5 GND 0.03fF
C90 a_11768_210.n0 GND 0.02fF
C91 a_11768_210.n1 GND 0.09fF
C92 a_11768_210.n2 GND 0.12fF
C93 a_11768_210.n3 GND 0.08fF
C94 a_11768_210.n4 GND 0.08fF
C95 a_11768_210.n5 GND 0.02fF
C96 a_11768_210.t1 GND 0.29fF
C97 a_11768_210.n6 GND 0.09fF
C98 a_11768_210.n7 GND 0.02fF
C99 a_11768_210.n8 GND 0.13fF
C100 a_11768_210.n9 GND 0.02fF
C101 a_11768_210.n10 GND 0.03fF
C102 a_11768_210.n11 GND 0.02fF
C103 a_14062_210.n0 GND 0.02fF
C104 a_14062_210.n1 GND 0.09fF
C105 a_14062_210.n2 GND 0.12fF
C106 a_14062_210.n3 GND 0.08fF
C107 a_14062_210.n4 GND 0.08fF
C108 a_14062_210.n5 GND 0.02fF
C109 a_14062_210.t1 GND 0.29fF
C110 a_14062_210.n6 GND 0.09fF
C111 a_14062_210.n7 GND 0.02fF
C112 a_14062_210.n8 GND 0.13fF
C113 a_14062_210.n9 GND 0.02fF
C114 a_14062_210.n10 GND 0.03fF
C115 a_14062_210.n11 GND 0.03fF
C116 a_1038_210.n0 GND 0.02fF
C117 a_1038_210.n1 GND 0.09fF
C118 a_1038_210.n2 GND 0.12fF
C119 a_1038_210.n3 GND 0.08fF
C120 a_1038_210.n4 GND 0.08fF
C121 a_1038_210.n5 GND 0.02fF
C122 a_1038_210.t1 GND 0.29fF
C123 a_1038_210.n6 GND 0.09fF
C124 a_1038_210.n7 GND 0.02fF
C125 a_1038_210.n8 GND 0.13fF
C126 a_1038_210.n9 GND 0.02fF
C127 a_1038_210.n10 GND 0.03fF
C128 a_1038_210.n11 GND 0.03fF
C129 a_15430_101.n0 GND 0.13fF
C130 a_15430_101.n1 GND 0.14fF
C131 a_15430_101.n2 GND 0.14fF
C132 a_12470_101.n0 GND 0.05fF
C133 a_12470_101.n1 GND 0.12fF
C134 a_12470_101.n2 GND 0.04fF
C135 a_12470_101.n3 GND 0.17fF
C136 a_10806_210.n0 GND 0.02fF
C137 a_10806_210.n1 GND 0.09fF
C138 a_10806_210.n2 GND 0.12fF
C139 a_10806_210.n3 GND 0.08fF
C140 a_10806_210.n4 GND 0.08fF
C141 a_10806_210.n5 GND 0.02fF
C142 a_10806_210.t1 GND 0.29fF
C143 a_10806_210.n6 GND 0.09fF
C144 a_10806_210.n7 GND 0.02fF
C145 a_10806_210.n8 GND 0.13fF
C146 a_10806_210.n9 GND 0.02fF
C147 a_10806_210.n10 GND 0.03fF
C148 a_10806_210.n11 GND 0.02fF
C149 a_2000_210.n0 GND 0.02fF
C150 a_2000_210.n1 GND 0.09fF
C151 a_2000_210.n2 GND 0.12fF
C152 a_2000_210.n3 GND 0.08fF
C153 a_2000_210.n4 GND 0.08fF
C154 a_2000_210.n5 GND 0.02fF
C155 a_2000_210.t1 GND 0.29fF
C156 a_2000_210.n6 GND 0.09fF
C157 a_2000_210.n7 GND 0.02fF
C158 a_2000_210.n8 GND 0.13fF
C159 a_2000_210.n9 GND 0.02fF
C160 a_2000_210.n10 GND 0.03fF
C161 a_2000_210.n11 GND 0.03fF
C162 a_3473_1050.n0 GND 0.29fF
C163 a_3473_1050.n1 GND 0.67fF
C164 a_3473_1050.n2 GND 0.04fF
C165 a_3473_1050.n3 GND 0.06fF
C166 a_3473_1050.n4 GND 0.04fF
C167 a_3473_1050.n5 GND 0.29fF
C168 a_3473_1050.n6 GND 0.70fF
C169 a_3473_1050.n7 GND 0.51fF
C170 a_3473_1050.n8 GND 0.53fF
C171 a_3473_1050.n9 GND 0.40fF
C172 a_11487_103.n0 GND 0.08fF
C173 a_11487_103.n1 GND 0.07fF
C174 a_11487_103.n2 GND 0.04fF
C175 a_11487_103.n3 GND 0.06fF
C176 a_11487_103.n4 GND 0.11fF
C177 a_11487_103.n5 GND 0.04fF
C178 a_11487_103.n7 GND 0.08fF
C179 a_343_411.n0 GND 0.57fF
C180 a_343_411.n1 GND 0.57fF
C181 a_343_411.n2 GND 0.41fF
C182 a_343_411.n3 GND 1.38fF
C183 a_343_411.n4 GND 0.40fF
C184 a_343_411.t11 GND 0.84fF
C185 a_343_411.n5 GND 0.89fF
C186 a_343_411.n6 GND 2.70fF
C187 a_343_411.n7 GND 0.06fF
C188 a_343_411.n8 GND 0.08fF
C189 a_343_411.n9 GND 0.05fF
C190 a_343_411.n10 GND 0.41fF
C191 a_343_411.n11 GND 0.77fF
C192 a_343_411.n12 GND 0.56fF
C193 a_343_411.n13 GND 0.69fF
C194 a_343_411.n14 GND 0.72fF
C195 a_4294_210.n0 GND 0.02fF
C196 a_4294_210.n1 GND 0.09fF
C197 a_4294_210.n2 GND 0.12fF
C198 a_4294_210.n3 GND 0.08fF
C199 a_4294_210.n4 GND 0.08fF
C200 a_4294_210.n5 GND 0.02fF
C201 a_4294_210.t1 GND 0.29fF
C202 a_4294_210.n6 GND 0.09fF
C203 a_4294_210.n7 GND 0.02fF
C204 a_4294_210.n8 GND 0.13fF
C205 a_4294_210.n9 GND 0.02fF
C206 a_4294_210.n10 GND 0.03fF
C207 a_4294_210.n11 GND 0.02fF
C208 a_4013_103.n0 GND 0.13fF
C209 a_4013_103.n1 GND 0.04fF
C210 a_4013_103.n2 GND 0.09fF
C211 a_4013_103.n3 GND 0.07fF
C212 a_4013_103.n4 GND 0.08fF
C213 a_4013_103.n5 GND 0.03fF
C214 a_13136_101.n0 GND 0.02fF
C215 a_13136_101.n1 GND 0.09fF
C216 a_13136_101.n2 GND 0.08fF
C217 a_13136_101.n3 GND 0.03fF
C218 a_13136_101.n4 GND 0.01fF
C219 a_13136_101.n5 GND 0.04fF
C220 a_13136_101.n6 GND 0.04fF
C221 a_13136_101.n7 GND 0.02fF
C222 a_13136_101.n8 GND 0.05fF
C223 a_13136_101.n9 GND 0.15fF
C224 a_13136_101.n10 GND 0.08fF
C225 a_13136_101.n11 GND 0.08fF
C226 a_13136_101.t1 GND 0.23fF
C227 a_13136_101.n12 GND 0.01fF
C228 a_6884_210.n0 GND 0.02fF
C229 a_6884_210.n1 GND 0.09fF
C230 a_6884_210.n2 GND 0.12fF
C231 a_6884_210.n3 GND 0.08fF
C232 a_6884_210.n4 GND 0.08fF
C233 a_6884_210.n5 GND 0.02fF
C234 a_6884_210.t1 GND 0.29fF
C235 a_6884_210.n6 GND 0.09fF
C236 a_6884_210.n7 GND 0.02fF
C237 a_6884_210.n8 GND 0.13fF
C238 a_6884_210.n9 GND 0.02fF
C239 a_6884_210.n10 GND 0.03fF
C240 a_6884_210.n11 GND 0.02fF
C241 a_6603_103.n0 GND 0.08fF
C242 a_6603_103.n1 GND 0.07fF
C243 a_6603_103.n2 GND 0.04fF
C244 a_6603_103.n3 GND 0.06fF
C245 a_6603_103.n4 GND 0.11fF
C246 a_6603_103.n5 GND 0.04fF
C247 a_6603_103.n7 GND 0.08fF
C248 SN.n0 GND 0.76fF
C249 SN.t11 GND 0.83fF
C250 SN.n1 GND 1.82fF
C251 SN.n2 GND 0.76fF
C252 SN.t5 GND 0.83fF
C253 SN.n3 GND 0.71fF
C254 SN.n4 GND 4.21fF
C255 SN.n5 GND 0.76fF
C256 SN.t6 GND 0.83fF
C257 SN.n6 GND 0.71fF
C258 SN.n7 GND 3.60fF
C259 SN.n8 GND 0.76fF
C260 SN.t0 GND 0.83fF
C261 SN.n9 GND 0.71fF
C262 SN.n10 GND 3.60fF
C263 SN.n11 GND 0.76fF
C264 SN.t1 GND 0.83fF
C265 SN.n12 GND 0.71fF
C266 SN.n13 GND 3.60fF
C267 SN.n14 GND 0.76fF
C268 SN.t14 GND 0.83fF
C269 SN.n15 GND 0.71fF
C270 SN.n16 GND 1.71fF
C271 a_13241_1050.n0 GND 0.36fF
C272 a_13241_1050.n1 GND 0.22fF
C273 a_13241_1050.n2 GND 0.70fF
C274 a_13241_1050.n3 GND 0.04fF
C275 a_13241_1050.n4 GND 0.05fF
C276 a_13241_1050.n5 GND 0.03fF
C277 a_13241_1050.n6 GND 0.30fF
C278 a_13241_1050.n7 GND 0.59fF
C279 a_13241_1050.n8 GND 0.46fF
C280 a_13241_1050.n9 GND 0.47fF
C281 a_8252_101.n0 GND 0.05fF
C282 a_8252_101.n1 GND 0.12fF
C283 a_8252_101.n2 GND 0.04fF
C284 a_8252_101.n3 GND 0.17fF
C285 a_9178_210.n0 GND 0.02fF
C286 a_9178_210.n1 GND 0.09fF
C287 a_9178_210.n2 GND 0.12fF
C288 a_9178_210.n3 GND 0.08fF
C289 a_9178_210.n4 GND 0.08fF
C290 a_9178_210.n5 GND 0.02fF
C291 a_9178_210.t1 GND 0.29fF
C292 a_9178_210.n6 GND 0.09fF
C293 a_9178_210.n7 GND 0.02fF
C294 a_9178_210.n8 GND 0.13fF
C295 a_9178_210.n9 GND 0.02fF
C296 a_9178_210.n10 GND 0.03fF
C297 a_9178_210.n11 GND 0.02fF
C298 a_2702_101.n0 GND 0.02fF
C299 a_2702_101.n1 GND 0.09fF
C300 a_2702_101.n2 GND 0.08fF
C301 a_2702_101.n3 GND 0.03fF
C302 a_2702_101.n4 GND 0.01fF
C303 a_2702_101.n5 GND 0.04fF
C304 a_2702_101.n6 GND 0.04fF
C305 a_2702_101.n7 GND 0.02fF
C306 a_2702_101.n8 GND 0.05fF
C307 a_2702_101.n9 GND 0.15fF
C308 a_2702_101.n10 GND 0.08fF
C309 a_2702_101.n11 GND 0.08fF
C310 a_2702_101.t1 GND 0.23fF
C311 a_2702_101.n12 GND 0.01fF
C312 a_11673_1050.n0 GND 0.39fF
C313 a_11673_1050.n1 GND 0.39fF
C314 a_11673_1050.n2 GND 0.38fF
C315 a_11673_1050.n3 GND 0.59fF
C316 a_11673_1050.n4 GND 0.04fF
C317 a_11673_1050.n5 GND 0.05fF
C318 a_11673_1050.n6 GND 0.03fF
C319 a_11673_1050.n7 GND 0.17fF
C320 a_11673_1050.n8 GND 0.69fF
C321 a_11673_1050.n9 GND 0.51fF
C322 a_11673_1050.n10 GND 0.47fF
C323 a_11673_1050.n11 GND 0.49fF
C324 a_11033_989.n0 GND 0.52fF
C325 a_11033_989.t8 GND 0.94fF
C326 a_11033_989.n1 GND 1.27fF
C327 a_11033_989.n2 GND 0.52fF
C328 a_11033_989.t12 GND 0.93fF
C329 a_11033_989.n3 GND 0.70fF
C330 a_11033_989.n4 GND 0.52fF
C331 a_11033_989.t10 GND 0.94fF
C332 a_11033_989.n5 GND 1.00fF
C333 a_11033_989.n6 GND 1.65fF
C334 a_11033_989.n7 GND 2.09fF
C335 a_11033_989.n8 GND 0.07fF
C336 a_11033_989.n9 GND 0.09fF
C337 a_11033_989.n10 GND 0.06fF
C338 a_11033_989.n11 GND 0.43fF
C339 a_11033_989.n12 GND 0.84fF
C340 a_11033_989.n13 GND 0.84fF
C341 a_11033_989.n14 GND 0.93fF
C342 a_11033_989.n15 GND 0.65fF
C343 a_6149_989.n0 GND 0.58fF
C344 a_6149_989.n1 GND 0.46fF
C345 a_6149_989.t6 GND 0.83fF
C346 a_6149_989.n2 GND 1.13fF
C347 a_6149_989.n3 GND 0.46fF
C348 a_6149_989.t11 GND 0.83fF
C349 a_6149_989.n4 GND 0.62fF
C350 a_6149_989.n5 GND 0.46fF
C351 a_6149_989.t9 GND 0.83fF
C352 a_6149_989.n6 GND 0.89fF
C353 a_6149_989.n7 GND 1.46fF
C354 a_6149_989.n8 GND 1.85fF
C355 a_6149_989.n9 GND 0.11fF
C356 a_6149_989.n10 GND 0.04fF
C357 a_6149_989.n11 GND 0.41fF
C358 a_6149_989.n12 GND 0.77fF
C359 a_6149_989.n13 GND 0.82fF
C360 a_6149_989.n14 GND 0.74fF
C361 QN.n0 GND 0.30fF
C362 QN.n1 GND 0.38fF
C363 QN.n2 GND 0.46fF
C364 QN.n3 GND 0.04fF
C365 QN.n4 GND 0.05fF
C366 QN.n5 GND 0.03fF
C367 QN.n6 GND 0.03fF
C368 QN.n7 GND 0.04fF
C369 QN.n8 GND 0.05fF
C370 QN.n9 GND 0.03fF
C371 QN.n10 GND 0.04fF
C372 QN.n11 GND 1.05fF
C373 QN.n12 GND 0.14fF
C374 QN.n13 GND 0.38fF
C375 QN.n14 GND 0.35fF
C376 QN.n15 GND 0.01fF
C377 a_13367_411.n0 GND 0.05fF
C378 a_13367_411.n1 GND 0.45fF
C379 a_13367_411.n2 GND 0.45fF
C380 a_13367_411.n3 GND 0.57fF
C381 a_13367_411.n4 GND 0.54fF
C382 a_13367_411.n5 GND 0.44fF
C383 a_13367_411.n6 GND 0.33fF
C384 a_13367_411.n7 GND 0.82fF
C385 a_13367_411.n8 GND 0.32fF
C386 a_13367_411.n9 GND 0.44fF
C387 a_13367_411.n10 GND 1.19fF
C388 a_13367_411.n11 GND 0.32fF
C389 a_13367_411.t8 GND 0.66fF
C390 a_13367_411.n12 GND 0.70fF
C391 a_13367_411.n13 GND 1.06fF
C392 a_13367_411.n14 GND 0.60fF
C393 a_13367_411.n15 GND 0.05fF
C394 a_13367_411.n16 GND 0.32fF
C395 a_13367_411.n17 GND 0.05fF
C396 a_4996_101.n0 GND 0.02fF
C397 a_4996_101.n1 GND 0.09fF
C398 a_4996_101.n2 GND 0.08fF
C399 a_4996_101.n3 GND 0.03fF
C400 a_4996_101.n4 GND 0.01fF
C401 a_4996_101.n5 GND 0.04fF
C402 a_4996_101.n6 GND 0.04fF
C403 a_4996_101.n7 GND 0.02fF
C404 a_4996_101.n8 GND 0.05fF
C405 a_4996_101.n9 GND 0.15fF
C406 a_4996_101.n10 GND 0.08fF
C407 a_4996_101.n11 GND 0.08fF
C408 a_4996_101.t1 GND 0.23fF
C409 a_4996_101.n12 GND 0.01fF
C410 a_16096_101.n0 GND 0.05fF
C411 a_16096_101.n1 GND 0.13fF
C412 a_16096_101.n2 GND 0.04fF
C413 a_16096_101.n3 GND 0.18fF
C414 a_10525_103.n0 GND 0.08fF
C415 a_10525_103.n1 GND 0.07fF
C416 a_10525_103.n2 GND 0.04fF
C417 a_10525_103.n3 GND 0.06fF
C418 a_10525_103.n4 GND 0.11fF
C419 a_10525_103.n5 GND 0.04fF
C420 a_10525_103.n7 GND 0.08fF
C421 a_9985_1050.n0 GND 0.49fF
C422 a_9985_1050.n1 GND 0.84fF
C423 a_9985_1050.n2 GND 0.49fF
C424 a_9985_1050.n3 GND 0.61fF
C425 a_9985_1050.n4 GND 1.21fF
C426 a_9985_1050.n5 GND 0.05fF
C427 a_9985_1050.n6 GND 0.07fF
C428 a_9985_1050.n7 GND 0.04fF
C429 a_9985_1050.n8 GND 0.22fF
C430 a_9985_1050.n9 GND 0.69fF
C431 a_9985_1050.n10 GND 0.64fF
C432 a_9985_1050.n11 GND 0.83fF
C433 a_9985_1050.n12 GND 0.50fF
C434 a_10111_411.n0 GND 0.67fF
C435 a_10111_411.n1 GND 0.48fF
C436 a_10111_411.n2 GND 1.62fF
C437 a_10111_411.n3 GND 0.48fF
C438 a_10111_411.t10 GND 0.99fF
C439 a_10111_411.n4 GND 1.05fF
C440 a_10111_411.n5 GND 3.19fF
C441 a_10111_411.n6 GND 0.07fF
C442 a_10111_411.n7 GND 0.09fF
C443 a_10111_411.n8 GND 0.52fF
C444 a_10111_411.n9 GND 0.93fF
C445 a_10111_411.n10 GND 0.66fF
C446 a_10111_411.n11 GND 0.85fF
C447 a_10111_411.n12 GND 0.81fF
C448 a_10111_411.n13 GND 0.67fF
C449 a_1905_1050.n0 GND 0.35fF
C450 a_1905_1050.n1 GND 0.35fF
C451 a_1905_1050.n2 GND 0.35fF
C452 a_1905_1050.n3 GND 0.54fF
C453 a_1905_1050.n4 GND 0.04fF
C454 a_1905_1050.n5 GND 0.05fF
C455 a_1905_1050.n6 GND 0.03fF
C456 a_1905_1050.n7 GND 0.15fF
C457 a_1905_1050.n8 GND 0.63fF
C458 a_1905_1050.n9 GND 0.46fF
C459 a_1905_1050.n10 GND 0.43fF
C460 a_1905_1050.n11 GND 0.45fF
C461 a_1265_989.n0 GND 0.39fF
C462 a_1265_989.t12 GND 0.71fF
C463 a_1265_989.n1 GND 0.96fF
C464 a_1265_989.n2 GND 0.39fF
C465 a_1265_989.t7 GND 0.70fF
C466 a_1265_989.n3 GND 0.53fF
C467 a_1265_989.n4 GND 0.39fF
C468 a_1265_989.t8 GND 0.71fF
C469 a_1265_989.n5 GND 0.76fF
C470 a_1265_989.n6 GND 1.24fF
C471 a_1265_989.n7 GND 1.58fF
C472 a_1265_989.n8 GND 0.05fF
C473 a_1265_989.n9 GND 0.07fF
C474 a_1265_989.n10 GND 0.04fF
C475 a_1265_989.n11 GND 0.32fF
C476 a_1265_989.n12 GND 0.64fF
C477 a_1265_989.n13 GND 0.63fF
C478 a_1265_989.n14 GND 0.70fF
C479 a_1265_989.n15 GND 0.49fF
C480 a_217_1050.n0 GND 0.32fF
C481 a_217_1050.n1 GND 0.32fF
C482 a_217_1050.n2 GND 0.55fF
C483 a_217_1050.n3 GND 0.32fF
C484 a_217_1050.n4 GND 0.39fF
C485 a_217_1050.n5 GND 0.79fF
C486 a_217_1050.n6 GND 0.23fF
C487 a_217_1050.n7 GND 0.46fF
C488 a_217_1050.n8 GND 0.54fF
C489 a_217_1050.n9 GND 0.42fF
C490 a_14869_1051.n0 GND 0.36fF
C491 a_14869_1051.n1 GND 0.32fF
C492 a_14869_1051.n2 GND 0.52fF
C493 a_14869_1051.n3 GND 0.30fF
C494 a_14869_1051.n4 GND 0.80fF
C495 a_14869_1051.n5 GND 0.43fF
C496 a_15533_1051.n0 GND 0.28fF
C497 a_15533_1051.n1 GND 0.36fF
C498 a_15533_1051.n2 GND 0.70fF
C499 a_15533_1051.n3 GND 0.27fF
C500 a_15533_1051.n4 GND 0.45fF
C501 a_15533_1051.n5 GND 0.28fF
C502 a_3599_411.n0 GND 0.08fF
C503 a_3599_411.n1 GND 0.75fF
C504 a_3599_411.n2 GND 0.75fF
C505 a_3599_411.n3 GND 0.96fF
C506 a_3599_411.n4 GND 0.91fF
C507 a_3599_411.n5 GND 0.92fF
C508 a_3599_411.n6 GND 0.70fF
C509 a_3599_411.n7 GND 0.85fF
C510 a_3599_411.n8 GND 1.18fF
C511 a_3599_411.n9 GND 0.70fF
C512 a_3599_411.n10 GND 8.46fF
C513 a_3599_411.n11 GND 0.65fF
C514 a_3599_411.t14 GND 0.98fF
C515 a_3599_411.n12 GND 1.19fF
C516 a_3599_411.n13 GND 10.95fF
C517 a_3599_411.n14 GND 1.00fF
C518 a_3599_411.n15 GND 0.08fF
C519 a_3599_411.n16 GND 0.38fF
C520 a_3599_411.n17 GND 0.09fF
C521 a_5227_411.n0 GND 0.65fF
C522 a_5227_411.n1 GND 0.65fF
C523 a_5227_411.n2 GND 0.47fF
C524 a_5227_411.n3 GND 1.57fF
C525 a_5227_411.n4 GND 0.46fF
C526 a_5227_411.t9 GND 0.96fF
C527 a_5227_411.n5 GND 1.02fF
C528 a_5227_411.n6 GND 3.09fF
C529 a_5227_411.n7 GND 0.07fF
C530 a_5227_411.n8 GND 0.09fF
C531 a_5227_411.n9 GND 0.50fF
C532 a_5227_411.n10 GND 0.90fF
C533 a_5227_411.n11 GND 0.64fF
C534 a_5227_411.n12 GND 0.78fF
C535 a_5227_411.n13 GND 0.83fF
C536 a_5101_1050.n0 GND 0.51fF
C537 a_5101_1050.n1 GND 0.49fF
C538 a_5101_1050.n2 GND 0.85fF
C539 a_5101_1050.n3 GND 0.49fF
C540 a_5101_1050.n4 GND 0.62fF
C541 a_5101_1050.n5 GND 1.22fF
C542 a_5101_1050.n6 GND 0.36fF
C543 a_5101_1050.n7 GND 0.72fF
C544 a_5101_1050.n8 GND 0.84fF
C545 a_5101_1050.n9 GND 0.65fF
C546 a_7586_101.n0 GND 0.05fF
C547 a_7586_101.n1 GND 0.02fF
C548 a_7586_101.n2 GND 0.12fF
C549 a_7586_101.n3 GND 0.04fF
C550 a_7586_101.n4 GND 0.17fF
C551 a_6789_1050.n0 GND 0.39fF
C552 a_6789_1050.n1 GND 0.39fF
C553 a_6789_1050.n2 GND 0.50fF
C554 a_6789_1050.n3 GND 0.47fF
C555 a_6789_1050.n4 GND 0.51fF
C556 a_6789_1050.n5 GND 0.38fF
C557 a_6789_1050.n6 GND 0.59fF
C558 a_6789_1050.n7 GND 0.70fF
C559 a_6789_1050.n8 GND 0.08fF
C560 a_6789_1050.n9 GND 0.16fF
C561 a_6789_1050.n10 GND 0.05fF
C562 VDD.n1 GND 0.03fF
C563 VDD.n2 GND 0.14fF
C564 VDD.n3 GND 0.03fF
C565 VDD.n4 GND 0.02fF
C566 VDD.n5 GND 0.06fF
C567 VDD.n6 GND 0.02fF
C568 VDD.n7 GND 0.02fF
C569 VDD.n8 GND 0.02fF
C570 VDD.n9 GND 0.02fF
C571 VDD.n10 GND 0.02fF
C572 VDD.n11 GND 0.02fF
C573 VDD.n12 GND 0.02fF
C574 VDD.n13 GND 0.02fF
C575 VDD.n14 GND 0.04fF
C576 VDD.n15 GND 0.01fF
C577 VDD.n20 GND 0.48fF
C578 VDD.n21 GND 0.29fF
C579 VDD.n22 GND 0.02fF
C580 VDD.n23 GND 0.04fF
C581 VDD.n24 GND 0.25fF
C582 VDD.n25 GND 0.01fF
C583 VDD.n26 GND 0.02fF
C584 VDD.n27 GND 0.01fF
C585 VDD.n28 GND 0.17fF
C586 VDD.n29 GND 0.01fF
C587 VDD.n30 GND 0.02fF
C588 VDD.n31 GND 0.08fF
C589 VDD.n32 GND 0.01fF
C590 VDD.n33 GND 0.03fF
C591 VDD.n34 GND 0.03fF
C592 VDD.n35 GND 0.15fF
C593 VDD.n36 GND 0.01fF
C594 VDD.n37 GND 0.03fF
C595 VDD.n38 GND 0.03fF
C596 VDD.n39 GND 0.17fF
C597 VDD.n40 GND 0.01fF
C598 VDD.n41 GND 0.02fF
C599 VDD.n42 GND 0.02fF
C600 VDD.n43 GND 0.26fF
C601 VDD.n44 GND 0.01fF
C602 VDD.n45 GND 0.02fF
C603 VDD.n46 GND 0.02fF
C604 VDD.n47 GND 0.29fF
C605 VDD.n48 GND 0.01fF
C606 VDD.n49 GND 0.02fF
C607 VDD.n50 GND 0.04fF
C608 VDD.n51 GND 0.06fF
C609 VDD.n52 GND 0.02fF
C610 VDD.n53 GND 0.02fF
C611 VDD.n54 GND 0.02fF
C612 VDD.n55 GND 0.02fF
C613 VDD.n56 GND 0.02fF
C614 VDD.n57 GND 0.02fF
C615 VDD.n58 GND 0.02fF
C616 VDD.n59 GND 0.02fF
C617 VDD.n60 GND 0.02fF
C618 VDD.n61 GND 0.02fF
C619 VDD.n62 GND 0.02fF
C620 VDD.n63 GND 0.03fF
C621 VDD.n64 GND 0.02fF
C622 VDD.n65 GND 0.23fF
C623 VDD.n66 GND 0.02fF
C624 VDD.n67 GND 0.02fF
C625 VDD.n69 GND 0.02fF
C626 VDD.n73 GND 0.29fF
C627 VDD.n74 GND 0.29fF
C628 VDD.n75 GND 0.01fF
C629 VDD.n76 GND 0.02fF
C630 VDD.n77 GND 0.04fF
C631 VDD.n78 GND 0.26fF
C632 VDD.n79 GND 0.01fF
C633 VDD.n80 GND 0.02fF
C634 VDD.n81 GND 0.02fF
C635 VDD.n82 GND 0.17fF
C636 VDD.n83 GND 0.01fF
C637 VDD.n84 GND 0.02fF
C638 VDD.n85 GND 0.02fF
C639 VDD.n86 GND 0.15fF
C640 VDD.n87 GND 0.01fF
C641 VDD.n88 GND 0.03fF
C642 VDD.n89 GND 0.03fF
C643 VDD.n90 GND 0.01fF
C644 VDD.n91 GND 0.03fF
C645 VDD.n92 GND 0.03fF
C646 VDD.n93 GND 0.17fF
C647 VDD.n94 GND 0.01fF
C648 VDD.n95 GND 0.02fF
C649 VDD.n96 GND 0.02fF
C650 VDD.n97 GND 0.25fF
C651 VDD.n98 GND 0.01fF
C652 VDD.n99 GND 0.02fF
C653 VDD.n100 GND 0.02fF
C654 VDD.n101 GND 0.29fF
C655 VDD.n102 GND 0.01fF
C656 VDD.n103 GND 0.02fF
C657 VDD.n104 GND 0.04fF
C658 VDD.n105 GND 0.22fF
C659 VDD.n106 GND 0.02fF
C660 VDD.n107 GND 0.02fF
C661 VDD.n108 GND 0.02fF
C662 VDD.n109 GND 0.06fF
C663 VDD.n110 GND 0.02fF
C664 VDD.n111 GND 0.02fF
C665 VDD.n112 GND 0.02fF
C666 VDD.n113 GND 0.02fF
C667 VDD.n114 GND 0.02fF
C668 VDD.n115 GND 0.02fF
C669 VDD.n116 GND 0.02fF
C670 VDD.n117 GND 0.02fF
C671 VDD.n118 GND 0.02fF
C672 VDD.n119 GND 0.02fF
C673 VDD.n120 GND 0.03fF
C674 VDD.n121 GND 0.02fF
C675 VDD.n122 GND 0.02fF
C676 VDD.n126 GND 0.29fF
C677 VDD.n127 GND 0.29fF
C678 VDD.n128 GND 0.01fF
C679 VDD.n129 GND 0.02fF
C680 VDD.n130 GND 0.04fF
C681 VDD.n131 GND 0.07fF
C682 VDD.n132 GND 0.25fF
C683 VDD.n133 GND 0.01fF
C684 VDD.n134 GND 0.01fF
C685 VDD.n135 GND 0.02fF
C686 VDD.n136 GND 0.17fF
C687 VDD.n137 GND 0.01fF
C688 VDD.n138 GND 0.02fF
C689 VDD.n139 GND 0.02fF
C690 VDD.n140 GND 0.08fF
C691 VDD.n141 GND 0.05fF
C692 VDD.n142 GND 0.01fF
C693 VDD.n143 GND 0.02fF
C694 VDD.n144 GND 0.03fF
C695 VDD.n145 GND 0.15fF
C696 VDD.n146 GND 0.01fF
C697 VDD.n147 GND 0.02fF
C698 VDD.n148 GND 0.03fF
C699 VDD.n149 GND 0.17fF
C700 VDD.n150 GND 0.01fF
C701 VDD.n151 GND 0.02fF
C702 VDD.n152 GND 0.02fF
C703 VDD.n153 GND 0.07fF
C704 VDD.n154 GND 0.26fF
C705 VDD.n155 GND 0.01fF
C706 VDD.n156 GND 0.01fF
C707 VDD.n157 GND 0.02fF
C708 VDD.n158 GND 0.29fF
C709 VDD.n159 GND 0.01fF
C710 VDD.n160 GND 0.02fF
C711 VDD.n161 GND 0.04fF
C712 VDD.n162 GND 0.27fF
C713 VDD.n163 GND 0.02fF
C714 VDD.n164 GND 0.02fF
C715 VDD.n165 GND 0.02fF
C716 VDD.n166 GND 0.06fF
C717 VDD.n167 GND 0.02fF
C718 VDD.n168 GND 0.02fF
C719 VDD.n169 GND 0.02fF
C720 VDD.n170 GND 0.02fF
C721 VDD.n171 GND 0.02fF
C722 VDD.n172 GND 0.02fF
C723 VDD.n173 GND 0.02fF
C724 VDD.n174 GND 0.02fF
C725 VDD.n175 GND 0.02fF
C726 VDD.n176 GND 0.02fF
C727 VDD.n177 GND 0.03fF
C728 VDD.n178 GND 0.02fF
C729 VDD.n179 GND 0.02fF
C730 VDD.n183 GND 0.29fF
C731 VDD.n184 GND 0.29fF
C732 VDD.n185 GND 0.01fF
C733 VDD.n186 GND 0.02fF
C734 VDD.n187 GND 0.04fF
C735 VDD.n188 GND 0.29fF
C736 VDD.n189 GND 0.01fF
C737 VDD.n190 GND 0.02fF
C738 VDD.n191 GND 0.02fF
C739 VDD.n192 GND 0.23fF
C740 VDD.n193 GND 0.01fF
C741 VDD.n194 GND 0.07fF
C742 VDD.n195 GND 0.02fF
C743 VDD.n196 GND 0.17fF
C744 VDD.n197 GND 0.01fF
C745 VDD.n198 GND 0.02fF
C746 VDD.n199 GND 0.02fF
C747 VDD.n200 GND 0.17fF
C748 VDD.n201 GND 0.01fF
C749 VDD.n202 GND 0.08fF
C750 VDD.n203 GND 0.05fF
C751 VDD.n204 GND 0.02fF
C752 VDD.n205 GND 0.02fF
C753 VDD.n206 GND 0.15fF
C754 VDD.n207 GND 0.02fF
C755 VDD.n208 GND 0.02fF
C756 VDD.n209 GND 0.03fF
C757 VDD.n210 GND 0.16fF
C758 VDD.n211 GND 0.02fF
C759 VDD.n212 GND 0.02fF
C760 VDD.n213 GND 0.03fF
C761 VDD.n214 GND 0.08fF
C762 VDD.n215 GND 0.05fF
C763 VDD.n216 GND 0.16fF
C764 VDD.n217 GND 0.01fF
C765 VDD.n218 GND 0.02fF
C766 VDD.n219 GND 0.02fF
C767 VDD.n220 GND 0.17fF
C768 VDD.n221 GND 0.01fF
C769 VDD.n222 GND 0.02fF
C770 VDD.n223 GND 0.02fF
C771 VDD.n224 GND 0.07fF
C772 VDD.n225 GND 0.23fF
C773 VDD.n226 GND 0.01fF
C774 VDD.n227 GND 0.01fF
C775 VDD.n228 GND 0.02fF
C776 VDD.n229 GND 0.29fF
C777 VDD.n230 GND 0.01fF
C778 VDD.n231 GND 0.02fF
C779 VDD.n232 GND 0.02fF
C780 VDD.n233 GND 0.29fF
C781 VDD.n234 GND 0.01fF
C782 VDD.n235 GND 0.02fF
C783 VDD.n236 GND 0.04fF
C784 VDD.n237 GND 0.27fF
C785 VDD.n238 GND 0.02fF
C786 VDD.n239 GND 0.02fF
C787 VDD.n240 GND 0.02fF
C788 VDD.n241 GND 0.06fF
C789 VDD.n242 GND 0.02fF
C790 VDD.n243 GND 0.02fF
C791 VDD.n244 GND 0.02fF
C792 VDD.n245 GND 0.02fF
C793 VDD.n246 GND 0.02fF
C794 VDD.n247 GND 0.02fF
C795 VDD.n248 GND 0.02fF
C796 VDD.n249 GND 0.02fF
C797 VDD.n250 GND 0.02fF
C798 VDD.n251 GND 0.02fF
C799 VDD.n252 GND 0.03fF
C800 VDD.n253 GND 0.02fF
C801 VDD.n254 GND 0.02fF
C802 VDD.n258 GND 0.29fF
C803 VDD.n259 GND 0.29fF
C804 VDD.n260 GND 0.01fF
C805 VDD.n261 GND 0.02fF
C806 VDD.n262 GND 0.04fF
C807 VDD.n263 GND 0.06fF
C808 VDD.n264 GND 0.25fF
C809 VDD.n265 GND 0.01fF
C810 VDD.n266 GND 0.01fF
C811 VDD.n267 GND 0.02fF
C812 VDD.n268 GND 0.17fF
C813 VDD.n269 GND 0.01fF
C814 VDD.n270 GND 0.02fF
C815 VDD.n271 GND 0.02fF
C816 VDD.n272 GND 0.08fF
C817 VDD.n273 GND 0.05fF
C818 VDD.n274 GND 0.01fF
C819 VDD.n275 GND 0.02fF
C820 VDD.n276 GND 0.03fF
C821 VDD.n277 GND 0.15fF
C822 VDD.n278 GND 0.01fF
C823 VDD.n279 GND 0.02fF
C824 VDD.n280 GND 0.03fF
C825 VDD.n281 GND 0.17fF
C826 VDD.n282 GND 0.01fF
C827 VDD.n283 GND 0.02fF
C828 VDD.n284 GND 0.02fF
C829 VDD.n285 GND 0.07fF
C830 VDD.n286 GND 0.26fF
C831 VDD.n287 GND 0.01fF
C832 VDD.n288 GND 0.01fF
C833 VDD.n289 GND 0.02fF
C834 VDD.n290 GND 0.29fF
C835 VDD.n291 GND 0.01fF
C836 VDD.n292 GND 0.02fF
C837 VDD.n293 GND 0.04fF
C838 VDD.n294 GND 0.22fF
C839 VDD.n295 GND 0.02fF
C840 VDD.n296 GND 0.02fF
C841 VDD.n297 GND 0.02fF
C842 VDD.n298 GND 0.06fF
C843 VDD.n299 GND 0.02fF
C844 VDD.n300 GND 0.02fF
C845 VDD.n301 GND 0.02fF
C846 VDD.n302 GND 0.02fF
C847 VDD.n303 GND 0.02fF
C848 VDD.n304 GND 0.02fF
C849 VDD.n305 GND 0.02fF
C850 VDD.n306 GND 0.02fF
C851 VDD.n307 GND 0.02fF
C852 VDD.n308 GND 0.02fF
C853 VDD.n309 GND 0.03fF
C854 VDD.n310 GND 0.02fF
C855 VDD.n311 GND 0.02fF
C856 VDD.n315 GND 0.29fF
C857 VDD.n316 GND 0.29fF
C858 VDD.n317 GND 0.01fF
C859 VDD.n318 GND 0.02fF
C860 VDD.n319 GND 0.04fF
C861 VDD.n320 GND 0.06fF
C862 VDD.n321 GND 0.25fF
C863 VDD.n322 GND 0.01fF
C864 VDD.n323 GND 0.01fF
C865 VDD.n324 GND 0.02fF
C866 VDD.n325 GND 0.17fF
C867 VDD.n326 GND 0.01fF
C868 VDD.n327 GND 0.02fF
C869 VDD.n328 GND 0.02fF
C870 VDD.n329 GND 0.08fF
C871 VDD.n330 GND 0.05fF
C872 VDD.n331 GND 0.01fF
C873 VDD.n332 GND 0.02fF
C874 VDD.n333 GND 0.03fF
C875 VDD.n334 GND 0.15fF
C876 VDD.n335 GND 0.01fF
C877 VDD.n336 GND 0.02fF
C878 VDD.n337 GND 0.03fF
C879 VDD.n338 GND 0.17fF
C880 VDD.n339 GND 0.01fF
C881 VDD.n340 GND 0.02fF
C882 VDD.n341 GND 0.02fF
C883 VDD.n342 GND 0.07fF
C884 VDD.n343 GND 0.26fF
C885 VDD.n344 GND 0.01fF
C886 VDD.n345 GND 0.01fF
C887 VDD.n346 GND 0.02fF
C888 VDD.n347 GND 0.29fF
C889 VDD.n348 GND 0.01fF
C890 VDD.n349 GND 0.02fF
C891 VDD.n350 GND 0.04fF
C892 VDD.n351 GND 0.27fF
C893 VDD.n352 GND 0.02fF
C894 VDD.n353 GND 0.02fF
C895 VDD.n354 GND 0.02fF
C896 VDD.n355 GND 0.06fF
C897 VDD.n356 GND 0.02fF
C898 VDD.n357 GND 0.02fF
C899 VDD.n358 GND 0.02fF
C900 VDD.n359 GND 0.02fF
C901 VDD.n360 GND 0.02fF
C902 VDD.n361 GND 0.02fF
C903 VDD.n362 GND 0.02fF
C904 VDD.n363 GND 0.02fF
C905 VDD.n364 GND 0.02fF
C906 VDD.n365 GND 0.02fF
C907 VDD.n366 GND 0.03fF
C908 VDD.n367 GND 0.02fF
C909 VDD.n368 GND 0.02fF
C910 VDD.n372 GND 0.29fF
C911 VDD.n373 GND 0.29fF
C912 VDD.n374 GND 0.01fF
C913 VDD.n375 GND 0.02fF
C914 VDD.n376 GND 0.04fF
C915 VDD.n377 GND 0.29fF
C916 VDD.n378 GND 0.01fF
C917 VDD.n379 GND 0.02fF
C918 VDD.n380 GND 0.02fF
C919 VDD.n381 GND 0.23fF
C920 VDD.n382 GND 0.01fF
C921 VDD.n383 GND 0.07fF
C922 VDD.n384 GND 0.02fF
C923 VDD.n385 GND 0.17fF
C924 VDD.n386 GND 0.01fF
C925 VDD.n387 GND 0.02fF
C926 VDD.n388 GND 0.02fF
C927 VDD.n389 GND 0.17fF
C928 VDD.n390 GND 0.01fF
C929 VDD.n391 GND 0.08fF
C930 VDD.n392 GND 0.05fF
C931 VDD.n393 GND 0.02fF
C932 VDD.n394 GND 0.02fF
C933 VDD.n395 GND 0.15fF
C934 VDD.n396 GND 0.02fF
C935 VDD.n397 GND 0.02fF
C936 VDD.n398 GND 0.03fF
C937 VDD.n399 GND 0.16fF
C938 VDD.n400 GND 0.02fF
C939 VDD.n401 GND 0.02fF
C940 VDD.n402 GND 0.03fF
C941 VDD.n403 GND 0.08fF
C942 VDD.n404 GND 0.05fF
C943 VDD.n405 GND 0.16fF
C944 VDD.n406 GND 0.01fF
C945 VDD.n407 GND 0.02fF
C946 VDD.n408 GND 0.02fF
C947 VDD.n409 GND 0.17fF
C948 VDD.n410 GND 0.01fF
C949 VDD.n411 GND 0.02fF
C950 VDD.n412 GND 0.02fF
C951 VDD.n413 GND 0.07fF
C952 VDD.n414 GND 0.23fF
C953 VDD.n415 GND 0.01fF
C954 VDD.n416 GND 0.01fF
C955 VDD.n417 GND 0.02fF
C956 VDD.n418 GND 0.29fF
C957 VDD.n419 GND 0.01fF
C958 VDD.n420 GND 0.02fF
C959 VDD.n421 GND 0.02fF
C960 VDD.n422 GND 0.29fF
C961 VDD.n423 GND 0.01fF
C962 VDD.n424 GND 0.02fF
C963 VDD.n425 GND 0.04fF
C964 VDD.n426 GND 0.32fF
C965 VDD.n427 GND 0.02fF
C966 VDD.n428 GND 0.02fF
C967 VDD.n429 GND 0.02fF
C968 VDD.n430 GND 0.06fF
C969 VDD.n431 GND 0.02fF
C970 VDD.n432 GND 0.02fF
C971 VDD.n433 GND 0.02fF
C972 VDD.n434 GND 0.02fF
C973 VDD.n435 GND 0.02fF
C974 VDD.n436 GND 0.02fF
C975 VDD.n437 GND 0.02fF
C976 VDD.n438 GND 0.02fF
C977 VDD.n439 GND 0.02fF
C978 VDD.n440 GND 0.02fF
C979 VDD.n441 GND 0.03fF
C980 VDD.n442 GND 0.02fF
C981 VDD.n443 GND 0.02fF
C982 VDD.n447 GND 0.29fF
C983 VDD.n448 GND 0.29fF
C984 VDD.n449 GND 0.01fF
C985 VDD.n450 GND 0.02fF
C986 VDD.n451 GND 0.04fF
C987 VDD.n452 GND 0.29fF
C988 VDD.n453 GND 0.01fF
C989 VDD.n454 GND 0.02fF
C990 VDD.n455 GND 0.02fF
C991 VDD.n456 GND 0.23fF
C992 VDD.n457 GND 0.01fF
C993 VDD.n458 GND 0.07fF
C994 VDD.n459 GND 0.02fF
C995 VDD.n460 GND 0.17fF
C996 VDD.n461 GND 0.01fF
C997 VDD.n462 GND 0.02fF
C998 VDD.n463 GND 0.02fF
C999 VDD.n464 GND 0.17fF
C1000 VDD.n465 GND 0.01fF
C1001 VDD.n466 GND 0.08fF
C1002 VDD.n467 GND 0.05fF
C1003 VDD.n468 GND 0.02fF
C1004 VDD.n469 GND 0.02fF
C1005 VDD.n470 GND 0.15fF
C1006 VDD.n471 GND 0.02fF
C1007 VDD.n472 GND 0.02fF
C1008 VDD.n473 GND 0.03fF
C1009 VDD.n474 GND 0.16fF
C1010 VDD.n475 GND 0.02fF
C1011 VDD.n476 GND 0.02fF
C1012 VDD.n477 GND 0.03fF
C1013 VDD.n478 GND 0.08fF
C1014 VDD.n479 GND 0.05fF
C1015 VDD.n480 GND 0.16fF
C1016 VDD.n481 GND 0.01fF
C1017 VDD.n482 GND 0.02fF
C1018 VDD.n483 GND 0.02fF
C1019 VDD.n484 GND 0.17fF
C1020 VDD.n485 GND 0.01fF
C1021 VDD.n486 GND 0.02fF
C1022 VDD.n487 GND 0.02fF
C1023 VDD.n488 GND 0.07fF
C1024 VDD.n489 GND 0.23fF
C1025 VDD.n490 GND 0.01fF
C1026 VDD.n491 GND 0.01fF
C1027 VDD.n492 GND 0.02fF
C1028 VDD.n493 GND 0.29fF
C1029 VDD.n494 GND 0.01fF
C1030 VDD.n495 GND 0.02fF
C1031 VDD.n496 GND 0.02fF
C1032 VDD.n497 GND 0.29fF
C1033 VDD.n498 GND 0.01fF
C1034 VDD.n499 GND 0.02fF
C1035 VDD.n500 GND 0.04fF
C1036 VDD.n501 GND 0.27fF
C1037 VDD.n502 GND 0.02fF
C1038 VDD.n503 GND 0.02fF
C1039 VDD.n504 GND 0.02fF
C1040 VDD.n505 GND 0.06fF
C1041 VDD.n506 GND 0.02fF
C1042 VDD.n507 GND 0.02fF
C1043 VDD.n508 GND 0.02fF
C1044 VDD.n509 GND 0.02fF
C1045 VDD.n510 GND 0.02fF
C1046 VDD.n511 GND 0.02fF
C1047 VDD.n512 GND 0.02fF
C1048 VDD.n513 GND 0.02fF
C1049 VDD.n514 GND 0.02fF
C1050 VDD.n515 GND 0.02fF
C1051 VDD.n516 GND 0.03fF
C1052 VDD.n517 GND 0.02fF
C1053 VDD.n518 GND 0.02fF
C1054 VDD.n522 GND 0.29fF
C1055 VDD.n523 GND 0.29fF
C1056 VDD.n524 GND 0.01fF
C1057 VDD.n525 GND 0.02fF
C1058 VDD.n526 GND 0.04fF
C1059 VDD.n527 GND 0.06fF
C1060 VDD.n528 GND 0.25fF
C1061 VDD.n529 GND 0.01fF
C1062 VDD.n530 GND 0.01fF
C1063 VDD.n531 GND 0.02fF
C1064 VDD.n532 GND 0.17fF
C1065 VDD.n533 GND 0.01fF
C1066 VDD.n534 GND 0.02fF
C1067 VDD.n535 GND 0.02fF
C1068 VDD.n536 GND 0.08fF
C1069 VDD.n537 GND 0.05fF
C1070 VDD.n538 GND 0.01fF
C1071 VDD.n539 GND 0.02fF
C1072 VDD.n540 GND 0.03fF
C1073 VDD.n541 GND 0.15fF
C1074 VDD.n542 GND 0.01fF
C1075 VDD.n543 GND 0.02fF
C1076 VDD.n544 GND 0.03fF
C1077 VDD.n545 GND 0.17fF
C1078 VDD.n546 GND 0.01fF
C1079 VDD.n547 GND 0.02fF
C1080 VDD.n548 GND 0.02fF
C1081 VDD.n549 GND 0.07fF
C1082 VDD.n550 GND 0.26fF
C1083 VDD.n551 GND 0.01fF
C1084 VDD.n552 GND 0.01fF
C1085 VDD.n553 GND 0.02fF
C1086 VDD.n554 GND 0.29fF
C1087 VDD.n555 GND 0.01fF
C1088 VDD.n556 GND 0.02fF
C1089 VDD.n557 GND 0.04fF
C1090 VDD.n558 GND 0.27fF
C1091 VDD.n559 GND 0.02fF
C1092 VDD.n560 GND 0.02fF
C1093 VDD.n561 GND 0.02fF
C1094 VDD.n562 GND 0.06fF
C1095 VDD.n563 GND 0.02fF
C1096 VDD.n564 GND 0.02fF
C1097 VDD.n565 GND 0.02fF
C1098 VDD.n566 GND 0.02fF
C1099 VDD.n567 GND 0.02fF
C1100 VDD.n568 GND 0.02fF
C1101 VDD.n569 GND 0.02fF
C1102 VDD.n570 GND 0.02fF
C1103 VDD.n571 GND 0.02fF
C1104 VDD.n572 GND 0.02fF
C1105 VDD.n573 GND 0.03fF
C1106 VDD.n574 GND 0.02fF
C1107 VDD.n575 GND 0.02fF
C1108 VDD.n579 GND 0.29fF
C1109 VDD.n580 GND 0.29fF
C1110 VDD.n581 GND 0.01fF
C1111 VDD.n582 GND 0.02fF
C1112 VDD.n583 GND 0.04fF
C1113 VDD.n584 GND 0.29fF
C1114 VDD.n585 GND 0.01fF
C1115 VDD.n586 GND 0.02fF
C1116 VDD.n587 GND 0.02fF
C1117 VDD.n588 GND 0.23fF
C1118 VDD.n589 GND 0.01fF
C1119 VDD.n590 GND 0.07fF
C1120 VDD.n591 GND 0.02fF
C1121 VDD.n592 GND 0.17fF
C1122 VDD.n593 GND 0.01fF
C1123 VDD.n594 GND 0.02fF
C1124 VDD.n595 GND 0.02fF
C1125 VDD.n596 GND 0.17fF
C1126 VDD.n597 GND 0.01fF
C1127 VDD.n598 GND 0.08fF
C1128 VDD.n599 GND 0.05fF
C1129 VDD.n600 GND 0.02fF
C1130 VDD.n601 GND 0.02fF
C1131 VDD.n602 GND 0.15fF
C1132 VDD.n603 GND 0.02fF
C1133 VDD.n604 GND 0.02fF
C1134 VDD.n605 GND 0.03fF
C1135 VDD.n606 GND 0.16fF
C1136 VDD.n607 GND 0.02fF
C1137 VDD.n608 GND 0.02fF
C1138 VDD.n609 GND 0.03fF
C1139 VDD.n610 GND 0.08fF
C1140 VDD.n611 GND 0.05fF
C1141 VDD.n612 GND 0.16fF
C1142 VDD.n613 GND 0.01fF
C1143 VDD.n614 GND 0.02fF
C1144 VDD.n615 GND 0.02fF
C1145 VDD.n616 GND 0.17fF
C1146 VDD.n617 GND 0.01fF
C1147 VDD.n618 GND 0.02fF
C1148 VDD.n619 GND 0.02fF
C1149 VDD.n620 GND 0.07fF
C1150 VDD.n621 GND 0.23fF
C1151 VDD.n622 GND 0.01fF
C1152 VDD.n623 GND 0.01fF
C1153 VDD.n624 GND 0.02fF
C1154 VDD.n625 GND 0.29fF
C1155 VDD.n626 GND 0.01fF
C1156 VDD.n627 GND 0.02fF
C1157 VDD.n628 GND 0.02fF
C1158 VDD.n629 GND 0.29fF
C1159 VDD.n630 GND 0.01fF
C1160 VDD.n631 GND 0.02fF
C1161 VDD.n632 GND 0.04fF
C1162 VDD.n633 GND 0.27fF
C1163 VDD.n634 GND 0.02fF
C1164 VDD.n635 GND 0.02fF
C1165 VDD.n636 GND 0.02fF
C1166 VDD.n637 GND 0.06fF
C1167 VDD.n638 GND 0.02fF
C1168 VDD.n639 GND 0.02fF
C1169 VDD.n640 GND 0.02fF
C1170 VDD.n641 GND 0.02fF
C1171 VDD.n642 GND 0.02fF
C1172 VDD.n643 GND 0.02fF
C1173 VDD.n644 GND 0.02fF
C1174 VDD.n645 GND 0.02fF
C1175 VDD.n646 GND 0.02fF
C1176 VDD.n647 GND 0.02fF
C1177 VDD.n648 GND 0.03fF
C1178 VDD.n649 GND 0.02fF
C1179 VDD.n650 GND 0.02fF
C1180 VDD.n654 GND 0.29fF
C1181 VDD.n655 GND 0.29fF
C1182 VDD.n656 GND 0.01fF
C1183 VDD.n657 GND 0.02fF
C1184 VDD.n658 GND 0.04fF
C1185 VDD.n659 GND 0.06fF
C1186 VDD.n660 GND 0.25fF
C1187 VDD.n661 GND 0.01fF
C1188 VDD.n662 GND 0.01fF
C1189 VDD.n663 GND 0.02fF
C1190 VDD.n664 GND 0.17fF
C1191 VDD.n665 GND 0.01fF
C1192 VDD.n666 GND 0.02fF
C1193 VDD.n667 GND 0.02fF
C1194 VDD.n668 GND 0.08fF
C1195 VDD.n669 GND 0.05fF
C1196 VDD.n670 GND 0.01fF
C1197 VDD.n671 GND 0.02fF
C1198 VDD.n672 GND 0.03fF
C1199 VDD.n673 GND 0.15fF
C1200 VDD.n674 GND 0.01fF
C1201 VDD.n675 GND 0.02fF
C1202 VDD.n676 GND 0.03fF
C1203 VDD.n677 GND 0.17fF
C1204 VDD.n678 GND 0.01fF
C1205 VDD.n679 GND 0.02fF
C1206 VDD.n680 GND 0.02fF
C1207 VDD.n681 GND 0.14fF
C1208 VDD.n682 GND 0.02fF
C1209 VDD.n683 GND 0.02fF
C1210 VDD.n684 GND 0.06fF
C1211 VDD.n685 GND 0.02fF
C1212 VDD.n686 GND 0.02fF
C1213 VDD.n687 GND 0.02fF
C1214 VDD.n688 GND 0.02fF
C1215 VDD.n689 GND 0.02fF
C1216 VDD.n690 GND 0.02fF
C1217 VDD.n691 GND 0.02fF
C1218 VDD.n692 GND 0.02fF
C1219 VDD.n693 GND 0.03fF
C1220 VDD.n694 GND 0.04fF
C1221 VDD.n695 GND 0.02fF
C1222 VDD.n699 GND 0.48fF
C1223 VDD.n700 GND 0.29fF
C1224 VDD.n701 GND 0.02fF
C1225 VDD.n702 GND 0.03fF
C1226 VDD.n703 GND 0.03fF
C1227 VDD.n704 GND 0.07fF
C1228 VDD.n705 GND 0.26fF
C1229 VDD.n706 GND 0.01fF
C1230 VDD.n707 GND 0.01fF
C1231 VDD.n708 GND 0.02fF
C1232 VDD.n709 GND 0.17fF
C1233 VDD.n710 GND 0.01fF
C1234 VDD.n711 GND 0.02fF
C1235 VDD.n712 GND 0.02fF
C1236 VDD.n713 GND 0.15fF
C1237 VDD.n714 GND 0.01fF
C1238 VDD.n715 GND 0.02fF
C1239 VDD.n716 GND 0.03fF
C1240 VDD.n717 GND 0.08fF
C1241 VDD.n718 GND 0.05fF
C1242 VDD.n719 GND 0.01fF
C1243 VDD.n720 GND 0.02fF
C1244 VDD.n721 GND 0.03fF
C1245 VDD.n722 GND 0.17fF
C1246 VDD.n723 GND 0.01fF
C1247 VDD.n724 GND 0.02fF
C1248 VDD.n725 GND 0.02fF
C1249 VDD.n726 GND 0.06fF
C1250 VDD.n727 GND 0.25fF
C1251 VDD.n728 GND 0.01fF
C1252 VDD.n729 GND 0.01fF
C1253 VDD.n730 GND 0.02fF
C1254 VDD.n731 GND 0.29fF
C1255 VDD.n732 GND 0.01fF
C1256 VDD.n733 GND 0.02fF
C1257 VDD.n734 GND 0.04fF
C1258 VDD.n735 GND 0.06fF
C1259 VDD.n736 GND 0.02fF
C1260 VDD.n737 GND 0.02fF
C1261 VDD.n738 GND 0.02fF
C1262 VDD.n739 GND 0.02fF
C1263 VDD.n740 GND 0.02fF
C1264 VDD.n741 GND 0.02fF
C1265 VDD.n742 GND 0.02fF
C1266 VDD.n743 GND 0.02fF
C1267 VDD.n744 GND 0.02fF
C1268 VDD.n745 GND 0.02fF
C1269 VDD.n746 GND 0.02fF
C1270 VDD.n747 GND 0.03fF
C1271 VDD.n748 GND 0.02fF
C1272 VDD.n751 GND 0.02fF
C1273 VDD.n753 GND 0.02fF
C1274 VDD.n754 GND 0.28fF
C1275 VDD.n755 GND 0.02fF
C1276 VDD.n757 GND 0.29fF
C1277 VDD.n758 GND 0.29fF
C1278 VDD.n759 GND 0.01fF
C1279 VDD.n760 GND 0.02fF
C1280 VDD.n761 GND 0.04fF
C1281 VDD.n762 GND 0.29fF
C1282 VDD.n763 GND 0.01fF
C1283 VDD.n764 GND 0.02fF
C1284 VDD.n765 GND 0.02fF
C1285 VDD.n766 GND 0.07fF
C1286 VDD.n767 GND 0.23fF
C1287 VDD.n768 GND 0.01fF
C1288 VDD.n769 GND 0.01fF
C1289 VDD.n770 GND 0.02fF
C1290 VDD.n771 GND 0.17fF
C1291 VDD.n772 GND 0.01fF
C1292 VDD.n773 GND 0.02fF
C1293 VDD.n774 GND 0.02fF
C1294 VDD.n775 GND 0.08fF
C1295 VDD.n776 GND 0.05fF
C1296 VDD.n777 GND 0.16fF
C1297 VDD.n778 GND 0.01fF
C1298 VDD.n779 GND 0.02fF
C1299 VDD.n780 GND 0.02fF
C1300 VDD.n781 GND 0.16fF
C1301 VDD.n782 GND 0.02fF
C1302 VDD.n783 GND 0.02fF
C1303 VDD.n784 GND 0.03fF
C1304 VDD.n785 GND 0.15fF
C1305 VDD.n786 GND 0.02fF
C1306 VDD.n787 GND 0.02fF
C1307 VDD.n788 GND 0.03fF
C1308 VDD.n789 GND 0.17fF
C1309 VDD.n790 GND 0.01fF
C1310 VDD.n791 GND 0.08fF
C1311 VDD.n792 GND 0.05fF
C1312 VDD.n793 GND 0.02fF
C1313 VDD.n794 GND 0.02fF
C1314 VDD.n795 GND 0.17fF
C1315 VDD.n796 GND 0.01fF
C1316 VDD.n797 GND 0.02fF
C1317 VDD.n798 GND 0.02fF
C1318 VDD.n799 GND 0.23fF
C1319 VDD.n800 GND 0.01fF
C1320 VDD.n801 GND 0.07fF
C1321 VDD.n802 GND 0.02fF
C1322 VDD.n803 GND 0.29fF
C1323 VDD.n804 GND 0.01fF
C1324 VDD.n805 GND 0.02fF
C1325 VDD.n806 GND 0.02fF
C1326 VDD.n807 GND 0.29fF
C1327 VDD.n808 GND 0.01fF
C1328 VDD.n809 GND 0.02fF
C1329 VDD.n810 GND 0.04fF
C1330 VDD.n811 GND 0.32fF
C1331 VDD.n812 GND 0.02fF
C1332 VDD.n813 GND 0.02fF
C1333 VDD.n814 GND 0.02fF
C1334 VDD.n815 GND 0.06fF
C1335 VDD.n816 GND 0.02fF
C1336 VDD.n817 GND 0.02fF
C1337 VDD.n818 GND 0.02fF
C1338 VDD.n819 GND 0.02fF
C1339 VDD.n820 GND 0.02fF
C1340 VDD.n821 GND 0.02fF
C1341 VDD.n822 GND 0.02fF
C1342 VDD.n823 GND 0.02fF
C1343 VDD.n824 GND 0.02fF
C1344 VDD.n825 GND 0.02fF
C1345 VDD.n826 GND 0.03fF
C1346 VDD.n827 GND 0.02fF
C1347 VDD.n828 GND 0.02fF
C1348 VDD.n832 GND 0.29fF
C1349 VDD.n833 GND 0.29fF
C1350 VDD.n834 GND 0.01fF
C1351 VDD.n835 GND 0.02fF
C1352 VDD.n836 GND 0.04fF
C1353 VDD.n837 GND 0.29fF
C1354 VDD.n838 GND 0.01fF
C1355 VDD.n839 GND 0.02fF
C1356 VDD.n840 GND 0.02fF
C1357 VDD.n841 GND 0.07fF
C1358 VDD.n842 GND 0.23fF
C1359 VDD.n843 GND 0.01fF
C1360 VDD.n844 GND 0.01fF
C1361 VDD.n845 GND 0.02fF
C1362 VDD.n846 GND 0.17fF
C1363 VDD.n847 GND 0.01fF
C1364 VDD.n848 GND 0.02fF
C1365 VDD.n849 GND 0.02fF
C1366 VDD.n850 GND 0.08fF
C1367 VDD.n851 GND 0.05fF
C1368 VDD.n852 GND 0.16fF
C1369 VDD.n853 GND 0.01fF
C1370 VDD.n854 GND 0.02fF
C1371 VDD.n855 GND 0.02fF
C1372 VDD.n856 GND 0.16fF
C1373 VDD.n857 GND 0.02fF
C1374 VDD.n858 GND 0.02fF
C1375 VDD.n859 GND 0.03fF
C1376 VDD.n860 GND 0.15fF
C1377 VDD.n861 GND 0.02fF
C1378 VDD.n862 GND 0.02fF
C1379 VDD.n863 GND 0.03fF
C1380 VDD.n864 GND 0.17fF
C1381 VDD.n865 GND 0.01fF
C1382 VDD.n866 GND 0.08fF
C1383 VDD.n867 GND 0.05fF
C1384 VDD.n868 GND 0.02fF
C1385 VDD.n869 GND 0.02fF
C1386 VDD.n870 GND 0.17fF
C1387 VDD.n871 GND 0.01fF
C1388 VDD.n872 GND 0.02fF
C1389 VDD.n873 GND 0.02fF
C1390 VDD.n874 GND 0.23fF
C1391 VDD.n875 GND 0.01fF
C1392 VDD.n876 GND 0.07fF
C1393 VDD.n877 GND 0.02fF
C1394 VDD.n878 GND 0.29fF
C1395 VDD.n879 GND 0.01fF
C1396 VDD.n880 GND 0.02fF
C1397 VDD.n881 GND 0.02fF
C1398 VDD.n882 GND 0.29fF
C1399 VDD.n883 GND 0.01fF
C1400 VDD.n884 GND 0.02fF
C1401 VDD.n885 GND 0.04fF
C1402 VDD.n886 GND 0.27fF
C1403 VDD.n887 GND 0.02fF
C1404 VDD.n888 GND 0.02fF
C1405 VDD.n889 GND 0.02fF
C1406 VDD.n890 GND 0.06fF
C1407 VDD.n891 GND 0.02fF
C1408 VDD.n892 GND 0.02fF
C1409 VDD.n893 GND 0.02fF
C1410 VDD.n894 GND 0.02fF
C1411 VDD.n895 GND 0.02fF
C1412 VDD.n896 GND 0.02fF
C1413 VDD.n897 GND 0.02fF
C1414 VDD.n898 GND 0.02fF
C1415 VDD.n899 GND 0.02fF
C1416 VDD.n900 GND 0.02fF
C1417 VDD.n901 GND 0.03fF
C1418 VDD.n902 GND 0.02fF
C1419 VDD.n903 GND 0.02fF
C1420 VDD.n907 GND 0.29fF
C1421 VDD.n908 GND 0.29fF
C1422 VDD.n909 GND 0.01fF
C1423 VDD.n910 GND 0.02fF
C1424 VDD.n911 GND 0.04fF
C1425 VDD.n912 GND 0.07fF
C1426 VDD.n913 GND 0.26fF
C1427 VDD.n914 GND 0.01fF
C1428 VDD.n915 GND 0.01fF
C1429 VDD.n916 GND 0.02fF
C1430 VDD.n917 GND 0.17fF
C1431 VDD.n918 GND 0.01fF
C1432 VDD.n919 GND 0.02fF
C1433 VDD.n920 GND 0.02fF
C1434 VDD.n921 GND 0.15fF
C1435 VDD.n922 GND 0.01fF
C1436 VDD.n923 GND 0.02fF
C1437 VDD.n924 GND 0.03fF
C1438 VDD.n925 GND 0.08fF
C1439 VDD.n926 GND 0.05fF
C1440 VDD.n927 GND 0.01fF
C1441 VDD.n928 GND 0.02fF
C1442 VDD.n929 GND 0.03fF
C1443 VDD.n930 GND 0.17fF
C1444 VDD.n931 GND 0.01fF
C1445 VDD.n932 GND 0.02fF
C1446 VDD.n933 GND 0.02fF
C1447 VDD.n934 GND 0.06fF
C1448 VDD.n935 GND 0.25fF
C1449 VDD.n936 GND 0.01fF
C1450 VDD.n937 GND 0.01fF
C1451 VDD.n938 GND 0.02fF
C1452 VDD.n939 GND 0.29fF
C1453 VDD.n940 GND 0.01fF
C1454 VDD.n941 GND 0.02fF
C1455 VDD.n942 GND 0.04fF
C1456 VDD.n943 GND 0.22fF
C1457 VDD.n944 GND 0.02fF
C1458 VDD.n945 GND 0.02fF
C1459 VDD.n946 GND 0.02fF
C1460 VDD.n947 GND 0.06fF
C1461 VDD.n948 GND 0.02fF
C1462 VDD.n949 GND 0.02fF
C1463 VDD.n950 GND 0.02fF
C1464 VDD.n951 GND 0.02fF
C1465 VDD.n952 GND 0.02fF
C1466 VDD.n953 GND 0.02fF
C1467 VDD.n954 GND 0.02fF
C1468 VDD.n955 GND 0.02fF
C1469 VDD.n956 GND 0.02fF
C1470 VDD.n957 GND 0.02fF
C1471 VDD.n958 GND 0.03fF
C1472 VDD.n959 GND 0.02fF
C1473 VDD.n960 GND 0.02fF
C1474 VDD.n964 GND 0.29fF
C1475 VDD.n965 GND 0.29fF
C1476 VDD.n966 GND 0.01fF
C1477 VDD.n967 GND 0.02fF
C1478 VDD.n968 GND 0.04fF
C1479 VDD.n969 GND 0.07fF
C1480 VDD.n970 GND 0.26fF
C1481 VDD.n971 GND 0.01fF
C1482 VDD.n972 GND 0.01fF
C1483 VDD.n973 GND 0.02fF
C1484 VDD.n974 GND 0.17fF
C1485 VDD.n975 GND 0.01fF
C1486 VDD.n976 GND 0.02fF
C1487 VDD.n977 GND 0.02fF
C1488 VDD.n978 GND 0.15fF
C1489 VDD.n979 GND 0.01fF
C1490 VDD.n980 GND 0.02fF
C1491 VDD.n981 GND 0.03fF
C1492 VDD.n982 GND 0.08fF
C1493 VDD.n983 GND 0.05fF
C1494 VDD.n984 GND 0.01fF
C1495 VDD.n985 GND 0.02fF
C1496 VDD.n986 GND 0.03fF
C1497 VDD.n987 GND 0.17fF
C1498 VDD.n988 GND 0.01fF
C1499 VDD.n989 GND 0.02fF
C1500 VDD.n990 GND 0.02fF
C1501 VDD.n991 GND 0.06fF
C1502 VDD.n992 GND 0.25fF
C1503 VDD.n993 GND 0.01fF
C1504 VDD.n994 GND 0.01fF
C1505 VDD.n995 GND 0.02fF
C1506 VDD.n996 GND 0.29fF
C1507 VDD.n997 GND 0.01fF
C1508 VDD.n998 GND 0.02fF
C1509 VDD.n999 GND 0.04fF
C1510 VDD.n1000 GND 0.27fF
C1511 VDD.n1001 GND 0.02fF
C1512 VDD.n1002 GND 0.02fF
C1513 VDD.n1003 GND 0.02fF
C1514 VDD.n1004 GND 0.06fF
C1515 VDD.n1005 GND 0.02fF
C1516 VDD.n1006 GND 0.02fF
C1517 VDD.n1007 GND 0.02fF
C1518 VDD.n1008 GND 0.02fF
C1519 VDD.n1009 GND 0.02fF
C1520 VDD.n1010 GND 0.02fF
C1521 VDD.n1011 GND 0.02fF
C1522 VDD.n1012 GND 0.02fF
C1523 VDD.n1013 GND 0.02fF
C1524 VDD.n1014 GND 0.02fF
C1525 VDD.n1015 GND 0.03fF
C1526 VDD.n1016 GND 0.02fF
C1527 VDD.n1017 GND 0.02fF
C1528 VDD.n1021 GND 0.29fF
C1529 VDD.n1022 GND 0.29fF
C1530 VDD.n1023 GND 0.01fF
C1531 VDD.n1024 GND 0.02fF
C1532 VDD.n1025 GND 0.04fF
C1533 VDD.n1026 GND 0.29fF
C1534 VDD.n1027 GND 0.01fF
C1535 VDD.n1028 GND 0.02fF
C1536 VDD.n1029 GND 0.02fF
C1537 VDD.n1030 GND 0.07fF
C1538 VDD.n1031 GND 0.23fF
C1539 VDD.n1032 GND 0.01fF
C1540 VDD.n1033 GND 0.01fF
C1541 VDD.n1034 GND 0.02fF
C1542 VDD.n1035 GND 0.17fF
C1543 VDD.n1036 GND 0.01fF
C1544 VDD.n1037 GND 0.02fF
C1545 VDD.n1038 GND 0.02fF
C1546 VDD.n1039 GND 0.08fF
C1547 VDD.n1040 GND 0.05fF
C1548 VDD.n1041 GND 0.16fF
C1549 VDD.n1042 GND 0.01fF
C1550 VDD.n1043 GND 0.02fF
C1551 VDD.n1044 GND 0.02fF
C1552 VDD.n1045 GND 0.16fF
C1553 VDD.n1046 GND 0.02fF
C1554 VDD.n1047 GND 0.02fF
C1555 VDD.n1048 GND 0.03fF
C1556 VDD.n1049 GND 0.15fF
C1557 VDD.n1050 GND 0.02fF
C1558 VDD.n1051 GND 0.02fF
C1559 VDD.n1052 GND 0.03fF
C1560 VDD.n1053 GND 0.17fF
C1561 VDD.n1054 GND 0.01fF
C1562 VDD.n1055 GND 0.08fF
C1563 VDD.n1056 GND 0.05fF
C1564 VDD.n1057 GND 0.02fF
C1565 VDD.n1058 GND 0.02fF
C1566 VDD.n1059 GND 0.17fF
C1567 VDD.n1060 GND 0.01fF
C1568 VDD.n1061 GND 0.02fF
C1569 VDD.n1062 GND 0.02fF
C1570 VDD.n1063 GND 0.23fF
C1571 VDD.n1064 GND 0.01fF
C1572 VDD.n1065 GND 0.07fF
C1573 VDD.n1066 GND 0.02fF
C1574 VDD.n1067 GND 0.29fF
C1575 VDD.n1068 GND 0.01fF
C1576 VDD.n1069 GND 0.02fF
C1577 VDD.n1070 GND 0.02fF
C1578 VDD.n1071 GND 0.29fF
C1579 VDD.n1072 GND 0.01fF
C1580 VDD.n1073 GND 0.02fF
C1581 VDD.n1074 GND 0.04fF
C1582 VDD.n1075 GND 0.27fF
C1583 VDD.n1076 GND 0.02fF
C1584 VDD.n1077 GND 0.02fF
C1585 VDD.n1078 GND 0.02fF
C1586 VDD.n1079 GND 0.06fF
C1587 VDD.n1080 GND 0.02fF
C1588 VDD.n1081 GND 0.02fF
C1589 VDD.n1082 GND 0.02fF
C1590 VDD.n1083 GND 0.02fF
C1591 VDD.n1084 GND 0.02fF
C1592 VDD.n1085 GND 0.02fF
C1593 VDD.n1086 GND 0.02fF
C1594 VDD.n1087 GND 0.02fF
C1595 VDD.n1088 GND 0.02fF
C1596 VDD.n1089 GND 0.02fF
C1597 VDD.n1090 GND 0.03fF
C1598 VDD.n1091 GND 0.02fF
C1599 VDD.n1092 GND 0.02fF
C1600 VDD.n1096 GND 0.29fF
C1601 VDD.n1097 GND 0.29fF
C1602 VDD.n1098 GND 0.01fF
C1603 VDD.n1099 GND 0.02fF
C1604 VDD.n1100 GND 0.04fF
C1605 VDD.n1101 GND 0.07fF
C1606 VDD.n1102 GND 0.26fF
C1607 VDD.n1103 GND 0.01fF
C1608 VDD.n1104 GND 0.01fF
C1609 VDD.n1105 GND 0.02fF
C1610 VDD.n1106 GND 0.17fF
C1611 VDD.n1107 GND 0.01fF
C1612 VDD.n1108 GND 0.02fF
C1613 VDD.n1109 GND 0.02fF
C1614 VDD.n1110 GND 0.15fF
C1615 VDD.n1111 GND 0.01fF
C1616 VDD.n1112 GND 0.02fF
C1617 VDD.n1113 GND 0.03fF
C1618 VDD.n1114 GND 0.08fF
C1619 VDD.n1115 GND 0.05fF
C1620 VDD.n1116 GND 0.01fF
C1621 VDD.n1117 GND 0.02fF
C1622 VDD.n1118 GND 0.03fF
C1623 VDD.n1119 GND 0.17fF
C1624 VDD.n1120 GND 0.01fF
C1625 VDD.n1121 GND 0.02fF
C1626 VDD.n1122 GND 0.02fF
C1627 VDD.n1123 GND 0.06fF
C1628 VDD.n1124 GND 0.25fF
C1629 VDD.n1125 GND 0.01fF
C1630 VDD.n1126 GND 0.01fF
C1631 VDD.n1127 GND 0.02fF
C1632 VDD.n1128 GND 0.29fF
C1633 VDD.n1129 GND 0.01fF
C1634 VDD.n1130 GND 0.02fF
C1635 VDD.n1131 GND 0.04fF
C1636 VDD.n1132 GND 0.27fF
C1637 VDD.n1133 GND 0.02fF
C1638 VDD.n1134 GND 0.02fF
C1639 VDD.n1135 GND 0.02fF
C1640 VDD.n1136 GND 0.06fF
C1641 VDD.n1137 GND 0.02fF
C1642 VDD.n1138 GND 0.02fF
C1643 VDD.n1139 GND 0.02fF
C1644 VDD.n1140 GND 0.02fF
C1645 VDD.n1141 GND 0.02fF
C1646 VDD.n1142 GND 0.02fF
C1647 VDD.n1143 GND 0.02fF
C1648 VDD.n1144 GND 0.02fF
C1649 VDD.n1145 GND 0.02fF
C1650 VDD.n1146 GND 0.02fF
C1651 VDD.n1147 GND 0.03fF
C1652 VDD.n1148 GND 0.02fF
C1653 VDD.n1149 GND 0.02fF
C1654 VDD.n1153 GND 0.29fF
C1655 VDD.n1154 GND 0.29fF
C1656 VDD.n1155 GND 0.01fF
C1657 VDD.n1156 GND 0.02fF
C1658 VDD.n1157 GND 0.04fF
C1659 VDD.n1158 GND 0.29fF
C1660 VDD.n1159 GND 0.01fF
C1661 VDD.n1160 GND 0.02fF
C1662 VDD.n1161 GND 0.02fF
C1663 VDD.n1162 GND 0.07fF
C1664 VDD.n1163 GND 0.23fF
C1665 VDD.n1164 GND 0.01fF
C1666 VDD.n1165 GND 0.01fF
C1667 VDD.n1166 GND 0.02fF
C1668 VDD.n1167 GND 0.17fF
C1669 VDD.n1168 GND 0.01fF
C1670 VDD.n1169 GND 0.02fF
C1671 VDD.n1170 GND 0.02fF
C1672 VDD.n1171 GND 0.08fF
C1673 VDD.n1172 GND 0.05fF
C1674 VDD.n1173 GND 0.16fF
C1675 VDD.n1174 GND 0.01fF
C1676 VDD.n1175 GND 0.02fF
C1677 VDD.n1176 GND 0.02fF
C1678 VDD.n1177 GND 0.16fF
C1679 VDD.n1178 GND 0.02fF
C1680 VDD.n1179 GND 0.02fF
C1681 VDD.n1180 GND 0.03fF
C1682 VDD.n1181 GND 0.15fF
C1683 VDD.n1182 GND 0.02fF
C1684 VDD.n1183 GND 0.02fF
C1685 VDD.n1184 GND 0.03fF
C1686 VDD.n1185 GND 0.17fF
C1687 VDD.n1186 GND 0.01fF
C1688 VDD.n1187 GND 0.08fF
C1689 VDD.n1188 GND 0.05fF
C1690 VDD.n1189 GND 0.02fF
C1691 VDD.n1190 GND 0.02fF
C1692 VDD.n1191 GND 0.17fF
C1693 VDD.n1192 GND 0.01fF
C1694 VDD.n1193 GND 0.02fF
C1695 VDD.n1194 GND 0.02fF
C1696 VDD.n1195 GND 0.23fF
C1697 VDD.n1196 GND 0.01fF
C1698 VDD.n1197 GND 0.07fF
C1699 VDD.n1198 GND 0.02fF
C1700 VDD.n1199 GND 0.29fF
C1701 VDD.n1200 GND 0.01fF
C1702 VDD.n1201 GND 0.02fF
C1703 VDD.n1202 GND 0.02fF
C1704 VDD.n1203 GND 0.29fF
C1705 VDD.n1204 GND 0.01fF
C1706 VDD.n1205 GND 0.02fF
C1707 VDD.n1206 GND 0.04fF
C1708 VDD.n1207 GND 0.32fF
C1709 VDD.n1208 GND 0.02fF
C1710 VDD.n1209 GND 0.02fF
C1711 VDD.n1210 GND 0.02fF
C1712 VDD.n1211 GND 0.06fF
C1713 VDD.n1212 GND 0.02fF
C1714 VDD.n1213 GND 0.02fF
C1715 VDD.n1214 GND 0.02fF
C1716 VDD.n1215 GND 0.02fF
C1717 VDD.n1216 GND 0.02fF
C1718 VDD.n1217 GND 0.02fF
C1719 VDD.n1218 GND 0.02fF
C1720 VDD.n1219 GND 0.02fF
C1721 VDD.n1220 GND 0.02fF
C1722 VDD.n1221 GND 0.02fF
C1723 VDD.n1222 GND 0.03fF
C1724 VDD.n1223 GND 0.02fF
C1725 VDD.n1224 GND 0.02fF
C1726 VDD.n1228 GND 0.29fF
C1727 VDD.n1229 GND 0.29fF
C1728 VDD.n1230 GND 0.01fF
C1729 VDD.n1231 GND 0.02fF
C1730 VDD.n1232 GND 0.04fF
C1731 VDD.n1233 GND 0.29fF
C1732 VDD.n1234 GND 0.01fF
C1733 VDD.n1235 GND 0.02fF
C1734 VDD.n1236 GND 0.02fF
C1735 VDD.n1237 GND 0.07fF
C1736 VDD.n1238 GND 0.23fF
C1737 VDD.n1239 GND 0.01fF
C1738 VDD.n1240 GND 0.01fF
C1739 VDD.n1241 GND 0.02fF
C1740 VDD.n1242 GND 0.17fF
C1741 VDD.n1243 GND 0.01fF
C1742 VDD.n1244 GND 0.02fF
C1743 VDD.n1245 GND 0.02fF
C1744 VDD.n1246 GND 0.08fF
C1745 VDD.n1247 GND 0.05fF
C1746 VDD.n1248 GND 0.16fF
C1747 VDD.n1249 GND 0.01fF
C1748 VDD.n1250 GND 0.02fF
C1749 VDD.n1251 GND 0.02fF
C1750 VDD.n1252 GND 0.16fF
C1751 VDD.n1253 GND 0.02fF
C1752 VDD.n1254 GND 0.02fF
C1753 VDD.n1255 GND 0.03fF
C1754 VDD.n1256 GND 0.15fF
C1755 VDD.n1257 GND 0.02fF
C1756 VDD.n1258 GND 0.02fF
C1757 VDD.n1259 GND 0.03fF
C1758 VDD.n1260 GND 0.17fF
C1759 VDD.n1261 GND 0.01fF
C1760 VDD.n1262 GND 0.08fF
C1761 VDD.n1263 GND 0.05fF
C1762 VDD.n1264 GND 0.02fF
C1763 VDD.n1265 GND 0.02fF
C1764 VDD.n1266 GND 0.17fF
C1765 VDD.n1267 GND 0.01fF
C1766 VDD.n1268 GND 0.02fF
C1767 VDD.n1269 GND 0.02fF
C1768 VDD.n1270 GND 0.23fF
C1769 VDD.n1271 GND 0.01fF
C1770 VDD.n1272 GND 0.07fF
C1771 VDD.n1273 GND 0.02fF
C1772 VDD.n1274 GND 0.29fF
C1773 VDD.n1275 GND 