magic
tech sky130A
magscale 1 2
timestamp 1648750605
<< locali >>
rect 15819 575 15853 609
<< metal1 >>
rect 55 1505 89 1539
rect 1378 945 14855 979
rect 171 871 11787 905
rect 11971 871 18230 905
rect 11971 831 12005 871
rect 11413 797 12005 831
rect 17185 797 17435 831
rect 19149 797 19183 831
rect 4679 723 4995 757
rect 10453 723 10766 757
rect 16224 723 16566 757
rect 4531 649 18515 683
rect 10314 575 11425 609
rect 16077 575 17184 609
rect 427 501 15854 535
rect 2344 427 14020 461
rect 55 13 89 47
use li1_M1_contact  li1_M1_contact_9 pcells
timestamp 1648061256
transform 1 0 5032 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_8
timestamp 1648061256
transform -1 0 4662 0 -1 740
box -53 -33 29 33
use dffsnrnx1_pcell  dffsnrnx1_pcell_0 pcells
timestamp 1648742386
transform 1 0 0 0 1 0
box -84 0 5856 1575
use dffsnrnx1_pcell  dffsnrnx1_pcell_1
timestamp 1648742386
transform 1 0 5772 0 1 0
box -84 0 5856 1575
use li1_M1_contact  li1_M1_contact_20
timestamp 1648061256
transform 1 0 5624 0 1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_15
timestamp 1648061256
transform -1 0 4514 0 -1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform 1 0 222 0 1 888
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_11
timestamp 1648061256
transform 1 0 10804 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_10
timestamp 1648061256
transform -1 0 10434 0 -1 740
box -53 -33 29 33
use dffsnrnx1_pcell  dffsnrnx1_pcell_2
timestamp 1648742386
transform 1 0 11544 0 1 0
box -84 0 5856 1575
use li1_M1_contact  li1_M1_contact_7
timestamp 1648061256
transform 1 0 11396 0 1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_5
timestamp 1648061256
transform -1 0 10286 0 -1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_3
timestamp 1648061256
transform -1 0 11396 0 -1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_2
timestamp 1648061256
transform -1 0 11766 0 -1 888
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform -1 0 5994 0 -1 888
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_17
timestamp 1648061256
transform 1 0 17464 0 -1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_14
timestamp 1648061256
transform 1 0 16576 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_13
timestamp 1648061256
transform -1 0 16206 0 -1 740
box -53 -33 29 33
use votern3x1_pcell  votern3x1_pcell_0 pcells
timestamp 1648740297
transform 1 0 17316 0 1 0
box -84 0 2082 1575
use li1_M1_contact  li1_M1_contact_19
timestamp 1648061256
transform -1 0 16058 0 -1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_4
timestamp 1648061256
transform 1 0 17168 0 1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_6
timestamp 1648061256
transform -1 0 17168 0 1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_16
timestamp 1648061256
transform -1 0 19166 0 -1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_12
timestamp 1648061256
transform 1 0 18500 0 -1 666
box -53 -33 29 33
<< labels >>
rlabel metal1 19149 797 19183 831 1 QN
port 1 n
rlabel metal1 205 871 239 905 1 D
port 2 n
rlabel metal1 1388 945 1422 979 1 CLK
port 3 n
rlabel metal1 2351 427 2385 461 1 SN
port 4 n
rlabel metal1 427 501 461 535 1 RN
port 5 n
rlabel metal1 55 1505 89 1539 1 VDD
port 6 n
rlabel metal1 55 13 89 47 1 VSS
port 7 n
<< end >>
