* SPICE3 file created from NOR2X1.ext - technology: sky130A

.subckt NOR2X1 Y A B VDD VSS
X0 a_131_1051# A VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8p ps=4.58u w=2u l=0.15u M=2
X1 Y A VSS VSS sky130_fd_pr__nfet_01v8 ad=3.582p pd=3.15u as=1.9366p ps=1.294u w=3u l=0.15u
X2 a_131_1051# B Y VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8p ps=4.58u w=2u l=0.15u M=2
X3 Y B VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
.ends
