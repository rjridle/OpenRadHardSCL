* SPICE3 file created from AND3X1.ext - technology: sky130A

.subckt AND3X1 Y A B C VDD VSS
X0 VDD B a_277_1050# VDD sky130_fd_pr__pfet_01v8 ad=3.36p pd=2.736u as=0p ps=0u w=2u l=0.15u M=2
X1 VDD C a_277_1050# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X2 Y a_277_1050# VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8p pd=4.58u as=0p ps=0u w=2u l=0.15u M=2
X3 a_277_1050# C a_372_210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X4 a_277_1050# A VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X5 VSS A a_91_103# VSS sky130_fd_pr__nfet_01v8 ad=1.3199p pd=9.67u as=0p ps=0u w=3u l=0.15u
X6 a_372_210# B a_91_103# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X7 Y a_277_1050# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=0p ps=0u w=3u l=0.15u
C0 a_277_1050# VDD 2.88fF
.ends
