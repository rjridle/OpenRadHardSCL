* NGSPICE file created from INVX1.ext - technology: sky130A

.subckt nmos_top a_85_108# a_55_92# a_n1_0# VSUBS
X0 a_85_108# a_55_92# a_n1_0# VSUBS sky130_fd_pr__nfet_01v8 ad=1.772e+11p pd=1.56e+06u as=1.15725e+12p ps=8.12e+06u w=3e+06u l=150000u
.ends

.subckt pmos2 a_144_n460# a_262_n399# a_88_n399# w_52_n435# a_174_n399#
X0 a_174_n399# a_144_n460# a_88_n399# w_52_n435# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.6e+11p ps=4.56e+06u w=2e+06u l=150000u
X1 a_262_n399# a_144_n460# a_174_n399# w_52_n435# sky130_fd_pr__pfet_01v8 ad=5.4e+11p pd=4.54e+06u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt invx1_pcell VSS VDD a_154_410# a_205_1105#
Xnmos_top_0 a_205_1105# a_154_410# VSS VSS nmos_top
Xpmos2_0 a_154_410# VDD VDD VDD a_205_1105# pmos2
.ends

.subckt INVX1 A Y VSS VDD
Xinvx1_pcell_0 VSS VDD A Y invx1_pcell
.ends

