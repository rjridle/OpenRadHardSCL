magic
tech sky130A
magscale 1 2
timestamp 1649361829
<< nwell >>
rect -84 832 2082 1575
<< nmos >>
rect 168 316 198 377
tri 198 316 214 332 sw
rect 362 324 392 377
tri 392 324 408 340 sw
rect 168 286 274 316
tri 274 286 304 316 sw
rect 362 294 468 324
tri 468 294 498 324 sw
rect 168 185 198 286
tri 198 270 214 286 nw
tri 258 270 274 286 ne
tri 198 185 214 201 sw
tri 258 185 274 201 se
rect 274 185 304 286
rect 362 193 392 294
tri 392 278 408 294 nw
tri 452 278 468 294 ne
tri 392 193 408 209 sw
tri 452 193 468 209 se
rect 468 193 498 294
tri 168 155 198 185 ne
rect 198 155 274 185
tri 274 155 304 185 nw
tri 362 163 392 193 ne
rect 392 163 468 193
tri 468 163 498 193 nw
rect 834 316 864 377
tri 864 316 880 332 sw
tri 1118 324 1134 340 se
rect 1134 324 1164 377
rect 834 286 940 316
tri 940 286 970 316 sw
tri 1028 294 1058 324 se
rect 1058 294 1164 324
rect 834 185 864 286
tri 864 270 880 286 nw
tri 924 270 940 286 ne
tri 864 185 880 201 sw
tri 924 185 940 201 se
rect 940 185 970 286
rect 1028 193 1058 294
tri 1058 278 1074 294 nw
tri 1118 278 1134 294 ne
tri 1058 193 1074 209 sw
tri 1118 193 1134 209 se
rect 1134 193 1164 294
tri 834 155 864 185 ne
rect 864 155 940 185
tri 940 155 970 185 nw
tri 1028 163 1058 193 ne
rect 1058 163 1134 193
tri 1134 163 1164 193 nw
rect 1500 316 1530 377
tri 1530 316 1546 332 sw
rect 1694 324 1724 377
tri 1724 324 1740 340 sw
rect 1500 286 1606 316
tri 1606 286 1636 316 sw
rect 1694 294 1800 324
tri 1800 294 1830 324 sw
rect 1500 185 1530 286
tri 1530 270 1546 286 nw
tri 1590 270 1606 286 ne
tri 1530 185 1546 201 sw
tri 1590 185 1606 201 se
rect 1606 185 1636 286
rect 1694 279 1725 294
tri 1725 279 1740 294 nw
tri 1784 279 1799 294 ne
rect 1799 279 1830 294
rect 1694 193 1724 279
tri 1724 193 1740 209 sw
tri 1784 193 1800 209 se
rect 1800 193 1830 279
tri 1500 155 1530 185 ne
rect 1530 155 1606 185
tri 1606 155 1636 185 nw
tri 1694 163 1724 193 ne
rect 1724 163 1800 193
tri 1800 163 1830 193 nw
<< pmos >>
rect 187 1051 217 1451
rect 275 1051 305 1451
rect 363 1051 393 1451
rect 451 1051 481 1451
rect 851 1051 881 1451
rect 939 1051 969 1451
rect 1027 1051 1057 1451
rect 1115 1051 1145 1451
rect 1519 1051 1549 1451
rect 1607 1051 1637 1451
rect 1695 1051 1725 1451
rect 1783 1051 1813 1451
<< ndiff >>
rect 112 361 168 377
rect 112 327 122 361
rect 156 327 168 361
rect 112 289 168 327
rect 198 361 362 377
rect 198 332 219 361
tri 198 316 214 332 ne
rect 214 327 219 332
rect 253 327 316 361
rect 350 327 362 361
rect 214 316 362 327
rect 392 361 552 377
rect 392 340 510 361
tri 392 324 408 340 ne
rect 408 327 510 340
rect 544 327 552 361
rect 408 324 552 327
rect 112 255 122 289
rect 156 255 168 289
tri 274 286 304 316 ne
rect 304 289 362 316
tri 468 294 498 324 ne
rect 112 221 168 255
rect 112 187 122 221
rect 156 187 168 221
rect 112 155 168 187
tri 198 270 214 286 se
rect 214 270 258 286
tri 258 270 274 286 sw
rect 198 236 274 270
rect 198 202 219 236
rect 253 202 274 236
rect 198 201 274 202
tri 198 185 214 201 ne
rect 214 185 258 201
tri 258 185 274 201 nw
rect 304 255 316 289
rect 350 255 362 289
rect 304 221 362 255
rect 304 187 316 221
rect 350 187 362 221
tri 392 278 408 294 se
rect 408 278 452 294
tri 452 278 468 294 sw
rect 392 245 468 278
rect 392 211 412 245
rect 446 211 468 245
rect 392 209 468 211
tri 392 193 408 209 ne
rect 408 193 452 209
tri 452 193 468 209 nw
rect 498 289 552 324
rect 498 255 510 289
rect 544 255 552 289
rect 498 221 552 255
tri 168 155 198 185 sw
tri 274 155 304 185 se
rect 304 163 362 187
tri 362 163 392 193 sw
tri 468 163 498 193 se
rect 498 187 510 221
rect 544 187 552 221
rect 498 163 552 187
rect 304 155 552 163
rect 112 151 552 155
rect 112 117 122 151
rect 156 117 316 151
rect 350 117 412 151
rect 446 117 510 151
rect 544 117 552 151
rect 112 101 552 117
rect 778 361 834 377
rect 778 327 788 361
rect 822 327 834 361
rect 778 289 834 327
rect 864 361 1134 377
rect 864 332 885 361
tri 864 316 880 332 ne
rect 880 327 885 332
rect 919 327 982 361
rect 1016 340 1134 361
rect 1016 327 1118 340
rect 880 324 1118 327
tri 1118 324 1134 340 nw
rect 1164 361 1220 377
rect 1164 327 1176 361
rect 1210 327 1220 361
rect 880 316 1028 324
rect 778 255 788 289
rect 822 255 834 289
tri 940 286 970 316 ne
rect 970 289 1028 316
tri 1028 294 1058 324 nw
rect 778 221 834 255
rect 778 187 788 221
rect 822 187 834 221
rect 778 155 834 187
tri 864 270 880 286 se
rect 880 270 924 286
tri 924 270 940 286 sw
rect 864 236 940 270
rect 864 202 885 236
rect 919 202 940 236
rect 864 201 940 202
tri 864 185 880 201 ne
rect 880 185 924 201
tri 924 185 940 201 nw
rect 970 255 982 289
rect 1016 255 1028 289
rect 970 221 1028 255
rect 970 187 982 221
rect 1016 187 1028 221
tri 1058 278 1074 294 se
rect 1074 278 1118 294
tri 1118 278 1134 294 sw
rect 1058 245 1134 278
rect 1058 211 1079 245
rect 1113 211 1134 245
rect 1058 209 1134 211
tri 1058 193 1074 209 ne
rect 1074 193 1118 209
tri 1118 193 1134 209 nw
rect 1164 289 1220 327
rect 1164 255 1176 289
rect 1210 255 1220 289
rect 1164 221 1220 255
tri 834 155 864 185 sw
tri 940 155 970 185 se
rect 970 163 1028 187
tri 1028 163 1058 193 sw
tri 1134 163 1164 193 se
rect 1164 187 1176 221
rect 1210 187 1220 221
rect 1164 163 1220 187
rect 970 155 1220 163
rect 778 151 1220 155
rect 778 117 788 151
rect 822 117 982 151
rect 1016 117 1079 151
rect 1113 117 1176 151
rect 1210 117 1220 151
rect 778 101 1220 117
rect 1444 361 1500 377
rect 1444 327 1454 361
rect 1488 327 1500 361
rect 1444 289 1500 327
rect 1530 361 1694 377
rect 1530 332 1551 361
tri 1530 316 1546 332 ne
rect 1546 327 1551 332
rect 1585 327 1648 361
rect 1682 327 1694 361
rect 1546 316 1694 327
rect 1724 340 1886 377
tri 1724 324 1740 340 ne
rect 1740 324 1886 340
rect 1444 255 1454 289
rect 1488 255 1500 289
tri 1606 286 1636 316 ne
rect 1636 289 1694 316
tri 1800 294 1830 324 ne
rect 1444 221 1500 255
rect 1444 187 1454 221
rect 1488 187 1500 221
rect 1444 155 1500 187
tri 1530 270 1546 286 se
rect 1546 270 1590 286
tri 1590 270 1606 286 sw
rect 1530 236 1606 270
rect 1530 202 1551 236
rect 1585 202 1606 236
rect 1530 201 1606 202
tri 1530 185 1546 201 ne
rect 1546 185 1590 201
tri 1590 185 1606 201 nw
rect 1636 255 1648 289
rect 1682 255 1694 289
tri 1725 279 1740 294 se
rect 1740 279 1784 294
tri 1784 279 1799 294 sw
rect 1830 289 1886 324
rect 1636 221 1694 255
rect 1636 187 1648 221
rect 1682 187 1694 221
rect 1724 245 1800 279
rect 1724 211 1745 245
rect 1779 211 1800 245
rect 1724 209 1800 211
tri 1724 193 1740 209 ne
rect 1740 193 1784 209
tri 1784 193 1800 209 nw
rect 1830 255 1842 289
rect 1876 255 1886 289
rect 1830 221 1886 255
tri 1500 155 1530 185 sw
tri 1606 155 1636 185 se
rect 1636 163 1694 187
tri 1694 163 1724 193 sw
tri 1800 163 1830 193 se
rect 1830 187 1842 221
rect 1876 187 1886 221
rect 1830 163 1886 187
rect 1636 155 1886 163
rect 1444 151 1886 155
rect 1444 117 1454 151
rect 1488 117 1648 151
rect 1682 117 1745 151
rect 1779 117 1842 151
rect 1876 117 1886 151
rect 1444 101 1886 117
<< pdiff >>
rect 131 1411 187 1451
rect 131 1377 141 1411
rect 175 1377 187 1411
rect 131 1343 187 1377
rect 131 1309 141 1343
rect 175 1309 187 1343
rect 131 1275 187 1309
rect 131 1241 141 1275
rect 175 1241 187 1275
rect 131 1207 187 1241
rect 131 1173 141 1207
rect 175 1173 187 1207
rect 131 1139 187 1173
rect 131 1105 141 1139
rect 175 1105 187 1139
rect 131 1051 187 1105
rect 217 1411 275 1451
rect 217 1377 229 1411
rect 263 1377 275 1411
rect 217 1343 275 1377
rect 217 1309 229 1343
rect 263 1309 275 1343
rect 217 1275 275 1309
rect 217 1241 229 1275
rect 263 1241 275 1275
rect 217 1207 275 1241
rect 217 1173 229 1207
rect 263 1173 275 1207
rect 217 1139 275 1173
rect 217 1105 229 1139
rect 263 1105 275 1139
rect 217 1051 275 1105
rect 305 1411 363 1451
rect 305 1377 317 1411
rect 351 1377 363 1411
rect 305 1343 363 1377
rect 305 1309 317 1343
rect 351 1309 363 1343
rect 305 1275 363 1309
rect 305 1241 317 1275
rect 351 1241 363 1275
rect 305 1207 363 1241
rect 305 1173 317 1207
rect 351 1173 363 1207
rect 305 1051 363 1173
rect 393 1411 451 1451
rect 393 1377 405 1411
rect 439 1377 451 1411
rect 393 1343 451 1377
rect 393 1309 405 1343
rect 439 1309 451 1343
rect 393 1275 451 1309
rect 393 1241 405 1275
rect 439 1241 451 1275
rect 393 1207 451 1241
rect 393 1173 405 1207
rect 439 1173 451 1207
rect 393 1051 451 1173
rect 481 1411 535 1451
rect 481 1377 493 1411
rect 527 1377 535 1411
rect 481 1343 535 1377
rect 481 1309 493 1343
rect 527 1309 535 1343
rect 481 1275 535 1309
rect 481 1241 493 1275
rect 527 1241 535 1275
rect 481 1207 535 1241
rect 481 1173 493 1207
rect 527 1173 535 1207
rect 481 1139 535 1173
rect 481 1105 493 1139
rect 527 1105 535 1139
rect 481 1051 535 1105
rect 797 1411 851 1451
rect 797 1377 805 1411
rect 839 1377 851 1411
rect 797 1343 851 1377
rect 797 1309 805 1343
rect 839 1309 851 1343
rect 797 1275 851 1309
rect 797 1241 805 1275
rect 839 1241 851 1275
rect 797 1207 851 1241
rect 797 1173 805 1207
rect 839 1173 851 1207
rect 797 1051 851 1173
rect 881 1343 939 1451
rect 881 1309 893 1343
rect 927 1309 939 1343
rect 881 1275 939 1309
rect 881 1241 893 1275
rect 927 1241 939 1275
rect 881 1207 939 1241
rect 881 1173 893 1207
rect 927 1173 939 1207
rect 881 1139 939 1173
rect 881 1105 893 1139
rect 927 1105 939 1139
rect 881 1051 939 1105
rect 969 1411 1027 1451
rect 969 1377 981 1411
rect 1015 1377 1027 1411
rect 969 1343 1027 1377
rect 969 1309 981 1343
rect 1015 1309 1027 1343
rect 969 1275 1027 1309
rect 969 1241 981 1275
rect 1015 1241 1027 1275
rect 969 1207 1027 1241
rect 969 1173 981 1207
rect 1015 1173 1027 1207
rect 969 1051 1027 1173
rect 1057 1343 1115 1451
rect 1057 1309 1069 1343
rect 1103 1309 1115 1343
rect 1057 1275 1115 1309
rect 1057 1241 1069 1275
rect 1103 1241 1115 1275
rect 1057 1207 1115 1241
rect 1057 1173 1069 1207
rect 1103 1173 1115 1207
rect 1057 1051 1115 1173
rect 1145 1411 1201 1451
rect 1145 1377 1157 1411
rect 1191 1377 1201 1411
rect 1145 1343 1201 1377
rect 1145 1309 1157 1343
rect 1191 1309 1201 1343
rect 1145 1275 1201 1309
rect 1145 1241 1157 1275
rect 1191 1241 1201 1275
rect 1145 1207 1201 1241
rect 1145 1173 1157 1207
rect 1191 1173 1201 1207
rect 1145 1051 1201 1173
rect 1463 1411 1519 1451
rect 1463 1377 1473 1411
rect 1507 1377 1519 1411
rect 1463 1343 1519 1377
rect 1463 1309 1473 1343
rect 1507 1309 1519 1343
rect 1463 1275 1519 1309
rect 1463 1241 1473 1275
rect 1507 1241 1519 1275
rect 1463 1207 1519 1241
rect 1463 1173 1473 1207
rect 1507 1173 1519 1207
rect 1463 1051 1519 1173
rect 1549 1343 1607 1451
rect 1549 1309 1561 1343
rect 1595 1309 1607 1343
rect 1549 1275 1607 1309
rect 1549 1241 1561 1275
rect 1595 1241 1607 1275
rect 1549 1207 1607 1241
rect 1549 1173 1561 1207
rect 1595 1173 1607 1207
rect 1549 1139 1607 1173
rect 1549 1105 1561 1139
rect 1595 1105 1607 1139
rect 1549 1051 1607 1105
rect 1637 1411 1695 1451
rect 1637 1377 1649 1411
rect 1683 1377 1695 1411
rect 1637 1343 1695 1377
rect 1637 1309 1649 1343
rect 1683 1309 1695 1343
rect 1637 1275 1695 1309
rect 1637 1241 1649 1275
rect 1683 1241 1695 1275
rect 1637 1207 1695 1241
rect 1637 1173 1649 1207
rect 1683 1173 1695 1207
rect 1637 1051 1695 1173
rect 1725 1343 1783 1451
rect 1725 1309 1737 1343
rect 1771 1309 1783 1343
rect 1725 1275 1783 1309
rect 1725 1241 1737 1275
rect 1771 1241 1783 1275
rect 1725 1207 1783 1241
rect 1725 1173 1737 1207
rect 1771 1173 1783 1207
rect 1725 1139 1783 1173
rect 1725 1105 1737 1139
rect 1771 1105 1783 1139
rect 1725 1051 1783 1105
rect 1813 1411 1867 1451
rect 1813 1377 1825 1411
rect 1859 1377 1867 1411
rect 1813 1343 1867 1377
rect 1813 1309 1825 1343
rect 1859 1309 1867 1343
rect 1813 1275 1867 1309
rect 1813 1241 1825 1275
rect 1859 1241 1867 1275
rect 1813 1207 1867 1241
rect 1813 1173 1825 1207
rect 1859 1173 1867 1207
rect 1813 1051 1867 1173
<< ndiffc >>
rect 122 327 156 361
rect 219 327 253 361
rect 316 327 350 361
rect 510 327 544 361
rect 122 255 156 289
rect 122 187 156 221
rect 219 202 253 236
rect 316 255 350 289
rect 316 187 350 221
rect 412 211 446 245
rect 510 255 544 289
rect 510 187 544 221
rect 122 117 156 151
rect 316 117 350 151
rect 412 117 446 151
rect 510 117 544 151
rect 788 327 822 361
rect 885 327 919 361
rect 982 327 1016 361
rect 1176 327 1210 361
rect 788 255 822 289
rect 788 187 822 221
rect 885 202 919 236
rect 982 255 1016 289
rect 982 187 1016 221
rect 1079 211 1113 245
rect 1176 255 1210 289
rect 1176 187 1210 221
rect 788 117 822 151
rect 982 117 1016 151
rect 1079 117 1113 151
rect 1176 117 1210 151
rect 1454 327 1488 361
rect 1551 327 1585 361
rect 1648 327 1682 361
rect 1454 255 1488 289
rect 1454 187 1488 221
rect 1551 202 1585 236
rect 1648 255 1682 289
rect 1648 187 1682 221
rect 1745 211 1779 245
rect 1842 255 1876 289
rect 1842 187 1876 221
rect 1454 117 1488 151
rect 1648 117 1682 151
rect 1745 117 1779 151
rect 1842 117 1876 151
<< pdiffc >>
rect 141 1377 175 1411
rect 141 1309 175 1343
rect 141 1241 175 1275
rect 141 1173 175 1207
rect 141 1105 175 1139
rect 229 1377 263 1411
rect 229 1309 263 1343
rect 229 1241 263 1275
rect 229 1173 263 1207
rect 229 1105 263 1139
rect 317 1377 351 1411
rect 317 1309 351 1343
rect 317 1241 351 1275
rect 317 1173 351 1207
rect 405 1377 439 1411
rect 405 1309 439 1343
rect 405 1241 439 1275
rect 405 1173 439 1207
rect 493 1377 527 1411
rect 493 1309 527 1343
rect 493 1241 527 1275
rect 493 1173 527 1207
rect 493 1105 527 1139
rect 805 1377 839 1411
rect 805 1309 839 1343
rect 805 1241 839 1275
rect 805 1173 839 1207
rect 893 1309 927 1343
rect 893 1241 927 1275
rect 893 1173 927 1207
rect 893 1105 927 1139
rect 981 1377 1015 1411
rect 981 1309 1015 1343
rect 981 1241 1015 1275
rect 981 1173 1015 1207
rect 1069 1309 1103 1343
rect 1069 1241 1103 1275
rect 1069 1173 1103 1207
rect 1157 1377 1191 1411
rect 1157 1309 1191 1343
rect 1157 1241 1191 1275
rect 1157 1173 1191 1207
rect 1473 1377 1507 1411
rect 1473 1309 1507 1343
rect 1473 1241 1507 1275
rect 1473 1173 1507 1207
rect 1561 1309 1595 1343
rect 1561 1241 1595 1275
rect 1561 1173 1595 1207
rect 1561 1105 1595 1139
rect 1649 1377 1683 1411
rect 1649 1309 1683 1343
rect 1649 1241 1683 1275
rect 1649 1173 1683 1207
rect 1737 1309 1771 1343
rect 1737 1241 1771 1275
rect 1737 1173 1771 1207
rect 1737 1105 1771 1139
rect 1825 1377 1859 1411
rect 1825 1309 1859 1343
rect 1825 1241 1859 1275
rect 1825 1173 1859 1207
<< psubdiff >>
rect -31 546 2029 572
rect -31 512 -17 546
rect 17 512 649 546
rect 683 512 1315 546
rect 1349 512 1981 546
rect 2015 512 2029 546
rect -31 510 2029 512
rect -31 474 31 510
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect 635 474 697 510
rect 635 440 649 474
rect 683 440 697 474
rect -31 368 -17 402
rect 17 368 31 402
rect 635 402 697 440
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect 635 368 649 402
rect 683 368 697 402
rect 1301 474 1363 510
rect 1301 440 1315 474
rect 1349 440 1363 474
rect 1301 402 1363 440
rect 1967 474 2029 510
rect 1967 440 1981 474
rect 2015 440 2029 474
rect 635 330 697 368
rect 635 296 649 330
rect 683 296 697 330
rect 635 258 697 296
rect 635 224 649 258
rect 683 224 697 258
rect 635 186 697 224
rect 635 152 649 186
rect 683 152 697 186
rect 635 114 697 152
rect -31 47 31 80
rect 635 80 649 114
rect 683 80 697 114
rect 1301 368 1315 402
rect 1349 368 1363 402
rect 1967 402 2029 440
rect 1301 330 1363 368
rect 1301 296 1315 330
rect 1349 296 1363 330
rect 1301 258 1363 296
rect 1301 224 1315 258
rect 1349 224 1363 258
rect 1301 186 1363 224
rect 1301 152 1315 186
rect 1349 152 1363 186
rect 1301 114 1363 152
rect 635 47 697 80
rect 1301 80 1315 114
rect 1349 80 1363 114
rect 1967 368 1981 402
rect 2015 368 2029 402
rect 1967 330 2029 368
rect 1967 296 1981 330
rect 2015 296 2029 330
rect 1967 258 2029 296
rect 1967 224 1981 258
rect 2015 224 2029 258
rect 1967 186 2029 224
rect 1967 152 1981 186
rect 2015 152 2029 186
rect 1967 114 2029 152
rect 1301 47 1363 80
rect 1967 80 1981 114
rect 2015 80 2029 114
rect 1967 47 2029 80
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 361 47
rect 395 13 433 47
rect 467 13 505 47
rect 539 13 577 47
rect 611 13 721 47
rect 755 13 793 47
rect 827 13 865 47
rect 899 13 937 47
rect 971 13 1027 47
rect 1061 13 1099 47
rect 1133 13 1171 47
rect 1205 13 1243 47
rect 1277 13 1387 47
rect 1421 13 1459 47
rect 1493 13 1531 47
rect 1565 13 1603 47
rect 1637 13 1693 47
rect 1727 13 1765 47
rect 1799 13 1837 47
rect 1871 13 1909 47
rect 1943 13 2029 47
rect -31 11 31 13
rect 635 11 697 13
rect 1301 11 1363 13
rect 1967 11 2029 13
<< nsubdiff >>
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 361 1539
rect 395 1505 433 1539
rect 467 1505 505 1539
rect 539 1505 577 1539
rect 611 1505 721 1539
rect 755 1505 793 1539
rect 827 1505 865 1539
rect 899 1505 937 1539
rect 971 1505 1027 1539
rect 1061 1505 1099 1539
rect 1133 1505 1171 1539
rect 1205 1505 1243 1539
rect 1277 1505 1387 1539
rect 1421 1505 1459 1539
rect 1493 1505 1531 1539
rect 1565 1505 1603 1539
rect 1637 1505 1693 1539
rect 1727 1505 1765 1539
rect 1799 1505 1837 1539
rect 1871 1505 1909 1539
rect 1943 1505 2029 1539
rect -31 1470 31 1505
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect 635 1470 697 1505
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect -31 1038 31 1076
rect 635 1436 649 1470
rect 683 1436 697 1470
rect 1301 1470 1363 1505
rect 635 1398 697 1436
rect 635 1364 649 1398
rect 683 1364 697 1398
rect 635 1326 697 1364
rect 635 1292 649 1326
rect 683 1292 697 1326
rect 635 1254 697 1292
rect 635 1220 649 1254
rect 683 1220 697 1254
rect 635 1182 697 1220
rect 635 1148 649 1182
rect 683 1148 697 1182
rect 635 1110 697 1148
rect 635 1076 649 1110
rect 683 1076 697 1110
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect 635 1038 697 1076
rect 1301 1436 1315 1470
rect 1349 1436 1363 1470
rect 1967 1470 2029 1505
rect 1301 1398 1363 1436
rect 1301 1364 1315 1398
rect 1349 1364 1363 1398
rect 1301 1326 1363 1364
rect 1301 1292 1315 1326
rect 1349 1292 1363 1326
rect 1301 1254 1363 1292
rect 1301 1220 1315 1254
rect 1349 1220 1363 1254
rect 1301 1182 1363 1220
rect 1301 1148 1315 1182
rect 1349 1148 1363 1182
rect 1301 1110 1363 1148
rect 1301 1076 1315 1110
rect 1349 1076 1363 1110
rect 635 1004 649 1038
rect 683 1004 697 1038
rect 635 966 697 1004
rect -31 930 31 932
rect 635 932 649 966
rect 683 932 697 966
rect 1301 1038 1363 1076
rect 1967 1436 1981 1470
rect 2015 1436 2029 1470
rect 1967 1398 2029 1436
rect 1967 1364 1981 1398
rect 2015 1364 2029 1398
rect 1967 1326 2029 1364
rect 1967 1292 1981 1326
rect 2015 1292 2029 1326
rect 1967 1254 2029 1292
rect 1967 1220 1981 1254
rect 2015 1220 2029 1254
rect 1967 1182 2029 1220
rect 1967 1148 1981 1182
rect 2015 1148 2029 1182
rect 1967 1110 2029 1148
rect 1967 1076 1981 1110
rect 2015 1076 2029 1110
rect 1301 1004 1315 1038
rect 1349 1004 1363 1038
rect 1301 966 1363 1004
rect 635 930 697 932
rect 1301 932 1315 966
rect 1349 932 1363 966
rect 1967 1038 2029 1076
rect 1967 1004 1981 1038
rect 2015 1004 2029 1038
rect 1967 966 2029 1004
rect 1301 930 1363 932
rect 1967 932 1981 966
rect 2015 932 2029 966
rect 1967 930 2029 932
rect -31 868 2029 930
<< psubdiffcont >>
rect -17 512 17 546
rect 649 512 683 546
rect 1315 512 1349 546
rect 1981 512 2015 546
rect -17 440 17 474
rect 649 440 683 474
rect -17 368 17 402
rect -17 296 17 330
rect -17 224 17 258
rect -17 152 17 186
rect -17 80 17 114
rect 649 368 683 402
rect 1315 440 1349 474
rect 1981 440 2015 474
rect 649 296 683 330
rect 649 224 683 258
rect 649 152 683 186
rect 649 80 683 114
rect 1315 368 1349 402
rect 1315 296 1349 330
rect 1315 224 1349 258
rect 1315 152 1349 186
rect 1315 80 1349 114
rect 1981 368 2015 402
rect 1981 296 2015 330
rect 1981 224 2015 258
rect 1981 152 2015 186
rect 1981 80 2015 114
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 361 13 395 47
rect 433 13 467 47
rect 505 13 539 47
rect 577 13 611 47
rect 721 13 755 47
rect 793 13 827 47
rect 865 13 899 47
rect 937 13 971 47
rect 1027 13 1061 47
rect 1099 13 1133 47
rect 1171 13 1205 47
rect 1243 13 1277 47
rect 1387 13 1421 47
rect 1459 13 1493 47
rect 1531 13 1565 47
rect 1603 13 1637 47
rect 1693 13 1727 47
rect 1765 13 1799 47
rect 1837 13 1871 47
rect 1909 13 1943 47
<< nsubdiffcont >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 361 1505 395 1539
rect 433 1505 467 1539
rect 505 1505 539 1539
rect 577 1505 611 1539
rect 721 1505 755 1539
rect 793 1505 827 1539
rect 865 1505 899 1539
rect 937 1505 971 1539
rect 1027 1505 1061 1539
rect 1099 1505 1133 1539
rect 1171 1505 1205 1539
rect 1243 1505 1277 1539
rect 1387 1505 1421 1539
rect 1459 1505 1493 1539
rect 1531 1505 1565 1539
rect 1603 1505 1637 1539
rect 1693 1505 1727 1539
rect 1765 1505 1799 1539
rect 1837 1505 1871 1539
rect 1909 1505 1943 1539
rect -17 1436 17 1470
rect -17 1364 17 1398
rect -17 1292 17 1326
rect -17 1220 17 1254
rect -17 1148 17 1182
rect -17 1076 17 1110
rect 649 1436 683 1470
rect 649 1364 683 1398
rect 649 1292 683 1326
rect 649 1220 683 1254
rect 649 1148 683 1182
rect 649 1076 683 1110
rect -17 1004 17 1038
rect -17 932 17 966
rect 1315 1436 1349 1470
rect 1315 1364 1349 1398
rect 1315 1292 1349 1326
rect 1315 1220 1349 1254
rect 1315 1148 1349 1182
rect 1315 1076 1349 1110
rect 649 1004 683 1038
rect 649 932 683 966
rect 1981 1436 2015 1470
rect 1981 1364 2015 1398
rect 1981 1292 2015 1326
rect 1981 1220 2015 1254
rect 1981 1148 2015 1182
rect 1981 1076 2015 1110
rect 1315 1004 1349 1038
rect 1315 932 1349 966
rect 1981 1004 2015 1038
rect 1981 932 2015 966
<< poly >>
rect 187 1451 217 1477
rect 275 1451 305 1477
rect 363 1451 393 1477
rect 451 1451 481 1477
rect 851 1451 881 1477
rect 939 1451 969 1477
rect 1027 1451 1057 1477
rect 1115 1451 1145 1477
rect 187 1020 217 1051
rect 275 1020 305 1051
rect 363 1020 393 1051
rect 451 1020 481 1051
rect 121 1004 305 1020
rect 121 970 131 1004
rect 165 990 305 1004
rect 351 1004 481 1020
rect 165 970 175 990
rect 121 954 175 970
rect 351 970 361 1004
rect 395 990 481 1004
rect 1519 1451 1549 1477
rect 1607 1451 1637 1477
rect 1695 1451 1725 1477
rect 1783 1451 1813 1477
rect 395 970 405 990
rect 351 954 405 970
rect 851 1020 881 1051
rect 939 1020 969 1051
rect 851 1004 969 1020
rect 851 990 871 1004
rect 861 970 871 990
rect 905 990 969 1004
rect 1027 1020 1057 1051
rect 1115 1020 1145 1051
rect 1027 1004 1211 1020
rect 1027 990 1167 1004
rect 905 970 915 990
rect 861 954 915 970
rect 1157 970 1167 990
rect 1201 970 1211 1004
rect 1157 954 1211 970
rect 1519 1020 1549 1051
rect 1607 1020 1637 1051
rect 1695 1020 1725 1051
rect 1783 1020 1813 1051
rect 1453 1004 1637 1020
rect 1453 970 1463 1004
rect 1497 990 1637 1004
rect 1679 1004 1813 1020
rect 1497 970 1507 990
rect 1453 954 1507 970
rect 1679 970 1689 1004
rect 1723 990 1813 1004
rect 1723 970 1733 990
rect 1679 954 1733 970
rect 121 461 175 477
rect 121 427 131 461
rect 165 441 175 461
rect 343 461 397 477
rect 165 427 198 441
rect 121 411 198 427
rect 343 427 353 461
rect 387 427 397 461
rect 343 411 397 427
rect 861 461 915 477
rect 861 441 871 461
rect 168 377 198 411
rect 362 377 392 411
rect 834 427 871 441
rect 905 427 915 461
rect 1157 461 1211 477
rect 1157 441 1167 461
rect 834 411 915 427
rect 1134 427 1167 441
rect 1201 427 1211 461
rect 1134 411 1211 427
rect 834 377 864 411
rect 1134 377 1164 411
rect 1453 461 1507 477
rect 1453 427 1463 461
rect 1497 441 1507 461
rect 1675 461 1729 477
rect 1497 427 1530 441
rect 1453 411 1530 427
rect 1675 427 1685 461
rect 1719 427 1729 461
rect 1675 411 1729 427
rect 1500 377 1530 411
rect 1694 377 1724 411
<< polycont >>
rect 131 970 165 1004
rect 361 970 395 1004
rect 871 970 905 1004
rect 1167 970 1201 1004
rect 1463 970 1497 1004
rect 1689 970 1723 1004
rect 131 427 165 461
rect 353 427 387 461
rect 871 427 905 461
rect 1167 427 1201 461
rect 1463 427 1497 461
rect 1685 427 1719 461
<< locali >>
rect -31 1539 2029 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 361 1539
rect 395 1505 433 1539
rect 467 1505 505 1539
rect 539 1505 577 1539
rect 611 1505 721 1539
rect 755 1505 793 1539
rect 827 1505 865 1539
rect 899 1505 937 1539
rect 971 1505 1027 1539
rect 1061 1505 1099 1539
rect 1133 1505 1171 1539
rect 1205 1505 1243 1539
rect 1277 1505 1387 1539
rect 1421 1505 1459 1539
rect 1493 1505 1531 1539
rect 1565 1505 1603 1539
rect 1637 1505 1693 1539
rect 1727 1505 1765 1539
rect 1799 1505 1837 1539
rect 1871 1505 1909 1539
rect 1943 1505 2029 1539
rect -31 1492 2029 1505
rect -31 1470 31 1492
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect -31 1038 31 1076
rect 141 1411 175 1492
rect 141 1343 175 1377
rect 141 1275 175 1309
rect 141 1207 175 1241
rect 141 1139 175 1173
rect 141 1071 175 1105
rect 229 1411 265 1445
rect 317 1411 351 1492
rect 229 1343 263 1377
rect 229 1275 263 1309
rect 229 1207 263 1241
rect 229 1139 263 1173
rect 317 1343 351 1377
rect 317 1275 351 1309
rect 317 1207 351 1241
rect 317 1157 351 1173
rect 405 1411 439 1445
rect 405 1343 439 1377
rect 405 1275 439 1309
rect 405 1207 439 1241
rect 405 1105 439 1173
rect 229 1071 405 1105
rect 493 1411 527 1492
rect 493 1343 527 1377
rect 493 1275 527 1309
rect 493 1207 527 1241
rect 493 1139 527 1173
rect 493 1071 527 1105
rect 635 1470 697 1492
rect 635 1436 649 1470
rect 683 1436 697 1470
rect 1301 1470 1363 1492
rect 635 1398 697 1436
rect 635 1364 649 1398
rect 683 1364 697 1398
rect 635 1326 697 1364
rect 635 1292 649 1326
rect 683 1292 697 1326
rect 635 1254 697 1292
rect 635 1220 649 1254
rect 683 1220 697 1254
rect 635 1182 697 1220
rect 635 1148 649 1182
rect 683 1148 697 1182
rect 635 1110 697 1148
rect 635 1076 649 1110
rect 683 1076 697 1110
rect 405 1055 439 1071
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect 635 1038 697 1076
rect 805 1411 1191 1445
rect 805 1343 839 1377
rect 805 1275 839 1309
rect 805 1207 839 1241
rect 805 1105 839 1173
rect 893 1343 927 1359
rect 893 1275 927 1309
rect 893 1207 927 1241
rect 893 1139 927 1173
rect 981 1343 1015 1377
rect 981 1275 1015 1309
rect 981 1207 1015 1241
rect 981 1157 1015 1173
rect 1069 1343 1103 1359
rect 1069 1275 1103 1309
rect 1069 1207 1103 1241
rect 1069 1105 1103 1173
rect 1157 1343 1191 1377
rect 1157 1275 1191 1309
rect 1157 1207 1191 1241
rect 1157 1121 1191 1173
rect 1301 1436 1315 1470
rect 1349 1436 1363 1470
rect 1967 1470 2029 1492
rect 1301 1398 1363 1436
rect 1301 1364 1315 1398
rect 1349 1364 1363 1398
rect 1301 1326 1363 1364
rect 1301 1292 1315 1326
rect 1349 1292 1363 1326
rect 1301 1254 1363 1292
rect 1301 1220 1315 1254
rect 1349 1220 1363 1254
rect 1301 1182 1363 1220
rect 1301 1148 1315 1182
rect 1349 1148 1363 1182
rect 893 1071 1069 1105
rect 805 1055 839 1071
rect 1069 1055 1103 1071
rect 1301 1110 1363 1148
rect 1301 1076 1315 1110
rect 1349 1076 1363 1110
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect -31 868 31 932
rect 131 1004 165 1020
rect 361 1004 395 1020
rect -31 546 31 572
rect -31 512 -17 546
rect 17 512 31 546
rect -31 474 31 512
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect 131 461 165 945
rect 131 411 165 427
rect 353 970 361 988
rect 353 954 395 970
rect 635 1004 649 1038
rect 683 1004 697 1038
rect 1301 1038 1363 1076
rect 1473 1411 1859 1445
rect 1473 1343 1507 1377
rect 1473 1275 1507 1309
rect 1473 1207 1507 1241
rect 1473 1105 1507 1173
rect 1561 1343 1595 1359
rect 1561 1275 1595 1309
rect 1561 1207 1595 1241
rect 1561 1139 1595 1173
rect 1649 1343 1683 1377
rect 1649 1275 1683 1309
rect 1649 1207 1683 1241
rect 1649 1157 1683 1173
rect 1737 1343 1771 1359
rect 1737 1275 1771 1309
rect 1737 1207 1771 1241
rect 1737 1139 1771 1173
rect 1825 1343 1859 1377
rect 1825 1275 1859 1309
rect 1825 1207 1859 1241
rect 1825 1157 1859 1173
rect 1967 1436 1981 1470
rect 2015 1436 2029 1470
rect 1967 1398 2029 1436
rect 1967 1364 1981 1398
rect 2015 1364 2029 1398
rect 1967 1326 2029 1364
rect 1967 1292 1981 1326
rect 2015 1292 2029 1326
rect 1967 1254 2029 1292
rect 1967 1220 1981 1254
rect 2015 1220 2029 1254
rect 1967 1182 2029 1220
rect 1967 1148 1981 1182
rect 2015 1148 2029 1182
rect 1967 1110 2029 1148
rect 1561 1071 1867 1105
rect 1473 1055 1507 1071
rect 635 966 697 1004
rect 353 905 387 954
rect 353 461 387 871
rect 635 932 649 966
rect 683 932 697 966
rect 635 868 697 932
rect 871 1004 905 1020
rect 353 411 387 427
rect 635 546 697 572
rect 635 512 649 546
rect 683 512 697 546
rect 635 474 697 512
rect 635 440 649 474
rect 683 440 697 474
rect -31 368 -17 402
rect 17 368 31 402
rect 635 402 697 440
rect 871 461 905 945
rect 871 411 905 427
rect 1167 1004 1201 1020
rect 1167 461 1201 970
rect 1301 1004 1315 1038
rect 1349 1004 1363 1038
rect 1301 966 1363 1004
rect 1301 932 1315 966
rect 1349 932 1363 966
rect 1301 868 1363 932
rect 1463 1004 1497 1020
rect 1167 411 1201 427
rect 1301 546 1363 572
rect 1301 512 1315 546
rect 1349 512 1363 546
rect 1301 474 1363 512
rect 1301 440 1315 474
rect 1349 440 1363 474
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect 122 361 156 377
rect 316 361 350 377
rect 156 327 219 361
rect 253 327 316 361
rect 122 289 156 327
rect 122 221 156 255
rect 316 289 350 327
rect 510 361 544 377
rect 413 281 447 297
rect 122 151 156 187
rect 122 101 156 117
rect 219 236 253 252
rect -31 62 31 80
rect 219 62 253 202
rect 316 221 350 255
rect 412 247 413 262
rect 412 245 447 247
rect 446 231 447 245
rect 510 289 544 327
rect 412 195 446 211
rect 510 221 544 255
rect 316 151 350 187
rect 510 151 544 187
rect 350 117 412 151
rect 446 117 510 151
rect 316 101 350 117
rect 510 101 544 117
rect 635 368 649 402
rect 683 368 697 402
rect 1301 402 1363 440
rect 1463 461 1497 970
rect 1463 411 1497 427
rect 1685 1004 1723 1020
rect 1685 970 1689 1004
rect 1685 954 1723 970
rect 1685 905 1719 954
rect 1685 461 1719 871
rect 1685 411 1719 427
rect 1833 831 1867 1071
rect 1967 1076 1981 1110
rect 2015 1076 2029 1110
rect 1967 1038 2029 1076
rect 1967 1004 1981 1038
rect 2015 1004 2029 1038
rect 1967 966 2029 1004
rect 1967 932 1981 966
rect 2015 932 2029 966
rect 1967 868 2029 932
rect 635 330 697 368
rect 635 296 649 330
rect 683 296 697 330
rect 635 258 697 296
rect 635 224 649 258
rect 683 224 697 258
rect 635 186 697 224
rect 635 152 649 186
rect 683 152 697 186
rect 635 114 697 152
rect 635 80 649 114
rect 683 80 697 114
rect 788 361 822 377
rect 982 361 1016 377
rect 822 327 885 361
rect 919 327 982 361
rect 788 289 822 327
rect 788 221 822 255
rect 982 289 1016 327
rect 1176 361 1210 377
rect 788 151 822 187
rect 788 101 822 117
rect 885 236 919 252
rect 635 62 697 80
rect 885 62 919 202
rect 982 221 1016 255
rect 1079 281 1113 297
rect 1079 245 1113 247
rect 1079 195 1113 211
rect 1176 289 1210 327
rect 1176 221 1210 255
rect 982 151 1016 187
rect 1176 151 1210 187
rect 1016 117 1079 151
rect 1113 117 1176 151
rect 982 101 1016 117
rect 1176 101 1210 117
rect 1301 368 1315 402
rect 1349 368 1363 402
rect 1301 330 1363 368
rect 1301 296 1315 330
rect 1349 296 1363 330
rect 1301 258 1363 296
rect 1301 224 1315 258
rect 1349 224 1363 258
rect 1301 186 1363 224
rect 1301 152 1315 186
rect 1349 152 1363 186
rect 1301 114 1363 152
rect 1301 80 1315 114
rect 1349 80 1363 114
rect 1454 361 1488 377
rect 1648 361 1682 377
rect 1833 374 1867 797
rect 1488 327 1551 361
rect 1585 327 1648 361
rect 1454 289 1488 327
rect 1454 221 1488 255
rect 1648 289 1682 327
rect 1454 151 1488 187
rect 1454 101 1488 117
rect 1551 236 1585 252
rect 1301 62 1363 80
rect 1551 62 1585 202
rect 1648 221 1682 255
rect 1745 340 1867 374
rect 1967 546 2029 572
rect 1967 512 1981 546
rect 2015 512 2029 546
rect 1967 474 2029 512
rect 1967 440 1981 474
rect 2015 440 2029 474
rect 1967 402 2029 440
rect 1967 368 1981 402
rect 2015 368 2029 402
rect 1745 281 1779 340
rect 1967 330 2029 368
rect 1745 245 1779 247
rect 1745 195 1779 211
rect 1842 289 1876 306
rect 1842 221 1876 255
rect 1648 151 1682 187
rect 1842 151 1876 187
rect 1682 117 1745 151
rect 1779 117 1842 151
rect 1648 101 1682 117
rect 1842 101 1876 117
rect 1967 296 1981 330
rect 2015 296 2029 330
rect 1967 258 2029 296
rect 1967 224 1981 258
rect 2015 224 2029 258
rect 1967 186 2029 224
rect 1967 152 1981 186
rect 2015 152 2029 186
rect 1967 114 2029 152
rect 1967 80 1981 114
rect 2015 80 2029 114
rect 1967 62 2029 80
rect -31 47 1079 62
rect 1113 47 2029 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 361 47
rect 395 13 433 47
rect 467 13 505 47
rect 539 13 577 47
rect 611 13 721 47
rect 755 13 793 47
rect 827 13 865 47
rect 899 13 937 47
rect 971 13 1027 47
rect 1061 13 1099 47
rect 1133 13 1171 47
rect 1205 13 1243 47
rect 1277 13 1387 47
rect 1421 13 1459 47
rect 1493 13 1531 47
rect 1565 13 1603 47
rect 1637 13 1693 47
rect 1727 13 1765 47
rect 1799 13 1837 47
rect 1871 13 1909 47
rect 1943 13 2029 47
rect -31 0 2029 13
<< viali >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 361 1505 395 1539
rect 433 1505 467 1539
rect 505 1505 539 1539
rect 577 1505 611 1539
rect 721 1505 755 1539
rect 793 1505 827 1539
rect 865 1505 899 1539
rect 937 1505 971 1539
rect 1027 1505 1061 1539
rect 1099 1505 1133 1539
rect 1171 1505 1205 1539
rect 1243 1505 1277 1539
rect 1387 1505 1421 1539
rect 1459 1505 1493 1539
rect 1531 1505 1565 1539
rect 1603 1505 1637 1539
rect 1693 1505 1727 1539
rect 1765 1505 1799 1539
rect 1837 1505 1871 1539
rect 1909 1505 1943 1539
rect 405 1071 439 1105
rect 805 1071 839 1105
rect 1069 1071 1103 1105
rect 131 970 165 979
rect 131 945 165 970
rect 1473 1071 1507 1105
rect 353 871 387 905
rect 871 970 905 979
rect 871 945 905 970
rect 1167 427 1201 461
rect 413 247 447 281
rect 1463 427 1497 461
rect 1685 871 1719 905
rect 1833 797 1867 831
rect 1079 247 1113 281
rect 1745 247 1779 281
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 361 13 395 47
rect 433 13 467 47
rect 505 13 539 47
rect 577 13 611 47
rect 721 13 755 47
rect 793 13 827 47
rect 865 13 899 47
rect 937 13 971 47
rect 1027 13 1061 47
rect 1099 13 1133 47
rect 1171 13 1205 47
rect 1243 13 1277 47
rect 1387 13 1421 47
rect 1459 13 1493 47
rect 1531 13 1565 47
rect 1603 13 1637 47
rect 1693 13 1727 47
rect 1765 13 1799 47
rect 1837 13 1871 47
rect 1909 13 1943 47
<< metal1 >>
rect -31 1539 2029 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 361 1539
rect 395 1505 433 1539
rect 467 1505 505 1539
rect 539 1505 577 1539
rect 611 1505 721 1539
rect 755 1505 793 1539
rect 827 1505 865 1539
rect 899 1505 937 1539
rect 971 1505 1027 1539
rect 1061 1505 1099 1539
rect 1133 1505 1171 1539
rect 1205 1505 1243 1539
rect 1277 1505 1387 1539
rect 1421 1505 1459 1539
rect 1493 1505 1531 1539
rect 1565 1505 1603 1539
rect 1637 1505 1693 1539
rect 1727 1505 1765 1539
rect 1799 1505 1837 1539
rect 1871 1505 1909 1539
rect 1943 1505 2029 1539
rect -31 1492 2029 1505
rect 399 1105 445 1111
rect 799 1105 845 1111
rect 1063 1105 1109 1111
rect 1467 1105 1513 1111
rect 393 1071 405 1105
rect 439 1071 805 1105
rect 839 1071 851 1105
rect 1057 1071 1069 1105
rect 1103 1071 1473 1105
rect 1507 1071 1519 1105
rect 399 1065 445 1071
rect 799 1065 845 1071
rect 1063 1065 1109 1071
rect 1467 1065 1513 1071
rect 125 979 171 985
rect 865 979 911 985
rect 119 945 131 979
rect 165 945 871 979
rect 905 945 917 979
rect 125 939 171 945
rect 865 939 911 945
rect 347 905 393 911
rect 1679 905 1725 911
rect 341 871 353 905
rect 387 871 1685 905
rect 1719 871 1731 905
rect 347 865 393 871
rect 1679 865 1725 871
rect 1827 831 1873 837
rect 1821 797 1833 831
rect 1867 797 1903 831
rect 1827 791 1873 797
rect 1161 461 1207 467
rect 1457 461 1503 467
rect 1155 427 1167 461
rect 1201 427 1463 461
rect 1497 427 1509 461
rect 1161 421 1207 427
rect 1457 421 1503 427
rect 407 281 453 287
rect 1073 281 1119 287
rect 1739 281 1785 287
rect 401 247 413 281
rect 447 247 1079 281
rect 1113 247 1745 281
rect 1779 247 1791 281
rect 407 241 453 247
rect 1073 241 1119 247
rect 1739 241 1785 247
rect -31 47 2029 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 361 47
rect 395 13 433 47
rect 467 13 505 47
rect 539 13 577 47
rect 611 13 721 47
rect 755 13 793 47
rect 827 13 865 47
rect 899 13 937 47
rect 971 13 1027 47
rect 1061 13 1099 47
rect 1133 13 1171 47
rect 1205 13 1243 47
rect 1277 13 1387 47
rect 1421 13 1459 47
rect 1493 13 1531 47
rect 1565 13 1603 47
rect 1637 13 1693 47
rect 1727 13 1765 47
rect 1799 13 1837 47
rect 1871 13 1909 47
rect 1943 13 2029 47
rect -31 0 2029 13
<< labels >>
rlabel metal1 1833 797 1867 831 1 YN
port 1 n
rlabel metal1 353 871 387 905 1 A
port 2 n
rlabel metal1 131 945 165 979 1 B
port 3 n
rlabel metal1 1167 427 1201 461 1 C
port 4 n
rlabel metal1 55 1505 89 1539 1 VDD
port 5 n
rlabel metal1 55 13 89 47 1 VSS
port 6 n
<< end >>
