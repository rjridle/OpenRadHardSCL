* SPICE3 file created from AND3X1.ext - technology: sky130A

.subckt AND3X1 Y A B C
X0 w_n84_832.t15 B.t0 a_277_1050.t6  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X1 w_n84_832.t1 C.t0 a_277_1050.t0 w_n84_832.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X2 Y.t2 a_277_1050.t7 w_n84_832.t11  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X3  饝 A.t1 a_91_103.t0  饝 sky130_fd_pr__nfet_01v8 ad=1.3199p pd=9.67u as=0p ps=0u w=0u l=0u
X4 a_277_1050.t1 A.t0 w_n84_832.t3 �饝 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X5 Y a_277_1050.t8  饝  饝 sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=0p ps=0u w=0u l=0u
X6 a_277_1050.t5 B.t1 w_n84_832.t13  饝 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X7 a_277_1050.t4 C.t2 w_n84_832.t7 �饝 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X8 w_n84_832.t9 a_277_1050.t9 Y.t1  饝 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X9 w_n84_832.t5 A.t2 a_277_1050.t2 �饝 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
C0 C A 0.02fF
C1 B C 0.18fF
C2 B A 0.18fF
R0 B.n0 B.t0 479.223
R1 B.n0 B.t1 375.52
R2 B.n1 B.t2 315.431
R3 B.n1 B.n0 168.611
R4 B B.n1 4.65
R5 a_277_1050.n5 a_277_1050.t9 512.525
R6 a_277_1050.n5 a_277_1050.t7 371.139
R7 a_277_1050.n9 a_277_1050.n7 286.879
R8 a_277_1050.n6 a_277_1050.t8 282.852
R9 a_277_1050.n6 a_277_1050.n5 247.347
R10 a_277_1050.n7 a_277_1050.n4 207.058
R11 a_277_1050.n3 a_277_1050.n2 161.352
R12 a_277_1050.n4 a_277_1050.n0 95.095
R13 a_277_1050.n3 a_277_1050.n1 95.095
R14 a_277_1050.n4 a_277_1050.n3 66.258
R15 a_277_1050.n9 a_277_1050.n8 15.218
R16 a_277_1050.n0 a_277_1050.t0 14.282
R17 a_277_1050.n0 a_277_1050.t4 14.282
R18 a_277_1050.n1 a_277_1050.t6 14.282
R19 a_277_1050.n1 a_277_1050.t5 14.282
R20 a_277_1050.n2 a_277_1050.t2 14.282
R21 a_277_1050.n2 a_277_1050.t1 14.282
R22 a_277_1050.n10 a_277_1050.n9 12.014
R23 a_277_1050.n7 a_277_1050.n6 10.343
R24 w_n84_832.n68 w_n84_832.n57 144.705
R25 w_n84_832.n77 w_n84_832.t1 143.754
R26 w_n84_832.n109 w_n84_832.t3 135.17
R27 w_n84_832.n37 w_n84_832.t11 135.17
R28 w_n84_832.n26 w_n84_832.t9 135.17
R29 w_n84_832.n135 w_n84_832.n134 129.475
R30 w_n84_832.n119 w_n84_832.n118 129.472
R31 w_n84_832.n53 w_n84_832.n52 92.5
R32 w_n84_832.n51 w_n84_832.n50 92.5
R33 w_n84_832.n49 w_n84_832.n48 92.5
R34 w_n84_832.n47 w_n84_832.n46 92.5
R35 w_n84_832.n55 w_n84_832.n54 92.5
R36 w_n84_832.n94 w_n84_832.n93 92.5
R37 w_n84_832.n92 w_n84_832.n91 92.5
R38 w_n84_832.n90 w_n84_832.n89 92.5
R39 w_n84_832.n88 w_n84_832.n87 92.5
R40 w_n84_832.n96 w_n84_832.n95 92.5
R41 w_n84_832.n16 w_n84_832.n3 92.5
R42 w_n84_832.n7 w_n84_832.n6 92.5
R43 w_n84_832.n9 w_n84_832.n8 92.5
R44 w_n84_832.n11 w_n84_832.n10 92.5
R45 w_n84_832.n13 w_n84_832.n12 92.5
R46 w_n84_832.n15 w_n84_832.n14 92.5
R47 w_n84_832.n23 w_n84_832.n22 92.059
R48 w_n84_832.n67 w_n84_832.n66 92.059
R49 w_n84_832.n102 w_n84_832.n101 92.059
R50 w_n84_832.n22 w_n84_832.n18 67.194
R51 w_n84_832.n22 w_n84_832.n19 67.194
R52 w_n84_832.n22 w_n84_832.n20 67.194
R53 w_n84_832.n22 w_n84_832.n21 67.194
R54 w_n84_832.n86 w_n84_832.n85 44.141
R55 w_n84_832.n7 w_n84_832.n5 44.141
R56 w_n84_832.n85 w_n84_832.n83 44.107
R57 w_n84_832.n5 w_n84_832.n4 44.107
R58 w_n84_832.n27  饝 43.472
R59 w_n84_832.n35  43.472
R60 w_n84_832.n22 w_n84_832.n17 41.052
R61 w_n84_832.n98 w_n84_832.n97 39.742
R62 w_n84_832.n65 w_n84_832.n62 39.742
R63 w_n84_832.n65 w_n84_832.n64 39.742
R64 w_n84_832.n61 w_n84_832.n60 39.742
R65 w_n84_832.n85 w_n84_832.n84 38
R66 w_n84_832.n64 w_n84_832.n63 36.774
R67 w_n84_832.n79 w_n84_832.t0 35.8
R68 w_n84_832.n114 �饝 33.243
R69 w_n84_832.n3 w_n84_832.n2 30.923
R70 w_n84_832.n101 w_n84_832.n99 26.38
R71 w_n84_832.n101 w_n84_832.n98 26.38
R72 w_n84_832.n101 w_n84_832.n100 26.38
R73 w_n84_832.n66 w_n84_832.n65 26.38
R74 w_n84_832.n66 w_n84_832.n61 26.38
R75 w_n84_832.n66 w_n84_832.n59 26.38
R76 w_n84_832.n66 w_n84_832.n58 26.38
R77 w_n84_832.n104 w_n84_832.n96 22.915
R78 w_n84_832.n25 w_n84_832.n16 22.915
R79 w_n84_832.n0 �饝 15.343
R80 w_n84_832.n96 w_n84_832.n94 14.864
R81 w_n84_832.n94 w_n84_832.n92 14.864
R82 w_n84_832.n92 w_n84_832.n90 14.864
R83 w_n84_832.n90 w_n84_832.n88 14.864
R84 w_n84_832.n88 w_n84_832.n86 14.864
R85 w_n84_832.n55 w_n84_832.n53 14.864
R86 w_n84_832.n53 w_n84_832.n51 14.864
R87 w_n84_832.n51 w_n84_832.n49 14.864
R88 w_n84_832.n49 w_n84_832.n47 14.864
R89 w_n84_832.n47 w_n84_832.n45 14.864
R90 w_n84_832.n45 w_n84_832.n44 14.864
R91 w_n84_832.n16 w_n84_832.n15 14.864
R92 w_n84_832.n15 w_n84_832.n13 14.864
R93 w_n84_832.n13 w_n84_832.n11 14.864
R94 w_n84_832.n11 w_n84_832.n9 14.864
R95 w_n84_832.n9 w_n84_832.n7 14.864
R96 w_n84_832.n69 w_n84_832.n56 14.864
R97 w_n84_832.n118 w_n84_832.t13 14.282
R98 w_n84_832.n118 w_n84_832.t5 14.282
R99 w_n84_832.n135 w_n84_832.t7 14.282
R100 w_n84_832.t15 w_n84_832.n135 14.282
R101 w_n84_832.n120 �饝 12.786
R102 w_n84_832.n25 w_n84_832.n24 8.855
R103 w_n84_832.n24 w_n84_832.n23 8.855
R104 w_n84_832.n29 w_n84_832.n28 8.855
R105 w_n84_832.n28 w_n84_832.n27 8.855
R106 w_n84_832.n33 w_n84_832.n32 8.855
R107 w_n84_832.n32 w_n84_832.n31 8.855
R108 w_n84_832.n38 w_n84_832.n36 8.855
R109 w_n84_832.n36 w_n84_832.n35 8.855
R110 w_n84_832.n42 w_n84_832.n41 8.855
R111 w_n84_832.n41 w_n84_832.n40 8.855
R112 w_n84_832.n69 w_n84_832.n68 8.855
R113 w_n84_832.n68 w_n84_832.n67 8.855
R114 w_n84_832.n73 w_n84_832.n72 8.855
R115 w_n84_832.n72 w_n84_832.n71 8.855
R116 w_n84_832.n77 w_n84_832.n76 8.855
R117 w_n84_832.n76 w_n84_832.n75 8.855
R118 w_n84_832.n81 w_n84_832.n80 8.855
R119 w_n84_832.n80 w_n84_832.n79 8.855
R120 w_n84_832.n130 w_n84_832.n1 8.855
R121 w_n84_832.n1 w_n84_832.n0 8.855
R122 w_n84_832.n133 w_n84_832.n132 8.855
R123 w_n84_832.n132 w_n84_832.n131 8.855
R124 w_n84_832.n126 w_n84_832.n125 8.855
R125 w_n84_832.n125 w_n84_832.n124 8.855
R126 w_n84_832.n122 w_n84_832.n121 8.855
R127 w_n84_832.n121 w_n84_832.n120 8.855
R128 w_n84_832.n116 w_n84_832.n115 8.855
R129 w_n84_832.n115 w_n84_832.n114 8.855
R130 w_n84_832.n112 w_n84_832.n111 8.855
R131 w_n84_832.n111 w_n84_832.n110 8.855
R132 w_n84_832.n107 w_n84_832.n106 8.855
R133 w_n84_832.n106 w_n84_832.n105 8.855
R134 w_n84_832.n104 w_n84_832.n103 8.855
R135 w_n84_832.n103 w_n84_832.n102 8.855
R136 w_n84_832.n134 w_n84_832.n133 8.258
R137 w_n84_832.n56 w_n84_832.n55 8.051
R138 w_n84_832.n124  饝 7.671
R139 w_n84_832.n122 w_n84_832.n119 7.019
R140 w_n84_832.n134 w_n84_832.n130 6.606
R141 w_n84_832.n131 ���i�U 5.114
R142 w_n84_832.n30 w_n84_832.n25 4.795
R143 w_n84_832.n30 w_n84_832.n29 4.65
R144 w_n84_832.n34 w_n84_832.n33 4.65
R145 w_n84_832.n39 w_n84_832.n38 4.65
R146 w_n84_832.n43 w_n84_832.n42 4.65
R147 w_n84_832.n70 w_n84_832.n69 4.65
R148 w_n84_832.n74 w_n84_832.n73 4.65
R149 w_n84_832.n78 w_n84_832.n77 4.65
R150 w_n84_832.n82 w_n84_832.n81 4.65
R151 w_n84_832.n130 w_n84_832.n129 4.65
R152 w_n84_832.n127 w_n84_832.n126 4.65
R153 w_n84_832.n123 w_n84_832.n122 4.65
R154 w_n84_832.n117 w_n84_832.n116 4.65
R155 w_n84_832.n113 w_n84_832.n112 4.65
R156 w_n84_832.n108 w_n84_832.n104 2.932
R157 w_n84_832.n108 w_n84_832.n107 2.844
R158 w_n84_832.n29 w_n84_832.n26 2.064
R159 w_n84_832.n38 w_n84_832.n37 2.064
R160 w_n84_832.n113 w_n84_832.n108 1.063
R161 w_n84_832.n112 w_n84_832.n109 0.412
R162 w_n84_832.n70 w_n84_832.n43 0.29
R163 w_n84_832.n128 w_n84_832.n127 0.197
R164 w_n84_832.n34 w_n84_832.n30 0.157
R165 w_n84_832.n39 w_n84_832.n34 0.157
R166 w_n84_832.n43 w_n84_832.n39 0.145
R167 w_n84_832.n74 w_n84_832.n70 0.145
R168 w_n84_832.n78 w_n84_832.n74 0.145
R169 w_n84_832.n82 w_n84_832.n78 0.145
R170 w_n84_832.n129 w_n84_832.n82 0.145
R171 w_n84_832.n129 w_n84_832.n128 0.145
R172 w_n84_832.n127 w_n84_832.n123 0.145
R173 w_n84_832.n123 w_n84_832.n117 0.145
R174 w_n84_832.n117 w_n84_832.n113 0.145
R175 C.n0 C.t2 454.685
R176 C.n0 C.t0 428.979
R177 C.n1 C.t1 283.824
R178 C.n1 C.n0 199.147
R179 C C.n1 4.65
R180 Y.n5 Y.n4 272.451
R181 Y.n5 Y.n0 271.281
R182 Y.n4 Y.n3 30
R183 Y.n2 Y.n1 24.383
R184 Y.n4 Y.n2 23.684
R185 Y.n0 Y.t1 14.282
R186 Y.n0 Y.t2 14.282
R187 Y Y.n5 4.65
R188 a_372_210.n9 a_372_210.n7 171.558
R189 a_372_210.t0 a_372_210.n9 75.765
R190 a_372_210.n3 a_372_210.n1 74.827
R191 a_372_210.n3 a_372_210.n2 27.476
R192 a_372_210.n7 a_372_210.n6 27.2
R193 a_372_210.n5 a_372_210.n4 23.498
R194 a_372_210.n7 a_372_210.n5 22.4
R195 a_372_210.t0 a_372_210.n11 20.241
R196 a_372_210.t0 a_372_210.n3 13.984
R197 a_372_210.n11 a_372_210.n10 13.494
R198 a_372_210.t0 a_372_210.n0 8.137
R199 a_372_210.n9 a_372_210.n8 1.505
R200 A.n0 A.t2 512.525
R201 A.n1 A.t1 389.251
R202 A.n0 A.t0 371.139
R203 A.n1 A.n0 207.695
R204 A A.n1 4.65
R205 a_91_103.t0 a_91_103.n7 59.616
R206 a_91_103.n4 a_91_103.n2 54.496
R207 a_91_103.n4 a_91_103.n3 54.496
R208 a_91_103.n1 a_91_103.n0 24.679
R209 a_91_103.t0 a_91_103.n1 7.505
R210 a_91_103.n6 a_91_103.n5 2.455
R211 a_91_103.n6 a_91_103.n4 0.636
R212 a_91_103.t0 a_91_103.n6 0.246
C3 C  饝 0.29fF
C4 B  饝 0.29fF
C5 A  饝 0.35fF
C6 a_91_103.n0  饝 0.08fF
C7 a_91_103.n1  饝 0.07fF
C8 a_91_103.n2  饝 0.04fF
C9 a_91_103.n3  饝 0.06fF
C10 a_91_103.n4  饝 0.03fF
C11 a_91_103.n5  饝 0.03fF
C12 a_91_103.n7  饝 0.08fF
C13 A.n0  饝 0.16fF
C14 A.n1  饝 0.25fF
C15 a_372_210.n0  饝 0.06fF
C16 a_372_210.n1  饝 0.09fF
C17 a_372_210.n2  饝 0.12fF
C18 a_372_210.n3  饝 0.08fF
C19 a_372_210.n4  饝 0.02fF
C20 a_372_210.n5  饝 0.03fF
C21 a_372_210.n6  饝 0.02fF
C22 a_372_210.n7  饝 0.03fF
C23 a_372_210.n8  饝 0.02fF
C24 a_372_210.n9  饝 0.13fF
C25 a_372_210.n10  饝 0.08fF
C26 a_372_210.n11  饝 0.02fF
C27 a_372_210.t0  饝 0.31fF
C28 Y.n0  饝 0.64fF
C29 Y.n1  饝 0.04fF
C30 Y.n2  饝 0.05fF
C31 Y.n3  饝 0.03fF
C32 Y.n4  饝 0.19fF
C33 Y.n5  饝 0.62fF
C34 C.n0  饝 0.22fF
C35 C.t1  饝 0.31fF
C36 C.n1  饝 0.25fF
C37 w_n84_832.n0  饝 0.12fF
C38 w_n84_832.n1  饝 0.01fF
C39 w_n84_832.n3  饝 0.02fF
C40 w_n84_832.n4  饝 0.07fF
C41 w_n84_832.n5  饝 0.02fF
C42 w_n84_832.n6  饝 0.02fF
C43 w_n84_832.n7  饝 0.04fF
C44 w_n84_832.n8  饝 0.02fF
C45 w_n84_832.n9  饝 0.02fF
C46 w_n84_832.n10  饝 0.02fF
C47 w_n84_832.n11  饝 0.02fF
C48 w_n84_832.n12  饝 0.02fF
C49 w_n84_832.n13  饝 0.02fF
C50 w_n84_832.n14  饝 0.02fF
C51 w_n84_832.n15  饝 0.02fF
C52 w_n84_832.n16  饝 0.03fF
C53 w_n84_832.n17  饝 0.01fF
C54 w_n84_832.n22  饝 0.34fF
C55 w_n84_832.n23  饝 0.21fF
C56 w_n84_832.n24  饝 0.01fF
C57 w_n84_832.n25  饝 0.02fF
C58 w_n84_832.n26  饝 0.05fF
C59 w_n84_832.n27  饝 0.15fF
C60 w_n84_832.n28  饝 0.01fF
C61 w_n84_832.n29  饝 0.01fF
C62 w_n84_832.n30  饝 0.05fF
C63 w_n84_832.n31  饝 0.13fF
C64 w_n84_832.n32  饝 0.01fF
C65 w_n84_832.n33  饝 0.02fF
C66 w_n84_832.n34  饝 0.02fF
C67 w_n84_832.n35  饝 0.15fF
C68 w_n84_832.n36  饝 0.01fF
C69 w_n84_832.n37  饝 0.05fF
C70 w_n84_832.n38  饝 0.01fF
C71 w_n84_832.n39  饝 0.02fF
C72 w_n84_832.n40  饝 0.21fF
C73 w_n84_832.n41  饝 0.01fF
C74 w_n84_832.n42  饝 0.02fF
C75 w_n84_832.n43  饝 0.03fF
C76 w_n84_832.n44  饝 0.04fF
C77 w_n84_832.n45  饝 0.02fF
C78 w_n84_832.n46  饝 0.02fF
C79 w_n84_832.n47  饝 0.02fF
C80 w_n84_832.n48  饝 0.02fF
C81 w_n84_832.n49  饝 0.02fF
C82 w_n84_832.n50  饝 0.02fF
C83 w_n84_832.n51  饝 0.02fF
C84 w_n84_832.n52  饝 0.02fF
C85 w_n84_832.n53  饝 0.02fF
C86 w_n84_832.n54  饝 0.02fF
C87 w_n84_832.n55  饝 0.01fF
C88 w_n84_832.n56  饝 0.02fF
C89 w_n84_832.n57  饝 0.02fF
C90 w_n84_832.n60  饝 0.02fF
C91 w_n84_832.n62  饝 0.02fF
C92 w_n84_832.n63  饝 0.17fF
C93 w_n84_832.n64  饝 0.01fF
C94 w_n84_832.n66  饝 0.21fF
C95 w_n84_832.n67  饝 0.21fF
C96 w_n84_832.n68  饝 0.01fF
C97 w_n84_832.n69  饝 0.02fF
C98 w_n84_832.n70  饝 0.03fF
C99 w_n84_832.n71  饝 0.21fF
C100 w_n84_832.n72  饝 0.01fF
C101 w_n84_832.n73  饝 0.02fF
C102 w_n84_832.n74  饝 0.02fF
C103 w_n84_832.n75  饝 0.17fF
C104 w_n84_832.n76  饝 0.01fF
C105 w_n84_832.n77  饝 0.05fF
C106 w_n84_832.n78  饝 0.02fF
C107 w_n84_832.n79  饝 0.13fF
C108 w_n84_832.n80  饝 0.01fF
C109 w_n84_832.n81  饝 0.02fF
C110 w_n84_83