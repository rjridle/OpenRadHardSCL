magic
tech sky130A
magscale 1 2
timestamp 1649945920
<< nwell >>
rect -84 832 2304 1575
<< nmos >>
rect 155 324 185 377
tri 185 324 201 340 sw
rect 155 294 261 324
tri 261 294 291 324 sw
rect 155 193 185 294
tri 185 278 201 294 nw
tri 245 278 261 294 ne
tri 185 193 201 209 sw
tri 245 193 261 209 se
rect 261 193 291 294
tri 155 163 185 193 ne
rect 185 163 261 193
tri 261 163 291 193 nw
rect 612 316 642 377
tri 642 316 658 332 sw
rect 806 324 836 377
tri 836 324 852 340 sw
rect 612 286 718 316
tri 718 286 748 316 sw
rect 806 294 912 324
tri 912 294 942 324 sw
rect 612 185 642 286
tri 642 270 658 286 nw
tri 702 270 718 286 ne
tri 642 185 658 201 sw
tri 702 185 718 201 se
rect 718 185 748 286
rect 806 193 836 294
tri 836 278 852 294 nw
tri 896 278 912 294 ne
tri 836 193 852 209 sw
tri 896 193 912 209 se
rect 912 193 942 294
tri 612 155 642 185 ne
rect 642 155 718 185
tri 718 155 748 185 nw
tri 806 163 836 193 ne
rect 836 163 912 193
tri 912 163 942 193 nw
rect 1278 316 1308 377
tri 1308 316 1324 332 sw
rect 1472 324 1502 377
tri 1502 324 1518 340 sw
rect 1278 286 1384 316
tri 1384 286 1414 316 sw
rect 1472 294 1578 324
tri 1578 294 1608 324 sw
rect 1278 185 1308 286
tri 1308 270 1324 286 nw
tri 1368 270 1384 286 ne
tri 1308 185 1324 201 sw
tri 1368 185 1384 201 se
rect 1384 185 1414 286
rect 1472 193 1502 294
tri 1502 278 1518 294 nw
tri 1562 278 1578 294 ne
tri 1502 193 1518 209 sw
tri 1562 193 1578 209 se
rect 1578 193 1608 294
tri 1278 155 1308 185 ne
rect 1308 155 1384 185
tri 1384 155 1414 185 nw
tri 1472 163 1502 193 ne
rect 1502 163 1578 193
tri 1578 163 1608 193 nw
tri 2019 324 2035 340 se
rect 2035 324 2065 377
tri 1929 294 1959 324 se
rect 1959 294 2065 324
rect 1929 193 1959 294
tri 1959 278 1975 294 nw
tri 2019 278 2035 294 ne
tri 1959 193 1975 209 sw
tri 2019 193 2035 209 se
rect 2035 193 2065 294
tri 1929 163 1959 193 ne
rect 1959 163 2035 193
tri 2035 163 2065 193 nw
<< pmos >>
rect 163 1050 193 1450
rect 251 1050 281 1450
rect 631 1051 661 1451
rect 719 1051 749 1451
rect 807 1051 837 1451
rect 895 1051 925 1451
rect 1297 1051 1327 1451
rect 1385 1051 1415 1451
rect 1473 1051 1503 1451
rect 1561 1051 1591 1451
rect 1939 1050 1969 1450
rect 2027 1050 2057 1450
<< ndiff >>
rect 99 361 155 377
rect 99 327 109 361
rect 143 327 155 361
rect 99 289 155 327
rect 185 361 345 377
rect 185 340 303 361
tri 185 324 201 340 ne
rect 201 327 303 340
rect 337 327 345 361
rect 201 324 345 327
tri 261 294 291 324 ne
rect 99 255 109 289
rect 143 255 155 289
rect 99 221 155 255
rect 99 187 109 221
rect 143 187 155 221
tri 185 278 201 294 se
rect 201 278 245 294
tri 245 278 261 294 sw
rect 185 245 261 278
rect 185 211 205 245
rect 239 211 261 245
rect 185 209 261 211
tri 185 193 201 209 ne
rect 201 193 245 209
tri 245 193 261 209 nw
rect 291 289 345 324
rect 291 255 303 289
rect 337 255 345 289
rect 291 221 345 255
rect 99 163 155 187
tri 155 163 185 193 sw
tri 261 163 291 193 se
rect 291 187 303 221
rect 337 187 345 221
rect 291 163 345 187
rect 99 151 345 163
rect 99 117 109 151
rect 143 117 205 151
rect 239 117 303 151
rect 337 117 345 151
rect 99 101 345 117
rect 556 361 612 377
rect 556 327 566 361
rect 600 327 612 361
rect 556 289 612 327
rect 642 361 806 377
rect 642 332 663 361
tri 642 316 658 332 ne
rect 658 327 663 332
rect 697 327 760 361
rect 794 327 806 361
rect 658 316 806 327
rect 836 340 998 377
tri 836 324 852 340 ne
rect 852 324 998 340
rect 556 255 566 289
rect 600 255 612 289
tri 718 286 748 316 ne
rect 748 289 806 316
tri 912 294 942 324 ne
rect 556 221 612 255
rect 556 187 566 221
rect 600 187 612 221
rect 556 155 612 187
tri 642 270 658 286 se
rect 658 270 702 286
tri 702 270 718 286 sw
rect 642 236 718 270
rect 642 202 663 236
rect 697 202 718 236
rect 642 201 718 202
tri 642 185 658 201 ne
rect 658 185 702 201
tri 702 185 718 201 nw
rect 748 255 760 289
rect 794 255 806 289
rect 748 221 806 255
rect 748 187 760 221
rect 794 187 806 221
tri 836 278 852 294 se
rect 852 278 896 294
tri 896 278 912 294 sw
rect 836 245 912 278
rect 836 211 857 245
rect 891 211 912 245
rect 836 209 912 211
tri 836 193 852 209 ne
rect 852 193 896 209
tri 896 193 912 209 nw
rect 942 289 998 324
rect 942 255 954 289
rect 988 255 998 289
rect 942 221 998 255
tri 612 155 642 185 sw
tri 718 155 748 185 se
rect 748 163 806 187
tri 806 163 836 193 sw
tri 912 163 942 193 se
rect 942 187 954 221
rect 988 187 998 221
rect 942 163 998 187
rect 748 155 998 163
rect 556 151 998 155
rect 556 117 566 151
rect 600 117 760 151
rect 794 117 857 151
rect 891 117 954 151
rect 988 117 998 151
rect 556 101 998 117
rect 1222 361 1278 377
rect 1222 327 1232 361
rect 1266 327 1278 361
rect 1222 289 1278 327
rect 1308 361 1472 377
rect 1308 332 1329 361
tri 1308 316 1324 332 ne
rect 1324 327 1329 332
rect 1363 327 1426 361
rect 1460 327 1472 361
rect 1324 316 1472 327
rect 1502 340 1664 377
tri 1502 324 1518 340 ne
rect 1518 324 1664 340
rect 1222 255 1232 289
rect 1266 255 1278 289
tri 1384 286 1414 316 ne
rect 1414 289 1472 316
tri 1578 294 1608 324 ne
rect 1222 221 1278 255
rect 1222 187 1232 221
rect 1266 187 1278 221
rect 1222 155 1278 187
tri 1308 270 1324 286 se
rect 1324 270 1368 286
tri 1368 270 1384 286 sw
rect 1308 236 1384 270
rect 1308 202 1329 236
rect 1363 202 1384 236
rect 1308 201 1384 202
tri 1308 185 1324 201 ne
rect 1324 185 1368 201
tri 1368 185 1384 201 nw
rect 1414 255 1426 289
rect 1460 255 1472 289
rect 1414 221 1472 255
rect 1414 187 1426 221
rect 1460 187 1472 221
tri 1502 278 1518 294 se
rect 1518 278 1562 294
tri 1562 278 1578 294 sw
rect 1502 245 1578 278
rect 1502 211 1523 245
rect 1557 211 1578 245
rect 1502 209 1578 211
tri 1502 193 1518 209 ne
rect 1518 193 1562 209
tri 1562 193 1578 209 nw
rect 1608 289 1664 324
rect 1608 255 1620 289
rect 1654 255 1664 289
rect 1608 221 1664 255
tri 1278 155 1308 185 sw
tri 1384 155 1414 185 se
rect 1414 163 1472 187
tri 1472 163 1502 193 sw
tri 1578 163 1608 193 se
rect 1608 187 1620 221
rect 1654 187 1664 221
rect 1608 163 1664 187
rect 1414 155 1664 163
rect 1222 151 1664 155
rect 1222 117 1232 151
rect 1266 117 1426 151
rect 1460 117 1523 151
rect 1557 117 1620 151
rect 1654 117 1664 151
rect 1222 101 1664 117
rect 1875 361 2035 377
rect 1875 327 1883 361
rect 1917 340 2035 361
rect 1917 327 2019 340
rect 1875 324 2019 327
tri 2019 324 2035 340 nw
rect 2065 361 2121 377
rect 2065 327 2077 361
rect 2111 327 2121 361
rect 1875 289 1929 324
tri 1929 294 1959 324 nw
rect 1875 255 1883 289
rect 1917 255 1929 289
rect 1875 221 1929 255
rect 1875 187 1883 221
rect 1917 187 1929 221
tri 1959 278 1975 294 se
rect 1975 278 2019 294
tri 2019 278 2035 294 sw
rect 1959 245 2035 278
rect 1959 211 1981 245
rect 2015 211 2035 245
rect 1959 209 2035 211
tri 1959 193 1975 209 ne
rect 1975 193 2019 209
tri 2019 193 2035 209 nw
rect 2065 289 2121 327
rect 2065 255 2077 289
rect 2111 255 2121 289
rect 2065 221 2121 255
rect 1875 163 1929 187
tri 1929 163 1959 193 sw
tri 2035 163 2065 193 se
rect 2065 187 2077 221
rect 2111 187 2121 221
rect 2065 163 2121 187
rect 1875 151 2121 163
rect 1875 117 1883 151
rect 1917 117 1981 151
rect 2015 117 2077 151
rect 2111 117 2121 151
rect 1875 101 2121 117
<< pdiff >>
rect 107 1412 163 1450
rect 107 1378 117 1412
rect 151 1378 163 1412
rect 107 1344 163 1378
rect 107 1310 117 1344
rect 151 1310 163 1344
rect 107 1276 163 1310
rect 107 1242 117 1276
rect 151 1242 163 1276
rect 107 1208 163 1242
rect 107 1174 117 1208
rect 151 1174 163 1208
rect 107 1139 163 1174
rect 107 1105 117 1139
rect 151 1105 163 1139
rect 107 1050 163 1105
rect 193 1412 251 1450
rect 193 1378 205 1412
rect 239 1378 251 1412
rect 193 1344 251 1378
rect 193 1310 205 1344
rect 239 1310 251 1344
rect 193 1276 251 1310
rect 193 1242 205 1276
rect 239 1242 251 1276
rect 193 1208 251 1242
rect 193 1174 205 1208
rect 239 1174 251 1208
rect 193 1139 251 1174
rect 193 1105 205 1139
rect 239 1105 251 1139
rect 193 1050 251 1105
rect 281 1412 335 1450
rect 281 1378 293 1412
rect 327 1378 335 1412
rect 281 1344 335 1378
rect 281 1310 293 1344
rect 327 1310 335 1344
rect 281 1276 335 1310
rect 281 1242 293 1276
rect 327 1242 335 1276
rect 281 1208 335 1242
rect 281 1174 293 1208
rect 327 1174 335 1208
rect 281 1139 335 1174
rect 281 1105 293 1139
rect 327 1105 335 1139
rect 281 1050 335 1105
rect 575 1411 631 1451
rect 575 1377 585 1411
rect 619 1377 631 1411
rect 575 1343 631 1377
rect 575 1309 585 1343
rect 619 1309 631 1343
rect 575 1275 631 1309
rect 575 1241 585 1275
rect 619 1241 631 1275
rect 575 1207 631 1241
rect 575 1173 585 1207
rect 619 1173 631 1207
rect 575 1139 631 1173
rect 575 1105 585 1139
rect 619 1105 631 1139
rect 575 1051 631 1105
rect 661 1343 719 1451
rect 661 1309 673 1343
rect 707 1309 719 1343
rect 661 1275 719 1309
rect 661 1241 673 1275
rect 707 1241 719 1275
rect 661 1207 719 1241
rect 661 1173 673 1207
rect 707 1173 719 1207
rect 661 1051 719 1173
rect 749 1411 807 1451
rect 749 1377 761 1411
rect 795 1377 807 1411
rect 749 1343 807 1377
rect 749 1309 761 1343
rect 795 1309 807 1343
rect 749 1275 807 1309
rect 749 1241 761 1275
rect 795 1241 807 1275
rect 749 1207 807 1241
rect 749 1173 761 1207
rect 795 1173 807 1207
rect 749 1139 807 1173
rect 749 1105 761 1139
rect 795 1105 807 1139
rect 749 1051 807 1105
rect 837 1343 895 1451
rect 837 1309 849 1343
rect 883 1309 895 1343
rect 837 1275 895 1309
rect 837 1241 849 1275
rect 883 1241 895 1275
rect 837 1207 895 1241
rect 837 1173 849 1207
rect 883 1173 895 1207
rect 837 1139 895 1173
rect 837 1105 849 1139
rect 883 1105 895 1139
rect 837 1051 895 1105
rect 925 1411 979 1451
rect 925 1377 937 1411
rect 971 1377 979 1411
rect 925 1343 979 1377
rect 925 1309 937 1343
rect 971 1309 979 1343
rect 925 1275 979 1309
rect 925 1241 937 1275
rect 971 1241 979 1275
rect 925 1207 979 1241
rect 925 1173 937 1207
rect 971 1173 979 1207
rect 925 1051 979 1173
rect 1241 1411 1297 1451
rect 1241 1377 1251 1411
rect 1285 1377 1297 1411
rect 1241 1343 1297 1377
rect 1241 1309 1251 1343
rect 1285 1309 1297 1343
rect 1241 1275 1297 1309
rect 1241 1241 1251 1275
rect 1285 1241 1297 1275
rect 1241 1207 1297 1241
rect 1241 1173 1251 1207
rect 1285 1173 1297 1207
rect 1241 1139 1297 1173
rect 1241 1105 1251 1139
rect 1285 1105 1297 1139
rect 1241 1051 1297 1105
rect 1327 1343 1385 1451
rect 1327 1309 1339 1343
rect 1373 1309 1385 1343
rect 1327 1275 1385 1309
rect 1327 1241 1339 1275
rect 1373 1241 1385 1275
rect 1327 1207 1385 1241
rect 1327 1173 1339 1207
rect 1373 1173 1385 1207
rect 1327 1051 1385 1173
rect 1415 1411 1473 1451
rect 1415 1377 1427 1411
rect 1461 1377 1473 1411
rect 1415 1343 1473 1377
rect 1415 1309 1427 1343
rect 1461 1309 1473 1343
rect 1415 1275 1473 1309
rect 1415 1241 1427 1275
rect 1461 1241 1473 1275
rect 1415 1207 1473 1241
rect 1415 1173 1427 1207
rect 1461 1173 1473 1207
rect 1415 1139 1473 1173
rect 1415 1105 1427 1139
rect 1461 1105 1473 1139
rect 1415 1051 1473 1105
rect 1503 1343 1561 1451
rect 1503 1309 1515 1343
rect 1549 1309 1561 1343
rect 1503 1275 1561 1309
rect 1503 1241 1515 1275
rect 1549 1241 1561 1275
rect 1503 1207 1561 1241
rect 1503 1173 1515 1207
rect 1549 1173 1561 1207
rect 1503 1139 1561 1173
rect 1503 1105 1515 1139
rect 1549 1105 1561 1139
rect 1503 1051 1561 1105
rect 1591 1411 1645 1451
rect 1591 1377 1603 1411
rect 1637 1377 1645 1411
rect 1591 1343 1645 1377
rect 1591 1309 1603 1343
rect 1637 1309 1645 1343
rect 1591 1275 1645 1309
rect 1591 1241 1603 1275
rect 1637 1241 1645 1275
rect 1591 1207 1645 1241
rect 1591 1173 1603 1207
rect 1637 1173 1645 1207
rect 1591 1051 1645 1173
rect 1885 1412 1939 1450
rect 1885 1378 1893 1412
rect 1927 1378 1939 1412
rect 1885 1344 1939 1378
rect 1885 1310 1893 1344
rect 1927 1310 1939 1344
rect 1885 1276 1939 1310
rect 1885 1242 1893 1276
rect 1927 1242 1939 1276
rect 1885 1208 1939 1242
rect 1885 1174 1893 1208
rect 1927 1174 1939 1208
rect 1885 1139 1939 1174
rect 1885 1105 1893 1139
rect 1927 1105 1939 1139
rect 1885 1050 1939 1105
rect 1969 1412 2027 1450
rect 1969 1378 1981 1412
rect 2015 1378 2027 1412
rect 1969 1344 2027 1378
rect 1969 1310 1981 1344
rect 2015 1310 2027 1344
rect 1969 1276 2027 1310
rect 1969 1242 1981 1276
rect 2015 1242 2027 1276
rect 1969 1208 2027 1242
rect 1969 1174 1981 1208
rect 2015 1174 2027 1208
rect 1969 1139 2027 1174
rect 1969 1105 1981 1139
rect 2015 1105 2027 1139
rect 1969 1050 2027 1105
rect 2057 1412 2113 1450
rect 2057 1378 2069 1412
rect 2103 1378 2113 1412
rect 2057 1344 2113 1378
rect 2057 1310 2069 1344
rect 2103 1310 2113 1344
rect 2057 1276 2113 1310
rect 2057 1242 2069 1276
rect 2103 1242 2113 1276
rect 2057 1208 2113 1242
rect 2057 1174 2069 1208
rect 2103 1174 2113 1208
rect 2057 1139 2113 1174
rect 2057 1105 2069 1139
rect 2103 1105 2113 1139
rect 2057 1050 2113 1105
<< ndiffc >>
rect 109 327 143 361
rect 303 327 337 361
rect 109 255 143 289
rect 109 187 143 221
rect 205 211 239 245
rect 303 255 337 289
rect 303 187 337 221
rect 109 117 143 151
rect 205 117 239 151
rect 303 117 337 151
rect 566 327 600 361
rect 663 327 697 361
rect 760 327 794 361
rect 566 255 600 289
rect 566 187 600 221
rect 663 202 697 236
rect 760 255 794 289
rect 760 187 794 221
rect 857 211 891 245
rect 954 255 988 289
rect 954 187 988 221
rect 566 117 600 151
rect 760 117 794 151
rect 857 117 891 151
rect 954 117 988 151
rect 1232 327 1266 361
rect 1329 327 1363 361
rect 1426 327 1460 361
rect 1232 255 1266 289
rect 1232 187 1266 221
rect 1329 202 1363 236
rect 1426 255 1460 289
rect 1426 187 1460 221
rect 1523 211 1557 245
rect 1620 255 1654 289
rect 1620 187 1654 221
rect 1232 117 1266 151
rect 1426 117 1460 151
rect 1523 117 1557 151
rect 1620 117 1654 151
rect 1883 327 1917 361
rect 2077 327 2111 361
rect 1883 255 1917 289
rect 1883 187 1917 221
rect 1981 211 2015 245
rect 2077 255 2111 289
rect 2077 187 2111 221
rect 1883 117 1917 151
rect 1981 117 2015 151
rect 2077 117 2111 151
<< pdiffc >>
rect 117 1378 151 1412
rect 117 1310 151 1344
rect 117 1242 151 1276
rect 117 1174 151 1208
rect 117 1105 151 1139
rect 205 1378 239 1412
rect 205 1310 239 1344
rect 205 1242 239 1276
rect 205 1174 239 1208
rect 205 1105 239 1139
rect 293 1378 327 1412
rect 293 1310 327 1344
rect 293 1242 327 1276
rect 293 1174 327 1208
rect 293 1105 327 1139
rect 585 1377 619 1411
rect 585 1309 619 1343
rect 585 1241 619 1275
rect 585 1173 619 1207
rect 585 1105 619 1139
rect 673 1309 707 1343
rect 673 1241 707 1275
rect 673 1173 707 1207
rect 761 1377 795 1411
rect 761 1309 795 1343
rect 761 1241 795 1275
rect 761 1173 795 1207
rect 761 1105 795 1139
rect 849 1309 883 1343
rect 849 1241 883 1275
rect 849 1173 883 1207
rect 849 1105 883 1139
rect 937 1377 971 1411
rect 937 1309 971 1343
rect 937 1241 971 1275
rect 937 1173 971 1207
rect 1251 1377 1285 1411
rect 1251 1309 1285 1343
rect 1251 1241 1285 1275
rect 1251 1173 1285 1207
rect 1251 1105 1285 1139
rect 1339 1309 1373 1343
rect 1339 1241 1373 1275
rect 1339 1173 1373 1207
rect 1427 1377 1461 1411
rect 1427 1309 1461 1343
rect 1427 1241 1461 1275
rect 1427 1173 1461 1207
rect 1427 1105 1461 1139
rect 1515 1309 1549 1343
rect 1515 1241 1549 1275
rect 1515 1173 1549 1207
rect 1515 1105 1549 1139
rect 1603 1377 1637 1411
rect 1603 1309 1637 1343
rect 1603 1241 1637 1275
rect 1603 1173 1637 1207
rect 1893 1378 1927 1412
rect 1893 1310 1927 1344
rect 1893 1242 1927 1276
rect 1893 1174 1927 1208
rect 1893 1105 1927 1139
rect 1981 1378 2015 1412
rect 1981 1310 2015 1344
rect 1981 1242 2015 1276
rect 1981 1174 2015 1208
rect 1981 1105 2015 1139
rect 2069 1378 2103 1412
rect 2069 1310 2103 1344
rect 2069 1242 2103 1276
rect 2069 1174 2103 1208
rect 2069 1105 2103 1139
<< psubdiff >>
rect -31 546 2251 572
rect -31 512 -17 546
rect 17 512 427 546
rect 461 512 1093 546
rect 1127 512 1759 546
rect 1793 512 2203 546
rect 2237 512 2251 546
rect -31 510 2251 512
rect -31 474 31 510
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect 413 474 475 510
rect -31 368 -17 402
rect 17 368 31 402
rect 413 440 427 474
rect 461 440 475 474
rect 413 402 475 440
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect 413 368 427 402
rect 461 368 475 402
rect 1079 474 1141 510
rect 1079 440 1093 474
rect 1127 440 1141 474
rect 1079 402 1141 440
rect 413 330 475 368
rect 413 296 427 330
rect 461 296 475 330
rect 413 258 475 296
rect 413 224 427 258
rect 461 224 475 258
rect 413 186 475 224
rect 413 152 427 186
rect 461 152 475 186
rect 413 114 475 152
rect -31 47 31 80
rect 413 80 427 114
rect 461 80 475 114
rect 1079 368 1093 402
rect 1127 368 1141 402
rect 1745 474 1807 510
rect 1745 440 1759 474
rect 1793 440 1807 474
rect 1745 402 1807 440
rect 1079 330 1141 368
rect 1079 296 1093 330
rect 1127 296 1141 330
rect 1079 258 1141 296
rect 1079 224 1093 258
rect 1127 224 1141 258
rect 1079 186 1141 224
rect 1079 152 1093 186
rect 1127 152 1141 186
rect 1079 114 1141 152
rect 413 47 475 80
rect 1079 80 1093 114
rect 1127 80 1141 114
rect 1745 368 1759 402
rect 1793 368 1807 402
rect 2189 474 2251 510
rect 2189 440 2203 474
rect 2237 440 2251 474
rect 2189 402 2251 440
rect 1745 330 1807 368
rect 1745 296 1759 330
rect 1793 296 1807 330
rect 1745 258 1807 296
rect 1745 224 1759 258
rect 1793 224 1807 258
rect 1745 186 1807 224
rect 1745 152 1759 186
rect 1793 152 1807 186
rect 1745 114 1807 152
rect 1079 47 1141 80
rect 1745 80 1759 114
rect 1793 80 1807 114
rect 2189 368 2203 402
rect 2237 368 2251 402
rect 2189 330 2251 368
rect 2189 296 2203 330
rect 2237 296 2251 330
rect 2189 258 2251 296
rect 2189 224 2203 258
rect 2237 224 2251 258
rect 2189 186 2251 224
rect 2189 152 2203 186
rect 2237 152 2251 186
rect 2189 114 2251 152
rect 1745 47 1807 80
rect 2189 80 2203 114
rect 2237 80 2251 114
rect 2189 47 2251 80
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 205 47
rect 239 13 283 47
rect 317 13 355 47
rect 389 13 499 47
rect 533 13 571 47
rect 605 13 643 47
rect 677 13 715 47
rect 749 13 805 47
rect 839 13 877 47
rect 911 13 949 47
rect 983 13 1021 47
rect 1055 13 1165 47
rect 1199 13 1237 47
rect 1271 13 1309 47
rect 1343 13 1381 47
rect 1415 13 1471 47
rect 1505 13 1543 47
rect 1577 13 1615 47
rect 1649 13 1687 47
rect 1721 13 1831 47
rect 1865 13 1903 47
rect 1937 13 1981 47
rect 2015 13 2059 47
rect 2093 13 2131 47
rect 2165 13 2251 47
rect -31 11 31 13
rect 413 11 475 13
rect 1079 11 1141 13
rect 1745 11 1807 13
rect 2189 11 2251 13
<< nsubdiff >>
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 205 1539
rect 239 1505 283 1539
rect 317 1505 355 1539
rect 389 1505 499 1539
rect 533 1505 571 1539
rect 605 1505 643 1539
rect 677 1505 715 1539
rect 749 1505 805 1539
rect 839 1505 877 1539
rect 911 1505 949 1539
rect 983 1505 1021 1539
rect 1055 1505 1165 1539
rect 1199 1505 1237 1539
rect 1271 1505 1309 1539
rect 1343 1505 1381 1539
rect 1415 1505 1471 1539
rect 1505 1505 1543 1539
rect 1577 1505 1615 1539
rect 1649 1505 1687 1539
rect 1721 1505 1831 1539
rect 1865 1505 1903 1539
rect 1937 1505 1981 1539
rect 2015 1505 2059 1539
rect 2093 1505 2131 1539
rect 2165 1505 2251 1539
rect -31 1470 31 1505
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect 413 1470 475 1505
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect -31 1038 31 1076
rect 413 1436 427 1470
rect 461 1436 475 1470
rect 1079 1470 1141 1505
rect 413 1398 475 1436
rect 413 1364 427 1398
rect 461 1364 475 1398
rect 413 1326 475 1364
rect 413 1292 427 1326
rect 461 1292 475 1326
rect 413 1254 475 1292
rect 413 1220 427 1254
rect 461 1220 475 1254
rect 413 1182 475 1220
rect 413 1148 427 1182
rect 461 1148 475 1182
rect 413 1110 475 1148
rect 413 1076 427 1110
rect 461 1076 475 1110
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect 413 1038 475 1076
rect 1079 1436 1093 1470
rect 1127 1436 1141 1470
rect 1745 1470 1807 1505
rect 1079 1398 1141 1436
rect 1079 1364 1093 1398
rect 1127 1364 1141 1398
rect 1079 1326 1141 1364
rect 1079 1292 1093 1326
rect 1127 1292 1141 1326
rect 1079 1254 1141 1292
rect 1079 1220 1093 1254
rect 1127 1220 1141 1254
rect 1079 1182 1141 1220
rect 1079 1148 1093 1182
rect 1127 1148 1141 1182
rect 1079 1110 1141 1148
rect 1079 1076 1093 1110
rect 1127 1076 1141 1110
rect 413 1004 427 1038
rect 461 1004 475 1038
rect 413 966 475 1004
rect -31 930 31 932
rect 413 932 427 966
rect 461 932 475 966
rect 1079 1038 1141 1076
rect 1745 1436 1759 1470
rect 1793 1436 1807 1470
rect 2189 1470 2251 1505
rect 1745 1398 1807 1436
rect 1745 1364 1759 1398
rect 1793 1364 1807 1398
rect 1745 1326 1807 1364
rect 1745 1292 1759 1326
rect 1793 1292 1807 1326
rect 1745 1254 1807 1292
rect 1745 1220 1759 1254
rect 1793 1220 1807 1254
rect 1745 1182 1807 1220
rect 1745 1148 1759 1182
rect 1793 1148 1807 1182
rect 1745 1110 1807 1148
rect 1745 1076 1759 1110
rect 1793 1076 1807 1110
rect 1079 1004 1093 1038
rect 1127 1004 1141 1038
rect 1079 966 1141 1004
rect 413 930 475 932
rect 1079 932 1093 966
rect 1127 932 1141 966
rect 1745 1038 1807 1076
rect 2189 1436 2203 1470
rect 2237 1436 2251 1470
rect 2189 1398 2251 1436
rect 2189 1364 2203 1398
rect 2237 1364 2251 1398
rect 2189 1326 2251 1364
rect 2189 1292 2203 1326
rect 2237 1292 2251 1326
rect 2189 1254 2251 1292
rect 2189 1220 2203 1254
rect 2237 1220 2251 1254
rect 2189 1182 2251 1220
rect 2189 1148 2203 1182
rect 2237 1148 2251 1182
rect 2189 1110 2251 1148
rect 2189 1076 2203 1110
rect 2237 1076 2251 1110
rect 1745 1004 1759 1038
rect 1793 1004 1807 1038
rect 1745 966 1807 1004
rect 2189 1038 2251 1076
rect 1079 930 1141 932
rect 1745 932 1759 966
rect 1793 932 1807 966
rect 2189 1004 2203 1038
rect 2237 1004 2251 1038
rect 2189 966 2251 1004
rect 1745 930 1807 932
rect 2189 932 2203 966
rect 2237 932 2251 966
rect 2189 930 2251 932
rect -31 868 2251 930
<< psubdiffcont >>
rect -17 512 17 546
rect 427 512 461 546
rect 1093 512 1127 546
rect 1759 512 1793 546
rect 2203 512 2237 546
rect -17 440 17 474
rect -17 368 17 402
rect 427 440 461 474
rect -17 296 17 330
rect -17 224 17 258
rect -17 152 17 186
rect -17 80 17 114
rect 427 368 461 402
rect 1093 440 1127 474
rect 427 296 461 330
rect 427 224 461 258
rect 427 152 461 186
rect 427 80 461 114
rect 1093 368 1127 402
rect 1759 440 1793 474
rect 1093 296 1127 330
rect 1093 224 1127 258
rect 1093 152 1127 186
rect 1093 80 1127 114
rect 1759 368 1793 402
rect 2203 440 2237 474
rect 1759 296 1793 330
rect 1759 224 1793 258
rect 1759 152 1793 186
rect 1759 80 1793 114
rect 2203 368 2237 402
rect 2203 296 2237 330
rect 2203 224 2237 258
rect 2203 152 2237 186
rect 2203 80 2237 114
rect 55 13 89 47
rect 127 13 161 47
rect 205 13 239 47
rect 283 13 317 47
rect 355 13 389 47
rect 499 13 533 47
rect 571 13 605 47
rect 643 13 677 47
rect 715 13 749 47
rect 805 13 839 47
rect 877 13 911 47
rect 949 13 983 47
rect 1021 13 1055 47
rect 1165 13 1199 47
rect 1237 13 1271 47
rect 1309 13 1343 47
rect 1381 13 1415 47
rect 1471 13 1505 47
rect 1543 13 1577 47
rect 1615 13 1649 47
rect 1687 13 1721 47
rect 1831 13 1865 47
rect 1903 13 1937 47
rect 1981 13 2015 47
rect 2059 13 2093 47
rect 2131 13 2165 47
<< nsubdiffcont >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 205 1505 239 1539
rect 283 1505 317 1539
rect 355 1505 389 1539
rect 499 1505 533 1539
rect 571 1505 605 1539
rect 643 1505 677 1539
rect 715 1505 749 1539
rect 805 1505 839 1539
rect 877 1505 911 1539
rect 949 1505 983 1539
rect 1021 1505 1055 1539
rect 1165 1505 1199 1539
rect 1237 1505 1271 1539
rect 1309 1505 1343 1539
rect 1381 1505 1415 1539
rect 1471 1505 1505 1539
rect 1543 1505 1577 1539
rect 1615 1505 1649 1539
rect 1687 1505 1721 1539
rect 1831 1505 1865 1539
rect 1903 1505 1937 1539
rect 1981 1505 2015 1539
rect 2059 1505 2093 1539
rect 2131 1505 2165 1539
rect -17 1436 17 1470
rect -17 1364 17 1398
rect -17 1292 17 1326
rect -17 1220 17 1254
rect -17 1148 17 1182
rect -17 1076 17 1110
rect 427 1436 461 1470
rect 427 1364 461 1398
rect 427 1292 461 1326
rect 427 1220 461 1254
rect 427 1148 461 1182
rect 427 1076 461 1110
rect -17 1004 17 1038
rect -17 932 17 966
rect 1093 1436 1127 1470
rect 1093 1364 1127 1398
rect 1093 1292 1127 1326
rect 1093 1220 1127 1254
rect 1093 1148 1127 1182
rect 1093 1076 1127 1110
rect 427 1004 461 1038
rect 427 932 461 966
rect 1759 1436 1793 1470
rect 1759 1364 1793 1398
rect 1759 1292 1793 1326
rect 1759 1220 1793 1254
rect 1759 1148 1793 1182
rect 1759 1076 1793 1110
rect 1093 1004 1127 1038
rect 1093 932 1127 966
rect 2203 1436 2237 1470
rect 2203 1364 2237 1398
rect 2203 1292 2237 1326
rect 2203 1220 2237 1254
rect 2203 1148 2237 1182
rect 2203 1076 2237 1110
rect 1759 1004 1793 1038
rect 1759 932 1793 966
rect 2203 1004 2237 1038
rect 2203 932 2237 966
<< poly >>
rect 163 1450 193 1476
rect 251 1450 281 1476
rect 631 1451 661 1477
rect 719 1451 749 1477
rect 807 1451 837 1477
rect 895 1451 925 1477
rect 163 1019 193 1050
rect 251 1019 281 1050
rect 121 1003 281 1019
rect 121 969 131 1003
rect 165 989 281 1003
rect 1297 1451 1327 1477
rect 1385 1451 1415 1477
rect 1473 1451 1503 1477
rect 1561 1451 1591 1477
rect 165 969 175 989
rect 121 953 175 969
rect 631 1020 661 1051
rect 719 1020 749 1051
rect 631 1004 749 1020
rect 631 990 649 1004
rect 639 970 649 990
rect 683 990 749 1004
rect 807 1020 837 1051
rect 895 1020 925 1051
rect 807 1004 925 1020
rect 807 990 871 1004
rect 683 970 693 990
rect 639 954 693 970
rect 861 970 871 990
rect 905 990 925 1004
rect 1939 1450 1969 1476
rect 2027 1450 2057 1476
rect 905 970 915 990
rect 861 954 915 970
rect 1297 1020 1327 1051
rect 1385 1020 1415 1051
rect 1297 1004 1415 1020
rect 1297 990 1315 1004
rect 1305 970 1315 990
rect 1349 990 1415 1004
rect 1473 1020 1503 1051
rect 1561 1020 1591 1051
rect 1473 1004 1591 1020
rect 1473 990 1537 1004
rect 1349 970 1359 990
rect 1305 954 1359 970
rect 1527 970 1537 990
rect 1571 990 1591 1004
rect 1571 970 1581 990
rect 1527 954 1581 970
rect 1939 1019 1969 1050
rect 2027 1019 2057 1050
rect 1939 1003 2099 1019
rect 1939 989 2055 1003
rect 2045 969 2055 989
rect 2089 969 2099 1003
rect 2045 953 2099 969
rect 121 461 175 477
rect 121 427 131 461
rect 165 441 175 461
rect 165 427 185 441
rect 121 411 185 427
rect 155 377 185 411
rect 639 461 693 477
rect 639 441 649 461
rect 612 427 649 441
rect 683 427 693 461
rect 861 461 915 477
rect 861 441 871 461
rect 612 411 693 427
rect 806 427 871 441
rect 905 427 915 461
rect 806 411 915 427
rect 1305 461 1359 477
rect 1305 441 1315 461
rect 612 377 642 411
rect 806 377 836 411
rect 1278 427 1315 441
rect 1349 427 1359 461
rect 1527 461 1581 477
rect 1527 441 1537 461
rect 1278 411 1359 427
rect 1472 427 1537 441
rect 1571 427 1581 461
rect 1472 411 1581 427
rect 2045 461 2099 477
rect 2045 441 2055 461
rect 1278 377 1308 411
rect 1472 377 1502 411
rect 2035 427 2055 441
rect 2089 427 2099 461
rect 2035 411 2099 427
rect 2035 377 2065 411
<< polycont >>
rect 131 969 165 1003
rect 649 970 683 1004
rect 871 970 905 1004
rect 1315 970 1349 1004
rect 1537 970 1571 1004
rect 2055 969 2089 1003
rect 131 427 165 461
rect 649 427 683 461
rect 871 427 905 461
rect 1315 427 1349 461
rect 1537 427 1571 461
rect 2055 427 2089 461
<< locali >>
rect -31 1539 2251 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 205 1539
rect 239 1505 283 1539
rect 317 1505 355 1539
rect 389 1505 499 1539
rect 533 1505 571 1539
rect 605 1505 643 1539
rect 677 1505 715 1539
rect 749 1505 805 1539
rect 839 1505 877 1539
rect 911 1505 949 1539
rect 983 1505 1021 1539
rect 1055 1505 1165 1539
rect 1199 1505 1237 1539
rect 1271 1505 1309 1539
rect 1343 1505 1381 1539
rect 1415 1505 1471 1539
rect 1505 1505 1543 1539
rect 1577 1505 1615 1539
rect 1649 1505 1687 1539
rect 1721 1505 1831 1539
rect 1865 1505 1903 1539
rect 1937 1505 1981 1539
rect 2015 1505 2059 1539
rect 2093 1505 2131 1539
rect 2165 1505 2251 1539
rect -31 1492 2251 1505
rect -31 1470 31 1492
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect 117 1412 151 1492
rect 117 1344 151 1378
rect 117 1276 151 1310
rect 117 1208 151 1242
rect 117 1139 151 1174
rect 117 1083 151 1105
rect 205 1412 239 1450
rect 205 1344 239 1378
rect 205 1276 239 1310
rect 205 1208 239 1242
rect 205 1139 239 1174
rect -31 1038 31 1076
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect -31 868 31 932
rect 131 1003 165 1019
rect 131 905 165 969
rect 205 979 239 1105
rect 293 1412 327 1492
rect 293 1344 327 1378
rect 293 1276 327 1310
rect 293 1208 327 1242
rect 293 1139 327 1174
rect 293 1083 327 1105
rect 413 1470 475 1492
rect 413 1436 427 1470
rect 461 1436 475 1470
rect 413 1398 475 1436
rect 413 1364 427 1398
rect 461 1364 475 1398
rect 413 1326 475 1364
rect 413 1292 427 1326
rect 461 1292 475 1326
rect 413 1254 475 1292
rect 413 1220 427 1254
rect 461 1220 475 1254
rect 413 1182 475 1220
rect 413 1148 427 1182
rect 461 1148 475 1182
rect 413 1110 475 1148
rect 413 1076 427 1110
rect 461 1076 475 1110
rect 413 1038 475 1076
rect 585 1411 619 1427
rect 585 1343 619 1377
rect 585 1275 619 1309
rect 585 1207 619 1241
rect 585 1139 619 1173
rect 673 1343 707 1492
rect 1079 1470 1141 1492
rect 673 1275 707 1309
rect 673 1207 707 1241
rect 673 1157 707 1173
rect 761 1411 971 1445
rect 761 1343 795 1377
rect 761 1275 795 1309
rect 761 1207 795 1241
rect 761 1139 795 1173
rect 585 1071 795 1105
rect 849 1343 883 1359
rect 849 1275 883 1309
rect 849 1207 883 1241
rect 849 1139 883 1173
rect 937 1343 971 1377
rect 937 1275 971 1309
rect 937 1207 971 1241
rect 937 1157 971 1173
rect 1079 1436 1093 1470
rect 1127 1436 1141 1470
rect 1079 1398 1141 1436
rect 1079 1364 1093 1398
rect 1127 1364 1141 1398
rect 1079 1326 1141 1364
rect 1079 1292 1093 1326
rect 1127 1292 1141 1326
rect 1079 1254 1141 1292
rect 1079 1220 1093 1254
rect 1127 1220 1141 1254
rect 1079 1182 1141 1220
rect 1079 1148 1093 1182
rect 1127 1148 1141 1182
rect 1079 1110 1141 1148
rect 849 1071 979 1105
rect 413 1004 427 1038
rect 461 1004 475 1038
rect 205 945 313 979
rect -31 546 31 572
rect -31 512 -17 546
rect 17 512 31 546
rect -31 474 31 512
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect 131 461 165 871
rect 279 535 313 945
rect 413 966 475 1004
rect 413 932 427 966
rect 461 932 475 966
rect 413 868 475 932
rect 649 1004 683 1020
rect 649 905 683 970
rect 279 461 313 501
rect 131 411 165 427
rect 205 427 313 461
rect 413 546 475 572
rect 413 512 427 546
rect 461 512 475 546
rect 413 474 475 512
rect 413 440 427 474
rect 461 440 475 474
rect -31 368 -17 402
rect 17 368 31 402
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect -31 62 31 80
rect 109 361 143 377
rect 109 289 143 327
rect 109 221 143 255
rect 205 245 239 427
rect 413 402 475 440
rect 649 461 683 871
rect 871 1004 905 1020
rect 871 831 905 970
rect 871 781 905 797
rect 945 757 979 1071
rect 1079 1076 1093 1110
rect 1127 1076 1141 1110
rect 1079 1038 1141 1076
rect 1251 1411 1285 1427
rect 1251 1343 1285 1377
rect 1251 1275 1285 1309
rect 1251 1207 1285 1241
rect 1251 1139 1285 1173
rect 1339 1343 1373 1492
rect 1745 1470 1807 1492
rect 1339 1275 1373 1309
rect 1339 1207 1373 1241
rect 1339 1157 1373 1173
rect 1427 1411 1637 1445
rect 1427 1343 1461 1377
rect 1427 1275 1461 1309
rect 1427 1207 1461 1241
rect 1427 1139 1461 1173
rect 1251 1071 1461 1105
rect 1515 1343 1549 1359
rect 1515 1275 1549 1309
rect 1515 1207 1549 1241
rect 1515 1139 1549 1173
rect 1603 1343 1637 1377
rect 1603 1275 1637 1309
rect 1603 1207 1637 1241
rect 1603 1157 1637 1173
rect 1745 1436 1759 1470
rect 1793 1436 1807 1470
rect 1745 1398 1807 1436
rect 1745 1364 1759 1398
rect 1793 1364 1807 1398
rect 1745 1326 1807 1364
rect 1745 1292 1759 1326
rect 1793 1292 1807 1326
rect 1745 1254 1807 1292
rect 1745 1220 1759 1254
rect 1793 1220 1807 1254
rect 1745 1182 1807 1220
rect 1745 1148 1759 1182
rect 1793 1148 1807 1182
rect 1745 1110 1807 1148
rect 1515 1071 1645 1105
rect 1079 1004 1093 1038
rect 1127 1004 1141 1038
rect 1079 966 1141 1004
rect 1079 932 1093 966
rect 1127 932 1141 966
rect 1079 868 1141 932
rect 1315 1004 1349 1020
rect 1315 905 1349 970
rect 1315 855 1349 871
rect 1537 1004 1571 1020
rect 649 411 683 427
rect 871 609 905 625
rect 871 461 905 575
rect 871 411 905 427
rect 205 195 239 211
rect 303 361 337 377
rect 303 289 337 327
rect 303 221 337 255
rect 109 151 143 187
rect 303 151 337 187
rect 143 117 205 151
rect 239 117 303 151
rect 109 62 143 117
rect 206 62 240 117
rect 303 62 337 117
rect 413 368 427 402
rect 461 368 475 402
rect 413 330 475 368
rect 413 296 427 330
rect 461 296 475 330
rect 413 258 475 296
rect 413 224 427 258
rect 461 224 475 258
rect 413 186 475 224
rect 413 152 427 186
rect 461 152 475 186
rect 413 114 475 152
rect 413 80 427 114
rect 461 80 475 114
rect 566 361 600 377
rect 760 361 794 377
rect 945 375 979 723
rect 1315 683 1349 699
rect 600 327 663 361
rect 697 327 760 361
rect 566 289 600 327
rect 566 221 600 255
rect 760 289 794 327
rect 566 151 600 187
rect 566 101 600 117
rect 663 236 697 252
rect 413 62 475 80
rect 663 62 697 202
rect 760 221 794 255
rect 857 341 979 375
rect 1079 546 1141 572
rect 1079 512 1093 546
rect 1127 512 1141 546
rect 1079 474 1141 512
rect 1079 440 1093 474
rect 1127 440 1141 474
rect 1079 402 1141 440
rect 1315 461 1349 649
rect 1315 411 1349 427
rect 1537 535 1571 970
rect 1537 461 1571 501
rect 1537 411 1571 427
rect 1611 757 1645 1071
rect 1745 1076 1759 1110
rect 1793 1076 1807 1110
rect 1893 1412 1927 1492
rect 1893 1344 1927 1378
rect 1893 1276 1927 1310
rect 1893 1208 1927 1242
rect 1893 1139 1927 1174
rect 1893 1083 1927 1105
rect 1981 1412 2015 1450
rect 1981 1344 2015 1378
rect 1981 1276 2015 1310
rect 1981 1208 2015 1242
rect 1981 1139 2015 1174
rect 1745 1038 1807 1076
rect 1745 1004 1759 1038
rect 1793 1004 1807 1038
rect 1745 966 1807 1004
rect 1981 979 2015 1105
rect 2069 1412 2103 1492
rect 2069 1344 2103 1378
rect 2069 1276 2103 1310
rect 2069 1208 2103 1242
rect 2069 1139 2103 1174
rect 2069 1083 2103 1105
rect 2189 1470 2251 1492
rect 2189 1436 2203 1470
rect 2237 1436 2251 1470
rect 2189 1398 2251 1436
rect 2189 1364 2203 1398
rect 2237 1364 2251 1398
rect 2189 1326 2251 1364
rect 2189 1292 2203 1326
rect 2237 1292 2251 1326
rect 2189 1254 2251 1292
rect 2189 1220 2203 1254
rect 2237 1220 2251 1254
rect 2189 1182 2251 1220
rect 2189 1148 2203 1182
rect 2237 1148 2251 1182
rect 2189 1110 2251 1148
rect 2189 1076 2203 1110
rect 2237 1076 2251 1110
rect 2189 1038 2251 1076
rect 1745 932 1759 966
rect 1793 932 1807 966
rect 1745 868 1807 932
rect 1907 945 2015 979
rect 2055 1003 2089 1019
rect 1907 905 1941 945
rect 1079 368 1093 402
rect 1127 368 1141 402
rect 857 245 891 341
rect 1079 330 1141 368
rect 857 195 891 211
rect 954 289 988 305
rect 954 221 988 255
rect 760 151 794 187
rect 954 151 988 187
rect 794 117 857 151
rect 891 117 954 151
rect 760 101 794 117
rect 954 101 988 117
rect 1079 296 1093 330
rect 1127 296 1141 330
rect 1079 258 1141 296
rect 1079 224 1093 258
rect 1127 224 1141 258
rect 1079 186 1141 224
rect 1079 152 1093 186
rect 1127 152 1141 186
rect 1079 114 1141 152
rect 1079 80 1093 114
rect 1127 80 1141 114
rect 1232 361 1266 377
rect 1426 361 1460 377
rect 1611 375 1645 723
rect 1907 609 1941 871
rect 1266 327 1329 361
rect 1363 327 1426 361
rect 1232 289 1266 327
rect 1232 221 1266 255
rect 1426 289 1460 327
rect 1232 151 1266 187
rect 1232 101 1266 117
rect 1329 236 1363 252
rect 1079 62 1141 80
rect 1329 62 1363 202
rect 1426 221 1460 255
rect 1523 341 1645 375
rect 1745 546 1807 572
rect 1745 512 1759 546
rect 1793 512 1807 546
rect 1745 474 1807 512
rect 1745 440 1759 474
rect 1793 440 1807 474
rect 1745 402 1807 440
rect 1907 461 1941 575
rect 2055 831 2089 969
rect 2189 1004 2203 1038
rect 2237 1004 2251 1038
rect 2189 966 2251 1004
rect 2189 932 2203 966
rect 2237 932 2251 966
rect 2189 868 2251 932
rect 2055 683 2089 797
rect 2055 609 2089 649
rect 2055 461 2089 575
rect 1907 427 2015 461
rect 1745 368 1759 402
rect 1793 368 1807 402
rect 1523 245 1557 341
rect 1745 330 1807 368
rect 1523 195 1557 211
rect 1620 289 1654 305
rect 1620 221 1654 255
rect 1426 151 1460 187
rect 1620 151 1654 187
rect 1460 117 1523 151
rect 1557 117 1620 151
rect 1426 101 1460 117
rect 1620 101 1654 117
rect 1745 296 1759 330
rect 1793 296 1807 330
rect 1745 258 1807 296
rect 1745 224 1759 258
rect 1793 224 1807 258
rect 1745 186 1807 224
rect 1745 152 1759 186
rect 1793 152 1807 186
rect 1745 114 1807 152
rect 1745 80 1759 114
rect 1793 80 1807 114
rect 1745 62 1807 80
rect 1883 361 1917 377
rect 1883 289 1917 327
rect 1883 221 1917 255
rect 1981 245 2015 427
rect 2055 411 2089 427
rect 2189 546 2251 572
rect 2189 512 2203 546
rect 2237 512 2251 546
rect 2189 474 2251 512
rect 2189 440 2203 474
rect 2237 440 2251 474
rect 2189 402 2251 440
rect 1981 195 2015 211
rect 2077 361 2111 377
rect 2077 289 2111 327
rect 2077 221 2111 255
rect 1883 151 1917 187
rect 2077 151 2111 187
rect 1917 117 1981 151
rect 2015 117 2077 151
rect 1883 62 1917 117
rect 1980 62 2014 117
rect 2077 62 2111 117
rect 2189 368 2203 402
rect 2237 368 2251 402
rect 2189 330 2251 368
rect 2189 296 2203 330
rect 2237 296 2251 330
rect 2189 258 2251 296
rect 2189 224 2203 258
rect 2237 224 2251 258
rect 2189 186 2251 224
rect 2189 152 2203 186
rect 2237 152 2251 186
rect 2189 114 2251 152
rect 2189 80 2203 114
rect 2237 80 2251 114
rect 2189 62 2251 80
rect -31 47 2251 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 205 47
rect 239 13 283 47
rect 317 13 355 47
rect 389 13 499 47
rect 533 13 571 47
rect 605 13 643 47
rect 677 13 715 47
rect 749 13 805 47
rect 839 13 877 47
rect 911 13 949 47
rect 983 13 1021 47
rect 1055 13 1165 47
rect 1199 13 1237 47
rect 1271 13 1309 47
rect 1343 13 1381 47
rect 1415 13 1471 47
rect 1505 13 1543 47
rect 1577 13 1615 47
rect 1649 13 1687 47
rect 1721 13 1831 47
rect 1865 13 1903 47
rect 1937 13 1981 47
rect 2015 13 2059 47
rect 2093 13 2131 47
rect 2165 13 2251 47
rect -31 0 2251 13
<< viali >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 205 1505 239 1539
rect 283 1505 317 1539
rect 355 1505 389 1539
rect 499 1505 533 1539
rect 571 1505 605 1539
rect 643 1505 677 1539
rect 715 1505 749 1539
rect 805 1505 839 1539
rect 877 1505 911 1539
rect 949 1505 983 1539
rect 1021 1505 1055 1539
rect 1165 1505 1199 1539
rect 1237 1505 1271 1539
rect 1309 1505 1343 1539
rect 1381 1505 1415 1539
rect 1471 1505 1505 1539
rect 1543 1505 1577 1539
rect 1615 1505 1649 1539
rect 1687 1505 1721 1539
rect 1831 1505 1865 1539
rect 1903 1505 1937 1539
rect 1981 1505 2015 1539
rect 2059 1505 2093 1539
rect 2131 1505 2165 1539
rect 131 871 165 905
rect 649 871 683 905
rect 279 501 313 535
rect 871 797 905 831
rect 1315 871 1349 905
rect 945 723 979 757
rect 871 575 905 609
rect 1315 649 1349 683
rect 1537 501 1571 535
rect 1907 871 1941 905
rect 1611 723 1645 757
rect 1907 575 1941 609
rect 2055 797 2089 831
rect 2055 649 2089 683
rect 2055 575 2089 609
rect 55 13 89 47
rect 127 13 161 47
rect 205 13 239 47
rect 283 13 317 47
rect 355 13 389 47
rect 499 13 533 47
rect 571 13 605 47
rect 643 13 677 47
rect 715 13 749 47
rect 805 13 839 47
rect 877 13 911 47
rect 949 13 983 47
rect 1021 13 1055 47
rect 1165 13 1199 47
rect 1237 13 1271 47
rect 1309 13 1343 47
rect 1381 13 1415 47
rect 1471 13 1505 47
rect 1543 13 1577 47
rect 1615 13 1649 47
rect 1687 13 1721 47
rect 1831 13 1865 47
rect 1903 13 1937 47
rect 1981 13 2015 47
rect 2059 13 2093 47
rect 2131 13 2165 47
<< metal1 >>
rect -31 1539 2251 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 205 1539
rect 239 1505 283 1539
rect 317 1505 355 1539
rect 389 1505 499 1539
rect 533 1505 571 1539
rect 605 1505 643 1539
rect 677 1505 715 1539
rect 749 1505 805 1539
rect 839 1505 877 1539
rect 911 1505 949 1539
rect 983 1505 1021 1539
rect 1055 1505 1165 1539
rect 1199 1505 1237 1539
rect 1271 1505 1309 1539
rect 1343 1505 1381 1539
rect 1415 1505 1471 1539
rect 1505 1505 1543 1539
rect 1577 1505 1615 1539
rect 1649 1505 1687 1539
rect 1721 1505 1831 1539
rect 1865 1505 1903 1539
rect 1937 1505 1981 1539
rect 2015 1505 2059 1539
rect 2093 1505 2131 1539
rect 2165 1505 2251 1539
rect -31 1492 2251 1505
rect 125 905 171 911
rect 643 905 689 911
rect 1309 905 1355 911
rect 1901 905 1947 911
rect 119 871 131 905
rect 165 871 649 905
rect 683 871 695 905
rect 1303 871 1315 905
rect 1349 871 1907 905
rect 1941 871 1953 905
rect 125 865 171 871
rect 643 865 689 871
rect 1309 865 1355 871
rect 1901 865 1947 871
rect 865 831 911 837
rect 2049 831 2095 837
rect 859 797 871 831
rect 905 797 2055 831
rect 2089 797 2101 831
rect 865 791 911 797
rect 2049 791 2095 797
rect 939 757 985 763
rect 1605 757 1651 763
rect 933 723 945 757
rect 979 723 1611 757
rect 1645 723 1657 757
rect 939 717 985 723
rect 1605 717 1651 723
rect 1309 683 1355 689
rect 2049 683 2095 689
rect 1303 649 1315 683
rect 1349 649 2055 683
rect 2089 649 2101 683
rect 1309 643 1355 649
rect 2049 643 2095 649
rect 865 609 911 615
rect 1901 609 1947 615
rect 2049 609 2095 615
rect 859 575 871 609
rect 905 575 1907 609
rect 1941 575 1953 609
rect 2019 575 2055 609
rect 2089 575 2101 609
rect 865 569 911 575
rect 1901 569 1947 575
rect 2049 569 2095 575
rect 273 535 319 541
rect 1531 535 1577 541
rect 267 501 279 535
rect 313 501 1537 535
rect 1571 501 1583 535
rect 273 495 319 501
rect 1531 495 1577 501
rect -31 47 2251 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 205 47
rect 239 13 283 47
rect 317 13 355 47
rect 389 13 499 47
rect 533 13 571 47
rect 605 13 643 47
rect 677 13 715 47
rect 749 13 805 47
rect 839 13 877 47
rect 911 13 949 47
rect 983 13 1021 47
rect 1055 13 1165 47
rect 1199 13 1237 47
rect 1271 13 1309 47
rect 1343 13 1381 47
rect 1415 13 1471 47
rect 1505 13 1543 47
rect 1577 13 1615 47
rect 1649 13 1687 47
rect 1721 13 1831 47
rect 1865 13 1903 47
rect 1937 13 1981 47
rect 2015 13 2059 47
rect 2093 13 2131 47
rect 2165 13 2251 47
rect -31 0 2251 13
<< labels >>
rlabel metal1 1611 723 1645 757 1 Y
port 1 n
rlabel metal1 131 871 165 905 1 A
port 2 n
rlabel metal1 2055 575 2089 609 1 B
port 3 n
rlabel metal1 55 1505 89 1539 1 VDD
port 4 n
rlabel metal1 55 13 89 47 1 VSS
port 5 n
<< end >>
