magic
tech sky130
magscale 1 2
timestamp 1652307457
<< error_p >>
rect -41 -17 -31 7
rect 31 -17 41 7
rect -17 -41 17 -31
<< nwell >>
rect -84 790 84 1533
<< pwell >>
rect -31 -31 31 541
<< psubdiff >>
rect -31 461 31 541
rect -31 427 -17 461
rect 17 427 31 461
rect -31 387 31 427
rect -31 353 -17 387
rect 17 353 31 387
rect -31 313 31 353
rect -31 279 -17 313
rect 17 279 31 313
rect -31 239 31 279
rect -31 205 -17 239
rect 17 205 31 239
rect -31 165 31 205
rect -31 131 -17 165
rect 17 131 31 165
rect -31 91 31 131
rect -31 57 -17 91
rect 17 57 31 91
rect -31 17 31 57
rect -31 -17 -17 17
rect 17 -17 31 17
rect -31 -31 31 -17
<< nsubdiff >>
rect -31 1423 31 1497
rect -31 1389 -17 1423
rect 17 1389 31 1423
rect -31 1349 31 1389
rect -31 1315 -17 1349
rect 17 1315 31 1349
rect -31 1275 31 1315
rect -31 1241 -17 1275
rect 17 1241 31 1275
rect -31 1201 31 1241
rect -31 1167 -17 1201
rect 17 1167 31 1201
rect -31 1127 31 1167
rect -31 1093 -17 1127
rect 17 1093 31 1127
rect -31 1053 31 1093
rect -31 1019 -17 1053
rect 17 1019 31 1053
rect -31 979 31 1019
rect -31 945 -17 979
rect 17 945 31 979
rect -31 905 31 945
rect -31 871 -17 905
rect 17 871 31 905
rect -31 826 31 871
<< psubdiffcont >>
rect -17 427 17 461
rect -17 353 17 387
rect -17 279 17 313
rect -17 205 17 239
rect -17 131 17 165
rect -17 57 17 91
rect -17 -17 17 17
<< nsubdiffcont >>
rect -17 1389 17 1423
rect -17 1315 17 1349
rect -17 1241 17 1275
rect -17 1167 17 1201
rect -17 1093 17 1127
rect -17 1019 17 1053
rect -17 945 17 979
rect -17 871 17 905
<< locali >>
rect -31 1497 31 1512
rect -31 1463 -17 1497
rect 17 1463 31 1497
rect -31 1423 31 1463
rect -31 1389 -17 1423
rect 17 1389 31 1423
rect -31 1349 31 1389
rect -31 1315 -17 1349
rect 17 1315 31 1349
rect -31 1275 31 1315
rect -31 1241 -17 1275
rect 17 1241 31 1275
rect -31 1201 31 1241
rect -31 1167 -17 1201
rect 17 1167 31 1201
rect -31 1127 31 1167
rect -31 1093 -17 1127
rect 17 1093 31 1127
rect -31 1053 31 1093
rect -31 1019 -17 1053
rect 17 1019 31 1053
rect -31 979 31 1019
rect -31 945 -17 979
rect 17 945 31 979
rect -31 905 31 945
rect -31 871 -17 905
rect 17 871 31 905
rect -31 826 31 871
rect -31 461 31 541
rect -31 427 -17 461
rect 17 427 31 461
rect -31 387 31 427
rect -31 353 -17 387
rect 17 353 31 387
rect -31 313 31 353
rect -31 279 -17 313
rect 17 279 31 313
rect -31 239 31 279
rect -31 205 -17 239
rect 17 205 31 239
rect -31 165 31 205
rect -31 131 -17 165
rect 17 131 31 165
rect -31 91 31 131
rect -31 57 -17 91
rect 17 57 31 91
rect -31 17 31 57
rect -31 -17 -17 17
rect 17 -17 31 17
rect -31 -31 31 -17
<< viali >>
rect -17 1463 17 1497
rect -17 -17 17 17
<< metal1 >>
rect -31 1497 31 1512
rect -31 1463 -17 1497
rect 17 1463 31 1497
rect -31 1450 31 1463
rect -31 17 31 31
rect -31 -17 -17 17
rect 17 -17 31 17
rect -31 -31 31 -17
<< end >>
