* SPICE3 file created from VOTERN3X1.ext - technology: sky130A

.subckt VOTERN3X1 YN A B C VDD VSS
X0 YN A a_112_102 VSS sky130_fd_pr__nfet_01v8 ad=5.373p pd=4.72u as=0p ps=0u w=3u l=0.15u
X1 a_217_1052 B VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.68p ps=1.368u w=2u l=0.15u M=2
X2 a_217_1052 B a_881_1052 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X3 YN C a_778_102 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X4 a_881_1052 A YN VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.16p ps=9.16u w=2u l=0.15u M=2
X5 a_217_1052 A VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X6 a_217_1052 C a_881_1052 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X7 YN C a_881_1052 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X8 VSS B a_778_102 VSS sky130_fd_pr__nfet_01v8 ad=5.373p pd=4.71u as=0p ps=0u w=3u l=0.15u
X9 VSS B a_112_102 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X10 VSS C a_1444_102 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X11 YN A a_1444_102 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u


.ends
