* SPICE3 file created from NOR2X1.ext - technology: sky130A

.subckt NOR2X1 Y A B VDD VSS
X0 a_131_1051 A VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=150000u M=2
X1 Y A VSS VSS sky130_fd_pr__nfet_01v8 ad=3.582e+11p pd=3.15e+06u as=1.9366e+12p ps=1.294e+07u w=3e+06u l=150000u
X2 a_131_1051 B Y VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=150000u M=2
X3 Y B VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
.ends
