* SPICE3 file created from INVX1.ext - technology: sky130A

.subckt INVX1 Y A VDD GND
X0 Y A.t1 GND.t0 GND sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=0p ps=0u w=0u l=0u
X1 Y.t1 A.t0 VDD.t3  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X2 Y A GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.1408p ps=8.1u w=3u l=0.15u
X3 VDD.t1 A.t2 Y.t0 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
C0 A VDD 0.38fF
C1 A Y 0.31fF
C2 VDD Y 1.04fF
R0 A.n0 A.t2 512.525
R1 A.n0 A.t0 371.139
R2 A.n1 A.t1 282.852
R3 A.n1 A.n0 247.347
R4 A.n2 A.n1 4.65
R5 A.n2 A 0.046
R6 VDD.n55 VDD.t3 135.17
R7 VDD.n24 VDD.t1 135.17
R8 VDD.n38 VDD.n37 92.5
R9 VDD.n36 VDD.n35 92.5
R10 VDD.n34 VDD.n33 92.5
R11 VDD.n32 VDD.n31 92.5
R12 VDD.n40 VDD.n39 92.5
R13 VDD.n14 VDD.n1 92.5
R14 VDD.n5 VDD.n4 92.5
R15 VDD.n7 VDD.n6 92.5
R16 VDD.n9 VDD.n8 92.5
R17 VDD.n11 VDD.n10 92.5
R18 VDD.n13 VDD.n12 92.5
R19 VDD.n21 VDD.n20 92.059
R20 VDD.n49 VDD.n48 92.059
R21 VDD.n20 VDD.n16 67.194
R22 VDD.n20 VDD.n17 67.194
R23 VDD.n20 VDD.n18 67.194
R24 VDD.n20 VDD.n19 67.194
R25 VDD.n5 VDD.n3 44.141
R26 VDD.n3 VDD.n2 44.107
R27 VDD.n25 VDD.t0 43.472
R28 VDD.n53  43.472
R29 VDD.n20 VDD.n15 41.052
R30 VDD.n47 VDD.n45 39.742
R31 VDD.n47 VDD.n46 39.742
R32 VDD.n44 VDD.n43 39.742
R33 VDD.n1 VDD.n0 30.923
R34 VDD.n48 VDD.n47 26.38
R35 VDD.n48 VDD.n44 26.38
R36 VDD.n48 VDD.n42 26.38
R37 VDD.n48 VDD.n41 26.38
R38 VDD.n51 VDD.n40 22.915
R39 VDD.n23 VDD.n14 22.915
R40 VDD.n40 VDD.n38 14.864
R41 VDD.n38 VDD.n36 14.864
R42 VDD.n36 VDD.n34 14.864
R43 VDD.n34 VDD.n32 14.864
R44 VDD.n32 VDD.n30 14.864
R45 VDD.n30 VDD.n29 14.864
R46 VDD.n14 VDD.n13 14.864
R47 VDD.n13 VDD.n11 14.864
R48 VDD.n11 VDD.n9 14.864
R49 VDD.n9 VDD.n7 14.864
R50 VDD.n7 VDD.n5 14.864
R51 VDD.n23 VDD.n22 8.855
R52 VDD.n22 VDD.n21 8.855
R53 VDD.n27 VDD.n26 8.855
R54 VDD.n26 VDD.n25 8.855
R55 VDD.n60 VDD.n59 8.855
R56 VDD.n59 VDD.n58 8.855
R57 VDD.n56 VDD.n54 8.855
R58 VDD.n54 VDD.n53 8.855
R59 VDD.n51 VDD.n50 8.855
R60 VDD.n50 VDD.n49 8.855
R61 VDD.n28 VDD.n23 4.795
R62 VDD.n28 VDD.n27 4.65
R63 VDD.n61 VDD.n60 4.65
R64 VDD.n57 VDD.n56 4.65
R65 VDD.n52 VDD.n51 4.65
R66 VDD.n27 VDD.n24 2.064
R67 VDD.n56 VDD.n55 2.064
R68 VDD.n52 VDD 0.207
R69 VDD.n61 VDD.n28 0.157
R70 VDD.n61 VDD.n57 0.157
R71 VDD.n57 VDD.n52 0.145
R72 Y.n5 Y.n4 272.451
R73 Y.n5 Y.n0 271.281
R74 Y.n4 Y.n3 30
R75 Y.n2 Y.n1 24.383
R76 Y.n4 Y.n2 23.684
R77 Y.n0 Y.t0 14.282
R78 Y.n0 Y.t1 14.282
R79 Y.n6 Y.n5 4.65
R80 Y.n6 Y 0.046
R81 GND.n18 GND.n17 37.582
R82 GND.t0 GND.n15 32.601
R83 GND.n15 GND.n14 21.734
R84 GND.n4 GND.n3 20.705
R85 GND.n24 GND.n23 20.705
R86 GND.n19 GND.n18 20.705
R87 GND.n3 GND.n2 19.952
R88 GND.n17 GND.t0 15.644
R89 GND.n17 GND.n16 13.541
R90 GND.n20 GND.n11 9.154
R91 GND.n26 GND.n25 9.154
R92 GND.n6 GND.n5 9.154
R93 GND.n7 GND.n1 4.795
R94 GND.n10 GND.n9 4.65
R95 GND.n7 GND.n6 4.65
R96 GND.n27 GND.n26 4.65
R97 GND.n21 GND.n20 4.65
R98 GND.n13 GND.n12 4.504
R99 GND.n6 GND.n4 4.129
R100 GND.n20 GND.n19 3.716
R101 GND.t0 GND.n13 2.452
R102 GND.n1 GND.n0 0.474
R103 GND.n9 GND.n8 0.474
R104 GND.n23 GND.n22 0.376
R105 GND.n10 GND 0.207
R106 GND.n26 GND.n24 0.206
R107 GND.n27 GND.n7 0.157
R108 GND.n27 GND.n21 0.157
R109 GND.n21 GND.n10 0.145
C3 VDD GND 0.98fF
C4 Y.n0 GND 0.63fF
C5 Y.n1 GND 0.04fF
C6 Y.n2 GND 0.05fF
C7 Y.n3 GND 0.03fF
C8 Y.n4 GND 0.18fF
C9 Y.n5 GND 0.61fF
C10 Y.n6 GND 0.01fF
C11 VDD.n1 GND 0.02fF
C12 VDD.n2 GND 0.06fF
C13 VDD.n3 GND 0.02fF
C14 VDD.n4 GND 0.01fF
C15 VDD.n5 GND 0.04fF
C16 VDD.n6 GND 0.01fF
C17 VDD.n7 GND 0.01fF
C18 VDD.n8 GND 0.01fF
C19 VDD.n9 GND 0.01fF
C20 VDD.n10 GND 0.01fF
C21 VDD.n11 GND 0.01fF
C22 VDD.n12 GND 0.01fF
C23 VDD.n13 GND 0.01fF
C24 VDD.n14 GND 0.02fF
C25 VDD.n15 GND 0.01fF
C26 VDD.n20 GND 0.27fF
C27 VDD.n21 GND 0.16fF
C28 VDD.n22 GND 0.01fF
C29 VDD.n23 GND 0.02fF
C30 VDD.n24 GND 0.04fF
C31 VDD.n25 GND 0.12fF
C32 VDD.n26 GND 0.01fF
C33 VDD.n27 GND 0.01fF
C34 VDD.n28 GND 0.04fF
C35 VDD.n29 GND 0.03fF
C36 VDD.n30 GND 0.01fF
C37 VDD.n31 GND 0.01fF
C38 VDD.n32 GND 0.01fF
C39 VDD.n33 GND 0.01fF
C40 VDD.n34 GND 0.01fF
C41 VDD.n35 GND 0.01fF
C42 VDD.n36 GND 0.01fF
C43 VDD.n37 GND 0.01fF
C44 VDD.n38 GND 0.01fF
C45 VDD.n39 GND 0.02fF
C46 VDD.n40 GND 0.02fF
C47 VDD.n43 GND 0.01fF
C48 VDD.n45 GND 0.01fF
C49 VDD.n46 GND 0.06fF
C50 VDD.n48 GND 0.27fF
C51 VDD.n49 GND 0.16fF
C52 VDD.n50 GND 0.01fF
C53 VDD.n51 GND 0.02fF
C54 VDD.n52 GND 0.02fF
C55 VDD.n53 GND 0.12fF
C56 VDD.n54 GND 0.01fF
C57 VDD.n55 GND 0.04fF
C58 VDD.n56 GND 0.01fF
C59 VDD.n57 GND 0.01fF
C60 VDD.n58 GND 0.10fF
C61 VDD.n59 GND 0.01fF
C62 VDD.n60 GND 0.01fF
C63 VDD.n61 GND 0.01fF
.ends
