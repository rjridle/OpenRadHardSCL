magic
tech sky130A
magscale 1 2
timestamp 1647328266
<< nwell >>
rect 84 1573 880 1575
rect 84 1556 878 1573
rect 84 1487 941 1556
rect 84 1145 878 1487
rect 84 1139 220 1145
rect 84 1105 205 1139
rect 229 1105 263 1139
rect 84 1102 220 1105
rect 279 1102 878 1145
rect 84 935 878 1102
rect 84 934 929 935
rect 84 859 931 934
rect 84 832 878 859
<< pdiffc >>
rect 201 1105 235 1139
rect 289 1105 323 1139
rect 465 1105 499 1139
rect 641 1105 675 1139
<< psubdiff >>
rect 31 510 931 572
rect 31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 343 47
rect 377 13 415 47
rect 449 13 513 47
rect 547 13 585 47
rect 619 13 657 47
rect 691 13 729 47
rect 763 13 801 47
rect 835 13 873 47
rect 907 13 931 47
<< nsubdiff >>
rect 31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 343 1539
rect 377 1505 415 1539
rect 449 1505 513 1539
rect 547 1505 585 1539
rect 619 1505 657 1539
rect 691 1505 729 1539
rect 763 1505 801 1539
rect 835 1505 873 1539
rect 907 1505 931 1539
rect 31 868 931 930
<< psubdiffcont >>
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 343 13 377 47
rect 415 13 449 47
rect 513 13 547 47
rect 585 13 619 47
rect 657 13 691 47
rect 729 13 763 47
rect 801 13 835 47
rect 873 13 907 47
<< nsubdiffcont >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 343 1505 377 1539
rect 415 1505 449 1539
rect 513 1505 547 1539
rect 585 1505 619 1539
rect 657 1505 691 1539
rect 729 1505 763 1539
rect 801 1505 835 1539
rect 873 1505 907 1539
<< poly >>
rect 147 411 195 441
rect 471 411 477 441
rect 147 405 177 411
rect 447 405 477 411
<< locali >>
rect 31 1539 931 1554
rect 31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 343 1539
rect 377 1505 415 1539
rect 449 1505 513 1539
rect 547 1505 585 1539
rect 619 1505 657 1539
rect 691 1505 729 1539
rect 763 1505 801 1539
rect 835 1505 873 1539
rect 907 1505 931 1539
rect 31 1492 931 1505
rect 201 1139 235 1162
rect 201 1089 235 1105
rect 289 1139 323 1157
rect 289 1094 323 1105
rect 465 1139 499 1157
rect 465 1094 499 1105
rect 641 1139 675 1157
rect 641 1094 675 1105
rect 289 1060 831 1094
rect 205 461 239 954
rect 427 461 461 954
rect 649 477 683 986
rect 797 378 831 1060
rect 700 344 831 378
rect 700 263 734 344
rect 393 210 603 244
rect 198 62 232 195
rect 31 47 931 62
rect 31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 343 47
rect 377 13 415 47
rect 449 13 513 47
rect 547 13 585 47
rect 619 13 657 47
rect 691 13 729 47
rect 763 13 801 47
rect 835 13 873 47
rect 907 13 931 47
rect 31 0 931 13
<< viali >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 343 1505 377 1539
rect 415 1505 449 1539
rect 513 1505 547 1539
rect 585 1505 619 1539
rect 657 1505 691 1539
rect 729 1505 763 1539
rect 801 1505 835 1539
rect 873 1505 907 1539
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 343 13 377 47
rect 415 13 449 47
rect 513 13 547 47
rect 585 13 619 47
rect 657 13 691 47
rect 729 13 763 47
rect 801 13 835 47
rect 873 13 907 47
<< metal1 >>
rect 31 1539 931 1554
rect 31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 343 1539
rect 377 1505 415 1539
rect 449 1505 513 1539
rect 547 1505 585 1539
rect 619 1505 657 1539
rect 691 1505 729 1539
rect 763 1505 801 1539
rect 835 1505 873 1539
rect 907 1505 931 1539
rect 31 1492 931 1505
rect 31 47 931 62
rect 31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 343 47
rect 377 13 415 47
rect 449 13 513 47
rect 547 13 585 47
rect 619 13 657 47
rect 691 13 729 47
rect 763 13 801 47
rect 835 13 873 47
rect 907 13 931 47
rect 31 0 931 13
use pmos2  pmos2_0
timestamp 1647328240
transform 1 0 103 0 1 1450
box 52 -460 352 42
use diff_ring_side  diff_ring_side_1
timestamp 1646086970
transform 1 0 0 0 1 0
box -84 0 84 1575
use nmos_bottom  nmos_bottom_0
timestamp 1646007130
transform -1 0 339 0 1 103
box 0 0 248 302
use poly_li1_contact  poly_li1_contact_0
timestamp 1645652543
transform 0 1 222 -1 0 987
box -33 -27 33 27
use poly_li1_contact  poly_li1_contact_1
timestamp 1645652543
transform 0 -1 222 1 0 444
box -33 -27 33 27
use pmos2  pmos2_2
timestamp 1647328240
transform 1 0 455 0 1 1450
box 52 -460 352 42
use pmos2  pmos2_1
timestamp 1647328240
transform 1 0 279 0 1 1450
box 52 -460 352 42
use poly_li1_contact  poly_li1_contact_2
timestamp 1645652543
transform 0 -1 444 1 0 444
box -33 -27 33 27
use poly_li1_contact  poly_li1_contact_3
timestamp 1645652543
transform 0 -1 444 1 0 987
box -33 -27 33 27
use nmos_side_left  nmos_side_left_0
timestamp 1645918720
transform 1 0 285 0 1 103
box 0 0 248 302
use nmos_top_trim1  nmos_top_trim1_0
timestamp 1646008046
transform -1 0 841 0 1 103
box 0 0 248 309
use poly_li1_contact  poly_li1_contact_4
timestamp 1645652543
transform 0 -1 666 1 0 444
box -33 -27 33 27
use poly_li1_contact  poly_li1_contact_5
timestamp 1645652543
transform 0 1 666 -1 0 987
box -33 -27 33 27
use diff_ring_side  diff_ring_side_0
timestamp 1646086970
transform 1 0 962 0 1 0
box -84 0 84 1575
<< end >>
