* NGSPICE file created from DFFX1.ext - technology: sky130A

.subckt nmos_bottom a_86_101# a_56_85# a_0_0# VSUBS
X0 a_86_101# a_56_85# a_0_0# VSUBS sky130_fd_pr__nfet_01v8 ad=1.772e+11p pd=1.56e+06u as=1.152e+12p ps=8.19e+06u w=3e+06u l=150000u
.ends

.subckt nmos_top_trim1 a_56_92# a_86_108# a_0_0# VSUBS
X0 a_86_108# a_56_92# a_0_0# VSUBS sky130_fd_pr__nfet_01v8 ad=1.772e+11p pd=1.56e+06u as=1.15725e+12p ps=8.12e+06u w=3e+06u l=150000u
.ends

.subckt pmos2 a_144_n460# a_262_n399# a_88_n399# w_52_n435# a_174_n399#
X0 a_174_n399# a_144_n460# a_88_n399# w_52_n435# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.6e+11p ps=4.56e+06u w=2e+06u l=150000u
X1 a_262_n399# a_144_n460# a_174_n399# w_52_n435# sky130_fd_pr__pfet_01v8 ad=5.4e+11p pd=4.54e+06u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt nand2x1_pcell VSS VDD a_229_1105# a_168_403# a_362_410#
Xnmos_bottom_0 VSS a_168_403# nmos_bottom_0/a_0_0# VSS nmos_bottom
Xnmos_top_trim1_0 a_362_410# a_229_1105# nmos_bottom_0/a_0_0# VSS nmos_top_trim1
Xpmos2_0 a_168_403# VDD VDD VDD a_229_1105# pmos2
Xpmos2_1 a_362_410# VDD VDD VDD a_229_1105# pmos2
.ends

.subckt nmos_side_left a_87_107# a_57_91# a_0_0# VSUBS
X0 a_87_107# a_57_91# a_0_0# VSUBS sky130_fd_pr__nfet_01v8 ad=1.6345e+11p pd=1.49e+06u as=1.17945e+12p ps=8.17e+06u w=3e+06u l=150000u
.ends

.subckt nand3x1_pcell VSS VDD a_289_1105# a_147_405# a_447_405# li_649_477# a_31_510#
Xnmos_bottom_0 VSS a_147_405# nmos_bottom_0/a_0_0# VSS nmos_bottom
Xnmos_top_trim1_0 li_649_477# a_289_1105# li_393_210# VSS nmos_top_trim1
Xnmos_side_left_0 li_393_210# a_447_405# nmos_bottom_0/a_0_0# VSS nmos_side_left
Xpmos2_0 a_147_405# VDD VDD VDD a_289_1105# pmos2
Xpmos2_1 a_447_405# VDD VDD VDD a_289_1105# pmos2
Xpmos2_2 li_649_477# VDD VDD VDD a_289_1105# pmos2
.ends

.subckt DFFX1 VSS VDD CLK D Q QN
Xnand2x1_pcell_2 VSS VDD m1_463_871# CLK m1_2165_723# nand2x1_pcell
Xnand2x1_pcell_3 VSS VDD QN m1_833_649# Q nand2x1_pcell
Xnand2x1_pcell_4 VSS VDD Q m1_463_871# QN nand2x1_pcell
Xnand3x1_pcell_0 VSS VDD m1_833_649# CLK m1_463_871# m1_685_723# VSS nand3x1_pcell
Xnand2x1_pcell_0 VSS VDD m1_685_723# m1_833_649# D nand2x1_pcell
Xnand2x1_pcell_1 VSS VDD m1_2165_723# m1_463_871# m1_685_723# nand2x1_pcell
.ends

