* SPICE3 file created from DFFRNQX1.ext - technology: sky130A

.subckt DFFRNQX1 Q D CLK RN VDD VSS
X0 a_599_989.t2 D.t0 VDD.t37 @��}�U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X1 VDD.t39 CLK.t0 a_277_1050.t5  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X2 VDD.t49 a_599_989.t7 a_2141_1050.t3 VDD.t48 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X3 VDD.t3 a_277_1050.t7 a_3829_1050.t2  \R. sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X4 a_599_989.t0 RN.t0 VDD.t33 �[R. sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X5 a_147_187.t3 CLK.t1 VDD.t11  \R. sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X6 a_3829_1050.t4 Q.t5 VDD.t47 �[R. sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X7 Q.t4 a_3829_1050.t7 VDD.t15  \R. sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X8 VDD.t25 a_599_989.t8 a_277_1050.t2 �[R. sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X9 VDD.t31 a_147_187.t9 a_2141_1050.t1  \R. sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X10 VDD.t9 a_2141_1050.t5 a_147_187.t1 �[R. sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X11 a_147_187.t4 RN.t1 VDD.t57  \R. sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X12 VSS a_147_187.t12 a_91_103.t0 VSS sky130_fd_pr__nfet_01v8 ad=1.0746p pd=9.42u as=0p ps=0u w=0u l=0u
X13 Q.t1 a_147_187.t10 VDD.t5 �[R. sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X14 a_277_1050.t0 a_147_187.t11 VDD.t29  \R. sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X15 VDD.t51 a_277_1050.t8 a_599_989.t3 �[R. sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X16 VDD.t59 RN.t3 a_599_989.t5  \R. sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X17 VDD.t43 Q.t6 a_3829_1050.t3 �[R. sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X18 VSS a_277_1050.t11 a_3643_103.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X19 a_277_1050.t4 CLK.t2 VDD.t1  \R. sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X20 a_2141_1050.t2 a_599_989.t10 VDD.t7 �[R. sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X21 a_3829_1050.t1 a_277_1050.t9 VDD.t19  \R. sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X22 VSS a_3829_1050.t8 a_4626_101.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X23 VDD.t55 RN.t4 a_3829_1050.t6 �[R. sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X24 VSS a_599_989.t12 a_2036_101.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X25 VDD.t35 D.t2 a_599_989.t1  \R. sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X26 VSS a_2141_1050.t7 a_2681_103.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X27 a_599_989.t6 a_277_1050.t10 VDD.t61 �[R. sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X28 a_277_1050.t1 a_599_989.t11 VDD.t23  \R. sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X29 a_2141_1050.t0 a_147_187.t13 VDD.t27 �[R. sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X30 a_3829_1050.t5 RN.t5 VDD.t53  \R. sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X31 a_147_187.t0 a_2141_1050.t6 VDD.t21 �[R. sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X32 VDD.t17 CLK.t4 a_147_187.t2  \R. sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X33 VDD.t41 a_3829_1050.t9 Q.t3 �[R. sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X34 VSS a_277_1050.t12 a_1053_103.t0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X35 VDD.t63 RN.t8 a_147_187.t6  \R. sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X36 VDD.t13 a_147_187.t14 Q.t0 �[R. sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X37 Q a_147_187.t7 a_4626_101.t0 VSS sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=0p ps=0u w=0u l=0u
X38 VDD.t45 a_147_187.t15 a_277_1050.t6  \R. sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
C0 D RN 0.18fF
C1 CLK VDD 1.98fF
C2 CLK RN 0.28fF
C3 CLK D 0.07fF
C4 Q VDD 2.14fF
C5 RN VDD 0.89fF
C6 Q RN 0.18fF
C7 D VDD 0.29fF
R0 D.n0 D.t2 479.223
R1 D.n0 D.t0 375.52
R2 D.n1 D.t1 287.572
R3 D.n1 D.n0 196.47
R4 D.n2 D.n1 4.65
R5 D.n2 D 0.046
R6 VDD.n286 VDD.n279 144.705
R7 VDD.n229 VDD.n222 144.705
R8 VDD.n154 VDD.n147 144.705
R9 VDD.n79 VDD.n68 144.705
R10 VDD.n362 VDD.n351 144.705
R11 VDD.n371 VDD.t25 143.754
R12 VDD.n295 VDD.t59 143.754
R13 VDD.n163 VDD.t63 143.754
R14 VDD.n88 VDD.t43 143.754
R15 VDD.n232 VDD.t31 143.754
R16 VDD.n24 VDD.t13 143.754
R17 VDD.n401 VDD.t29 135.17
R18 VDD.n325 VDD.t61 135.17
R19 VDD.n254 VDD.t7 135.17
R20 VDD.n193 VDD.t21 135.17
R21 VDD.n118 VDD.t19 135.17
R22 VDD.n46 VDD.t15 135.17
R23 VDD.n392 VDD.n391 129.472
R24 VDD.n380 VDD.n379 129.472
R25 VDD.n316 VDD.n315 129.472
R26 VDD.n304 VDD.n303 129.472
R27 VDD.n242 VDD.n241 129.472
R28 VDD.n184 VDD.n183 129.472
R29 VDD.n172 VDD.n171 129.472
R30 VDD.n109 VDD.n108 129.472
R31 VDD.n97 VDD.n96 129.472
R32 VDD.n34 VDD.n33 129.472
R33 VDD.n64 VDD.n63 92.5
R34 VDD.n62 VDD.n61 92.5
R35 VDD.n60 VDD.n59 92.5
R36 VDD.n58 VDD.n57 92.5
R37 VDD.n66 VDD.n65 92.5
R38 VDD.n143 VDD.n142 92.5
R39 VDD.n141 VDD.n140 92.5
R40 VDD.n139 VDD.n138 92.5
R41 VDD.n137 VDD.n136 92.5
R42 VDD.n145 VDD.n144 92.5
R43 VDD.n218 VDD.n217 92.5
R44 VDD.n216 VDD.n215 92.5
R45 VDD.n214 VDD.n213 92.5
R46 VDD.n212 VDD.n211 92.5
R47 VDD.n220 VDD.n219 92.5
R48 VDD.n275 VDD.n274 92.5
R49 VDD.n273 VDD.n272 92.5
R50 VDD.n271 VDD.n270 92.5
R51 VDD.n269 VDD.n268 92.5
R52 VDD.n277 VDD.n276 92.5
R53 VDD.n347 VDD.n346 92.5
R54 VDD.n345 VDD.n344 92.5
R55 VDD.n343 VDD.n342 92.5
R56 VDD.n341 VDD.n340 92.5
R57 VDD.n349 VDD.n348 92.5
R58 VDD.n421 VDD.n420 92.5
R59 VDD.n419 VDD.n418 92.5
R60 VDD.n417 VDD.n416 92.5
R61 VDD.n415 VDD.n414 92.5
R62 VDD.n423 VDD.n422 92.5
R63 VDD.n14 VDD.n1 92.5
R64 VDD.n5 VDD.n4 92.5
R65 VDD.n7 VDD.n6 92.5
R66 VDD.n9 VDD.n8 92.5
R67 VDD.n11 VDD.n10 92.5
R68 VDD.n13 VDD.n12 92.5
R69 VDD.n21 VDD.n20 92.059
R70 VDD.n78 VDD.n77 92.059
R71 VDD.n153 VDD.n152 92.059
R72 VDD.n228 VDD.n227 92.059
R73 VDD.n285 VDD.n284 92.059
R74 VDD.n361 VDD.n360 92.059
R75 VDD.n429 VDD.n428 92.059
R76 VDD.n20 VDD.n16 67.194
R77 VDD.n20 VDD.n17 67.194
R78 VDD.n20 VDD.n18 67.194
R79 VDD.n20 VDD.n19 67.194
R80 VDD.n413 VDD.n412 44.141
R81 VDD.n267 VDD.n266 44.141
R82 VDD.n210 VDD.n209 44.141
R83 VDD.n135 VDD.n134 44.141
R84 VDD.n5 VDD.n3 44.141
R85 VDD.n266 VDD.n264 44.107
R86 VDD.n209 VDD.n207 44.107
R87 VDD.n134 VDD.n132 44.107
R88 VDD.n412 VDD.n410 44.107
R89 VDD.n3 VDD.n2 44.107
R90 VDD.n20 VDD.n15 41.052
R91 VDD.n72 VDD.n70 39.742
R92 VDD.n72 VDD.n71 39.742
R93 VDD.n74 VDD.n73 39.742
R94 VDD.n149 VDD.n148 39.742
R95 VDD.n224 VDD.n223 39.742
R96 VDD.n281 VDD.n280 39.742
R97 VDD.n425 VDD.n424 39.742
R98 VDD.n359 VDD.n356 39.742
R99 VDD.n359 VDD.n358 39.742
R100 VDD.n355 VDD.n354 39.742
R101 VDD.n134 VDD.n133 38
R102 VDD.n209 VDD.n208 38
R103 VDD.n266 VDD.n265 38
R104 VDD.n412 VDD.n411 38
R105 VDD.n264 VDD.n263 36.774
R106 VDD.n207 VDD.n206 36.774
R107 VDD.n132 VDD.n131 36.774
R108 VDD.n70 VDD.n69 36.774
R109 VDD.n358 VDD.n357 36.774
R110 VDD.n90 �[R. 35.8
R111 VDD.n165  \R. 35.8
R112 VDD.n297  \R. 35.8
R113 VDD.n373 �[R. 35.8
R114 VDD.n114  \R. 33.243
R115 VDD.n189 �[R. 33.243
R116 VDD.n321 �[R. 33.243
R117 VDD.n397  \R. 33.243
R118 VDD.n1 VDD.n0 30.923
R119 VDD.n77 VDD.n75 26.38
R120 VDD.n77 VDD.n74 26.38
R121 VDD.n77 VDD.n72 26.38
R122 VDD.n77 VDD.n76 26.38
R123 VDD.n152 VDD.n150 26.38
R124 VDD.n152 VDD.n149 26.38
R125 VDD.n152 VDD.n151 26.38
R126 VDD.n227 VDD.n225 26.38
R127 VDD.n227 VDD.n224 26.38
R128 VDD.n227 VDD.n226 26.38
R129 VDD.n284 VDD.n282 26.38
R130 VDD.n284 VDD.n281 26.38
R131 VDD.n284 VDD.n283 26.38
R132 VDD.n428 VDD.n426 26.38
R133 VDD.n428 VDD.n425 26.38
R134 VDD.n428 VDD.n427 26.38
R135 VDD.n360 VDD.n359 26.38
R136 VDD.n360 VDD.n355 26.38
R137 VDD.n360 VDD.n353 26.38
R138 VDD.n360 VDD.n352 26.38
R139 VDD.n431 VDD.n423 22.915
R140 VDD.n23 VDD.n14 22.915
R141 VDD.n29 �[R. 20.457
R142 VDD.n237  \R. 20.457
R143 VDD.n42  \R. 17.9
R144 VDD.n250 �[R. 17.9
R145 VDD.n94 �[R. 15.343
R146 VDD.n169  \R. 15.343
R147 VDD.n301 �[R. 15.343
R148 VDD.n377  \R. 15.343
R149 VDD.n423 VDD.n421 14.864
R150 VDD.n421 VDD.n419 14.864
R151 VDD.n419 VDD.n417 14.864
R152 VDD.n417 VDD.n415 14.864
R153 VDD.n415 VDD.n413 14.864
R154 VDD.n277 VDD.n275 14.864
R155 VDD.n275 VDD.n273 14.864
R156 VDD.n273 VDD.n271 14.864
R157 VDD.n271 VDD.n269 14.864
R158 VDD.n269 VDD.n267 14.864
R159 VDD.n220 VDD.n218 14.864
R160 VDD.n218 VDD.n216 14.864
R161 VDD.n216 VDD.n214 14.864
R162 VDD.n214 VDD.n212 14.864
R163 VDD.n212 VDD.n210 14.864
R164 VDD.n145 VDD.n143 14.864
R165 VDD.n143 VDD.n141 14.864
R166 VDD.n141 VDD.n139 14.864
R167 VDD.n139 VDD.n137 14.864
R168 VDD.n137 VDD.n135 14.864
R169 VDD.n66 VDD.n64 14.864
R170 VDD.n64 VDD.n62 14.864
R171 VDD.n62 VDD.n60 14.864
R172 VDD.n60 VDD.n58 14.864
R173 VDD.n58 VDD.n56 14.864
R174 VDD.n56 VDD.n55 14.864
R175 VDD.n349 VDD.n347 14.864
R176 VDD.n347 VDD.n345 14.864
R177 VDD.n345 VDD.n343 14.864
R178 VDD.n343 VDD.n341 14.864
R179 VDD.n341 VDD.n339 14.864
R180 VDD.n339 VDD.n338 14.864
R181 VDD.n14 VDD.n13 14.864
R182 VDD.n13 VDD.n11 14.864
R183 VDD.n11 VDD.n9 14.864
R184 VDD.n9 VDD.n7 14.864
R185 VDD.n7 VDD.n5 14.864
R186 VDD.n80 VDD.n67 14.864
R187 VDD.n155 VDD.n146 14.864
R188 VDD.n230 VDD.n221 14.864
R189 VDD.n287 VDD.n278 14.864
R190 VDD.n363 VDD.n350 14.864
R191 VDD.n391 VDD.t1 14.282
R192 VDD.n391 VDD.t45 14.282
R193 VDD.n379 VDD.t23 14.282
R194 VDD.n379 VDD.t39 14.282
R195 VDD.n315 VDD.t37 14.282
R196 VDD.n315 VDD.t51 14.282
R197 VDD.n303 VDD.t33 14.282
R198 VDD.n303 VDD.t35 14.282
R199 VDD.n241 VDD.t27 14.282
R200 VDD.n241 VDD.t49 14.282
R201 VDD.n183 VDD.t11 14.282
R202 VDD.n183 VDD.t9 14.282
R203 VDD.n171 VDD.t57 14.282
R204 VDD.n171 VDD.t17 14.282
R205 VDD.n108 VDD.t53 14.282
R206 VDD.n108 VDD.t3 14.282
R207 VDD.n96 VDD.t47 14.282
R208 VDD.n96 VDD.t55 14.282
R209 VDD.n33 VDD.t5 14.282
R210 VDD.n33 VDD.t41 14.282
R211 VDD.n110  \R. 12.786
R212 VDD.n185 �[R. 12.786
R213 VDD.n317 �[R. 12.786
R214 VDD.n393  \R. 12.786
R215 VDD.n36 VDD.n34 9.083
R216 VDD.n244 VDD.n242 9.083
R217 VDD.n23 VDD.n22 8.855
R218 VDD.n22 VDD.n21 8.855
R219 VDD.n27 VDD.n26 8.855
R220 VDD.n26 VDD.n25 8.855
R221 VDD.n31 VDD.n30 8.855
R222 VDD.n30 VDD.n29 8.855
R223 VDD.n36 VDD.n35 8.855
R224 VDD.n35 �[R. 8.855
R225 VDD.n40 VDD.n39 8.855
R226 VDD.n39 VDD.n38 8.855
R227 VDD.n44 VDD.n43 8.855
R228 VDD.n43 VDD.n42 8.855
R229 VDD.n49 VDD.n48 8.855
R230 VDD.n48 VDD.n47 8.855
R231 VDD.n53 VDD.n52 8.855
R232 VDD.n52 VDD.n51 8.855
R233 VDD.n80 VDD.n79 8.855
R234 VDD.n79 VDD.n78 8.855
R235 VDD.n84 VDD.n83 8.855
R236 VDD.n83 VDD.n82 8.855
R237 VDD.n88 VDD.n87 8.855
R238 VDD.n87 VDD.n86 8.855
R239 VDD.n92 VDD.n91 8.855
R240 VDD.n91 VDD.n90 8.855
R241 VDD.n98 VDD.n95 8.855
R242 VDD.n95 VDD.n94 8.855
R243 VDD.n102 VDD.n101 8.855
R244 VDD.n101 VDD.n100 8.855
R245 VDD.n106 VDD.n105 8.855
R246 VDD.n105 VDD.n104 8.855
R247 VDD.n112 VDD.n111 8.855
R248 VDD.n111 VDD.n110 8.855
R249 VDD.n116 VDD.n115 8.855
R250 VDD.n115 VDD.n114 8.855
R251 VDD.n121 VDD.n120 8.855
R252 VDD.n120 VDD.n119 8.855
R253 VDD.n125 VDD.n124 8.855
R254 VDD.n124 VDD.n123 8.855
R255 VDD.n129 VDD.n128 8.855
R256 VDD.n128 VDD.n127 8.855
R257 VDD.n155 VDD.n154 8.855
R258 VDD.n154 VDD.n153 8.855
R259 VDD.n159 VDD.n158 8.855
R260 VDD.n158 VDD.n157 8.855
R261 VDD.n163 VDD.n162 8.855
R262 VDD.n162 VDD.n161 8.855
R263 VDD.n167 VDD.n166 8.855
R264 VDD.n166 VDD.n165 8.855
R265 VDD.n173 VDD.n170 8.855
R266 VDD.n170 VDD.n169 8.855
R267 VDD.n177 VDD.n176 8.855
R268 VDD.n176 VDD.n175 8.855
R269 VDD.n181 VDD.n180 8.855
R270 VDD.n180 VDD.n179 8.855
R271 VDD.n187 VDD.n186 8.855
R272 VDD.n186 VDD.n185 8.855
R273 VDD.n191 VDD.n190 8.855
R274 VDD.n190 VDD.n189 8.855
R275 VDD.n196 VDD.n195 8.855
R276 VDD.n195 VDD.n194 8.855
R277 VDD.n200 VDD.n199 8.855
R278 VDD.n199 VDD.n198 8.855
R279 VDD.n204 VDD.n203 8.855
R280 VDD.n203 VDD.n202 8.855
R281 VDD.n230 VDD.n229 8.855
R282 VDD.n229 VDD.n228 8.855
R283 VDD.n235 VDD.n234 8.855
R284 VDD.n234 VDD.n233 8.855
R285 VDD.n239 VDD.n238 8.855
R286 VDD.n238 VDD.n237 8.855
R287 VDD.n244 VDD.n243 8.855
R288 VDD.n243 �[R. 8.855
R289 VDD.n248 VDD.n247 8.855
R290 VDD.n247 VDD.n246 8.855
R291 VDD.n252 VDD.n251 8.855
R292 VDD.n251 VDD.n250 8.855
R293 VDD.n257 VDD.n256 8.855
R294 VDD.n256 VDD.n255 8.855
R295 VDD.n261 VDD.n260 8.855
R296 VDD.n260 VDD.n259 8.855
R297 VDD.n287 VDD.n286 8.855
R298 VDD.n286 VDD.n285 8.855
R299 VDD.n291 VDD.n290 8.855
R300 VDD.n290 VDD.n289 8.855
R301 VDD.n295 VDD.n294 8.855
R302 VDD.n294 VDD.n293 8.855
R303 VDD.n299 VDD.n298 8.855
R304 VDD.n298 VDD.n297 8.855
R305 VDD.n305 VDD.n302 8.855
R306 VDD.n302 VDD.n301 8.855
R307 VDD.n309 VDD.n308 8.855
R308 VDD.n308 VDD.n307 8.855
R309 VDD.n313 VDD.n312 8.855
R310 VDD.n312 VDD.n311 8.855
R311 VDD.n319 VDD.n318 8.855
R312 VDD.n318 VDD.n317 8.855
R313 VDD.n323 VDD.n322 8.855
R314 VDD.n322 VDD.n321 8.855
R315 VDD.n328 VDD.n327 8.855
R316 VDD.n327 VDD.n326 8.855
R317 VDD.n332 VDD.n331 8.855
R318 VDD.n331 VDD.n330 8.855
R319 VDD.n336 VDD.n335 8.855
R320 VDD.n335 VDD.n334 8.855
R321 VDD.n363 VDD.n362 8.855
R322 VDD.n362 VDD.n361 8.855
R323 VDD.n367 VDD.n366 8.855
R324 VDD.n366 VDD.n365 8.855
R325 VDD.n371 VDD.n370 8.855
R326 VDD.n370 VDD.n369 8.855
R327 VDD.n375 VDD.n374 8.855
R328 VDD.n374 VDD.n373 8.855
R329 VDD.n381 VDD.n378 8.855
R330 VDD.n378 VDD.n377 8.855
R331 VDD.n385 VDD.n384 8.855
R332 VDD.n384 VDD.n383 8.855
R333 VDD.n389 VDD.n388 8.855
R334 VDD.n388 VDD.n387 8.855
R335 VDD.n395 VDD.n394 8.855
R336 VDD.n394 VDD.n393 8.855
R337 VDD.n399 VDD.n398 8.855
R338 VDD.n398 VDD.n397 8.855
R339 VDD.n404 VDD.n403 8.855
R340 VDD.n403 VDD.n402 8.855
R341 VDD.n408 VDD.n407 8.855
R342 VDD.n407 VDD.n406 8.855
R343 VDD.n431 VDD.n430 8.855
R344 VDD.n430 VDD.n429 8.855
R345 VDD.n278 VDD.n277 8.051
R346 VDD.n221 VDD.n220 8.051
R347 VDD.n146 VDD.n145 8.051
R348 VDD.n67 VDD.n66 8.051
R349 VDD.n350 VDD.n349 8.051
R350 VDD.n104  \R. 7.671
R351 VDD.n179  \R. 7.671
R352 VDD.n311 @��}�U 7.671
R353 VDD.n387  \R. 7.671
R354 VDD.n112 VDD.n109 7.019
R355 VDD.n187 VDD.n184 7.019
R356 VDD.n319 VDD.n316 7.019
R357 VDD.n395 VDD.n392 7.019
R358 VDD.n98 VDD.n97 6.606
R359 VDD.n173 VDD.n172 6.606
R360 VDD.n305 VDD.n304 6.606
R361 VDD.n381 VDD.n380 6.606
R362 VDD.n100 �[R. 5.114
R363 VDD.n175  \R. 5.114
R364 VDD.n307  \R. 5.114
R365 VDD.n383 @{o}�U 5.114
R366 VDD.n32 VDD.n31 4.65
R367 VDD.n37 VDD.n36 4.65
R368 VDD.n41 VDD.n40 4.65
R369 VDD.n45 VDD.n44 4.65
R370 VDD.n50 VDD.n49 4.65
R371 VDD.n54 VDD.n53 4.65
R372 VDD.n81 VDD.n80 4.65
R373 VDD.n85 VDD.n84 4.65
R374 VDD.n89 VDD.n88 4.65
R375 VDD.n93 VDD.n92 4.65
R376 VDD.n99 VDD.n98 4.65
R377 VDD.n103 VDD.n102 4.65
R378 VDD.n107 VDD.n106 4.65
R379 VDD.n113 VDD.n112 4.65
R380 VDD.n117 VDD.n116 4.65
R381 VDD.n122 VDD.n121 4.65
R382 VDD.n126 VDD.n125 4.65
R383 VDD.n130 VDD.n129 4.65
R384 VDD.n156 VDD.n155 4.65
R385 VDD.n160 VDD.n159 4.65
R386 VDD.n164 VDD.n163 4.65
R387 VDD.n168 VDD.n167 4.65
R388 VDD.n174 VDD.n173 4.65
R389 VDD.n178 VDD.n177 4.65
R390 VDD.n182 VDD.n181 4.65
R391 VDD.n188 VDD.n187 4.65
R392 VDD.n192 VDD.n191 4.65
R393 VDD.n197 VDD.n196 4.65
R394 VDD.n201 VDD.n200 4.65
R395 VDD.n205 VDD.n204 4.65
R396 VDD.n231 VDD.n230 4.65
R397 VDD.n236 VDD.n235 4.65
R398 VDD.n240 VDD.n239 4.65
R399 VDD.n245 VDD.n244 4.65
R400 VDD.n249 VDD.n248 4.65
R401 VDD.n253 VDD.n252 4.65
R402 VDD.n258 VDD.n257 4.65
R403 VDD.n262 VDD.n261 4.65
R404 VDD.n288 VDD.n287 4.65
R405 VDD.n292 VDD.n291 4.65
R406 VDD.n296 VDD.n295 4.65
R407 VDD.n300 VDD.n299 4.65
R408 VDD.n306 VDD.n305 4.65
R409 VDD.n310 VDD.n309 4.65
R410 VDD.n314 VDD.n313 4.65
R411 VDD.n320 VDD.n319 4.65
R412 VDD.n324 VDD.n323 4.65
R413 VDD.n329 VDD.n328 4.65
R414 VDD.n333 VDD.n332 4.65
R415 VDD.n337 VDD.n336 4.65
R416 VDD.n364 VDD.n363 4.65
R417 VDD.n368 VDD.n367 4.65
R418 VDD.n372 VDD.n371 4.65
R419 VDD.n376 VDD.n375 4.65
R420 VDD.n382 VDD.n381 4.65
R421 VDD.n386 VDD.n385 4.65
R422 VDD.n390 VDD.n389 4.65
R423 VDD.n396 VDD.n395 4.65
R424 VDD.n400 VDD.n399 4.65
R425 VDD.n405 VDD.n404 4.65
R426 VDD.n409 VDD.n408 4.65
R427 VDD.n432 VDD.n431 4.65
R428 VDD.n28 VDD.n23 2.933
R429 VDD.n49 VDD.n46 2.89
R430 VDD.n257 VDD.n254 2.89
R431 VDD.n28 VDD.n27 2.844
R432 VDD.n38 �[R. 2.557
R433 VDD.n246 VDD.t48 2.557
R434 VDD.n27 VDD.n24 2.477
R435 VDD.n235 VDD.n232 2.477
R436 VDD.n32 VDD.n28 1.063
R437 VDD.n121 VDD.n118 0.412
R438 VDD.n196 VDD.n193 0.412
R439 VDD.n328 VDD.n325 0.412
R440 VDD.n404 VDD.n401 0.412
R441 VDD.n81 VDD.n54 0.29
R442 VDD.n156 VDD.n130 0.29
R443 VDD.n231 VDD.n205 0.29
R444 VDD.n288 VDD.n262 0.29
R445 VDD.n364 VDD.n337 0.29
R446 VDD.n107 VDD.n103 0.197
R447 VDD.n182 VDD.n178 0.197
R448 VDD.n314 VDD.n310 0.197
R449 VDD.n390 VDD.n386 0.197
R450 VDD.n41 VDD.n37 0.181
R451 VDD.n249 VDD.n245 0.181
R452 VDD.n37 VDD.n32 0.145
R453 VDD.n45 VDD.n41 0.145
R454 VDD.n50 VDD.n45 0.145
R455 VDD.n54 VDD.n50 0.145
R456 VDD.n85 VDD.n81 0.145
R457 VDD.n89 VDD.n85 0.145
R458 VDD.n93 VDD.n89 0.145
R459 VDD.n99 VDD.n93 0.145
R460 VDD.n103 VDD.n99 0.145
R461 VDD.n113 VDD.n107 0.145
R462 VDD.n117 VDD.n113 0.145
R463 VDD.n122 VDD.n117 0.145
R464 VDD.n126 VDD.n122 0.145
R465 VDD.n130 VDD.n126 0.145
R466 VDD.n160 VDD.n156 0.145
R467 VDD.n164 VDD.n160 0.145
R468 VDD.n168 VDD.n164 0.145
R469 VDD.n174 VDD.n168 0.145
R470 VDD.n178 VDD.n174 0.145
R471 VDD.n188 VDD.n182 0.145
R472 VDD.n192 VDD.n188 0.145
R473 VDD.n197 VDD.n192 0.145
R474 VDD.n201 VDD.n197 0.145
R475 VDD.n205 VDD.n201 0.145
R476 VDD.n236 VDD.n231 0.145
R477 VDD.n240 VDD.n236 0.145
R478 VDD.n245 VDD.n240 0.145
R479 VDD.n253 VDD.n249 0.145
R480 VDD.n258 VDD.n253 0.145
R481 VDD.n262 VDD.n258 0.145
R482 VDD.n292 VDD.n288 0.145
R483 VDD.n296 VDD.n292 0.145
R484 VDD.n300 VDD.n296 0.145
R485 VDD.n306 VDD.n300 0.145
R486 VDD.n310 VDD.n306 0.145
R487 VDD.n320 VDD.n314 0.145
R488 VDD.n324 VDD.n320 0.145
R489 VDD.n329 VDD.n324 0.145
R490 VDD.n333 VDD.n329 0.145
R491 VDD.n337 VDD.n333 0.145
R492 VDD.n368 VDD.n364 0.145
R493 VDD.n372 VDD.n368 0.145
R494 VDD.n376 VDD.n372 0.145
R495 VDD.n382 VDD.n376 0.145
R496 VDD.n386 VDD.n382 0.145
R497 VDD.n396 VDD.n390 0.145
R498 VDD.n400 VDD.n396 0.145
R499 VDD.n405 VDD.n400 0.145
R500 VDD.n409 VDD.n405 0.145
R501 VDD.n432 VDD.n409 0.145
R502 VDD.n432 VDD 0.034
R503 a_599_989.n1 a_599_989.t7 480.392
R504 a_599_989.n3 a_599_989.t11 454.685
R505 a_599_989.n3 a_599_989.t8 428.979
R506 a_599_989.n1 a_599_989.t10 403.272
R507 a_599_989.n2 a_599_989.t12 357.204
R508 a_599_989.n4 a_599_989.t9 311.683
R509 a_599_989.n10 a_599_989.n9 308.216
R510 a_599_989.n11 a_599_989.n10 179.199
R511 a_599_989.n4 a_599_989.n3 171.288
R512 a_599_989.n2 a_599_989.n1 171.288
R513 a_599_989.n13 a_599_989.n12 161.352
R514 a_599_989.n11 a_599_989.n0 95.095
R515 a_599_989.n14 a_599_989.n13 95.094
R516 a_599_989.n13 a_599_989.n11 66.258
R517 a_599_989.n9 a_599_989.n8 30
R518 a_599_989.n7 a_599_989.n6 24.383
R519 a_599_989.n9 a_599_989.n7 23.684
R520 a_599_989.n0 a_599_989.t5 14.282
R521 a_599_989.n0 a_599_989.t0 14.282
R522 a_599_989.n12 a_599_989.t3 14.282
R523 a_599_989.n12 a_599_989.t6 14.282
R524 a_599_989.n14 a_599_989.t1 14.282
R525 a_599_989.t2 a_599_989.n14 14.282
R526 a_599_989.n5 a_599_989.n4 8.685
R527 a_599_989.n5 a_599_989.n2 5.965
R528 a_599_989.n10 a_599_989.n5 4.65
R529 CLK.n2 CLK.t0 459.505
R530 CLK.n0 CLK.t4 459.505
R531 CLK.n3 CLK.t3 399.181
R532 CLK.n1 CLK.t5 399.181
R533 CLK.n2 CLK.t2 384.527
R534 CLK.n0 CLK.t1 384.527
R535 CLK.n3 CLK.n2 33.832
R536 CLK.n1 CLK.n0 33.832
R537 CLK.n4 CLK.n1 11.555
R538 CLK.n4 CLK.n3 2.079
R539 CLK.n4 CLK 0.046
R540 a_277_1050.n2 a_277_1050.t8 512.525
R541 a_277_1050.n0 a_277_1050.t7 512.525
R542 a_277_1050.n3 a_277_1050.t12 389.251
R543 a_277_1050.n1 a_277_1050.t11 389.251
R544 a_277_1050.n2 a_277_1050.t10 371.139
R545 a_277_1050.n0 a_277_1050.t9 371.139
R546 a_277_1050.n9 a_277_1050.n8 336.075
R547 a_277_1050.n3 a_277_1050.n2 207.695
R548 a_277_1050.n1 a_277_1050.n0 207.695
R549 a_277_1050.n12 a_277_1050.n11 161.352
R550 a_277_1050.n13 a_277_1050.n9 151.34
R551 a_277_1050.n12 a_277_1050.n10 95.095
R552 a_277_1050.n14 a_277_1050.n13 95.094
R553 a_277_1050.n13 a_277_1050.n12 66.258
R554 a_277_1050.n8 a_277_1050.n7 30
R555 a_277_1050.n6 a_277_1050.n5 24.383
R556 a_277_1050.n8 a_277_1050.n6 23.684
R557 a_277_1050.n10 a_277_1050.t5 14.282
R558 a_277_1050.n10 a_277_1050.t4 14.282
R559 a_277_1050.n11 a_277_1050.t6 14.282
R560 a_277_1050.n11 a_277_1050.t0 14.282
R561 a_277_1050.t2 a_277_1050.n14 14.282
R562 a_277_1050.n14 a_277_1050.t1 14.282
R563 a_277_1050.n4 a_277_1050.n1 14.126
R564 a_277_1050.n9 a_277_1050.n4 5.965
R565 a_277_1050.n4 a_277_1050.n3 4.65
R566 a_2141_1050.n1 a_2141_1050.t5 512.525
R567 a_2141_1050.n1 a_2141_1050.t6 371.139
R568 a_2141_1050.n2 a_2141_1050.t7 361.392
R569 a_2141_1050.n4 a_2141_1050.n3 327.32
R570 a_2141_1050.n2 a_2141_1050.n1 235.554
R571 a_2141_1050.n5 a_2141_1050.n4 159.999
R572 a_2141_1050.n6 a_2141_1050.n5 157.963
R573 a_2141_1050.n5 a_2141_1050.n0 91.706
R574 a_2141_1050.n0 a_2141_1050.t1 14.282
R575 a_2141_1050.n0 a_2141_1050.t0 14.282
R576 a_2141_1050.t3 a_2141_1050.n6 14.282
R577 a_2141_1050.n6 a_2141_1050.t2 14.282
R578 a_2141_1050.n4 a_2141_1050.n2 10.615
R579 a_3829_1050.n2 a_3829_1050.t9 480.392
R580 a_3829_1050.n2 a_3829_1050.t7 403.272
R581 a_3829_1050.n3 a_3829_1050.t8 357.204
R582 a_3829_1050.n5 a_3829_1050.n4 329.955
R583 a_3829_1050.n6 a_3829_1050.n5 179.199
R584 a_3829_1050.n3 a_3829_1050.n2 171.288
R585 a_3829_1050.n8 a_3829_1050.n7 161.352
R586 a_3829_1050.n6 a_3829_1050.n1 95.095
R587 a_3829_1050.n7 a_3829_1050.n0 95.095
R588 a_3829_1050.n7 a_3829_1050.n6 66.258
R589 a_3829_1050.n1 a_3829_1050.t3 14.282
R590 a_3829_1050.n1 a_3829_1050.t4 14.282
R591 a_3829_1050.n0 a_3829_1050.t6 14.282
R592 a_3829_1050.n0 a_3829_1050.t5 14.282
R593 a_3829_1050.t2 a_3829_1050.n8 14.282
R594 a_3829_1050.n8 a_3829_1050.t1 14.282
R595 a_3829_1050.n5 a_3829_1050.n3 10.615
R596 a_1053_103.t0 a_1053_103.n3 117.777
R597 a_1053_103.n6 a_1053_103.n4 55.785
R598 a_1053_103.n6 a_1053_103.n5 51.696
R599 a_1053_103.t0 a_1053_103.n6 39.361
R600 a_1053_103.n2 a_1053_103.n0 32.662
R601 a_1053_103.t0 a_1053_103.n2 3.034
R602 a_1053_103.n2 a_1053_103.n1 0.443
R603 a_1334_210.n10 a_1334_210.n8 171.558
R604 a_1334_210.n8 a_1334_210.t1 75.764
R605 a_1334_210.n11 a_1334_210.n0 49.6
R606 a_1334_210.n3 a_1334_210.n2 27.476
R607 a_1334_210.n10 a_1334_210.n9 27.2
R608 a_1334_210.n11 a_1334_210.n10 22.4
R609 a_1334_210.t1 a_1334_210.n5 20.241
R610 a_1334_210.n7 a_1334_210.n6 19.952
R611 a_1334_210.t1 a_1334_210.n3 13.984
R612 a_1334_210.n5 a_1334_210.n4 13.494
R613 a_1334_210.t1 a_1334_210.n1 7.04
R614 a_1334_210.n8 a_1334_210.n7 1.505
R615 VSS.n196 VSS.n195 237.558
R616 VSS.n154 VSS.n153 237.558
R617 VSS.n121 VSS.n120 237.558
R618 VSS.n76 VSS.n75 237.558
R619 VSS.n31 VSS.n30 237.558
R620 VSS.n28 VSS.n27 210.82
R621 VSS.n193 VSS.n192 210.82
R622 VSS.n151 VSS.n150 210.82
R623 VSS.n118 VSS.n117 210.82
R624 VSS.n73 VSS.n72 210.82
R625 VSS.n183 VSS.n182 173.365
R626 VSS.n225 VSS.n224 173.365
R627 VSS.n63 VSS.n62 152.358
R628 VSS.n108 VSS.n107 152.358
R629 VSS.n17 VSS.n16 151.605
R630 VSS.n140 VSS.n139 151.605
R631 VSS.n16 VSS.n15 28.421
R632 VSS.n62 VSS.n61 28.421
R633 VSS.n107 VSS.n106 28.421
R634 VSS.n139 VSS.n138 28.421
R635 VSS.n16 VSS.n14 25.263
R636 VSS.n62 VSS.n60 25.263
R637 VSS.n107 VSS.n105 25.263
R638 VSS.n139 VSS.n137 25.263
R639 VSS.n14 VSS.n13 24.383
R640 VSS.n60 VSS.n59 24.383
R641 VSS.n105 VSS.n104 24.383
R642 VSS.n137 VSS.n136 24.383
R643 VSS.n29 VSS.n28 18.953
R644 VSS.n194 VSS.n193 18.953
R645 VSS.n152 VSS.n151 18.953
R646 VSS.n119 VSS.n118 18.953
R647 VSS.n74 VSS.n73 18.953
R648 VSS.n32 VSS.n29 14.864
R649 VSS.n77 VSS.n74 14.864
R650 VSS.n122 VSS.n119 14.864
R651 VSS.n155 VSS.n152 14.864
R652 VSS.n197 VSS.n194 14.864
R653 VSS.n229 VSS.n228 9.154
R654 VSS.n226 VSS.n223 9.154
R655 VSS.n221 VSS.n220 9.154
R656 VSS.n218 VSS.n217 9.154
R657 VSS.n215 VSS.n214 9.154
R658 VSS.n212 VSS.n211 9.154
R659 VSS.n209 VSS.n208 9.154
R660 VSS.n206 VSS.n205 9.154
R661 VSS.n203 VSS.n202 9.154
R662 VSS.n200 VSS.n199 9.154
R663 VSS.n197 VSS.n196 9.154
R664 VSS.n190 VSS.n189 9.154
R665 VSS.n187 VSS.n186 9.154
R666 VSS.n184 VSS.n181 9.154
R667 VSS.n179 VSS.n178 9.154
R668 VSS.n176 VSS.n175 9.154
R669 VSS.n173 VSS.n172 9.154
R670 VSS.n170 VSS.n169 9.154
R671 VSS.n167 VSS.n166 9.154
R672 VSS.n164 VSS.n163 9.154
R673 VSS.n161 VSS.n160 9.154
R674 VSS.n158 VSS.n157 9.154
R675 VSS.n155 VSS.n154 9.154
R676 VSS.n148 VSS.n147 9.154
R677 VSS.n145 VSS.n144 9.154
R678 VSS.n142 VSS.n141 9.154
R679 VSS.n134 VSS.n133 9.154
R680 VSS.n131 VSS.n130 9.154
R681 VSS.n128 VSS.n127 9.154
R682 VSS.n125 VSS.n124 9.154
R683 VSS.n122 VSS.n121 9.154
R684 VSS.n115 VSS.n114 9.154
R685 VSS.n112 VSS.n111 9.154
R686 VSS.n109 VSS.n103 9.154
R687 VSS.n101 VSS.n100 9.154
R688 VSS.n98 VSS.n97 9.154
R689 VSS.n95 VSS.n94 9.154
R690 VSS.n92 VSS.n91 9.154
R691 VSS.n89 VSS.n88 9.154
R692 VSS.n86 VSS.n85 9.154
R693 VSS.n83 VSS.n82 9.154
R694 VSS.n80 VSS.n79 9.154
R695 VSS.n77 VSS.n76 9.154
R696 VSS.n70 VSS.n69 9.154
R697 VSS.n67 VSS.n66 9.154
R698 VSS.n64 VSS.n58 9.154
R699 VSS.n56 VSS.n55 9.154
R700 VSS.n53 VSS.n52 9.154
R701 VSS.n50 VSS.n49 9.154
R702 VSS.n47 VSS.n46 9.154
R703 VSS.n44 VSS.n43 9.154
R704 VSS.n41 VSS.n40 9.154
R705 VSS.n38 VSS.n37 9.154
R706 VSS.n35 VSS.n34 9.154
R707 VSS.n32 VSS.n31 9.154
R708 VSS.n25 VSS.n24 9.154
R709 VSS.n22 VSS.n21 9.154
R710 VSS.n19 VSS.n18 9.154
R711 VSS.n11 VSS.n10 9.154
R712 VSS.n8 VSS.n7 9.154
R713 VSS.n5 VSS.n4 9.154
R714 VSS.n2 VSS.n1 9.154
R715 VSS.n233 VSS.n232 4.65
R716 VSS.n6 VSS.n5 4.65
R717 VSS.n9 VSS.n8 4.65
R718 VSS.n12 VSS.n11 4.65
R719 VSS.n20 VSS.n19 4.65
R720 VSS.n23 VSS.n22 4.65
R721 VSS.n26 VSS.n25 4.65
R722 VSS.n33 VSS.n32 4.65
R723 VSS.n36 VSS.n35 4.65
R724 VSS.n39 VSS.n38 4.65
R725 VSS.n42 VSS.n41 4.65
R726 VSS.n45 VSS.n44 4.65
R727 VSS.n48 VSS.n47 4.65
R728 VSS.n51 VSS.n50 4.65
R729 VSS.n54 VSS.n53 4.65
R730 VSS.n57 VSS.n56 4.65
R731 VSS.n65 VSS.n64 4.65
R732 VSS.n68 VSS.n67 4.65
R733 VSS.n71 VSS.n70 4.65
R734 VSS.n78 VSS.n77 4.65
R735 VSS.n81 VSS.n80 4.65
R736 VSS.n84 VSS.n83 4.65
R737 VSS.n87 VSS.n86 4.65
R738 VSS.n90 VSS.n89 4.65
R739 VSS.n93 VSS.n92 4.65
R740 VSS.n96 VSS.n95 4.65
R741 VSS.n99 VSS.n98 4.65
R742 VSS.n102 VSS.n101 4.65
R743 VSS.n110 VSS.n109 4.65
R744 VSS.n113 VSS.n112 4.65
R745 VSS.n116 VSS.n115 4.65
R746 VSS.n123 VSS.n122 4.65
R747 VSS.n126 VSS.n125 4.65
R748 VSS.n129 VSS.n128 4.65
R749 VSS.n132 VSS.n131 4.65
R750 VSS.n135 VSS.n134 4.65
R751 VSS.n143 VSS.n142 4.65
R752 VSS.n146 VSS.n145 4.65
R753 VSS.n149 VSS.n148 4.65
R754 VSS.n156 VSS.n155 4.65
R755 VSS.n159 VSS.n158 4.65
R756 VSS.n162 VSS.n161 4.65
R757 VSS.n165 VSS.n164 4.65
R758 VSS.n168 VSS.n167 4.65
R759 VSS.n171 VSS.n170 4.65
R760 VSS.n174 VSS.n173 4.65
R761 VSS.n177 VSS.n176 4.65
R762 VSS.n180 VSS.n179 4.65
R763 VSS.n185 VSS.n184 4.65
R764 VSS.n188 VSS.n187 4.65
R765 VSS.n191 VSS.n190 4.65
R766 VSS.n198 VSS.n197 4.65
R767 VSS.n201 VSS.n200 4.65
R768 VSS.n204 VSS.n203 4.65
R769 VSS.n207 VSS.n206 4.65
R770 VSS.n210 VSS.n209 4.65
R771 VSS.n213 VSS.n212 4.65
R772 VSS.n216 VSS.n215 4.65
R773 VSS.n219 VSS.n218 4.65
R774 VSS.n222 VSS.n221 4.65
R775 VSS.n227 VSS.n226 4.65
R776 VSS.n230 VSS.n229 4.65
R777 VSS.n19 VSS.n17 4.129
R778 VSS.n142 VSS.n140 4.129
R779 VSS.n3 VSS.n0 3.407
R780 VSS.n3 VSS.n2 2.844
R781 VSS.n6 VSS.n3 1.063
R782 VSS.n232 VSS.n231 0.474
R783 VSS.n33 VSS.n26 0.29
R784 VSS.n78 VSS.n71 0.29
R785 VSS.n123 VSS.n116 0.29
R786 VSS.n156 VSS.n149 0.29
R787 VSS.n198 VSS.n191 0.29
R788 VSS.n64 VSS.n63 0.206
R789 VSS.n109 VSS.n108 0.206
R790 VSS.n184 VSS.n183 0.206
R791 VSS.n226 VSS.n225 0.206
R792 VSS.n51 VSS.n48 0.197
R793 VSS.n96 VSS.n93 0.197
R794 VSS.n174 VSS.n171 0.197
R795 VSS.n216 VSS.n213 0.197
R796 VSS.n12 VSS.n9 0.181
R797 VSS.n135 VSS.n132 0.181
R798 VSS.n9 VSS.n6 0.145
R799 VSS.n20 VSS.n12 0.145
R800 VSS.n23 VSS.n20 0.145
R801 VSS.n26 VSS.n23 0.145
R802 VSS.n36 VSS.n33 0.145
R803 VSS.n39 VSS.n36 0.145
R804 VSS.n42 VSS.n39 0.145
R805 VSS.n45 VSS.n42 0.145
R806 VSS.n48 VSS.n45 0.145
R807 VSS.n54 VSS.n51 0.145
R808 VSS.n57 VSS.n54 0.145
R809 VSS.n65 VSS.n57 0.145
R810 VSS.n68 VSS.n65 0.145
R811 VSS.n71 VSS.n68 0.145
R812 VSS.n81 VSS.n78 0.145
R813 VSS.n84 VSS.n81 0.145
R814 VSS.n87 VSS.n84 0.145
R815 VSS.n90 VSS.n87 0.145
R816 VSS.n93 VSS.n90 0.145
R817 VSS.n99 VSS.n96 0.145
R818 VSS.n102 VSS.n99 0.145
R819 VSS.n110 VSS.n102 0.145
R820 VSS.n113 VSS.n110 0.145
R821 VSS.n116 VSS.n113 0.145
R822 VSS.n126 VSS.n123 0.145
R823 VSS.n129 VSS.n126 0.145
R824 VSS.n132 VSS.n129 0.145
R825 VSS.n143 VSS.n135 0.145
R826 VSS.n146 VSS.n143 0.145
R827 VSS.n149 VSS.n146 0.145
R828 VSS.n159 VSS.n156 0.145
R829 VSS.n162 VSS.n159 0.145
R830 VSS.n165 VSS.n162 0.145
R831 VSS.n168 VSS.n165 0.145
R832 VSS.n171 VSS.n168 0.145
R833 VSS.n177 VSS.n174 0.145
R834 VSS.n180 VSS.n177 0.145
R835 VSS.n185 VSS.n180 0.145
R836 VSS.n188 VSS.n185 0.145
R837 VSS.n191 VSS.n188 0.145
R838 VSS.n201 VSS.n198 0.145
R839 VSS.n204 VSS.n201 0.145
R840 VSS.n207 VSS.n204 0.145
R841 VSS.n210 VSS.n207 0.145
R842 VSS.n213 VSS.n210 0.145
R843 VSS.n219 VSS.n216 0.145
R844 VSS.n222 VSS.n219 0.145
R845 VSS.n227 VSS.n222 0.145
R846 VSS.n230 VSS.n227 0.145
R847 VSS.n233 VSS.n230 0.145
R848 VSS.n233 VSS 0.034
R849 a_147_187.n6 a_147_187.t15 512.525
R850 a_147_187.n4 a_147_187.t9 472.359
R851 a_147_187.n2 a_147_187.t14 472.359
R852 a_147_187.n7 a_147_187.t12 417.109
R853 a_147_187.n4 a_147_187.t13 384.527
R854 a_147_187.n2 a_147_187.t10 384.527
R855 a_147_187.n13 a_147_187.n12 379.457
R856 a_147_187.n6 a_147_187.t11 371.139
R857 a_147_187.n5 a_147_187.t8 370.613
R858 a_147_187.n3 a_147_187.t7 370.613
R859 a_147_187.n7 a_147_187.n6 179.837
R860 a_147_187.n16 a_147_187.n15 161.352
R861 a_147_187.n5 a_147_187.n4 127.096
R862 a_147_187.n3 a_147_187.n2 127.096
R863 a_147_187.n14 a_147_187.n13 123.481
R864 a_147_187.n14 a_147_187.n1 95.095
R865 a_147_187.n15 a_147_187.n0 95.095
R866 a_147_187.n15 a_147_187.n14 66.258
R867 a_147_187.n12 a_147_187.n11 22.578
R868 a_147_187.n1 a_147_187.t6 14.282
R869 a_147_187.n1 a_147_187.t4 14.282
R870 a_147_187.n0 a_147_187.t2 14.282
R871 a_147_187.n0 a_147_187.t3 14.282
R872 a_147_187.t1 a_147_187.n16 14.282
R873 a_147_187.n16 a_147_187.t0 14.282
R874 a_147_187.n8 a_147_187.n7 12.222
R875 a_147_187.n9 a_147_187.n3 10.046
R876 a_147_187.n12 a_147_187.n10 8.58
R877 a_147_187.n8 a_147_187.n5 4.65
R878 a_147_187.n13 a_147_187.n9 4.65
R879 a_147_187.n9 a_147_187.n8 4.035
R880 a_4626_101.n3 a_4626_101.n1 42.788
R881 a_4626_101.t0 a_4626_101.n0 8.137
R882 a_4626_101.n3 a_4626_101.n2 4.665
R883 a_4626_101.t0 a_4626_101.n3 0.06
R884 Q.n5 Q.t5 454.685
R885 Q.n5 Q.t6 428.979
R886 Q.n4 Q.n3 355.179
R887 Q.n6 Q.t7 339.542
R888 Q.n2 Q.n1 157.964
R889 Q.n6 Q.n5 143.429
R890 Q.n4 Q.n2 132.141
R891 Q.n2 Q.n0 91.706
R892 Q.n0 Q.t0 14.282
R893 Q.n0 Q.t1 14.282
R894 Q.n1 Q.t3 14.282
R895 Q.n1 Q.t4 14.282
R896 Q Q.n6 7.551
R897 Q.n7 Q.n4 4.65
R898 Q.n7 Q 0.046
R899 a_2036_101.n11 a_2036_101.n10 68.43
R900 a_2036_101.n3 a_2036_101.n2 62.817
R901 a_2036_101.n7 a_2036_101.n6 38.626
R902 a_2036_101.n6 a_2036_101.n5 35.955
R903 a_2036_101.n3 a_2036_101.n1 26.202
R904 a_2036_101.t0 a_2036_101.n3 19.737
R905 a_2036_101.t1 a_2036_101.n8 8.137
R906 a_2036_101.t0 a_2036_101.n4 7.273
R907 a_2036_101.t0 a_2036_101.n0 6.109
R908 a_2036_101.t1 a_2036_101.n7 4.864
R909 a_2036_101.t0 a_2036_101.n12 2.074
R910 a_2036_101.n12 a_2036_101.t1 0.937
R911 a_2036_101.t1 a_2036_101.n11 0.763
R912 a_2036_101.n11 a_2036_101.n9 0.185
R913 RN.n0 RN.t4 479.223
R914 RN.n5 RN.t0 454.685
R915 RN.n2 RN.t1 454.685
R916 RN.n5 RN.t3 428.979
R917 RN.n2 RN.t8 428.979
R918 RN.n0 RN.t5 375.52
R919 RN.n6 RN.n5 254.865
R920 RN.n3 RN.n2 254.865
R921 RN.n1 RN.n0 252.188
R922 RN.n1 RN.t7 231.854
R923 RN.n6 RN.t6 228.106
R924 RN.n3 RN.t2 228.106
R925 RN.n4 RN.n1 7.325
R926 RN.n7 RN.n4 5.94
R927 RN.n4 RN.n3 4.65
R928 RN.n7 RN.n6 4.65
R929 RN.n7 RN 0.046
R930 a_372_210.n9 a_372_210.n7 171.558
R931 a_372_210.t0 a_372_210.n9 75.765
R932 a_372_210.n3 a_372_210.n1 74.827
R933 a_372_210.n3 a_372_210.n2 27.476
R934 a_372_210.n7 a_372_210.n6 27.2
R935 a_372_210.n5 a_372_210.n4 23.498
R936 a_372_210.n7 a_372_210.n5 22.4
R937 a_372_210.t0 a_372_210.n11 20.241
R938 a_372_210.t0 a_372_210.n3 13.984
R939 a_372_210.n11 a_372_210.n10 13.494
R940 a_372_210.t0 a_372_210.n0 8.137
R941 a_372_210.n9 a_372_210.n8 1.505
R942 a_2962_210.n9 a_2962_210.n7 171.558
R943 a_2962_210.t0 a_2962_210.n9 75.765
R944 a_2962_210.n3 a_2962_210.n1 74.827
R945 a_2962_210.n3 a_2962_210.n2 27.476
R946 a_2962_210.n7 a_2962_210.n6 27.2
R947 a_2962_210.n5 a_2962_210.n4 23.498
R948 a_2962_210.n7 a_2962_210.n5 22.4
R949 a_2962_210.t0 a_2962_210.n11 20.241
R950 a_2962_210.t0 a_2962_210.n3 13.984
R951 a_2962_210.n11 a_2962_210.n10 13.494
R952 a_2962_210.t0 a_2962_210.n0 8.137
R953 a_2962_210.n9 a_2962_210.n8 1.505
R954 a_91_103.t0 a_91_103.n7 59.616
R955 a_91_103.n4 a_91_103.n2 54.496
R956 a_91_103.n4 a_91_103.n3 54.496
R957 a_91_103.n1 a_91_103.n0 24.679
R958 a_91_103.t0 a_91_103.n1 7.505
R959 a_91_103.n6 a_91_103.n5 2.455
R960 a_91_103.n6 a_91_103.n4 0.636
R961 a_91_103.t0 a_91_103.n6 0.246
R962 a_3924_210.n9 a_3924_210.n7 171.558
R963 a_3924_210.t0 a_3924_210.n9 75.765
R964 a_3924_210.n3 a_3924_210.n1 74.827
R965 a_3924_210.n3 a_3924_210.n2 27.476
R966 a_3924_210.n7 a_3924_210.n6 27.2
R967 a_3924_210.n5 a_3924_210.n4 23.498
R968 a_3924_210.n7 a_3924_210.n5 22.4
R969 a_3924_210.t0 a_3924_210.n11 20.241
R970 a_3924_210.t0 a_3924_210.n3 13.984
R971 a_3924_210.n11 a_3924_210.n10 13.494
R972 a_3924_210.t0 a_3924_210.n0 8.137
R973 a_3924_210.n9 a_3924_210.n8 1.505
R974 a_3643_103.t0 a_3643_103.n7 59.616
R975 a_3643_103.n4 a_3643_103.n2 54.496
R976 a_3643_103.n4 a_3643_103.n3 54.496
R977 a_3643_103.n1 a_3643_103.n0 24.679
R978 a_3643_103.t0 a_3643_103.n1 7.505
R979 a_3643_103.n6 a_3643_103.n5 2.455
R980 a_3643_103.n6 a_3643_103.n4 0.636
R981 a_3643_103.t0 a_3643_103.n6 0.246
R982 a_2681_103.n5 a_2681_103.n4 66.708
R983 a_2681_103.n2 a_2681_103.n0 25.439
R984 a_2681_103.n5 a_2681_103.n3 19.496
R985 a_2681_103.t0 a_2681_103.n5 13.756
R986 a_2681_103.n2 a_2681_103.n1 2.455
R987 a_2681_103.t0 a_2681_103.n2 0.246
C8 RN VSS 1.72fF
C9 VDD VSS 8.54fF
C10 a_2681_103.n0 VSS 0.11fF
C11 a_2681_103.n1 VSS 0.04fF
C12 a_2681_103.n2 VSS 0.03fF
C13 a_2681_103.n3 VSS 0.07fF
C14 a_2681_103.n4 VSS 0.08fF
C15 a_2681_103.n5 VSS 0.03fF
C16 a_3643_103.n0 VSS 0.08fF
C17 a_3643_103.n1 VSS 0.07fF
C18 a_3643_103.n2 VSS 0.04fF
C19 a_3643_103.n3 VSS 0.06fF
C20 a_3643_103.n4 VSS 0.03fF
C21 a_3643_103.n5 VSS 0.04fF
C22 a_3643_103.n7 VSS 0.08fF
C23 a_3924_210.n0 VSS 0.07fF
C24 a_3924_210.n1 VSS 0.09fF
C25 a_3924_210.n2 VSS 0.12fF
C26 a_3924_210.n3 VSS 0.08fF
C27 a_3924_210.n4 VSS 0.02fF
C28 a_3924_210.n5 VSS 0.03fF
C29 a_3924_210.n6 VSS 0.02fF
C30 a_3924_210.n7 VSS 0.03fF
C31 a_3924_210.n8 VSS 0.02fF
C32 a_3924_210.n9 VSS 0.13fF
C33 a_3924_210.n10 VSS 0.08fF
C34 a_3924_210.n11 VSS 0.02fF
C35 a_3924_210.t0 VSS 0.31fF
C36 a_91_103.n0 VSS 0.08fF
C37 a_91_103.n1 VSS 0.07fF
C38 a_91_103.n2 VSS 0.04fF
C39 a_91_103.n3 VSS 0.06fF
C40 a_91_103.n4 VSS 0.03fF
C41 a_91_103.n5 VSS 0.03fF
C42 a_91_103.n7 VSS 0.08fF
C43 a_2962_210.n0 VSS 0.07fF
C44 a_2962_210.n1 VSS 0.09fF
C45 a_2962_210.n2 VSS 0.12fF
C46 a_2962_210.n3 VSS 0.08fF
C47 a_2962_210.n4 VSS 0.02fF
C48 a_2962_210.n5 VSS 0.03fF
C49 a_2962_210.n6 VSS 0.02fF
C50 a_2962_210.n7 VSS 0.03fF
C51 a_2962_210.n8 VSS 0.02fF
C52 a_2962_210.n9 VSS 0.13fF
C53 a_2962_210.n10 VSS 0.08fF
C54 a_2962_210.n11 VSS 0.02fF
C55 a_2962_210.t0 VSS 0.31fF
C56 a_372_210.n0 VSS 0.07fF
C57 a_372_210.n1 VSS 0.09fF
C58 a_372_210.n2 VSS 0.12fF
C59 a_372_210.n3 VSS 0.08fF
C60 a_372_210.n4 VSS 0.02fF
C61 a_372_210.n5 VSS 0.03fF
C62 a_372_210.n6 VSS 0.02fF
C63 a_372_210.n7 VSS 0.03fF
C64 a_372_210.n8 VSS 0.02fF
C65 a_372_210.n9 VSS 0.13fF
C66 a_372_210.n10 VSS 0.08fF
C67 a_372_210.n11 VSS 0.02fF
C68 a_372_210.t0 VSS 0.31fF
C69 RN.n0 VSS 0.33fF
C70 RN.t7 VSS 0.36fF
C71 RN.n1 VSS 0.40fF
C72 RN.n2 VSS 0.32fF
C73 RN.t2 VSS 0.36fF
C74 RN.n3 VSS 0.30fF
C75 RN.n4 VSS 0.92fF
C76 RN.n5 VSS 0.32fF
C77 RN.t6 VSS 0.37fF
C78 RN.n6 VSS 0.30fF
C79 RN.n7 VSS 0.53fF
C80 a_2036_101.n0 VSS 0.02fF
C81 a_2036_101.n1 VSS 0.09fF
C82 a_2036_101.n2 VSS 0.08fF
C83 a_2036_101.n3 VSS 0.03fF
C84 a_2036_101.n4 VSS 0.01fF
C85 a_2036_101.n5 VSS 0.04fF
C86 a_2036_101.n6 VSS 0.04fF
C87 a_2036_101.n7 VSS 0.02fF
C88 a_2036_101.n8 VSS 0.05fF
C89 a_2036_101.n9 VSS 0.15fF
C90 a_2036_101.n10 VSS 0.08fF
C91 a_2036_101.n11 VSS 0.08fF
C92 a_2036_101.t1 VSS 0.23fF
C93 a_2036_101.n12 VSS 0.01fF
C94 Q.n0 VSS 0.38fF
C95 Q.n1 VSS 0.48fF
C96 Q.n2 VSS 0.54fF
C97 Q.n3 VSS 0.36fF
C98 Q.n4 VSS 0.51fF
C99 Q.n5 VSS 0.30fF
C100 Q.t7 VSS 0.54fF
C101 Q.n6 VSS 0.54fF
C102 Q.n7 VSS 0.03fF
C103 a_4626_101.n0 VSS 0.05fF
C104 a_4626_101.n1 VSS 0.12fF
C105 a_4626_101.n2 VSS 0.04fF
C106 a_4626_101.n3 VSS 0.16fF
C107 a_147_187.n0 VSS 0.58fF
C108 a_147_187.n1 VSS 0.58fF
C109 a_147_187.n2 VSS 0.41fF
C110 a_147_187.n3 VSS 1.08fF
C111 a_147_187.n4 VSS 0.41fF
C112 a_147_187.t8 VSS 0.86fF
C113 a_147_187.n5 VSS 0.58fF
C114 a_147_187.n6 VSS 0.42fF
C115 a_147_187.n7 VSS 1.51fF
C116 a_147_187.n8 VSS 2.43fF
C117 a_147_187.n9 VSS 2.02fF
C118 a_147_187.n10 VSS 0.06fF
C119 a_147_187.n11 VSS 0.08fF
C120 a_147_187.n12 VSS 0.45fF
C121 a_147_187.n13 VSS 0.80fF
C122 a_147_187.n14 VSS 0.58fF
C123 a_147_187.n15 VSS 0.70fF
C124 a_147_187.n16 VSS 0.74fF
C125 a_1334_210.n0 VSS 0.02fF
C126 a_1334_210.n1 VSS 0.09fF
C127 a_1334_210.n2 VSS 0.12fF
C128 a_1334_210.n3 VSS 0.08fF
C129 a_1334_210.n4 VSS 0.08fF
C130 a_1334_210.n5 VSS 0.02fF
C131 a_1334_210.t1 VSS 0.29fF
C132 a_1334_210.n6 VSS 0.09fF
C133 a_1334_210.n7 VSS 0.02fF
C134 a_1334_210.n8 VSS 0.13fF
C135 a_1334_210.n9 VSS 0.02fF
C136 a_1334_210.n10 VSS 0.03fF
C137 a_1334_210.n11 VSS 0.02fF
C138 a_1053_103.n0 VSS 0.13fF
C139 a_1053_103.n1 VSS 0.04fF
C140 a_1053_103.n2 VSS 0.09fF
C141 a_1053_103.n3 VSS 0.03fF
C142 a_1053_103.n4 VSS 0.08fF
C143 a_1053_103.n5 VSS 0.07fF
C144 a_1053_103.n6 VSS 0.04fF
C145 a_3829_1050.n0 VSS 0.32fF
C146 a_3829_1050.n1 VSS 0.32fF
C147 a_3829_1050.n2 VSS 0.27fF
C148 a_3829_1050.n3 VSS 0.50fF
C149 a_3829_1050.n4 VSS 0.28fF
C150 a_3829_1050.n5 VSS 0.59fF
C151 a_3829_1050.n6 VSS 0.37fF
C152 a_3829_1050.n7 VSS 0.39fF
C153 a_3829_1050.n8 VSS 0.41fF
C154 a_2141_1050.n0 VSS 0.36fF
C155 a_2141_1050.n1 VSS 0.31fF
C156 a_2141_1050.n2 VSS 0.62fF
C157 a_2141_1050.n3 VSS 0.31fF
C158 a_2141_1050.n4 VSS 0.65fF
C159 a_2141_1050.n5 VSS 0.54fF
C160 a_2141_1050.n6 VSS 0.46fF
C161 a_277_1050.n0 VSS 0.41fF
C162 a_277_1050.n1 VSS 1.62fF
C163 a_277_1050.n2 VSS 0.41fF
C164 a_277_1050.n3 VSS 0.65fF
C165 a_277_1050.n4 VSS 2.31fF
C166 a_277_1050.n5 VSS 0.05fF
C167 a_277_1050.n6 VSS 0.07fF
C168 a_277_1050.n7 VSS 0.05fF
C169 a_277_1050.n8 VSS 0.35fF
C170 a_277_1050.n9 VSS 0.76fF
C171 a_277_1050.n10 VSS 0.53fF
C172 a_277_1050.n11 VSS 0.67fF
C173 a_277_1050.n12 VSS 0.64fF
C174 a_277_1050.n13 VSS 0.56fF
C175 a_277_1050.n14 VSS 0.53fF
C176 a_599_989.n0 VSS 0.40fF
C177 a_599_989.n1 VSS 0.34fF
C178 a_599_989.n2 VSS 0.48fF
C179 a_599_989.n3 VSS 0.34fF
C180 a_599_989.t9 VSS 0.55fF
C181 a_599_989.n4 VSS 0.65fF
C182 a_599_989.n5 VSS 1.04fF
C183 a_599_989.n6 VSS 0.04fF
C184 a_599_989.n7 VSS 0.06fF
C185 a_599_989.n8 VSS 0.04fF
C186 a_599_989.n9 VSS 0.23fF
C187 a_599_989.n10 VSS 0.54fF
C188 a_599_989.n11 VSS 0.46fF
C189 a_599_989.n12 VSS 0.51fF
C190 a_599_989.n13 VSS 0.49fF
C191 a_599_989.n14 VSS 0.40fF
C192 VDD.n1 VSS 0.03fF
C193 VDD.n2 VSS 0.14fF
C194 VDD.n3 VSS 0.03fF
C195 VDD.n4 VSS 0.02fF
C196 VDD.n5 VSS 0.06fF
C197 VDD.n6 VSS 0.02fF
C198 VDD.n7 VSS 0.02fF
C199 VDD.n8 VSS 0.02fF
C200 VDD.n9 VSS 0.02fF
C201 VDD.n10 VSS 0.02fF
C202 VDD.n11 VSS 0.02fF
C203 VDD.n12 VSS 0.02fF
C204 VDD.n13 VSS 0.02fF
C205 VDD.n14 VSS 0.04fF
C206 VDD.n15 VSS 0.01fF
C207 VDD.n20 VSS 0.46fF
C208 VDD.n21 VSS 0.27fF
C209 VDD.n22 VSS 0.02fF
C210 VDD.n23 VSS 0.03fF
C211 VDD.n24 VSS 0.06fF
C212 VDD.n25 VSS 0.24fF
C213 VDD.n26 VSS 0.01fF
C214 VDD.n27 VSS 0.01fF
C215 VDD.n28 VSS 0.01fF
C216 VDD.n29 VSS 0.17fF
C217 VDD.n30 VSS 0.01fF
C218 VDD.n31 VSS 0.02fF
C219 VDD.n32 VSS 0.08fF
C220 VDD.n33 VSS 0.08fF
C221 VDD.n34 VSS 0.05fF
C222 VDD.n35 VSS 0.01fF
C223 VDD.n36 VSS 0.02fF
C224 VDD.n37 VSS 0.03fF
C225 VDD.n38 VSS 0.14fF
C226 VDD.n39 VSS 0.01fF
C227 VDD.n40 VSS 0.02fF
C228 VDD.n41 VSS 0.03fF
C229 VDD.n42 VSS 0.16fF
C230 VDD.n43 VSS 0.01fF
C231 VDD.n44 VSS 0.02fF
C232 VDD.n45 VSS 0.02fF
C233 VDD.n46 VSS 0.06fF
C234 VDD.n47 VSS 0.25fF
C235 VDD.n48 VSS 0.01fF
C236 VDD.n49 VSS 0.01fF
C237 VDD.n50 VSS 0.02fF
C238 VDD.n51 VSS 0.27fF
C239 VDD.n52 VSS 0.01fF
C240 VDD.n53 VSS 0.02fF
C241 VDD.n54 VSS 0.03fF
C242 VDD.n55 VSS 0.05fF
C243 VDD.n56 VSS 0.02fF
C244 VDD.n57 VSS 0.02fF
C245 VDD.n58 VSS 0.02fF
C246 VDD.n59 VSS 0.02fF
C247 VDD.n60 VSS 0.02fF
C248 VDD.n61 VSS 0.02fF
C249 VDD.n62 VSS 0.02fF
C250 VDD.n63 VSS 0.02fF
C251 VDD.n64 VSS 0.02fF
C252 VDD.n65 VSS 0.02fF
C253 VDD.n66 VSS 0.02fF
C254 VDD.n67 VSS 0.03fF
C255 VDD.n68 VSS 0.02fF
C256 VDD.n69 VSS 0.27fF
C257 VDD.n70 VSS 0.02fF
C258 VDD.n71 VSS 0.02fF
C259 VDD.n73 VSS 0.02fF
C260 VDD.n77 VSS 0.27fF
C261 VDD.n78 VSS 0.27fF
C262 VDD.n79 VSS 0.01fF
C263 VDD.n80 VSS 0.02fF
C264 VDD.n81 VSS 0.03fF
C265 VDD.n82 VSS 0.27fF
C266 VDD.n83 VSS 0.01fF
C267 VDD.n84 VSS 0.02fF
C268 VDD.n85 VSS 0.02fF
C269 VDD.n86 VSS 0.22fF
C270 VDD.n87 VSS 0.01fF
C271 VDD.n88 VSS 0.07fF
C272 VDD.n89 VSS 0.02fF
C273 VDD.n90 VSS 0.17fF
C274 VDD.n91 VSS 0.01fF
C275 VDD.n92 VSS 0.02fF
C276 VDD.n93 VSS 0.02fF
C277 VDD.n94 VSS 0.16fF
C278 VDD.n95 VSS 0.01fF
C279 VDD.n96 VSS 0.08fF
C280 VDD.n97 VSS 0.05fF
C281 VDD.n98 VSS 0.02fF
C282 VDD.n99 VSS 0.02fF
C283 VDD.n100 VSS 0.14fF
C284 VDD.n101 VSS 0.01fF
C285 VDD.n102 VSS 0.02fF
C286 VDD.n103 VSS 0.03fF
C287 VDD.n104 VSS 0.15fF
C288 VDD.n105 VSS 0.01fF
C289 VDD.n106 VSS 0.02fF
C290 VDD.n107 VSS 0.03fF
C291 VDD.n108 VSS 0.08fF
C292 VDD.n109 VSS 0.05fF
C293 VDD.n110 VSS 0.16fF
C294 VDD.n111 VSS 0.01fF
C295 VDD.n112 VSS 0.02fF
C296 VDD.n113 VSS 0.02fF
C297 VDD.n114 VSS 0.17fF
C298 VDD.n115 VSS 0.01fF
C299 VDD.n116 VSS 0.02fF
C300 VDD.n117 VSS 0.02fF
C301 VDD.n118 VSS 0.06fF
C302 VDD.n119 VSS 0.22fF
C303 VDD.n120 VSS 0.01fF
C304 VDD.n121 VSS 0.01fF
C305 VDD.n122 VSS 0.02fF
C306 VDD.n123 VSS 0.27fF
C307 VDD.n124 VSS 0.01fF
C308 VDD.n125 VSS 0.02fF
C309 VDD.n126 VSS 0.02fF
C310 VDD.n127 VSS 0.27fF
C311 VDD.n128 VSS 0.01fF
C312 VDD.n129 VSS 0.02fF
C313 VDD.n130 VSS 0.03fF
C314 VDD.n131 VSS 0.31fF
C315 VDD.n132 VSS 0.02fF
C316 VDD.n133 VSS 0.02fF
C317 VDD.n134 VSS 0.02fF
C318 VDD.n135 VSS 0.06fF
C319 VDD.n136 VSS 0.02fF
C320 VDD.n137 VSS 0.02fF
C321 VDD.n138 VSS 0.02fF
C322 VDD.n139 VSS 0.02fF
C323 VDD.n140 VSS 0.02fF
C324 VDD.n141 VSS 0.02fF
C325 VDD.n142 VSS 0.02fF
C326 VDD.n143 VSS 0.02fF
C327 VDD.n144 VSS 0.02fF
C328 VDD.n145 VSS 0.02fF
C329 VDD.n146 VSS 0.03fF
C330 VDD.n147 VSS 0.02fF
C331 VDD.n148 VSS 0.02fF
C332 VDD.n152 VSS 0.27fF
C333 VDD.n153 VSS 0.27fF
C334 VDD.n154 VSS 0.01fF
C335 VDD.n155 VSS 0.02fF
C336 VDD.n156 VSS 0.03fF
C337 VDD.n157 VSS 0.27fF
C338 VDD.n158 VSS 0.01fF
C339 VDD.n159 VSS 0.02fF
C340 VDD.n160 VSS 0.02fF
C341 VDD.n161 VSS 0.22fF
C342 VDD.n162 VSS 0.01fF
C343 VDD.n163 VSS 0.07fF
C344 VDD.n164 VSS 0.02fF
C345 VDD.n165 VSS 0.17fF
C346 VDD.n166 VSS 0.01fF
C347 VDD.n167 VSS 0.02fF
C348 VDD.n168 VSS 0.02fF
C349 VDD.n169 VSS 0.16fF
C350 VDD.n170 VSS 0.01fF
C351 VDD.n171 VSS 0.08fF
C352 VDD.n172 VSS 0.05fF
C353 VDD.n173 VSS 0.02fF
C354 VDD.n174 VSS 0.02fF
C355 VDD.n175 VSS 0.14fF
C356 VDD.n176 VSS 0.01fF
C357 VDD.n177 VSS 0.02fF
C358 VDD.n178 VSS 0.03fF
C359 VDD.n179 VSS 0.15fF
C360 VDD.n180 VSS 0.01fF
C361 VDD.n181 VSS 0.02fF
C362 VDD.n182 VSS 0.03fF
C363 VDD.n183 VSS 0.08fF
C364 VDD.n184 VSS 0.05fF
C365 VDD.n185 VSS 0.16fF
C366 VDD.n186 VSS 0.01fF
C367 VDD.n187 VSS 0.02fF
C368 VDD.n188 VSS 0.02fF
C369 VDD.n189 VSS 0.17fF
C370 VDD.n190 VSS 0.01fF
C371 VDD.n191 VSS 0.02fF
C372 VDD.n192 VSS 0.02fF
C373 VDD.n193 VSS 0.06fF
C374 VDD.n194 VSS 0.22fF
C375 VDD.n195 VSS 0.01fF
C376 VDD.n196 VSS 0.01fF
C377 VDD.n197 VSS 0.02fF
C378 VDD.n198 VSS 0.27fF
C379 VDD.n199 VSS 0.01fF
C380 VDD.n200 VSS 0.02fF
C381 VDD.n201 VSS 0.02fF
C382 VDD.n202 VSS 0.27fF
C383 VDD.n203 VSS 0.01fF
C384 VDD.n204 VSS 0.02fF
C385 VDD.n205 VSS 0.03fF
C386 VDD.n206 VSS 0.26fF
C387 VDD.n207 VSS 0.02fF
C388 VDD.n208 VSS 0.02fF
C389 VDD.n209 VSS 0.02fF
C390 VDD.n210 VSS 0.06fF
C391 VDD.n211 VSS 0.02fF
C392 VDD.n212 VSS 0.02fF
C393 VDD.n213 VSS 0.02fF
C394 VDD.n214 VSS 0.02fF
C395 VDD.n215 VSS 0.02fF
C396 VDD.n216 VSS 0.02fF
C397 VDD.n217 VSS 0.02fF
C398 VDD.n218 VSS 0.02fF
C399 VDD.n219 VSS 0.02fF
C400 VDD.n220 VSS 0.02fF
C401 VDD.n221 VSS 0.03fF
C402 VDD.n222 VSS 0.02fF
C403 VDD.n223 VSS 0.02fF
C404 VDD.n227 VSS 0.27fF
C405 VDD.n228 VSS 0.27fF
C406 VDD.n229 VSS 0.01fF
C407 VDD.n230 VSS 0.02fF
C408 VDD.n231 VSS 0.03fF
C409 VDD.n232 VSS 0.06fF
C410 VDD.n233 VSS 0.24fF
C411 VDD.n234 VSS 0.01fF
C412 VDD.n235 VSS 0.01fF
C413 VDD.n236 VSS 0.02fF
C414 VDD.n237 VSS 0.17fF
C415 VDD.n238 VSS 0.01fF
C416 VDD.n239 VSS 0.02fF
C417 VDD.n240 VSS 0.02fF
C418 VDD.n241 VSS 0.08fF
C419 VDD.n242 VSS 0.05fF
C420 VDD.n243 VSS 0.01fF
C421 VDD.n244 VSS 0.02fF
C422 VDD.n245 VSS 0.03fF
C423 VDD.n246 VSS 0.14fF
C424 VDD.n247 VSS 0.01fF
C425 VDD.n248 VSS 0.02fF
C426 VDD.n249 VSS 0.03fF
C427 VDD.n250 VSS 0.16fF
C428 VDD.n251 VSS 0.01fF
C429 VDD.n252 VSS 0.02fF
C430 VDD.n253 VSS 0.02fF
C431 VDD.n254 VSS 0.06fF
C432 VDD.n255 VSS 0.25fF
C433 VDD.n256 VSS 0.01fF
C434 VDD.n257 VSS 0.01fF
C435 VDD.n258 VSS 0.02fF
C436 VDD.n259 VSS 0.27fF
C437 VDD.n260 VSS 0.01fF
C438 VDD.n261 VSS 0.02fF
C439 VDD.n262 VSS 0.03fF
C440 VDD.n263 VSS 0.26fF
C441 VDD.n264 VSS 0.02fF
C442 VDD.n265 VSS 0.02fF
C443 VDD.n266 VSS 0.02fF
C444 VDD.n267 VSS 0.06fF
C445 VDD.n268 VSS 0.02fF
C446 VDD.n269 VSS 0.02fF
C447 VDD.n270 VSS 0.02fF
C448 VDD.n271 VSS 0.02fF
C449 VDD.n272 VSS 0.02fF
C450 VDD.n273 VSS 0.02fF
C451 VDD.n274 VSS 0.02fF
C452 VDD.n275 VSS 0.02fF
C453 VDD.n276 VSS 0.02fF
C454 VDD.n277 VSS 0.02fF
C455 VDD.n278 VSS 0.03fF
C456 VDD.n279 VSS 0.02fF
C457 VDD.n280 VSS 0.02fF
C458 VDD.n284 VSS 0.27fF
C459 VDD.n285 VSS 0.27fF
C460 VDD.n286 VSS 0.01fF
C461 VDD.n287 VSS 0.02fF
C462 VDD.n288 VSS 0.03fF
C463 VDD.n289 VSS 0.27fF
C464 VDD.n290 VSS 0.01fF
C465 VDD.n291 VSS 0.02fF
C466 VDD.n292 VSS 0.02fF
C467 VDD.n293 VSS 0.22fF
C468 VDD.n294 VSS 0.01fF
C469 VDD.n295 VSS 0.07fF
C470 VDD.n296 VSS 0.02fF
C471 VDD.n297 VSS 0.17fF
C472 VDD.n298 VSS 0.01fF
C473 VDD.n299 VSS 0.02fF
C474 VDD.n300 VSS 0.02fF
C475 VDD.n301 VSS 0.16fF
C476 VDD.n302 VSS 0.01fF
C477 VDD.n303 VSS 0.08fF
C478 VDD.n304 VSS 0.05fF
C479 VDD.n305 VSS 0.02fF
C480 VDD.n306 VSS 0.02fF
C481 VDD.n307 VSS 0.14fF
C482 VDD.n308 VSS 0.01fF
C483 VDD.n309 VSS 0.02fF
C484 VDD.n310 VSS 0.03fF
C485 VDD.n311 VSS 0.15fF
C486 VDD.n312 VSS 0.01fF
C487 VDD.n313 VSS 0.02fF
C488 VDD.n314 VSS 0.03fF
C489 VDD.n315 VSS 0.08fF
C490 VDD.n316 VSS 0.05fF
C491 VDD.n317 VSS 0.16fF
C492 VDD.n318 VSS 0.01fF
C493 VDD.n319 VSS 0.02fF
C494 VDD.n320 VSS 0.02fF
C495 VDD.n321 VSS 0.17fF
C496 VDD.n322 VSS 0.01fF
C497 VDD.n323 VSS 0.02fF
C498 VDD.n324 VSS 0.02fF
C499 VDD.n325 VSS 0.06fF
C500 VDD.n326 VSS 0.22fF
C501 VDD.n327 VSS 0.01fF
C502 VDD.n328 VSS 0.01fF
C503 VDD.n329 VSS 0.02fF
C504 VDD.n330 VSS 0.27fF
C505 VDD.n331 VSS 0.01fF
C506 VDD.n332 VSS 0.02fF
C507 VDD.n333 VSS 0.02fF
C508 VDD.n334 VSS 0.27fF
C509 VDD.n335 VSS 0.01fF
C510 VDD.n336 VSS 0.02fF
C511 VDD.n337 VSS 0.03fF
C512 VDD.n338 VSS 0.05fF
C513 VDD.n339 VSS 0.02fF
C514 VDD.n340 VSS 0.02fF
C515 VDD.n341 VSS 0.02fF
C516 VDD.n342 VSS 0.02fF
C517 VDD.n343 VSS 0.02fF
C518 VDD.n344 VSS 0.02fF
C519 VDD.n345 VSS 0.02fF
C520 VDD.n346 VSS 0.02fF
C521 VDD.n347 VSS 0.02fF
C522 VDD.n348 VSS 0.02fF
C523 VDD.n349 VSS 0.02fF
C524 VDD.n350 VSS 0.03fF
C525 VDD.n351 VSS 0.02fF
C526 VDD.n354 VSS 0.02fF
C527 VDD.n356 VSS 0.02fF
C528 VDD.n357 VSS 0.31fF
C529 VDD.n358 VSS 0.02fF
C530 VDD.n360 VSS 0.27fF
C531 VDD.n361 VSS 0.27fF
C532 VDD.n362 VSS 0.01fF
C533 VDD.n363 VSS 0.02fF
C534 VDD.n364 VSS 0.03fF
C535 VDD.n365 VSS 0.27fF
C536 VDD.n366 VSS 0.01fF
C537 VDD.n367 VSS 0.02fF
C538 VDD.n368 VSS 0.02fF
C539 VDD.n369 VSS 0.22fF
C540 VDD.n370 VSS 0.01fF
C541 VDD.n371 VSS 0.07fF
C542 VDD.n372 VSS 0.02fF
C543 VDD.n373 VSS 0.17fF
C544 VDD.n374 VSS 0.01fF
C545 VDD.n375 VSS 0.02fF
C546 VDD.n376 VSS 0.02fF
C547 VDD.n377 VSS 0.16fF
C548 VDD.n378 VSS 0.01fF
C549 VDD.n379 VSS 0.08fF
C550 VDD.n380 VSS 0.05fF
C551 VDD.n381 VSS 0.02fF
C552 VDD.n382 VSS 0.02fF
C553 VDD.n383 VSS 0.14fF
C554 VDD.n384 VSS 0.01fF
C555 VDD.n385 VSS 0.02fF
C556 VDD.n386 VSS 0.03fF
C557 VDD.n387 VSS 0.15fF
C558 VDD.n388 VSS 0.01fF
C559 VDD.n389 VSS 0.02fF
C560 VDD.n390 VSS 0.03fF
C561 VDD.n391 VSS 0.08fF
C562 VDD.n392 VSS 0.05fF
C563 VDD.n393 VSS 0.16fF
C564 VDD.n394 VSS 0.01fF
C565 VDD.n395 VSS 0.02fF
C566 VDD.n396 VSS 0.02fF
C567 VDD.n397 VSS 0.17fF
C568 VDD.n398 VSS 0.01fF
C569 VDD.n399 VSS 0.02fF
C570 VDD.n400 VSS 0.02fF
C571 VDD.n401 VSS 0.06fF
C572 VDD.n402 VSS 0.22fF
C573 VDD.n403 VSS 0.01fF
C574 VDD.n404 VSS 0.01fF
C575 VDD.n405 VSS 0.02fF
C576 VDD.n406 VSS 0.27fF
C577 VDD.n