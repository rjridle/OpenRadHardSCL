magic
tech sky130A
magscale 1 2
timestamp 1643656459
<< nmos >>
rect 152 226 182 288
tri 56 196 86 226 se
rect 86 196 182 226
rect 56 92 86 196
tri 86 180 102 196 nw
tri 136 180 152 196 ne
tri 86 92 102 108 sw
tri 136 92 152 108 se
rect 152 92 182 196
tri 56 62 86 92 ne
rect 86 62 152 92
tri 152 62 182 92 nw
<< ndiff >>
rect 0 260 152 288
rect 0 226 10 260
rect 44 226 152 260
rect 182 260 238 288
rect 182 226 194 260
rect 228 226 238 260
rect 0 189 56 226
tri 56 196 86 226 nw
rect 0 155 10 189
rect 44 155 56 189
rect 0 121 56 155
rect 0 87 10 121
rect 44 87 56 121
tri 86 180 102 196 se
rect 102 180 136 196
tri 136 180 152 196 sw
rect 86 155 152 180
rect 86 121 102 155
rect 136 121 152 155
rect 86 108 152 121
tri 86 92 102 108 ne
rect 102 92 136 108
tri 136 92 152 108 nw
rect 182 189 238 226
rect 182 155 194 189
rect 228 155 238 189
rect 182 121 238 155
rect 0 62 56 87
tri 56 62 86 92 sw
tri 152 62 182 92 se
rect 182 87 194 121
rect 228 87 238 121
rect 182 62 238 87
rect 0 50 238 62
rect 0 16 10 50
rect 44 16 102 50
rect 136 16 194 50
rect 228 16 238 50
rect 0 0 238 16
<< ndiffc >>
rect 10 226 44 260
rect 194 226 228 260
rect 10 155 44 189
rect 10 87 44 121
rect 102 121 136 155
rect 194 155 228 189
rect 194 87 228 121
rect 10 16 44 50
rect 102 16 136 50
rect 194 16 228 50
<< poly >>
rect 152 288 182 314
<< locali >>
rect 10 260 44 288
rect 10 189 44 226
rect 194 260 228 288
rect 194 189 228 226
rect 10 121 44 155
rect 102 155 136 171
rect 102 105 136 121
rect 194 121 228 155
rect 10 50 44 87
rect 194 50 228 87
rect 44 16 102 50
rect 136 16 194 50
rect 10 0 44 16
rect 194 0 228 16
<< end >>
