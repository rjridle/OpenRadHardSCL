magic
tech sky130A
magscale 1 2
timestamp 1649549310
<< nwell >>
rect -528 832 4080 1575
<< nmos >>
rect -289 324 -259 377
tri -259 324 -243 340 sw
rect -289 294 -183 324
tri -183 294 -153 324 sw
rect -289 193 -259 294
tri -259 278 -243 294 nw
tri -199 278 -183 294 ne
tri -259 193 -243 209 sw
tri -199 193 -183 209 se
rect -183 193 -153 294
tri -289 163 -259 193 ne
rect -259 163 -183 193
tri -183 163 -153 193 nw
rect 155 324 185 377
tri 185 324 201 340 sw
rect 155 294 261 324
tri 261 294 291 324 sw
rect 155 193 185 294
tri 185 278 201 294 nw
tri 245 278 261 294 ne
tri 185 193 201 209 sw
tri 245 193 261 209 se
rect 261 193 291 294
tri 155 163 185 193 ne
rect 185 163 261 193
tri 261 163 291 193 nw
rect 612 316 642 377
tri 642 316 658 332 sw
rect 806 324 836 377
tri 836 324 852 340 sw
rect 612 286 718 316
tri 718 286 748 316 sw
rect 806 294 912 324
tri 912 294 942 324 sw
rect 612 185 642 286
tri 642 270 658 286 nw
tri 702 270 718 286 ne
tri 642 185 658 201 sw
tri 702 185 718 201 se
rect 718 185 748 286
rect 806 193 836 294
tri 836 278 852 294 nw
tri 896 278 912 294 ne
tri 836 193 852 209 sw
tri 896 193 912 209 se
rect 912 193 942 294
tri 612 155 642 185 ne
rect 642 155 718 185
tri 718 155 748 185 nw
tri 806 163 836 193 ne
rect 836 163 912 193
tri 912 163 942 193 nw
rect 1265 324 1295 377
tri 1295 324 1311 340 sw
rect 1265 294 1371 324
tri 1371 294 1401 324 sw
rect 1265 193 1295 294
tri 1295 278 1311 294 nw
tri 1355 278 1371 294 ne
tri 1295 193 1311 209 sw
tri 1355 193 1371 209 se
rect 1371 193 1401 294
tri 1265 163 1295 193 ne
rect 1295 163 1371 193
tri 1371 163 1401 193 nw
rect 1722 316 1752 377
tri 1752 316 1768 332 sw
rect 1916 324 1946 377
tri 1946 324 1962 340 sw
rect 1722 286 1828 316
tri 1828 286 1858 316 sw
rect 1916 294 2022 324
tri 2022 294 2052 324 sw
rect 1722 185 1752 286
tri 1752 270 1768 286 nw
tri 1812 270 1828 286 ne
tri 1752 185 1768 201 sw
tri 1812 185 1828 201 se
rect 1828 185 1858 286
rect 1916 193 1946 294
tri 1946 278 1962 294 nw
tri 2006 278 2022 294 ne
tri 1946 193 1962 209 sw
tri 2006 193 2022 209 se
rect 2022 193 2052 294
tri 1722 155 1752 185 ne
rect 1752 155 1828 185
tri 1828 155 1858 185 nw
tri 1916 163 1946 193 ne
rect 1946 163 2022 193
tri 2022 163 2052 193 nw
rect 2375 324 2405 377
tri 2405 324 2421 340 sw
rect 2375 294 2481 324
tri 2481 294 2511 324 sw
rect 2375 193 2405 294
tri 2405 278 2421 294 nw
tri 2465 278 2481 294 ne
tri 2405 193 2421 209 sw
tri 2465 193 2481 209 se
rect 2481 193 2511 294
tri 2375 163 2405 193 ne
rect 2405 163 2481 193
tri 2481 163 2511 193 nw
rect 2832 324 2862 377
tri 2862 324 2878 340 sw
rect 3026 324 3056 377
tri 3056 324 3072 340 sw
rect 2832 294 2938 324
tri 2938 294 2968 324 sw
rect 2832 193 2862 294
tri 2862 278 2878 294 nw
tri 2922 278 2938 294 ne
tri 2862 193 2878 209 sw
tri 2922 193 2938 209 se
rect 2938 193 2968 294
rect 3026 294 3132 324
tri 3132 294 3162 324 sw
rect 3026 279 3057 294
tri 3057 279 3072 294 nw
tri 3116 279 3131 294 ne
rect 3131 279 3162 294
tri 2832 163 2862 193 ne
rect 2862 163 2938 193
tri 2938 163 2968 193 nw
rect 3026 193 3056 279
tri 3056 193 3072 209 sw
tri 3116 193 3132 209 se
rect 3132 193 3162 279
tri 3026 163 3056 193 ne
rect 3056 163 3132 193
tri 3132 163 3162 193 nw
rect 3498 324 3528 377
tri 3528 324 3544 340 sw
rect 3692 324 3722 377
tri 3722 324 3738 340 sw
rect 3498 294 3604 324
tri 3604 294 3634 324 sw
rect 3498 193 3528 294
tri 3528 278 3544 294 nw
tri 3588 278 3604 294 ne
tri 3528 193 3544 209 sw
tri 3588 193 3604 209 se
rect 3604 193 3634 294
rect 3692 294 3798 324
tri 3798 294 3828 324 sw
rect 3692 279 3723 294
tri 3723 279 3738 294 nw
tri 3782 279 3797 294 ne
rect 3797 279 3828 294
tri 3498 163 3528 193 ne
rect 3528 163 3604 193
tri 3604 163 3634 193 nw
rect 3692 193 3722 279
tri 3722 193 3738 209 sw
tri 3782 193 3798 209 se
rect 3798 193 3828 279
tri 3692 163 3722 193 ne
rect 3722 163 3798 193
tri 3798 163 3828 193 nw
<< pmos >>
rect -281 1050 -251 1450
rect -193 1050 -163 1450
rect 163 1050 193 1450
rect 251 1050 281 1450
rect 631 1050 661 1450
rect 719 1050 749 1450
rect 807 1050 837 1450
rect 895 1050 925 1450
rect 1273 1050 1303 1450
rect 1361 1050 1391 1450
rect 1741 1050 1771 1450
rect 1829 1050 1859 1450
rect 1917 1050 1947 1450
rect 2005 1050 2035 1450
rect 2383 1050 2413 1450
rect 2471 1050 2501 1450
rect 2851 1051 2881 1451
rect 2939 1051 2969 1451
rect 3027 1051 3057 1451
rect 3115 1051 3145 1451
rect 3517 1051 3547 1451
rect 3605 1051 3635 1451
rect 3693 1051 3723 1451
rect 3781 1051 3811 1451
<< ndiff >>
rect -345 361 -289 377
rect -345 327 -335 361
rect -301 327 -289 361
rect -345 289 -289 327
rect -259 361 -99 377
rect -259 340 -141 361
tri -259 324 -243 340 ne
rect -243 327 -141 340
rect -107 327 -99 361
rect -243 324 -99 327
tri -183 294 -153 324 ne
rect -345 255 -335 289
rect -301 255 -289 289
rect -345 221 -289 255
rect -345 187 -335 221
rect -301 187 -289 221
tri -259 278 -243 294 se
rect -243 278 -199 294
tri -199 278 -183 294 sw
rect -259 245 -183 278
rect -259 211 -239 245
rect -205 211 -183 245
rect -259 209 -183 211
tri -259 193 -243 209 ne
rect -243 193 -199 209
tri -199 193 -183 209 nw
rect -153 289 -99 324
rect -153 255 -141 289
rect -107 255 -99 289
rect -153 221 -99 255
rect -345 163 -289 187
tri -289 163 -259 193 sw
tri -183 163 -153 193 se
rect -153 187 -141 221
rect -107 187 -99 221
rect -153 163 -99 187
rect -345 151 -99 163
rect -345 117 -335 151
rect -301 117 -239 151
rect -205 117 -141 151
rect -107 117 -99 151
rect -345 101 -99 117
rect 99 361 155 377
rect 99 327 109 361
rect 143 327 155 361
rect 99 289 155 327
rect 185 361 345 377
rect 185 340 303 361
tri 185 324 201 340 ne
rect 201 327 303 340
rect 337 327 345 361
rect 201 324 345 327
tri 261 294 291 324 ne
rect 99 255 109 289
rect 143 255 155 289
rect 99 221 155 255
rect 99 187 109 221
rect 143 187 155 221
tri 185 278 201 294 se
rect 201 278 245 294
tri 245 278 261 294 sw
rect 185 245 261 278
rect 185 211 205 245
rect 239 211 261 245
rect 185 209 261 211
tri 185 193 201 209 ne
rect 201 193 245 209
tri 245 193 261 209 nw
rect 291 289 345 324
rect 291 255 303 289
rect 337 255 345 289
rect 291 221 345 255
rect 99 163 155 187
tri 155 163 185 193 sw
tri 261 163 291 193 se
rect 291 187 303 221
rect 337 187 345 221
rect 291 163 345 187
rect 99 151 345 163
rect 99 117 109 151
rect 143 117 205 151
rect 239 117 303 151
rect 337 117 345 151
rect 99 101 345 117
rect 556 361 612 377
rect 556 327 566 361
rect 600 327 612 361
rect 556 289 612 327
rect 642 361 806 377
rect 642 332 663 361
tri 642 316 658 332 ne
rect 658 327 663 332
rect 697 327 760 361
rect 794 327 806 361
rect 658 316 806 327
rect 836 340 998 377
tri 836 324 852 340 ne
rect 852 324 998 340
rect 556 255 566 289
rect 600 255 612 289
tri 718 286 748 316 ne
rect 748 289 806 316
tri 912 294 942 324 ne
rect 556 221 612 255
rect 556 187 566 221
rect 600 187 612 221
rect 556 155 612 187
tri 642 270 658 286 se
rect 658 270 702 286
tri 702 270 718 286 sw
rect 642 236 718 270
rect 642 202 663 236
rect 697 202 718 236
rect 642 201 718 202
tri 642 185 658 201 ne
rect 658 185 702 201
tri 702 185 718 201 nw
rect 748 255 760 289
rect 794 255 806 289
rect 748 221 806 255
rect 748 187 760 221
rect 794 187 806 221
tri 836 278 852 294 se
rect 852 278 896 294
tri 896 278 912 294 sw
rect 836 245 912 278
rect 836 211 857 245
rect 891 211 912 245
rect 836 209 912 211
tri 836 193 852 209 ne
rect 852 193 896 209
tri 896 193 912 209 nw
rect 942 289 998 324
rect 942 255 954 289
rect 988 255 998 289
rect 942 221 998 255
tri 612 155 642 185 sw
tri 718 155 748 185 se
rect 748 163 806 187
tri 806 163 836 193 sw
tri 912 163 942 193 se
rect 942 187 954 221
rect 988 187 998 221
rect 942 163 998 187
rect 748 155 998 163
rect 556 151 998 155
rect 556 117 566 151
rect 600 117 760 151
rect 794 117 857 151
rect 891 117 954 151
rect 988 117 998 151
rect 556 101 998 117
rect 1209 361 1265 377
rect 1209 327 1219 361
rect 1253 327 1265 361
rect 1209 289 1265 327
rect 1295 361 1455 377
rect 1295 340 1413 361
tri 1295 324 1311 340 ne
rect 1311 327 1413 340
rect 1447 327 1455 361
rect 1311 324 1455 327
tri 1371 294 1401 324 ne
rect 1209 255 1219 289
rect 1253 255 1265 289
rect 1209 221 1265 255
rect 1209 187 1219 221
rect 1253 187 1265 221
tri 1295 278 1311 294 se
rect 1311 278 1355 294
tri 1355 278 1371 294 sw
rect 1295 245 1371 278
rect 1295 211 1315 245
rect 1349 211 1371 245
rect 1295 209 1371 211
tri 1295 193 1311 209 ne
rect 1311 193 1355 209
tri 1355 193 1371 209 nw
rect 1401 289 1455 324
rect 1401 255 1413 289
rect 1447 255 1455 289
rect 1401 221 1455 255
rect 1209 163 1265 187
tri 1265 163 1295 193 sw
tri 1371 163 1401 193 se
rect 1401 187 1413 221
rect 1447 187 1455 221
rect 1401 163 1455 187
rect 1209 151 1455 163
rect 1209 117 1219 151
rect 1253 117 1315 151
rect 1349 117 1413 151
rect 1447 117 1455 151
rect 1209 101 1455 117
rect 1666 361 1722 377
rect 1666 327 1676 361
rect 1710 327 1722 361
rect 1666 289 1722 327
rect 1752 361 1916 377
rect 1752 332 1773 361
tri 1752 316 1768 332 ne
rect 1768 327 1773 332
rect 1807 327 1870 361
rect 1904 327 1916 361
rect 1768 316 1916 327
rect 1946 340 2108 377
tri 1946 324 1962 340 ne
rect 1962 324 2108 340
rect 1666 255 1676 289
rect 1710 255 1722 289
tri 1828 286 1858 316 ne
rect 1858 289 1916 316
tri 2022 294 2052 324 ne
rect 1666 221 1722 255
rect 1666 187 1676 221
rect 1710 187 1722 221
rect 1666 155 1722 187
tri 1752 270 1768 286 se
rect 1768 270 1812 286
tri 1812 270 1828 286 sw
rect 1752 236 1828 270
rect 1752 202 1773 236
rect 1807 202 1828 236
rect 1752 201 1828 202
tri 1752 185 1768 201 ne
rect 1768 185 1812 201
tri 1812 185 1828 201 nw
rect 1858 255 1870 289
rect 1904 255 1916 289
rect 1858 221 1916 255
rect 1858 187 1870 221
rect 1904 187 1916 221
tri 1946 278 1962 294 se
rect 1962 278 2006 294
tri 2006 278 2022 294 sw
rect 1946 245 2022 278
rect 1946 211 1967 245
rect 2001 211 2022 245
rect 1946 209 2022 211
tri 1946 193 1962 209 ne
rect 1962 193 2006 209
tri 2006 193 2022 209 nw
rect 2052 289 2108 324
rect 2052 255 2064 289
rect 2098 255 2108 289
rect 2052 221 2108 255
tri 1722 155 1752 185 sw
tri 1828 155 1858 185 se
rect 1858 163 1916 187
tri 1916 163 1946 193 sw
tri 2022 163 2052 193 se
rect 2052 187 2064 221
rect 2098 187 2108 221
rect 2052 163 2108 187
rect 1858 155 2108 163
rect 1666 151 2108 155
rect 1666 117 1676 151
rect 1710 117 1870 151
rect 1904 117 1967 151
rect 2001 117 2064 151
rect 2098 117 2108 151
rect 1666 101 2108 117
rect 2319 361 2375 377
rect 2319 327 2329 361
rect 2363 327 2375 361
rect 2319 289 2375 327
rect 2405 361 2565 377
rect 2405 340 2523 361
tri 2405 324 2421 340 ne
rect 2421 327 2523 340
rect 2557 327 2565 361
rect 2421 324 2565 327
tri 2481 294 2511 324 ne
rect 2319 255 2329 289
rect 2363 255 2375 289
rect 2319 221 2375 255
rect 2319 187 2329 221
rect 2363 187 2375 221
tri 2405 278 2421 294 se
rect 2421 278 2465 294
tri 2465 278 2481 294 sw
rect 2405 245 2481 278
rect 2405 211 2425 245
rect 2459 211 2481 245
rect 2405 209 2481 211
tri 2405 193 2421 209 ne
rect 2421 193 2465 209
tri 2465 193 2481 209 nw
rect 2511 289 2565 324
rect 2511 255 2523 289
rect 2557 255 2565 289
rect 2511 221 2565 255
rect 2319 163 2375 187
tri 2375 163 2405 193 sw
tri 2481 163 2511 193 se
rect 2511 187 2523 221
rect 2557 187 2565 221
rect 2511 163 2565 187
rect 2319 151 2565 163
rect 2319 117 2329 151
rect 2363 117 2425 151
rect 2459 117 2523 151
rect 2557 117 2565 151
rect 2319 101 2565 117
rect 2776 361 2832 377
rect 2776 327 2786 361
rect 2820 327 2832 361
rect 2776 289 2832 327
rect 2862 340 3026 377
tri 2862 324 2878 340 ne
rect 2878 324 3026 340
rect 3056 340 3218 377
tri 3056 324 3072 340 ne
rect 3072 324 3218 340
tri 2938 294 2968 324 ne
rect 2776 255 2786 289
rect 2820 255 2832 289
rect 2776 221 2832 255
rect 2776 187 2786 221
rect 2820 187 2832 221
tri 2862 278 2878 294 se
rect 2878 278 2922 294
tri 2922 278 2938 294 sw
rect 2862 245 2938 278
rect 2862 211 2883 245
rect 2917 211 2938 245
rect 2862 209 2938 211
tri 2862 193 2878 209 ne
rect 2878 193 2922 209
tri 2922 193 2938 209 nw
rect 2968 289 3026 324
tri 3132 294 3162 324 ne
rect 2968 255 2980 289
rect 3014 255 3026 289
tri 3057 279 3072 294 se
rect 3072 279 3116 294
tri 3116 279 3131 294 sw
rect 3162 289 3218 324
rect 2968 221 3026 255
rect 2776 163 2832 187
tri 2832 163 2862 193 sw
tri 2938 163 2968 193 se
rect 2968 187 2980 221
rect 3014 187 3026 221
rect 3056 245 3132 279
rect 3056 211 3077 245
rect 3111 211 3132 245
rect 3056 209 3132 211
tri 3056 193 3072 209 ne
rect 3072 193 3116 209
tri 3116 193 3132 209 nw
rect 3162 255 3174 289
rect 3208 255 3218 289
rect 3162 221 3218 255
rect 2968 163 3026 187
tri 3026 163 3056 193 sw
tri 3132 163 3162 193 se
rect 3162 187 3174 221
rect 3208 187 3218 221
rect 3162 163 3218 187
rect 2776 151 3218 163
rect 2776 117 2786 151
rect 2820 117 2883 151
rect 2917 117 2980 151
rect 3014 117 3077 151
rect 3111 117 3174 151
rect 3208 117 3218 151
rect 2776 101 3218 117
rect 3442 361 3498 377
rect 3442 327 3452 361
rect 3486 327 3498 361
rect 3442 289 3498 327
rect 3528 340 3692 377
tri 3528 324 3544 340 ne
rect 3544 324 3692 340
rect 3722 340 3884 377
tri 3722 324 3738 340 ne
rect 3738 324 3884 340
tri 3604 294 3634 324 ne
rect 3442 255 3452 289
rect 3486 255 3498 289
rect 3442 221 3498 255
rect 3442 187 3452 221
rect 3486 187 3498 221
tri 3528 278 3544 294 se
rect 3544 278 3588 294
tri 3588 278 3604 294 sw
rect 3528 245 3604 278
rect 3528 211 3549 245
rect 3583 211 3604 245
rect 3528 209 3604 211
tri 3528 193 3544 209 ne
rect 3544 193 3588 209
tri 3588 193 3604 209 nw
rect 3634 289 3692 324
tri 3798 294 3828 324 ne
rect 3634 255 3646 289
rect 3680 255 3692 289
tri 3723 279 3738 294 se
rect 3738 279 3782 294
tri 3782 279 3797 294 sw
rect 3828 289 3884 324
rect 3634 221 3692 255
rect 3442 163 3498 187
tri 3498 163 3528 193 sw
tri 3604 163 3634 193 se
rect 3634 187 3646 221
rect 3680 187 3692 221
rect 3722 245 3798 279
rect 3722 211 3743 245
rect 3777 211 3798 245
rect 3722 209 3798 211
tri 3722 193 3738 209 ne
rect 3738 193 3782 209
tri 3782 193 3798 209 nw
rect 3828 255 3840 289
rect 3874 255 3884 289
rect 3828 221 3884 255
rect 3634 163 3692 187
tri 3692 163 3722 193 sw
tri 3798 163 3828 193 se
rect 3828 187 3840 221
rect 3874 187 3884 221
rect 3828 163 3884 187
rect 3442 151 3884 163
rect 3442 117 3452 151
rect 3486 117 3549 151
rect 3583 117 3646 151
rect 3680 117 3743 151
rect 3777 117 3840 151
rect 3874 117 3884 151
rect 3442 101 3884 117
<< pdiff >>
rect -337 1412 -281 1450
rect -337 1378 -327 1412
rect -293 1378 -281 1412
rect -337 1344 -281 1378
rect -337 1310 -327 1344
rect -293 1310 -281 1344
rect -337 1276 -281 1310
rect -337 1242 -327 1276
rect -293 1242 -281 1276
rect -337 1208 -281 1242
rect -337 1174 -327 1208
rect -293 1174 -281 1208
rect -337 1139 -281 1174
rect -337 1105 -327 1139
rect -293 1105 -281 1139
rect -337 1050 -281 1105
rect -251 1412 -193 1450
rect -251 1378 -239 1412
rect -205 1378 -193 1412
rect -251 1344 -193 1378
rect -251 1310 -239 1344
rect -205 1310 -193 1344
rect -251 1276 -193 1310
rect -251 1242 -239 1276
rect -205 1242 -193 1276
rect -251 1208 -193 1242
rect -251 1174 -239 1208
rect -205 1174 -193 1208
rect -251 1139 -193 1174
rect -251 1105 -239 1139
rect -205 1105 -193 1139
rect -251 1050 -193 1105
rect -163 1412 -109 1450
rect -163 1378 -151 1412
rect -117 1378 -109 1412
rect -163 1344 -109 1378
rect -163 1310 -151 1344
rect -117 1310 -109 1344
rect -163 1276 -109 1310
rect -163 1242 -151 1276
rect -117 1242 -109 1276
rect -163 1208 -109 1242
rect -163 1174 -151 1208
rect -117 1174 -109 1208
rect -163 1139 -109 1174
rect -163 1105 -151 1139
rect -117 1105 -109 1139
rect -163 1050 -109 1105
rect 107 1412 163 1450
rect 107 1378 117 1412
rect 151 1378 163 1412
rect 107 1344 163 1378
rect 107 1310 117 1344
rect 151 1310 163 1344
rect 107 1276 163 1310
rect 107 1242 117 1276
rect 151 1242 163 1276
rect 107 1208 163 1242
rect 107 1174 117 1208
rect 151 1174 163 1208
rect 107 1139 163 1174
rect 107 1105 117 1139
rect 151 1105 163 1139
rect 107 1050 163 1105
rect 193 1412 251 1450
rect 193 1378 205 1412
rect 239 1378 251 1412
rect 193 1344 251 1378
rect 193 1310 205 1344
rect 239 1310 251 1344
rect 193 1276 251 1310
rect 193 1242 205 1276
rect 239 1242 251 1276
rect 193 1208 251 1242
rect 193 1174 205 1208
rect 239 1174 251 1208
rect 193 1139 251 1174
rect 193 1105 205 1139
rect 239 1105 251 1139
rect 193 1050 251 1105
rect 281 1412 335 1450
rect 281 1378 293 1412
rect 327 1378 335 1412
rect 281 1344 335 1378
rect 281 1310 293 1344
rect 327 1310 335 1344
rect 281 1276 335 1310
rect 281 1242 293 1276
rect 327 1242 335 1276
rect 281 1208 335 1242
rect 281 1174 293 1208
rect 327 1174 335 1208
rect 281 1139 335 1174
rect 281 1105 293 1139
rect 327 1105 335 1139
rect 281 1050 335 1105
rect 575 1412 631 1450
rect 575 1378 585 1412
rect 619 1378 631 1412
rect 575 1344 631 1378
rect 575 1310 585 1344
rect 619 1310 631 1344
rect 575 1276 631 1310
rect 575 1242 585 1276
rect 619 1242 631 1276
rect 575 1208 631 1242
rect 575 1174 585 1208
rect 619 1174 631 1208
rect 575 1139 631 1174
rect 575 1105 585 1139
rect 619 1105 631 1139
rect 575 1050 631 1105
rect 661 1412 719 1450
rect 661 1378 673 1412
rect 707 1378 719 1412
rect 661 1344 719 1378
rect 661 1310 673 1344
rect 707 1310 719 1344
rect 661 1276 719 1310
rect 661 1242 673 1276
rect 707 1242 719 1276
rect 661 1208 719 1242
rect 661 1174 673 1208
rect 707 1174 719 1208
rect 661 1139 719 1174
rect 661 1105 673 1139
rect 707 1105 719 1139
rect 661 1050 719 1105
rect 749 1412 807 1450
rect 749 1378 761 1412
rect 795 1378 807 1412
rect 749 1344 807 1378
rect 749 1310 761 1344
rect 795 1310 807 1344
rect 749 1276 807 1310
rect 749 1242 761 1276
rect 795 1242 807 1276
rect 749 1208 807 1242
rect 749 1174 761 1208
rect 795 1174 807 1208
rect 749 1050 807 1174
rect 837 1412 895 1450
rect 837 1378 849 1412
rect 883 1378 895 1412
rect 837 1344 895 1378
rect 837 1310 849 1344
rect 883 1310 895 1344
rect 837 1276 895 1310
rect 837 1242 849 1276
rect 883 1242 895 1276
rect 837 1208 895 1242
rect 837 1174 849 1208
rect 883 1174 895 1208
rect 837 1139 895 1174
rect 837 1105 849 1139
rect 883 1105 895 1139
rect 837 1050 895 1105
rect 925 1412 979 1450
rect 925 1378 937 1412
rect 971 1378 979 1412
rect 925 1344 979 1378
rect 925 1310 937 1344
rect 971 1310 979 1344
rect 925 1276 979 1310
rect 925 1242 937 1276
rect 971 1242 979 1276
rect 925 1208 979 1242
rect 925 1174 937 1208
rect 971 1174 979 1208
rect 925 1050 979 1174
rect 1217 1412 1273 1450
rect 1217 1378 1227 1412
rect 1261 1378 1273 1412
rect 1217 1344 1273 1378
rect 1217 1310 1227 1344
rect 1261 1310 1273 1344
rect 1217 1276 1273 1310
rect 1217 1242 1227 1276
rect 1261 1242 1273 1276
rect 1217 1208 1273 1242
rect 1217 1174 1227 1208
rect 1261 1174 1273 1208
rect 1217 1139 1273 1174
rect 1217 1105 1227 1139
rect 1261 1105 1273 1139
rect 1217 1050 1273 1105
rect 1303 1412 1361 1450
rect 1303 1378 1315 1412
rect 1349 1378 1361 1412
rect 1303 1344 1361 1378
rect 1303 1310 1315 1344
rect 1349 1310 1361 1344
rect 1303 1276 1361 1310
rect 1303 1242 1315 1276
rect 1349 1242 1361 1276
rect 1303 1208 1361 1242
rect 1303 1174 1315 1208
rect 1349 1174 1361 1208
rect 1303 1139 1361 1174
rect 1303 1105 1315 1139
rect 1349 1105 1361 1139
rect 1303 1050 1361 1105
rect 1391 1412 1445 1450
rect 1391 1378 1403 1412
rect 1437 1378 1445 1412
rect 1391 1344 1445 1378
rect 1391 1310 1403 1344
rect 1437 1310 1445 1344
rect 1391 1276 1445 1310
rect 1391 1242 1403 1276
rect 1437 1242 1445 1276
rect 1391 1208 1445 1242
rect 1391 1174 1403 1208
rect 1437 1174 1445 1208
rect 1391 1139 1445 1174
rect 1391 1105 1403 1139
rect 1437 1105 1445 1139
rect 1391 1050 1445 1105
rect 1685 1412 1741 1450
rect 1685 1378 1695 1412
rect 1729 1378 1741 1412
rect 1685 1344 1741 1378
rect 1685 1310 1695 1344
rect 1729 1310 1741 1344
rect 1685 1276 1741 1310
rect 1685 1242 1695 1276
rect 1729 1242 1741 1276
rect 1685 1208 1741 1242
rect 1685 1174 1695 1208
rect 1729 1174 1741 1208
rect 1685 1139 1741 1174
rect 1685 1105 1695 1139
rect 1729 1105 1741 1139
rect 1685 1050 1741 1105
rect 1771 1412 1829 1450
rect 1771 1378 1783 1412
rect 1817 1378 1829 1412
rect 1771 1344 1829 1378
rect 1771 1310 1783 1344
rect 1817 1310 1829 1344
rect 1771 1276 1829 1310
rect 1771 1242 1783 1276
rect 1817 1242 1829 1276
rect 1771 1208 1829 1242
rect 1771 1174 1783 1208
rect 1817 1174 1829 1208
rect 1771 1139 1829 1174
rect 1771 1105 1783 1139
rect 1817 1105 1829 1139
rect 1771 1050 1829 1105
rect 1859 1412 1917 1450
rect 1859 1378 1871 1412
rect 1905 1378 1917 1412
rect 1859 1344 1917 1378
rect 1859 1310 1871 1344
rect 1905 1310 1917 1344
rect 1859 1276 1917 1310
rect 1859 1242 1871 1276
rect 1905 1242 1917 1276
rect 1859 1208 1917 1242
rect 1859 1174 1871 1208
rect 1905 1174 1917 1208
rect 1859 1050 1917 1174
rect 1947 1412 2005 1450
rect 1947 1378 1959 1412
rect 1993 1378 2005 1412
rect 1947 1344 2005 1378
rect 1947 1310 1959 1344
rect 1993 1310 2005 1344
rect 1947 1276 2005 1310
rect 1947 1242 1959 1276
rect 1993 1242 2005 1276
rect 1947 1208 2005 1242
rect 1947 1174 1959 1208
rect 1993 1174 2005 1208
rect 1947 1139 2005 1174
rect 1947 1105 1959 1139
rect 1993 1105 2005 1139
rect 1947 1050 2005 1105
rect 2035 1412 2089 1450
rect 2035 1378 2047 1412
rect 2081 1378 2089 1412
rect 2035 1344 2089 1378
rect 2035 1310 2047 1344
rect 2081 1310 2089 1344
rect 2035 1276 2089 1310
rect 2035 1242 2047 1276
rect 2081 1242 2089 1276
rect 2035 1208 2089 1242
rect 2035 1174 2047 1208
rect 2081 1174 2089 1208
rect 2035 1050 2089 1174
rect 2327 1412 2383 1450
rect 2327 1378 2337 1412
rect 2371 1378 2383 1412
rect 2327 1344 2383 1378
rect 2327 1310 2337 1344
rect 2371 1310 2383 1344
rect 2327 1276 2383 1310
rect 2327 1242 2337 1276
rect 2371 1242 2383 1276
rect 2327 1208 2383 1242
rect 2327 1174 2337 1208
rect 2371 1174 2383 1208
rect 2327 1139 2383 1174
rect 2327 1105 2337 1139
rect 2371 1105 2383 1139
rect 2327 1050 2383 1105
rect 2413 1412 2471 1450
rect 2413 1378 2425 1412
rect 2459 1378 2471 1412
rect 2413 1344 2471 1378
rect 2413 1310 2425 1344
rect 2459 1310 2471 1344
rect 2413 1276 2471 1310
rect 2413 1242 2425 1276
rect 2459 1242 2471 1276
rect 2413 1208 2471 1242
rect 2413 1174 2425 1208
rect 2459 1174 2471 1208
rect 2413 1139 2471 1174
rect 2413 1105 2425 1139
rect 2459 1105 2471 1139
rect 2413 1050 2471 1105
rect 2501 1412 2555 1450
rect 2501 1378 2513 1412
rect 2547 1378 2555 1412
rect 2501 1344 2555 1378
rect 2501 1310 2513 1344
rect 2547 1310 2555 1344
rect 2501 1276 2555 1310
rect 2501 1242 2513 1276
rect 2547 1242 2555 1276
rect 2501 1208 2555 1242
rect 2501 1174 2513 1208
rect 2547 1174 2555 1208
rect 2501 1139 2555 1174
rect 2501 1105 2513 1139
rect 2547 1105 2555 1139
rect 2501 1050 2555 1105
rect 2795 1411 2851 1451
rect 2795 1377 2805 1411
rect 2839 1377 2851 1411
rect 2795 1343 2851 1377
rect 2795 1309 2805 1343
rect 2839 1309 2851 1343
rect 2795 1275 2851 1309
rect 2795 1241 2805 1275
rect 2839 1241 2851 1275
rect 2795 1207 2851 1241
rect 2795 1173 2805 1207
rect 2839 1173 2851 1207
rect 2795 1139 2851 1173
rect 2795 1105 2805 1139
rect 2839 1105 2851 1139
rect 2795 1051 2851 1105
rect 2881 1411 2939 1451
rect 2881 1377 2893 1411
rect 2927 1377 2939 1411
rect 2881 1343 2939 1377
rect 2881 1309 2893 1343
rect 2927 1309 2939 1343
rect 2881 1275 2939 1309
rect 2881 1241 2893 1275
rect 2927 1241 2939 1275
rect 2881 1207 2939 1241
rect 2881 1173 2893 1207
rect 2927 1173 2939 1207
rect 2881 1051 2939 1173
rect 2969 1411 3027 1451
rect 2969 1377 2981 1411
rect 3015 1377 3027 1411
rect 2969 1343 3027 1377
rect 2969 1309 2981 1343
rect 3015 1309 3027 1343
rect 2969 1275 3027 1309
rect 2969 1241 2981 1275
rect 3015 1241 3027 1275
rect 2969 1207 3027 1241
rect 2969 1173 2981 1207
rect 3015 1173 3027 1207
rect 2969 1139 3027 1173
rect 2969 1105 2981 1139
rect 3015 1105 3027 1139
rect 2969 1051 3027 1105
rect 3057 1343 3115 1451
rect 3057 1309 3069 1343
rect 3103 1309 3115 1343
rect 3057 1275 3115 1309
rect 3057 1241 3069 1275
rect 3103 1241 3115 1275
rect 3057 1207 3115 1241
rect 3057 1173 3069 1207
rect 3103 1173 3115 1207
rect 3057 1139 3115 1173
rect 3057 1105 3069 1139
rect 3103 1105 3115 1139
rect 3057 1051 3115 1105
rect 3145 1411 3199 1451
rect 3145 1377 3157 1411
rect 3191 1377 3199 1411
rect 3145 1343 3199 1377
rect 3145 1309 3157 1343
rect 3191 1309 3199 1343
rect 3145 1275 3199 1309
rect 3145 1241 3157 1275
rect 3191 1241 3199 1275
rect 3145 1207 3199 1241
rect 3145 1173 3157 1207
rect 3191 1173 3199 1207
rect 3145 1051 3199 1173
rect 3461 1411 3517 1451
rect 3461 1377 3471 1411
rect 3505 1377 3517 1411
rect 3461 1343 3517 1377
rect 3461 1309 3471 1343
rect 3505 1309 3517 1343
rect 3461 1275 3517 1309
rect 3461 1241 3471 1275
rect 3505 1241 3517 1275
rect 3461 1207 3517 1241
rect 3461 1173 3471 1207
rect 3505 1173 3517 1207
rect 3461 1139 3517 1173
rect 3461 1105 3471 1139
rect 3505 1105 3517 1139
rect 3461 1051 3517 1105
rect 3547 1411 3605 1451
rect 3547 1377 3559 1411
rect 3593 1377 3605 1411
rect 3547 1343 3605 1377
rect 3547 1309 3559 1343
rect 3593 1309 3605 1343
rect 3547 1275 3605 1309
rect 3547 1241 3559 1275
rect 3593 1241 3605 1275
rect 3547 1207 3605 1241
rect 3547 1173 3559 1207
rect 3593 1173 3605 1207
rect 3547 1051 3605 1173
rect 3635 1411 3693 1451
rect 3635 1377 3647 1411
rect 3681 1377 3693 1411
rect 3635 1343 3693 1377
rect 3635 1309 3647 1343
rect 3681 1309 3693 1343
rect 3635 1275 3693 1309
rect 3635 1241 3647 1275
rect 3681 1241 3693 1275
rect 3635 1207 3693 1241
rect 3635 1173 3647 1207
rect 3681 1173 3693 1207
rect 3635 1139 3693 1173
rect 3635 1105 3647 1139
rect 3681 1105 3693 1139
rect 3635 1051 3693 1105
rect 3723 1343 3781 1451
rect 3723 1309 3735 1343
rect 3769 1309 3781 1343
rect 3723 1275 3781 1309
rect 3723 1241 3735 1275
rect 3769 1241 3781 1275
rect 3723 1207 3781 1241
rect 3723 1173 3735 1207
rect 3769 1173 3781 1207
rect 3723 1139 3781 1173
rect 3723 1105 3735 1139
rect 3769 1105 3781 1139
rect 3723 1051 3781 1105
rect 3811 1411 3865 1451
rect 3811 1377 3823 1411
rect 3857 1377 3865 1411
rect 3811 1343 3865 1377
rect 3811 1309 3823 1343
rect 3857 1309 3865 1343
rect 3811 1275 3865 1309
rect 3811 1241 3823 1275
rect 3857 1241 3865 1275
rect 3811 1207 3865 1241
rect 3811 1173 3823 1207
rect 3857 1173 3865 1207
rect 3811 1051 3865 1173
<< ndiffc >>
rect -335 327 -301 361
rect -141 327 -107 361
rect -335 255 -301 289
rect -335 187 -301 221
rect -239 211 -205 245
rect -141 255 -107 289
rect -141 187 -107 221
rect -335 117 -301 151
rect -239 117 -205 151
rect -141 117 -107 151
rect 109 327 143 361
rect 303 327 337 361
rect 109 255 143 289
rect 109 187 143 221
rect 205 211 239 245
rect 303 255 337 289
rect 303 187 337 221
rect 109 117 143 151
rect 205 117 239 151
rect 303 117 337 151
rect 566 327 600 361
rect 663 327 697 361
rect 760 327 794 361
rect 566 255 600 289
rect 566 187 600 221
rect 663 202 697 236
rect 760 255 794 289
rect 760 187 794 221
rect 857 211 891 245
rect 954 255 988 289
rect 954 187 988 221
rect 566 117 600 151
rect 760 117 794 151
rect 857 117 891 151
rect 954 117 988 151
rect 1219 327 1253 361
rect 1413 327 1447 361
rect 1219 255 1253 289
rect 1219 187 1253 221
rect 1315 211 1349 245
rect 1413 255 1447 289
rect 1413 187 1447 221
rect 1219 117 1253 151
rect 1315 117 1349 151
rect 1413 117 1447 151
rect 1676 327 1710 361
rect 1773 327 1807 361
rect 1870 327 1904 361
rect 1676 255 1710 289
rect 1676 187 1710 221
rect 1773 202 1807 236
rect 1870 255 1904 289
rect 1870 187 1904 221
rect 1967 211 2001 245
rect 2064 255 2098 289
rect 2064 187 2098 221
rect 1676 117 1710 151
rect 1870 117 1904 151
rect 1967 117 2001 151
rect 2064 117 2098 151
rect 2329 327 2363 361
rect 2523 327 2557 361
rect 2329 255 2363 289
rect 2329 187 2363 221
rect 2425 211 2459 245
rect 2523 255 2557 289
rect 2523 187 2557 221
rect 2329 117 2363 151
rect 2425 117 2459 151
rect 2523 117 2557 151
rect 2786 327 2820 361
rect 2786 255 2820 289
rect 2786 187 2820 221
rect 2883 211 2917 245
rect 2980 255 3014 289
rect 2980 187 3014 221
rect 3077 211 3111 245
rect 3174 255 3208 289
rect 3174 187 3208 221
rect 2786 117 2820 151
rect 2883 117 2917 151
rect 2980 117 3014 151
rect 3077 117 3111 151
rect 3174 117 3208 151
rect 3452 327 3486 361
rect 3452 255 3486 289
rect 3452 187 3486 221
rect 3549 211 3583 245
rect 3646 255 3680 289
rect 3646 187 3680 221
rect 3743 211 3777 245
rect 3840 255 3874 289
rect 3840 187 3874 221
rect 3452 117 3486 151
rect 3549 117 3583 151
rect 3646 117 3680 151
rect 3743 117 3777 151
rect 3840 117 3874 151
<< pdiffc >>
rect -327 1378 -293 1412
rect -327 1310 -293 1344
rect -327 1242 -293 1276
rect -327 1174 -293 1208
rect -327 1105 -293 1139
rect -239 1378 -205 1412
rect -239 1310 -205 1344
rect -239 1242 -205 1276
rect -239 1174 -205 1208
rect -239 1105 -205 1139
rect -151 1378 -117 1412
rect -151 1310 -117 1344
rect -151 1242 -117 1276
rect -151 1174 -117 1208
rect -151 1105 -117 1139
rect 117 1378 151 1412
rect 117 1310 151 1344
rect 117 1242 151 1276
rect 117 1174 151 1208
rect 117 1105 151 1139
rect 205 1378 239 1412
rect 205 1310 239 1344
rect 205 1242 239 1276
rect 205 1174 239 1208
rect 205 1105 239 1139
rect 293 1378 327 1412
rect 293 1310 327 1344
rect 293 1242 327 1276
rect 293 1174 327 1208
rect 293 1105 327 1139
rect 585 1378 619 1412
rect 585 1310 619 1344
rect 585 1242 619 1276
rect 585 1174 619 1208
rect 585 1105 619 1139
rect 673 1378 707 1412
rect 673 1310 707 1344
rect 673 1242 707 1276
rect 673 1174 707 1208
rect 673 1105 707 1139
rect 761 1378 795 1412
rect 761 1310 795 1344
rect 761 1242 795 1276
rect 761 1174 795 1208
rect 849 1378 883 1412
rect 849 1310 883 1344
rect 849 1242 883 1276
rect 849 1174 883 1208
rect 849 1105 883 1139
rect 937 1378 971 1412
rect 937 1310 971 1344
rect 937 1242 971 1276
rect 937 1174 971 1208
rect 1227 1378 1261 1412
rect 1227 1310 1261 1344
rect 1227 1242 1261 1276
rect 1227 1174 1261 1208
rect 1227 1105 1261 1139
rect 1315 1378 1349 1412
rect 1315 1310 1349 1344
rect 1315 1242 1349 1276
rect 1315 1174 1349 1208
rect 1315 1105 1349 1139
rect 1403 1378 1437 1412
rect 1403 1310 1437 1344
rect 1403 1242 1437 1276
rect 1403 1174 1437 1208
rect 1403 1105 1437 1139
rect 1695 1378 1729 1412
rect 1695 1310 1729 1344
rect 1695 1242 1729 1276
rect 1695 1174 1729 1208
rect 1695 1105 1729 1139
rect 1783 1378 1817 1412
rect 1783 1310 1817 1344
rect 1783 1242 1817 1276
rect 1783 1174 1817 1208
rect 1783 1105 1817 1139
rect 1871 1378 1905 1412
rect 1871 1310 1905 1344
rect 1871 1242 1905 1276
rect 1871 1174 1905 1208
rect 1959 1378 1993 1412
rect 1959 1310 1993 1344
rect 1959 1242 1993 1276
rect 1959 1174 1993 1208
rect 1959 1105 1993 1139
rect 2047 1378 2081 1412
rect 2047 1310 2081 1344
rect 2047 1242 2081 1276
rect 2047 1174 2081 1208
rect 2337 1378 2371 1412
rect 2337 1310 2371 1344
rect 2337 1242 2371 1276
rect 2337 1174 2371 1208
rect 2337 1105 2371 1139
rect 2425 1378 2459 1412
rect 2425 1310 2459 1344
rect 2425 1242 2459 1276
rect 2425 1174 2459 1208
rect 2425 1105 2459 1139
rect 2513 1378 2547 1412
rect 2513 1310 2547 1344
rect 2513 1242 2547 1276
rect 2513 1174 2547 1208
rect 2513 1105 2547 1139
rect 2805 1377 2839 1411
rect 2805 1309 2839 1343
rect 2805 1241 2839 1275
rect 2805 1173 2839 1207
rect 2805 1105 2839 1139
rect 2893 1377 2927 1411
rect 2893 1309 2927 1343
rect 2893 1241 2927 1275
rect 2893 1173 2927 1207
rect 2981 1377 3015 1411
rect 2981 1309 3015 1343
rect 2981 1241 3015 1275
rect 2981 1173 3015 1207
rect 2981 1105 3015 1139
rect 3069 1309 3103 1343
rect 3069 1241 3103 1275
rect 3069 1173 3103 1207
rect 3069 1105 3103 1139
rect 3157 1377 3191 1411
rect 3157 1309 3191 1343
rect 3157 1241 3191 1275
rect 3157 1173 3191 1207
rect 3471 1377 3505 1411
rect 3471 1309 3505 1343
rect 3471 1241 3505 1275
rect 3471 1173 3505 1207
rect 3471 1105 3505 1139
rect 3559 1377 3593 1411
rect 3559 1309 3593 1343
rect 3559 1241 3593 1275
rect 3559 1173 3593 1207
rect 3647 1377 3681 1411
rect 3647 1309 3681 1343
rect 3647 1241 3681 1275
rect 3647 1173 3681 1207
rect 3647 1105 3681 1139
rect 3735 1309 3769 1343
rect 3735 1241 3769 1275
rect 3735 1173 3769 1207
rect 3735 1105 3769 1139
rect 3823 1377 3857 1411
rect 3823 1309 3857 1343
rect 3823 1241 3857 1275
rect 3823 1173 3857 1207
<< psubdiff >>
rect -475 546 4027 572
rect -475 512 -461 546
rect -427 512 -17 546
rect 17 512 427 546
rect 461 512 1093 546
rect 1127 512 1537 546
rect 1571 512 2203 546
rect 2237 512 2647 546
rect 2681 512 3313 546
rect 3347 512 3979 546
rect 4013 512 4027 546
rect -475 510 4027 512
rect -475 474 -413 510
rect -475 440 -461 474
rect -427 440 -413 474
rect -475 402 -413 440
rect -31 474 31 510
rect -475 368 -461 402
rect -427 368 -413 402
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect 413 474 475 510
rect -475 330 -413 368
rect -475 296 -461 330
rect -427 296 -413 330
rect -475 258 -413 296
rect -475 224 -461 258
rect -427 224 -413 258
rect -475 186 -413 224
rect -475 152 -461 186
rect -427 152 -413 186
rect -475 114 -413 152
rect -475 80 -461 114
rect -427 80 -413 114
rect -31 368 -17 402
rect 17 368 31 402
rect 413 440 427 474
rect 461 440 475 474
rect 413 402 475 440
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -475 47 -413 80
rect -31 80 -17 114
rect 17 80 31 114
rect 413 368 427 402
rect 461 368 475 402
rect 1079 474 1141 510
rect 1079 440 1093 474
rect 1127 440 1141 474
rect 1079 402 1141 440
rect 1523 474 1585 510
rect 413 330 475 368
rect 413 296 427 330
rect 461 296 475 330
rect 413 258 475 296
rect 413 224 427 258
rect 461 224 475 258
rect 413 186 475 224
rect 413 152 427 186
rect 461 152 475 186
rect 413 114 475 152
rect -31 47 31 80
rect 413 80 427 114
rect 461 80 475 114
rect 1079 368 1093 402
rect 1127 368 1141 402
rect 1523 440 1537 474
rect 1571 440 1585 474
rect 1523 402 1585 440
rect 1079 330 1141 368
rect 1079 296 1093 330
rect 1127 296 1141 330
rect 1079 258 1141 296
rect 1079 224 1093 258
rect 1127 224 1141 258
rect 1079 186 1141 224
rect 1079 152 1093 186
rect 1127 152 1141 186
rect 1079 114 1141 152
rect 413 47 475 80
rect 1079 80 1093 114
rect 1127 80 1141 114
rect 1523 368 1537 402
rect 1571 368 1585 402
rect 2189 474 2251 510
rect 2189 440 2203 474
rect 2237 440 2251 474
rect 2189 402 2251 440
rect 2633 474 2695 510
rect 1523 330 1585 368
rect 1523 296 1537 330
rect 1571 296 1585 330
rect 1523 258 1585 296
rect 1523 224 1537 258
rect 1571 224 1585 258
rect 1523 186 1585 224
rect 1523 152 1537 186
rect 1571 152 1585 186
rect 1523 114 1585 152
rect 1079 47 1141 80
rect 1523 80 1537 114
rect 1571 80 1585 114
rect 2189 368 2203 402
rect 2237 368 2251 402
rect 2633 440 2647 474
rect 2681 440 2695 474
rect 2633 402 2695 440
rect 2189 330 2251 368
rect 2189 296 2203 330
rect 2237 296 2251 330
rect 2189 258 2251 296
rect 2189 224 2203 258
rect 2237 224 2251 258
rect 2189 186 2251 224
rect 2189 152 2203 186
rect 2237 152 2251 186
rect 2189 114 2251 152
rect 1523 47 1585 80
rect 2189 80 2203 114
rect 2237 80 2251 114
rect 2633 368 2647 402
rect 2681 368 2695 402
rect 3299 474 3361 510
rect 3299 440 3313 474
rect 3347 440 3361 474
rect 3299 402 3361 440
rect 2633 330 2695 368
rect 2633 296 2647 330
rect 2681 296 2695 330
rect 2633 258 2695 296
rect 2633 224 2647 258
rect 2681 224 2695 258
rect 2633 186 2695 224
rect 2633 152 2647 186
rect 2681 152 2695 186
rect 2633 114 2695 152
rect 2189 47 2251 80
rect 2633 80 2647 114
rect 2681 80 2695 114
rect 3299 368 3313 402
rect 3347 368 3361 402
rect 3965 474 4027 510
rect 3965 440 3979 474
rect 4013 440 4027 474
rect 3965 402 4027 440
rect 3299 330 3361 368
rect 3299 296 3313 330
rect 3347 296 3361 330
rect 3299 258 3361 296
rect 3299 224 3313 258
rect 3347 224 3361 258
rect 3299 186 3361 224
rect 3299 152 3313 186
rect 3347 152 3361 186
rect 3299 114 3361 152
rect 2633 47 2695 80
rect 3299 80 3313 114
rect 3347 80 3361 114
rect 3965 368 3979 402
rect 4013 368 4027 402
rect 3965 330 4027 368
rect 3965 296 3979 330
rect 4013 296 4027 330
rect 3965 258 4027 296
rect 3965 224 3979 258
rect 4013 224 4027 258
rect 3965 186 4027 224
rect 3965 152 3979 186
rect 4013 152 4027 186
rect 3965 114 4027 152
rect 3299 47 3361 80
rect 3965 80 3979 114
rect 4013 80 4027 114
rect 3965 47 4027 80
rect -475 13 -389 47
rect -355 13 -317 47
rect -283 13 -239 47
rect -205 13 -161 47
rect -127 13 -89 47
rect -55 13 55 47
rect 89 13 127 47
rect 161 13 205 47
rect 239 13 283 47
rect 317 13 355 47
rect 389 13 499 47
rect 533 13 571 47
rect 605 13 643 47
rect 677 13 715 47
rect 749 13 805 47
rect 839 13 877 47
rect 911 13 949 47
rect 983 13 1021 47
rect 1055 13 1165 47
rect 1199 13 1237 47
rect 1271 13 1315 47
rect 1349 13 1393 47
rect 1427 13 1465 47
rect 1499 13 1609 47
rect 1643 13 1681 47
rect 1715 13 1753 47
rect 1787 13 1825 47
rect 1859 13 1915 47
rect 1949 13 1987 47
rect 2021 13 2059 47
rect 2093 13 2131 47
rect 2165 13 2275 47
rect 2309 13 2347 47
rect 2381 13 2425 47
rect 2459 13 2503 47
rect 2537 13 2575 47
rect 2609 13 2719 47
rect 2753 13 2791 47
rect 2825 13 2863 47
rect 2897 13 2935 47
rect 2969 13 3025 47
rect 3059 13 3097 47
rect 3131 13 3169 47
rect 3203 13 3241 47
rect 3275 13 3385 47
rect 3419 13 3457 47
rect 3491 13 3529 47
rect 3563 13 3601 47
rect 3635 13 3691 47
rect 3725 13 3763 47
rect 3797 13 3835 47
rect 3869 13 3907 47
rect 3941 13 4027 47
rect -475 11 -413 13
rect -31 11 31 13
rect 413 11 475 13
rect 1079 11 1141 13
rect 1523 11 1585 13
rect 2189 11 2251 13
rect 2633 11 2695 13
rect 3299 11 3361 13
rect 3965 11 4027 13
<< nsubdiff >>
rect -475 1505 -389 1539
rect -355 1505 -317 1539
rect -283 1505 -239 1539
rect -205 1505 -161 1539
rect -127 1505 -89 1539
rect -55 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 205 1539
rect 239 1505 283 1539
rect 317 1505 355 1539
rect 389 1505 499 1539
rect 533 1505 571 1539
rect 605 1505 643 1539
rect 677 1505 715 1539
rect 749 1505 805 1539
rect 839 1505 877 1539
rect 911 1505 949 1539
rect 983 1505 1021 1539
rect 1055 1505 1165 1539
rect 1199 1505 1237 1539
rect 1271 1505 1315 1539
rect 1349 1505 1393 1539
rect 1427 1505 1465 1539
rect 1499 1505 1609 1539
rect 1643 1505 1681 1539
rect 1715 1505 1753 1539
rect 1787 1505 1825 1539
rect 1859 1505 1915 1539
rect 1949 1505 1987 1539
rect 2021 1505 2059 1539
rect 2093 1505 2131 1539
rect 2165 1505 2275 1539
rect 2309 1505 2347 1539
rect 2381 1505 2425 1539
rect 2459 1505 2503 1539
rect 2537 1505 2575 1539
rect 2609 1505 2719 1539
rect 2753 1505 2791 1539
rect 2825 1505 2863 1539
rect 2897 1505 2935 1539
rect 2969 1505 3025 1539
rect 3059 1505 3097 1539
rect 3131 1505 3169 1539
rect 3203 1505 3241 1539
rect 3275 1505 3385 1539
rect 3419 1505 3457 1539
rect 3491 1505 3529 1539
rect 3563 1505 3601 1539
rect 3635 1505 3691 1539
rect 3725 1505 3763 1539
rect 3797 1505 3835 1539
rect 3869 1505 3907 1539
rect 3941 1505 4027 1539
rect -475 1470 -413 1505
rect -475 1436 -461 1470
rect -427 1436 -413 1470
rect -31 1470 31 1505
rect -475 1398 -413 1436
rect -475 1364 -461 1398
rect -427 1364 -413 1398
rect -475 1326 -413 1364
rect -475 1292 -461 1326
rect -427 1292 -413 1326
rect -475 1254 -413 1292
rect -475 1220 -461 1254
rect -427 1220 -413 1254
rect -475 1182 -413 1220
rect -475 1148 -461 1182
rect -427 1148 -413 1182
rect -475 1110 -413 1148
rect -475 1076 -461 1110
rect -427 1076 -413 1110
rect -475 1038 -413 1076
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect 413 1470 475 1505
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect -475 1004 -461 1038
rect -427 1004 -413 1038
rect -475 966 -413 1004
rect -475 932 -461 966
rect -427 932 -413 966
rect -31 1038 31 1076
rect 413 1436 427 1470
rect 461 1436 475 1470
rect 1079 1470 1141 1505
rect 413 1398 475 1436
rect 413 1364 427 1398
rect 461 1364 475 1398
rect 413 1326 475 1364
rect 413 1292 427 1326
rect 461 1292 475 1326
rect 413 1254 475 1292
rect 413 1220 427 1254
rect 461 1220 475 1254
rect 413 1182 475 1220
rect 413 1148 427 1182
rect 461 1148 475 1182
rect 413 1110 475 1148
rect 413 1076 427 1110
rect 461 1076 475 1110
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -475 930 -413 932
rect -31 932 -17 966
rect 17 932 31 966
rect 413 1038 475 1076
rect 1079 1436 1093 1470
rect 1127 1436 1141 1470
rect 1523 1470 1585 1505
rect 1079 1398 1141 1436
rect 1079 1364 1093 1398
rect 1127 1364 1141 1398
rect 1079 1326 1141 1364
rect 1079 1292 1093 1326
rect 1127 1292 1141 1326
rect 1079 1254 1141 1292
rect 1079 1220 1093 1254
rect 1127 1220 1141 1254
rect 1079 1182 1141 1220
rect 1079 1148 1093 1182
rect 1127 1148 1141 1182
rect 1079 1110 1141 1148
rect 1079 1076 1093 1110
rect 1127 1076 1141 1110
rect 413 1004 427 1038
rect 461 1004 475 1038
rect 413 966 475 1004
rect -31 930 31 932
rect 413 932 427 966
rect 461 932 475 966
rect 1079 1038 1141 1076
rect 1523 1436 1537 1470
rect 1571 1436 1585 1470
rect 2189 1470 2251 1505
rect 1523 1398 1585 1436
rect 1523 1364 1537 1398
rect 1571 1364 1585 1398
rect 1523 1326 1585 1364
rect 1523 1292 1537 1326
rect 1571 1292 1585 1326
rect 1523 1254 1585 1292
rect 1523 1220 1537 1254
rect 1571 1220 1585 1254
rect 1523 1182 1585 1220
rect 1523 1148 1537 1182
rect 1571 1148 1585 1182
rect 1523 1110 1585 1148
rect 1523 1076 1537 1110
rect 1571 1076 1585 1110
rect 1079 1004 1093 1038
rect 1127 1004 1141 1038
rect 1079 966 1141 1004
rect 413 930 475 932
rect 1079 932 1093 966
rect 1127 932 1141 966
rect 1523 1038 1585 1076
rect 2189 1436 2203 1470
rect 2237 1436 2251 1470
rect 2633 1470 2695 1505
rect 2189 1398 2251 1436
rect 2189 1364 2203 1398
rect 2237 1364 2251 1398
rect 2189 1326 2251 1364
rect 2189 1292 2203 1326
rect 2237 1292 2251 1326
rect 2189 1254 2251 1292
rect 2189 1220 2203 1254
rect 2237 1220 2251 1254
rect 2189 1182 2251 1220
rect 2189 1148 2203 1182
rect 2237 1148 2251 1182
rect 2189 1110 2251 1148
rect 2189 1076 2203 1110
rect 2237 1076 2251 1110
rect 1523 1004 1537 1038
rect 1571 1004 1585 1038
rect 1523 966 1585 1004
rect 1079 930 1141 932
rect 1523 932 1537 966
rect 1571 932 1585 966
rect 2189 1038 2251 1076
rect 2633 1436 2647 1470
rect 2681 1436 2695 1470
rect 3299 1470 3361 1505
rect 2633 1398 2695 1436
rect 2633 1364 2647 1398
rect 2681 1364 2695 1398
rect 2633 1326 2695 1364
rect 2633 1292 2647 1326
rect 2681 1292 2695 1326
rect 2633 1254 2695 1292
rect 2633 1220 2647 1254
rect 2681 1220 2695 1254
rect 2633 1182 2695 1220
rect 2633 1148 2647 1182
rect 2681 1148 2695 1182
rect 2633 1110 2695 1148
rect 2633 1076 2647 1110
rect 2681 1076 2695 1110
rect 2189 1004 2203 1038
rect 2237 1004 2251 1038
rect 2189 966 2251 1004
rect 1523 930 1585 932
rect 2189 932 2203 966
rect 2237 932 2251 966
rect 2633 1038 2695 1076
rect 3299 1436 3313 1470
rect 3347 1436 3361 1470
rect 3965 1470 4027 1505
rect 3299 1398 3361 1436
rect 3299 1364 3313 1398
rect 3347 1364 3361 1398
rect 3299 1326 3361 1364
rect 3299 1292 3313 1326
rect 3347 1292 3361 1326
rect 3299 1254 3361 1292
rect 3299 1220 3313 1254
rect 3347 1220 3361 1254
rect 3299 1182 3361 1220
rect 3299 1148 3313 1182
rect 3347 1148 3361 1182
rect 3299 1110 3361 1148
rect 3299 1076 3313 1110
rect 3347 1076 3361 1110
rect 2633 1004 2647 1038
rect 2681 1004 2695 1038
rect 2633 966 2695 1004
rect 2189 930 2251 932
rect 2633 932 2647 966
rect 2681 932 2695 966
rect 3299 1038 3361 1076
rect 3965 1436 3979 1470
rect 4013 1436 4027 1470
rect 3965 1398 4027 1436
rect 3965 1364 3979 1398
rect 4013 1364 4027 1398
rect 3965 1326 4027 1364
rect 3965 1292 3979 1326
rect 4013 1292 4027 1326
rect 3965 1254 4027 1292
rect 3965 1220 3979 1254
rect 4013 1220 4027 1254
rect 3965 1182 4027 1220
rect 3965 1148 3979 1182
rect 4013 1148 4027 1182
rect 3965 1110 4027 1148
rect 3965 1076 3979 1110
rect 4013 1076 4027 1110
rect 3299 1004 3313 1038
rect 3347 1004 3361 1038
rect 3299 966 3361 1004
rect 2633 930 2695 932
rect 3299 932 3313 966
rect 3347 932 3361 966
rect 3965 1038 4027 1076
rect 3965 1004 3979 1038
rect 4013 1004 4027 1038
rect 3965 966 4027 1004
rect 3299 930 3361 932
rect 3965 932 3979 966
rect 4013 932 4027 966
rect 3965 930 4027 932
rect -475 868 4027 930
<< psubdiffcont >>
rect -461 512 -427 546
rect -17 512 17 546
rect 427 512 461 546
rect 1093 512 1127 546
rect 1537 512 1571 546
rect 2203 512 2237 546
rect 2647 512 2681 546
rect 3313 512 3347 546
rect 3979 512 4013 546
rect -461 440 -427 474
rect -461 368 -427 402
rect -17 440 17 474
rect -461 296 -427 330
rect -461 224 -427 258
rect -461 152 -427 186
rect -461 80 -427 114
rect -17 368 17 402
rect 427 440 461 474
rect -17 296 17 330
rect -17 224 17 258
rect -17 152 17 186
rect -17 80 17 114
rect 427 368 461 402
rect 1093 440 1127 474
rect 427 296 461 330
rect 427 224 461 258
rect 427 152 461 186
rect 427 80 461 114
rect 1093 368 1127 402
rect 1537 440 1571 474
rect 1093 296 1127 330
rect 1093 224 1127 258
rect 1093 152 1127 186
rect 1093 80 1127 114
rect 1537 368 1571 402
rect 2203 440 2237 474
rect 1537 296 1571 330
rect 1537 224 1571 258
rect 1537 152 1571 186
rect 1537 80 1571 114
rect 2203 368 2237 402
rect 2647 440 2681 474
rect 2203 296 2237 330
rect 2203 224 2237 258
rect 2203 152 2237 186
rect 2203 80 2237 114
rect 2647 368 2681 402
rect 3313 440 3347 474
rect 2647 296 2681 330
rect 2647 224 2681 258
rect 2647 152 2681 186
rect 2647 80 2681 114
rect 3313 368 3347 402
rect 3979 440 4013 474
rect 3313 296 3347 330
rect 3313 224 3347 258
rect 3313 152 3347 186
rect 3313 80 3347 114
rect 3979 368 4013 402
rect 3979 296 4013 330
rect 3979 224 4013 258
rect 3979 152 4013 186
rect 3979 80 4013 114
rect -389 13 -355 47
rect -317 13 -283 47
rect -239 13 -205 47
rect -161 13 -127 47
rect -89 13 -55 47
rect 55 13 89 47
rect 127 13 161 47
rect 205 13 239 47
rect 283 13 317 47
rect 355 13 389 47
rect 499 13 533 47
rect 571 13 605 47
rect 643 13 677 47
rect 715 13 749 47
rect 805 13 839 47
rect 877 13 911 47
rect 949 13 983 47
rect 1021 13 1055 47
rect 1165 13 1199 47
rect 1237 13 1271 47
rect 1315 13 1349 47
rect 1393 13 1427 47
rect 1465 13 1499 47
rect 1609 13 1643 47
rect 1681 13 1715 47
rect 1753 13 1787 47
rect 1825 13 1859 47
rect 1915 13 1949 47
rect 1987 13 2021 47
rect 2059 13 2093 47
rect 2131 13 2165 47
rect 2275 13 2309 47
rect 2347 13 2381 47
rect 2425 13 2459 47
rect 2503 13 2537 47
rect 2575 13 2609 47
rect 2719 13 2753 47
rect 2791 13 2825 47
rect 2863 13 2897 47
rect 2935 13 2969 47
rect 3025 13 3059 47
rect 3097 13 3131 47
rect 3169 13 3203 47
rect 3241 13 3275 47
rect 3385 13 3419 47
rect 3457 13 3491 47
rect 3529 13 3563 47
rect 3601 13 3635 47
rect 3691 13 3725 47
rect 3763 13 3797 47
rect 3835 13 3869 47
rect 3907 13 3941 47
<< nsubdiffcont >>
rect -389 1505 -355 1539
rect -317 1505 -283 1539
rect -239 1505 -205 1539
rect -161 1505 -127 1539
rect -89 1505 -55 1539
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 205 1505 239 1539
rect 283 1505 317 1539
rect 355 1505 389 1539
rect 499 1505 533 1539
rect 571 1505 605 1539
rect 643 1505 677 1539
rect 715 1505 749 1539
rect 805 1505 839 1539
rect 877 1505 911 1539
rect 949 1505 983 1539
rect 1021 1505 1055 1539
rect 1165 1505 1199 1539
rect 1237 1505 1271 1539
rect 1315 1505 1349 1539
rect 1393 1505 1427 1539
rect 1465 1505 1499 1539
rect 1609 1505 1643 1539
rect 1681 1505 1715 1539
rect 1753 1505 1787 1539
rect 1825 1505 1859 1539
rect 1915 1505 1949 1539
rect 1987 1505 2021 1539
rect 2059 1505 2093 1539
rect 2131 1505 2165 1539
rect 2275 1505 2309 1539
rect 2347 1505 2381 1539
rect 2425 1505 2459 1539
rect 2503 1505 2537 1539
rect 2575 1505 2609 1539
rect 2719 1505 2753 1539
rect 2791 1505 2825 1539
rect 2863 1505 2897 1539
rect 2935 1505 2969 1539
rect 3025 1505 3059 1539
rect 3097 1505 3131 1539
rect 3169 1505 3203 1539
rect 3241 1505 3275 1539
rect 3385 1505 3419 1539
rect 3457 1505 3491 1539
rect 3529 1505 3563 1539
rect 3601 1505 3635 1539
rect 3691 1505 3725 1539
rect 3763 1505 3797 1539
rect 3835 1505 3869 1539
rect 3907 1505 3941 1539
rect -461 1436 -427 1470
rect -461 1364 -427 1398
rect -461 1292 -427 1326
rect -461 1220 -427 1254
rect -461 1148 -427 1182
rect -461 1076 -427 1110
rect -17 1436 17 1470
rect -17 1364 17 1398
rect -17 1292 17 1326
rect -17 1220 17 1254
rect -17 1148 17 1182
rect -17 1076 17 1110
rect -461 1004 -427 1038
rect -461 932 -427 966
rect 427 1436 461 1470
rect 427 1364 461 1398
rect 427 1292 461 1326
rect 427 1220 461 1254
rect 427 1148 461 1182
rect 427 1076 461 1110
rect -17 1004 17 1038
rect -17 932 17 966
rect 1093 1436 1127 1470
rect 1093 1364 1127 1398
rect 1093 1292 1127 1326
rect 1093 1220 1127 1254
rect 1093 1148 1127 1182
rect 1093 1076 1127 1110
rect 427 1004 461 1038
rect 427 932 461 966
rect 1537 1436 1571 1470
rect 1537 1364 1571 1398
rect 1537 1292 1571 1326
rect 1537 1220 1571 1254
rect 1537 1148 1571 1182
rect 1537 1076 1571 1110
rect 1093 1004 1127 1038
rect 1093 932 1127 966
rect 2203 1436 2237 1470
rect 2203 1364 2237 1398
rect 2203 1292 2237 1326
rect 2203 1220 2237 1254
rect 2203 1148 2237 1182
rect 2203 1076 2237 1110
rect 1537 1004 1571 1038
rect 1537 932 1571 966
rect 2647 1436 2681 1470
rect 2647 1364 2681 1398
rect 2647 1292 2681 1326
rect 2647 1220 2681 1254
rect 2647 1148 2681 1182
rect 2647 1076 2681 1110
rect 2203 1004 2237 1038
rect 2203 932 2237 966
rect 3313 1436 3347 1470
rect 3313 1364 3347 1398
rect 3313 1292 3347 1326
rect 3313 1220 3347 1254
rect 3313 1148 3347 1182
rect 3313 1076 3347 1110
rect 2647 1004 2681 1038
rect 2647 932 2681 966
rect 3979 1436 4013 1470
rect 3979 1364 4013 1398
rect 3979 1292 4013 1326
rect 3979 1220 4013 1254
rect 3979 1148 4013 1182
rect 3979 1076 4013 1110
rect 3313 1004 3347 1038
rect 3313 932 3347 966
rect 3979 1004 4013 1038
rect 3979 932 4013 966
<< poly >>
rect -281 1450 -251 1476
rect -193 1450 -163 1476
rect 163 1450 193 1476
rect 251 1450 281 1476
rect -281 1019 -251 1050
rect -193 1019 -163 1050
rect -323 1003 -163 1019
rect -323 969 -313 1003
rect -279 989 -163 1003
rect 631 1450 661 1476
rect 719 1450 749 1476
rect 807 1450 837 1476
rect 895 1450 925 1476
rect 163 1019 193 1050
rect 251 1019 281 1050
rect -279 969 -269 989
rect -323 953 -269 969
rect 121 1003 281 1019
rect 121 969 131 1003
rect 165 989 281 1003
rect 1273 1450 1303 1476
rect 1361 1450 1391 1476
rect 165 969 175 989
rect 121 953 175 969
rect 631 1019 661 1050
rect 719 1019 749 1050
rect 807 1019 837 1050
rect 895 1019 925 1050
rect 631 1003 749 1019
rect 631 989 649 1003
rect 639 969 649 989
rect 683 989 749 1003
rect 793 1003 925 1019
rect 683 969 693 989
rect 639 953 693 969
rect 793 969 803 1003
rect 837 989 925 1003
rect 1741 1450 1771 1476
rect 1829 1450 1859 1476
rect 1917 1450 1947 1476
rect 2005 1450 2035 1476
rect 1273 1019 1303 1050
rect 1361 1019 1391 1050
rect 837 969 847 989
rect 793 953 847 969
rect 1231 1003 1391 1019
rect 1231 969 1241 1003
rect 1275 989 1391 1003
rect 2383 1450 2413 1476
rect 2471 1450 2501 1476
rect 1275 969 1285 989
rect 1231 953 1285 969
rect 1741 1019 1771 1050
rect 1829 1019 1859 1050
rect 1917 1019 1947 1050
rect 2005 1019 2035 1050
rect 1741 1003 1859 1019
rect 1741 989 1759 1003
rect 1749 969 1759 989
rect 1793 989 1859 1003
rect 1903 1003 2035 1019
rect 1793 969 1803 989
rect 1749 953 1803 969
rect 1903 969 1913 1003
rect 1947 989 2035 1003
rect 2851 1451 2881 1477
rect 2939 1451 2969 1477
rect 3027 1451 3057 1477
rect 3115 1451 3145 1477
rect 2383 1019 2413 1050
rect 2471 1019 2501 1050
rect 1947 969 1957 989
rect 1903 953 1957 969
rect 2341 1003 2501 1019
rect 2341 969 2351 1003
rect 2385 989 2501 1003
rect 3517 1451 3547 1477
rect 3605 1451 3635 1477
rect 3693 1451 3723 1477
rect 3781 1451 3811 1477
rect 2851 1020 2881 1051
rect 2939 1020 2969 1051
rect 3027 1020 3057 1051
rect 3115 1020 3145 1051
rect 2385 969 2395 989
rect 2341 953 2395 969
rect 2828 1004 2969 1020
rect 2828 970 2838 1004
rect 2872 990 2969 1004
rect 3014 1004 3145 1020
rect 2872 970 2882 990
rect 2828 954 2882 970
rect 3014 970 3024 1004
rect 3058 990 3145 1004
rect 3517 1020 3547 1051
rect 3605 1020 3635 1051
rect 3693 1020 3723 1051
rect 3781 1020 3811 1051
rect 3058 970 3068 990
rect 3014 954 3068 970
rect 3494 1004 3635 1020
rect 3494 970 3504 1004
rect 3538 990 3635 1004
rect 3680 1004 3811 1020
rect 3538 970 3548 990
rect 3494 954 3548 970
rect 3680 970 3690 1004
rect 3724 990 3811 1004
rect 3724 970 3734 990
rect 3680 954 3734 970
rect -323 461 -269 477
rect -323 427 -313 461
rect -279 441 -269 461
rect -279 427 -259 441
rect -323 411 -259 427
rect -289 377 -259 411
rect 121 461 175 477
rect 121 427 131 461
rect 165 441 175 461
rect 165 427 185 441
rect 121 411 185 427
rect 155 377 185 411
rect 639 461 693 477
rect 639 441 649 461
rect 612 427 649 441
rect 683 427 693 461
rect 612 411 693 427
rect 787 461 841 477
rect 787 427 797 461
rect 831 427 841 461
rect 787 411 841 427
rect 612 377 642 411
rect 806 377 836 411
rect 1231 461 1285 477
rect 1231 427 1241 461
rect 1275 441 1285 461
rect 1275 427 1295 441
rect 1231 411 1295 427
rect 1265 377 1295 411
rect 1749 461 1803 477
rect 1749 441 1759 461
rect 1722 427 1759 441
rect 1793 427 1803 461
rect 1722 411 1803 427
rect 1897 461 1951 477
rect 1897 427 1907 461
rect 1941 427 1951 461
rect 1897 411 1951 427
rect 1722 377 1752 411
rect 1916 377 1946 411
rect 2341 461 2395 477
rect 2341 427 2351 461
rect 2385 441 2395 461
rect 2385 427 2405 441
rect 2341 411 2405 427
rect 2375 377 2405 411
rect 2859 461 2913 477
rect 2859 441 2869 461
rect 2832 427 2869 441
rect 2903 427 2913 461
rect 2832 411 2913 427
rect 3007 461 3061 477
rect 3007 427 3017 461
rect 3051 427 3061 461
rect 3007 411 3061 427
rect 3525 461 3579 477
rect 3525 441 3535 461
rect 2832 377 2862 411
rect 3026 377 3056 411
rect 3498 427 3535 441
rect 3569 427 3579 461
rect 3498 411 3579 427
rect 3673 461 3727 477
rect 3673 427 3683 461
rect 3717 427 3727 461
rect 3673 411 3727 427
rect 3498 377 3528 411
rect 3692 377 3722 411
<< polycont >>
rect -313 969 -279 1003
rect 131 969 165 1003
rect 649 969 683 1003
rect 803 969 837 1003
rect 1241 969 1275 1003
rect 1759 969 1793 1003
rect 1913 969 1947 1003
rect 2351 969 2385 1003
rect 2838 970 2872 1004
rect 3024 970 3058 1004
rect 3504 970 3538 1004
rect 3690 970 3724 1004
rect -313 427 -279 461
rect 131 427 165 461
rect 649 427 683 461
rect 797 427 831 461
rect 1241 427 1275 461
rect 1759 427 1793 461
rect 1907 427 1941 461
rect 2351 427 2385 461
rect 2869 427 2903 461
rect 3017 427 3051 461
rect 3535 427 3569 461
rect 3683 427 3717 461
<< locali >>
rect -475 1539 4027 1554
rect -475 1505 -389 1539
rect -355 1505 -317 1539
rect -283 1505 -239 1539
rect -205 1505 -161 1539
rect -127 1505 -89 1539
rect -55 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 205 1539
rect 239 1505 283 1539
rect 317 1505 355 1539
rect 389 1505 499 1539
rect 533 1505 571 1539
rect 605 1505 643 1539
rect 677 1505 715 1539
rect 749 1505 805 1539
rect 839 1505 877 1539
rect 911 1505 949 1539
rect 983 1505 1021 1539
rect 1055 1505 1165 1539
rect 1199 1505 1237 1539
rect 1271 1505 1315 1539
rect 1349 1505 1393 1539
rect 1427 1505 1465 1539
rect 1499 1505 1609 1539
rect 1643 1505 1681 1539
rect 1715 1505 1753 1539
rect 1787 1505 1825 1539
rect 1859 1505 1915 1539
rect 1949 1505 1987 1539
rect 2021 1505 2059 1539
rect 2093 1505 2131 1539
rect 2165 1505 2275 1539
rect 2309 1505 2347 1539
rect 2381 1505 2425 1539
rect 2459 1505 2503 1539
rect 2537 1505 2575 1539
rect 2609 1505 2719 1539
rect 2753 1505 2791 1539
rect 2825 1505 2863 1539
rect 2897 1505 2935 1539
rect 2969 1505 3025 1539
rect 3059 1505 3097 1539
rect 3131 1505 3169 1539
rect 3203 1505 3241 1539
rect 3275 1505 3385 1539
rect 3419 1505 3457 1539
rect 3491 1505 3529 1539
rect 3563 1505 3601 1539
rect 3635 1505 3691 1539
rect 3725 1505 3763 1539
rect 3797 1505 3835 1539
rect 3869 1505 3907 1539
rect 3941 1505 4027 1539
rect -475 1492 4027 1505
rect -475 1470 -413 1492
rect -475 1436 -461 1470
rect -427 1436 -413 1470
rect -475 1398 -413 1436
rect -475 1364 -461 1398
rect -427 1364 -413 1398
rect -475 1326 -413 1364
rect -475 1292 -461 1326
rect -427 1292 -413 1326
rect -475 1254 -413 1292
rect -475 1220 -461 1254
rect -427 1220 -413 1254
rect -475 1182 -413 1220
rect -475 1148 -461 1182
rect -427 1148 -413 1182
rect -475 1110 -413 1148
rect -475 1076 -461 1110
rect -427 1076 -413 1110
rect -327 1412 -293 1492
rect -327 1344 -293 1378
rect -327 1276 -293 1310
rect -327 1208 -293 1242
rect -327 1139 -293 1174
rect -327 1083 -293 1105
rect -239 1412 -205 1450
rect -239 1344 -205 1378
rect -239 1276 -205 1310
rect -239 1208 -205 1242
rect -239 1139 -205 1174
rect -475 1038 -413 1076
rect -475 1004 -461 1038
rect -427 1004 -413 1038
rect -475 966 -413 1004
rect -475 932 -461 966
rect -427 932 -413 966
rect -475 868 -413 932
rect -313 1003 -279 1019
rect -313 609 -279 969
rect -239 979 -205 1105
rect -151 1412 -117 1492
rect -151 1344 -117 1378
rect -151 1276 -117 1310
rect -151 1208 -117 1242
rect -151 1139 -117 1174
rect -151 1083 -117 1105
rect -31 1470 31 1492
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect 117 1412 151 1492
rect 117 1344 151 1378
rect 117 1276 151 1310
rect 117 1208 151 1242
rect 117 1139 151 1174
rect 117 1083 151 1105
rect 205 1412 239 1450
rect 205 1344 239 1378
rect 205 1276 239 1310
rect 205 1208 239 1242
rect 205 1139 239 1174
rect -31 1038 31 1076
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -239 945 -131 979
rect -475 546 -413 572
rect -475 512 -461 546
rect -427 512 -413 546
rect -475 474 -413 512
rect -475 440 -461 474
rect -427 440 -413 474
rect -475 402 -413 440
rect -313 461 -279 575
rect -165 609 -131 945
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect -31 868 31 932
rect 131 1003 165 1019
rect -165 461 -131 575
rect 131 831 165 969
rect 205 979 239 1105
rect 293 1412 327 1492
rect 293 1344 327 1378
rect 293 1276 327 1310
rect 293 1208 327 1242
rect 293 1139 327 1174
rect 293 1083 327 1105
rect 413 1470 475 1492
rect 413 1436 427 1470
rect 461 1436 475 1470
rect 413 1398 475 1436
rect 413 1364 427 1398
rect 461 1364 475 1398
rect 413 1326 475 1364
rect 413 1292 427 1326
rect 461 1292 475 1326
rect 413 1254 475 1292
rect 413 1220 427 1254
rect 461 1220 475 1254
rect 413 1182 475 1220
rect 413 1148 427 1182
rect 461 1148 475 1182
rect 413 1110 475 1148
rect 413 1076 427 1110
rect 461 1076 475 1110
rect 413 1038 475 1076
rect 585 1412 619 1492
rect 585 1344 619 1378
rect 585 1276 619 1310
rect 585 1208 619 1242
rect 585 1139 619 1174
rect 585 1073 619 1105
rect 673 1412 707 1450
rect 673 1344 707 1378
rect 673 1276 707 1310
rect 673 1208 707 1242
rect 673 1139 707 1174
rect 761 1412 795 1492
rect 761 1344 795 1378
rect 761 1276 795 1310
rect 761 1208 795 1242
rect 761 1157 795 1174
rect 849 1412 883 1450
rect 849 1344 883 1378
rect 849 1276 883 1310
rect 849 1208 883 1242
rect 673 1103 707 1105
rect 849 1139 883 1174
rect 937 1412 971 1492
rect 937 1344 971 1378
rect 937 1276 971 1310
rect 937 1208 971 1242
rect 937 1157 971 1174
rect 1079 1470 1141 1492
rect 1079 1436 1093 1470
rect 1127 1436 1141 1470
rect 1079 1398 1141 1436
rect 1079 1364 1093 1398
rect 1127 1364 1141 1398
rect 1079 1326 1141 1364
rect 1079 1292 1093 1326
rect 1127 1292 1141 1326
rect 1079 1254 1141 1292
rect 1079 1220 1093 1254
rect 1127 1220 1141 1254
rect 1079 1182 1141 1220
rect 849 1103 883 1105
rect 1079 1148 1093 1182
rect 1127 1148 1141 1182
rect 1079 1110 1141 1148
rect 673 1069 979 1103
rect 413 1004 427 1038
rect 461 1004 475 1038
rect 205 945 313 979
rect -313 411 -279 427
rect -239 427 -131 461
rect -31 546 31 572
rect -31 512 -17 546
rect 17 512 31 546
rect -31 474 31 512
rect -31 440 -17 474
rect 17 440 31 474
rect -475 368 -461 402
rect -427 368 -413 402
rect -475 330 -413 368
rect -475 296 -461 330
rect -427 296 -413 330
rect -475 258 -413 296
rect -475 224 -461 258
rect -427 224 -413 258
rect -475 186 -413 224
rect -475 152 -461 186
rect -427 152 -413 186
rect -475 114 -413 152
rect -475 80 -461 114
rect -427 80 -413 114
rect -475 62 -413 80
rect -335 361 -301 377
rect -335 289 -301 327
rect -335 221 -301 255
rect -239 245 -205 427
rect -31 402 31 440
rect 131 461 165 797
rect 279 757 313 945
rect 413 966 475 1004
rect 413 932 427 966
rect 461 932 475 966
rect 413 868 475 932
rect 649 1003 683 1019
rect 803 1003 837 1019
rect 279 461 313 723
rect 649 757 683 969
rect 131 411 165 427
rect 205 427 313 461
rect 413 546 475 572
rect 413 512 427 546
rect 461 512 475 546
rect 413 474 475 512
rect 413 440 427 474
rect 461 440 475 474
rect -239 195 -205 211
rect -141 361 -107 377
rect -141 289 -107 327
rect -141 221 -107 255
rect -335 151 -301 187
rect -141 151 -107 187
rect -301 117 -239 151
rect -205 117 -141 151
rect -335 62 -301 117
rect -238 62 -204 117
rect -141 62 -107 117
rect -31 368 -17 402
rect 17 368 31 402
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect -31 62 31 80
rect 109 361 143 377
rect 109 289 143 327
rect 109 221 143 255
rect 205 245 239 427
rect 413 402 475 440
rect 649 461 683 723
rect 649 411 683 427
rect 797 969 803 988
rect 797 953 837 969
rect 797 609 831 953
rect 797 461 831 575
rect 797 411 831 427
rect 945 683 979 1069
rect 1079 1076 1093 1110
rect 1127 1076 1141 1110
rect 1227 1412 1261 1492
rect 1227 1344 1261 1378
rect 1227 1276 1261 1310
rect 1227 1208 1261 1242
rect 1227 1139 1261 1174
rect 1227 1083 1261 1105
rect 1315 1412 1349 1450
rect 1315 1344 1349 1378
rect 1315 1276 1349 1310
rect 1315 1208 1349 1242
rect 1315 1139 1349 1174
rect 1079 1038 1141 1076
rect 1079 1004 1093 1038
rect 1127 1004 1141 1038
rect 1079 966 1141 1004
rect 1079 932 1093 966
rect 1127 932 1141 966
rect 1079 868 1141 932
rect 1241 1003 1275 1019
rect 205 195 239 211
rect 303 361 337 377
rect 303 289 337 327
rect 303 221 337 255
rect 109 151 143 187
rect 303 151 337 187
rect 143 117 205 151
rect 239 117 303 151
rect 109 62 143 117
rect 206 62 240 117
rect 303 62 337 117
rect 413 368 427 402
rect 461 368 475 402
rect 413 330 475 368
rect 413 296 427 330
rect 461 296 475 330
rect 413 258 475 296
rect 413 224 427 258
rect 461 224 475 258
rect 413 186 475 224
rect 413 152 427 186
rect 461 152 475 186
rect 413 114 475 152
rect 413 80 427 114
rect 461 80 475 114
rect 566 361 600 377
rect 760 361 794 377
rect 945 376 979 649
rect 1241 683 1275 969
rect 1315 979 1349 1105
rect 1403 1412 1437 1492
rect 1403 1344 1437 1378
rect 1403 1276 1437 1310
rect 1403 1208 1437 1242
rect 1403 1139 1437 1174
rect 1403 1083 1437 1105
rect 1523 1470 1585 1492
rect 1523 1436 1537 1470
rect 1571 1436 1585 1470
rect 1523 1398 1585 1436
rect 1523 1364 1537 1398
rect 1571 1364 1585 1398
rect 1523 1326 1585 1364
rect 1523 1292 1537 1326
rect 1571 1292 1585 1326
rect 1523 1254 1585 1292
rect 1523 1220 1537 1254
rect 1571 1220 1585 1254
rect 1523 1182 1585 1220
rect 1523 1148 1537 1182
rect 1571 1148 1585 1182
rect 1523 1110 1585 1148
rect 1523 1076 1537 1110
rect 1571 1076 1585 1110
rect 1523 1038 1585 1076
rect 1695 1412 1729 1492
rect 1695 1344 1729 1378
rect 1695 1276 1729 1310
rect 1695 1208 1729 1242
rect 1695 1139 1729 1174
rect 1695 1073 1729 1105
rect 1783 1412 1817 1450
rect 1783 1344 1817 1378
rect 1783 1276 1817 1310
rect 1783 1208 1817 1242
rect 1783 1139 1817 1174
rect 1871 1412 1905 1492
rect 1871 1344 1905 1378
rect 1871 1276 1905 1310
rect 1871 1208 1905 1242
rect 1871 1157 1905 1174
rect 1959 1412 1993 1450
rect 1959 1344 1993 1378
rect 1959 1276 1993 1310
rect 1959 1208 1993 1242
rect 1783 1103 1817 1105
rect 1959 1139 1993 1174
rect 2047 1412 2081 1492
rect 2047 1344 2081 1378
rect 2047 1276 2081 1310
rect 2047 1208 2081 1242
rect 2047 1157 2081 1174
rect 2189 1470 2251 1492
rect 2189 1436 2203 1470
rect 2237 1436 2251 1470
rect 2189 1398 2251 1436
rect 2189 1364 2203 1398
rect 2237 1364 2251 1398
rect 2189 1326 2251 1364
rect 2189 1292 2203 1326
rect 2237 1292 2251 1326
rect 2189 1254 2251 1292
rect 2189 1220 2203 1254
rect 2237 1220 2251 1254
rect 2189 1182 2251 1220
rect 1959 1103 1993 1105
rect 2189 1148 2203 1182
rect 2237 1148 2251 1182
rect 2189 1110 2251 1148
rect 1783 1069 2089 1103
rect 1523 1004 1537 1038
rect 1571 1004 1585 1038
rect 1315 945 1423 979
rect 600 327 663 361
rect 697 327 760 361
rect 566 289 600 327
rect 566 221 600 255
rect 760 289 794 327
rect 566 151 600 187
rect 566 101 600 117
rect 663 236 697 252
rect 413 62 475 80
rect 663 62 697 202
rect 760 221 794 255
rect 857 342 979 376
rect 1079 546 1141 572
rect 1079 512 1093 546
rect 1127 512 1141 546
rect 1079 474 1141 512
rect 1079 440 1093 474
rect 1127 440 1141 474
rect 1079 402 1141 440
rect 1241 461 1275 649
rect 1389 757 1423 945
rect 1523 966 1585 1004
rect 1523 932 1537 966
rect 1571 932 1585 966
rect 1523 868 1585 932
rect 1759 1003 1793 1019
rect 1913 1003 1947 1019
rect 1389 461 1423 723
rect 1759 609 1793 969
rect 1241 411 1275 427
rect 1315 427 1423 461
rect 1523 546 1585 572
rect 1523 512 1537 546
rect 1571 512 1585 546
rect 1523 474 1585 512
rect 1523 440 1537 474
rect 1571 440 1585 474
rect 1079 368 1093 402
rect 1127 368 1141 402
rect 857 245 891 342
rect 1079 330 1141 368
rect 857 195 891 211
rect 954 289 988 305
rect 954 221 988 255
rect 760 151 794 187
rect 954 151 988 187
rect 794 117 857 151
rect 891 117 954 151
rect 760 101 794 117
rect 954 101 988 117
rect 1079 296 1093 330
rect 1127 296 1141 330
rect 1079 258 1141 296
rect 1079 224 1093 258
rect 1127 224 1141 258
rect 1079 186 1141 224
rect 1079 152 1093 186
rect 1127 152 1141 186
rect 1079 114 1141 152
rect 1079 80 1093 114
rect 1127 80 1141 114
rect 1079 62 1141 80
rect 1219 361 1253 377
rect 1219 289 1253 327
rect 1219 221 1253 255
rect 1315 245 1349 427
rect 1523 402 1585 440
rect 1759 461 1793 575
rect 1759 411 1793 427
rect 1907 969 1913 988
rect 1907 953 1947 969
rect 1907 831 1941 953
rect 1907 461 1941 797
rect 1907 411 1941 427
rect 2055 683 2089 1069
rect 2189 1076 2203 1110
rect 2237 1076 2251 1110
rect 2337 1412 2371 1492
rect 2337 1344 2371 1378
rect 2337 1276 2371 1310
rect 2337 1208 2371 1242
rect 2337 1139 2371 1174
rect 2337 1083 2371 1105
rect 2425 1412 2459 1450
rect 2425 1344 2459 1378
rect 2425 1276 2459 1310
rect 2425 1208 2459 1242
rect 2425 1139 2459 1174
rect 2189 1038 2251 1076
rect 2189 1004 2203 1038
rect 2237 1004 2251 1038
rect 2189 966 2251 1004
rect 2189 932 2203 966
rect 2237 932 2251 966
rect 2189 868 2251 932
rect 2351 1003 2385 1019
rect 1315 195 1349 211
rect 1413 361 1447 377
rect 1413 289 1447 327
rect 1413 221 1447 255
rect 1219 151 1253 187
rect 1413 151 1447 187
rect 1253 117 1315 151
rect 1349 117 1413 151
rect 1219 62 1253 117
rect 1316 62 1350 117
rect 1413 62 1447 117
rect 1523 368 1537 402
rect 1571 368 1585 402
rect 1523 330 1585 368
rect 1523 296 1537 330
rect 1571 296 1585 330
rect 1523 258 1585 296
rect 1523 224 1537 258
rect 1571 224 1585 258
rect 1523 186 1585 224
rect 1523 152 1537 186
rect 1571 152 1585 186
rect 1523 114 1585 152
rect 1523 80 1537 114
rect 1571 80 1585 114
rect 1676 361 1710 377
rect 1870 361 1904 377
rect 2055 376 2089 649
rect 2351 683 2385 969
rect 2425 979 2459 1105
rect 2513 1412 2547 1492
rect 2513 1344 2547 1378
rect 2513 1276 2547 1310
rect 2513 1208 2547 1242
rect 2513 1139 2547 1174
rect 2513 1083 2547 1105
rect 2633 1470 2695 1492
rect 2633 1436 2647 1470
rect 2681 1436 2695 1470
rect 2633 1398 2695 1436
rect 2633 1364 2647 1398
rect 2681 1364 2695 1398
rect 2633 1326 2695 1364
rect 2633 1292 2647 1326
rect 2681 1292 2695 1326
rect 2633 1254 2695 1292
rect 2633 1220 2647 1254
rect 2681 1220 2695 1254
rect 2633 1182 2695 1220
rect 2633 1148 2647 1182
rect 2681 1148 2695 1182
rect 2633 1110 2695 1148
rect 2633 1076 2647 1110
rect 2681 1076 2695 1110
rect 2633 1038 2695 1076
rect 2805 1411 2839 1451
rect 2805 1343 2839 1377
rect 2805 1275 2839 1309
rect 2805 1207 2839 1241
rect 2805 1139 2839 1173
rect 2893 1411 2927 1492
rect 3299 1470 3361 1492
rect 2893 1343 2927 1377
rect 2893 1275 2927 1309
rect 2893 1207 2927 1241
rect 2893 1157 2927 1173
rect 2981 1411 3191 1445
rect 2981 1343 3015 1377
rect 2981 1275 3015 1309
rect 2981 1207 3015 1241
rect 2981 1139 3015 1173
rect 2805 1071 3015 1105
rect 3069 1343 3103 1359
rect 3069 1275 3103 1309
rect 3069 1207 3103 1241
rect 3069 1139 3103 1173
rect 3157 1343 3191 1377
rect 3157 1275 3191 1309
rect 3157 1207 3191 1241
rect 3157 1157 3191 1173
rect 3299 1436 3313 1470
rect 3347 1436 3361 1470
rect 3299 1398 3361 1436
rect 3299 1364 3313 1398
rect 3347 1364 3361 1398
rect 3299 1326 3361 1364
rect 3299 1292 3313 1326
rect 3347 1292 3361 1326
rect 3299 1254 3361 1292
rect 3299 1220 3313 1254
rect 3347 1220 3361 1254
rect 3299 1182 3361 1220
rect 3299 1148 3313 1182
rect 3347 1148 3361 1182
rect 3299 1110 3361 1148
rect 3069 1071 3199 1105
rect 2633 1004 2647 1038
rect 2681 1004 2695 1038
rect 2425 945 2533 979
rect 1710 327 1773 361
rect 1807 327 1870 361
rect 1676 289 1710 327
rect 1676 221 1710 255
rect 1870 289 1904 327
rect 1676 151 1710 187
rect 1676 101 1710 117
rect 1773 236 1807 252
rect 1523 62 1585 80
rect 1773 62 1807 202
rect 1870 221 1904 255
rect 1967 342 2089 376
rect 2189 546 2251 572
rect 2189 512 2203 546
rect 2237 512 2251 546
rect 2189 474 2251 512
rect 2189 440 2203 474
rect 2237 440 2251 474
rect 2189 402 2251 440
rect 2351 461 2385 649
rect 2499 831 2533 945
rect 2633 966 2695 1004
rect 2633 932 2647 966
rect 2681 932 2695 966
rect 2838 1004 2872 1020
rect 3024 1004 3058 1020
rect 2872 970 2903 988
rect 2838 954 2903 970
rect 2633 868 2695 932
rect 2499 461 2533 797
rect 2869 757 2903 954
rect 2351 411 2385 427
rect 2425 427 2533 461
rect 2633 546 2695 572
rect 2633 512 2647 546
rect 2681 512 2695 546
rect 2633 474 2695 512
rect 2633 440 2647 474
rect 2681 440 2695 474
rect 2189 368 2203 402
rect 2237 368 2251 402
rect 1967 245 2001 342
rect 2189 330 2251 368
rect 1967 195 2001 211
rect 2064 289 2098 305
rect 2064 221 2098 255
rect 1870 151 1904 187
rect 2064 151 2098 187
rect 1904 117 1967 151
rect 2001 117 2064 151
rect 1870 101 1904 117
rect 2064 101 2098 117
rect 2189 296 2203 330
rect 2237 296 2251 330
rect 2189 258 2251 296
rect 2189 224 2203 258
rect 2237 224 2251 258
rect 2189 186 2251 224
rect 2189 152 2203 186
rect 2237 152 2251 186
rect 2189 114 2251 152
rect 2189 80 2203 114
rect 2237 80 2251 114
rect 2189 62 2251 80
rect 2329 361 2363 377
rect 2329 289 2363 327
rect 2329 221 2363 255
rect 2425 245 2459 427
rect 2633 402 2695 440
rect 2869 461 2903 723
rect 2869 411 2903 427
rect 3017 970 3024 988
rect 3017 954 3058 970
rect 3017 757 3051 954
rect 3017 461 3051 723
rect 3017 411 3051 427
rect 3165 683 3199 1071
rect 3299 1076 3313 1110
rect 3347 1076 3361 1110
rect 3299 1038 3361 1076
rect 3471 1411 3505 1451
rect 3471 1343 3505 1377
rect 3471 1275 3505 1309
rect 3471 1207 3505 1241
rect 3471 1139 3505 1173
rect 3559 1411 3593 1492
rect 3965 1470 4027 1492
rect 3559 1343 3593 1377
rect 3559 1275 3593 1309
rect 3559 1207 3593 1241
rect 3559 1157 3593 1173
rect 3647 1411 3857 1445
rect 3647 1343 3681 1377
rect 3647 1275 3681 1309
rect 3647 1207 3681 1241
rect 3647 1139 3681 1173
rect 3471 1071 3681 1105
rect 3735 1343 3769 1359
rect 3735 1275 3769 1309
rect 3735 1207 3769 1241
rect 3735 1139 3769 1173
rect 3823 1343 3857 1377
rect 3823 1275 3857 1309
rect 3823 1207 3857 1241
rect 3823 1157 3857 1173
rect 3965 1436 3979 1470
rect 4013 1436 4027 1470
rect 3965 1398 4027 1436
rect 3965 1364 3979 1398
rect 4013 1364 4027 1398
rect 3965 1326 4027 1364
rect 3965 1292 3979 1326
rect 4013 1292 4027 1326
rect 3965 1254 4027 1292
rect 3965 1220 3979 1254
rect 4013 1220 4027 1254
rect 3965 1182 4027 1220
rect 3965 1148 3979 1182
rect 4013 1148 4027 1182
rect 3965 1110 4027 1148
rect 3735 1071 3865 1105
rect 3299 1004 3313 1038
rect 3347 1004 3361 1038
rect 3299 966 3361 1004
rect 3299 932 3313 966
rect 3347 932 3361 966
rect 3504 1004 3538 1020
rect 3690 1004 3724 1020
rect 3538 970 3569 988
rect 3504 954 3569 970
rect 3299 868 3361 932
rect 2425 195 2459 211
rect 2523 361 2557 377
rect 2523 289 2557 327
rect 2523 221 2557 255
rect 2329 151 2363 187
rect 2523 151 2557 187
rect 2363 117 2425 151
rect 2459 117 2523 151
rect 2329 62 2363 117
rect 2426 62 2460 117
rect 2523 62 2557 117
rect 2633 368 2647 402
rect 2681 368 2695 402
rect 2633 330 2695 368
rect 2633 296 2647 330
rect 2681 296 2695 330
rect 2633 258 2695 296
rect 2633 224 2647 258
rect 2681 224 2695 258
rect 2633 186 2695 224
rect 2633 152 2647 186
rect 2681 152 2695 186
rect 2633 114 2695 152
rect 2633 80 2647 114
rect 2681 80 2695 114
rect 2633 62 2695 80
rect 2786 361 2820 377
rect 3165 376 3199 649
rect 3535 683 3569 954
rect 2786 289 2820 327
rect 2786 221 2820 255
rect 2883 342 3199 376
rect 3299 546 3361 572
rect 3299 512 3313 546
rect 3347 512 3361 546
rect 3299 474 3361 512
rect 3299 440 3313 474
rect 3347 440 3361 474
rect 3299 402 3361 440
rect 3535 461 3569 649
rect 3535 411 3569 427
rect 3683 970 3690 988
rect 3683 954 3724 970
rect 3683 831 3717 954
rect 3683 461 3717 797
rect 3683 411 3717 427
rect 3831 757 3865 1071
rect 3965 1076 3979 1110
rect 4013 1076 4027 1110
rect 3965 1038 4027 1076
rect 3965 1004 3979 1038
rect 4013 1004 4027 1038
rect 3965 966 4027 1004
rect 3965 932 3979 966
rect 4013 932 4027 966
rect 3965 868 4027 932
rect 3299 368 3313 402
rect 3347 368 3361 402
rect 2883 245 2917 342
rect 2883 195 2917 211
rect 2980 289 3014 306
rect 2980 221 3014 255
rect 2786 151 2820 187
rect 3077 245 3111 342
rect 3299 330 3361 368
rect 3077 195 3111 211
rect 3174 289 3208 306
rect 3174 221 3208 255
rect 2980 151 3014 187
rect 3174 151 3208 187
rect 2820 117 2883 151
rect 2917 117 2980 151
rect 3014 117 3077 151
rect 3111 117 3174 151
rect 2786 62 2820 117
rect 2883 62 2917 117
rect 2980 62 3014 117
rect 3077 62 3111 117
rect 3174 62 3208 117
rect 3299 296 3313 330
rect 3347 296 3361 330
rect 3299 258 3361 296
rect 3299 224 3313 258
rect 3347 224 3361 258
rect 3299 186 3361 224
rect 3299 152 3313 186
rect 3347 152 3361 186
rect 3299 114 3361 152
rect 3299 80 3313 114
rect 3347 80 3361 114
rect 3299 62 3361 80
rect 3452 361 3486 377
rect 3831 376 3865 723
rect 3452 289 3486 327
rect 3452 221 3486 255
rect 3549 342 3865 376
rect 3965 546 4027 572
rect 3965 512 3979 546
rect 4013 512 4027 546
rect 3965 474 4027 512
rect 3965 440 3979 474
rect 4013 440 4027 474
rect 3965 402 4027 440
rect 3965 368 3979 402
rect 4013 368 4027 402
rect 3549 245 3583 342
rect 3549 195 3583 211
rect 3646 289 3680 306
rect 3646 221 3680 255
rect 3452 151 3486 187
rect 3743 245 3777 342
rect 3965 330 4027 368
rect 3743 195 3777 211
rect 3840 289 3874 306
rect 3840 221 3874 255
rect 3646 151 3680 187
rect 3840 151 3874 187
rect 3486 117 3549 151
rect 3583 117 3646 151
rect 3680 117 3743 151
rect 3777 117 3840 151
rect 3452 62 3486 117
rect 3549 62 3583 117
rect 3646 62 3680 117
rect 3743 62 3777 117
rect 3840 62 3874 117
rect 3965 296 3979 330
rect 4013 296 4027 330
rect 3965 258 4027 296
rect 3965 224 3979 258
rect 4013 224 4027 258
rect 3965 186 4027 224
rect 3965 152 3979 186
rect 4013 152 4027 186
rect 3965 114 4027 152
rect 3965 80 3979 114
rect 4013 80 4027 114
rect 3965 62 4027 80
rect -475 47 4027 62
rect -475 13 -389 47
rect -355 13 -317 47
rect -283 13 -239 47
rect -205 13 -161 47
rect -127 13 -89 47
rect -55 13 55 47
rect 89 13 127 47
rect 161 13 205 47
rect 239 13 283 47
rect 317 13 355 47
rect 389 13 499 47
rect 533 13 571 47
rect 605 13 643 47
rect 677 13 715 47
rect 749 13 805 47
rect 839 13 877 47
rect 911 13 949 47
rect 983 13 1021 47
rect 1055 13 1165 47
rect 1199 13 1237 47
rect 1271 13 1315 47
rect 1349 13 1393 47
rect 1427 13 1465 47
rect 1499 13 1609 47
rect 1643 13 1681 47
rect 1715 13 1753 47
rect 1787 13 1825 47
rect 1859 13 1915 47
rect 1949 13 1987 47
rect 2021 13 2059 47
rect 2093 13 2131 47
rect 2165 13 2275 47
rect 2309 13 2347 47
rect 2381 13 2425 47
rect 2459 13 2503 47
rect 2537 13 2575 47
rect 2609 13 2719 47
rect 2753 13 2791 47
rect 2825 13 2863 47
rect 2897 13 2935 47
rect 2969 13 3025 47
rect 3059 13 3097 47
rect 3131 13 3169 47
rect 3203 13 3241 47
rect 3275 13 3385 47
rect 3419 13 3457 47
rect 3491 13 3529 47
rect 3563 13 3601 47
rect 3635 13 3691 47
rect 3725 13 3763 47
rect 3797 13 3835 47
rect 3869 13 3907 47
rect 3941 13 4027 47
rect -475 0 4027 13
<< viali >>
rect -389 1505 -355 1539
rect -317 1505 -283 1539
rect -239 1505 -205 1539
rect -161 1505 -127 1539
rect -89 1505 -55 1539
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 205 1505 239 1539
rect 283 1505 317 1539
rect 355 1505 389 1539
rect 499 1505 533 1539
rect 571 1505 605 1539
rect 643 1505 677 1539
rect 715 1505 749 1539
rect 805 1505 839 1539
rect 877 1505 911 1539
rect 949 1505 983 1539
rect 1021 1505 1055 1539
rect 1165 1505 1199 1539
rect 1237 1505 1271 1539
rect 1315 1505 1349 1539
rect 1393 1505 1427 1539
rect 1465 1505 1499 1539
rect 1609 1505 1643 1539
rect 1681 1505 1715 1539
rect 1753 1505 1787 1539
rect 1825 1505 1859 1539
rect 1915 1505 1949 1539
rect 1987 1505 2021 1539
rect 2059 1505 2093 1539
rect 2131 1505 2165 1539
rect 2275 1505 2309 1539
rect 2347 1505 2381 1539
rect 2425 1505 2459 1539
rect 2503 1505 2537 1539
rect 2575 1505 2609 1539
rect 2719 1505 2753 1539
rect 2791 1505 2825 1539
rect 2863 1505 2897 1539
rect 2935 1505 2969 1539
rect 3025 1505 3059 1539
rect 3097 1505 3131 1539
rect 3169 1505 3203 1539
rect 3241 1505 3275 1539
rect 3385 1505 3419 1539
rect 3457 1505 3491 1539
rect 3529 1505 3563 1539
rect 3601 1505 3635 1539
rect 3691 1505 3725 1539
rect 3763 1505 3797 1539
rect 3835 1505 3869 1539
rect 3907 1505 3941 1539
rect -313 575 -279 609
rect -165 575 -131 609
rect 131 797 165 831
rect 279 723 313 757
rect 649 723 683 757
rect 797 575 831 609
rect 945 649 979 683
rect 1241 649 1275 683
rect 1389 723 1423 757
rect 1759 575 1793 609
rect 1907 797 1941 831
rect 2055 649 2089 683
rect 2351 649 2385 683
rect 2499 797 2533 831
rect 2869 723 2903 757
rect 3017 723 3051 757
rect 3165 649 3199 683
rect 3535 649 3569 683
rect 3683 797 3717 831
rect 3831 723 3865 757
rect -389 13 -355 47
rect -317 13 -283 47
rect -239 13 -205 47
rect -161 13 -127 47
rect -89 13 -55 47
rect 55 13 89 47
rect 127 13 161 47
rect 205 13 239 47
rect 283 13 317 47
rect 355 13 389 47
rect 499 13 533 47
rect 571 13 605 47
rect 643 13 677 47
rect 715 13 749 47
rect 805 13 839 47
rect 877 13 911 47
rect 949 13 983 47
rect 1021 13 1055 47
rect 1165 13 1199 47
rect 1237 13 1271 47
rect 1315 13 1349 47
rect 1393 13 1427 47
rect 1465 13 1499 47
rect 1609 13 1643 47
rect 1681 13 1715 47
rect 1753 13 1787 47
rect 1825 13 1859 47
rect 1915 13 1949 47
rect 1987 13 2021 47
rect 2059 13 2093 47
rect 2131 13 2165 47
rect 2275 13 2309 47
rect 2347 13 2381 47
rect 2425 13 2459 47
rect 2503 13 2537 47
rect 2575 13 2609 47
rect 2719 13 2753 47
rect 2791 13 2825 47
rect 2863 13 2897 47
rect 2935 13 2969 47
rect 3025 13 3059 47
rect 3097 13 3131 47
rect 3169 13 3203 47
rect 3241 13 3275 47
rect 3385 13 3419 47
rect 3457 13 3491 47
rect 3529 13 3563 47
rect 3601 13 3635 47
rect 3691 13 3725 47
rect 3763 13 3797 47
rect 3835 13 3869 47
rect 3907 13 3941 47
<< metal1 >>
rect -475 1539 4027 1554
rect -475 1505 -389 1539
rect -355 1505 -317 1539
rect -283 1505 -239 1539
rect -205 1505 -161 1539
rect -127 1505 -89 1539
rect -55 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 205 1539
rect 239 1505 283 1539
rect 317 1505 355 1539
rect 389 1505 499 1539
rect 533 1505 571 1539
rect 605 1505 643 1539
rect 677 1505 715 1539
rect 749 1505 805 1539
rect 839 1505 877 1539
rect 911 1505 949 1539
rect 983 1505 1021 1539
rect 1055 1505 1165 1539
rect 1199 1505 1237 1539
rect 1271 1505 1315 1539
rect 1349 1505 1393 1539
rect 1427 1505 1465 1539
rect 1499 1505 1609 1539
rect 1643 1505 1681 1539
rect 1715 1505 1753 1539
rect 1787 1505 1825 1539
rect 1859 1505 1915 1539
rect 1949 1505 1987 1539
rect 2021 1505 2059 1539
rect 2093 1505 2131 1539
rect 2165 1505 2275 1539
rect 2309 1505 2347 1539
rect 2381 1505 2425 1539
rect 2459 1505 2503 1539
rect 2537 1505 2575 1539
rect 2609 1505 2719 1539
rect 2753 1505 2791 1539
rect 2825 1505 2863 1539
rect 2897 1505 2935 1539
rect 2969 1505 3025 1539
rect 3059 1505 3097 1539
rect 3131 1505 3169 1539
rect 3203 1505 3241 1539
rect 3275 1505 3385 1539
rect 3419 1505 3457 1539
rect 3491 1505 3529 1539
rect 3563 1505 3601 1539
rect 3635 1505 3691 1539
rect 3725 1505 3763 1539
rect 3797 1505 3835 1539
rect 3869 1505 3907 1539
rect 3941 1505 4027 1539
rect -475 1492 4027 1505
rect 125 831 171 837
rect 1901 831 1947 837
rect 2493 831 2539 837
rect 3677 831 3723 837
rect 119 797 131 831
rect 165 797 1907 831
rect 1941 797 1953 831
rect 2487 797 2499 831
rect 2533 797 3683 831
rect 3717 797 3729 831
rect 125 791 171 797
rect 1901 791 1947 797
rect 2493 791 2539 797
rect 3677 791 3723 797
rect 273 757 319 763
rect 643 757 689 763
rect 1383 757 1429 763
rect 2863 757 2909 763
rect 3011 757 3057 763
rect 3825 757 3871 763
rect 267 723 279 757
rect 313 723 649 757
rect 683 723 695 757
rect 1377 723 1389 757
rect 1423 723 2869 757
rect 2903 723 2915 757
rect 3005 723 3017 757
rect 3051 723 3831 757
rect 3865 723 3877 757
rect 273 717 319 723
rect 643 717 689 723
rect 1383 717 1429 723
rect 2863 717 2909 723
rect 3011 717 3057 723
rect 3825 717 3871 723
rect 939 683 985 689
rect 1235 683 1281 689
rect 2049 683 2095 689
rect 2345 683 2391 689
rect 3159 683 3205 689
rect 3529 683 3575 689
rect 933 649 945 683
rect 979 649 1241 683
rect 1275 649 1287 683
rect 2043 649 2055 683
rect 2089 649 2351 683
rect 2385 649 2397 683
rect 3153 649 3165 683
rect 3199 649 3535 683
rect 3569 649 3581 683
rect 939 643 985 649
rect 1235 643 1281 649
rect 2049 643 2095 649
rect 2345 643 2391 649
rect 3159 643 3205 649
rect 3529 643 3575 649
rect -319 609 -273 615
rect -171 609 -125 615
rect 791 609 837 615
rect 1753 609 1799 615
rect -349 575 -313 609
rect -279 575 -267 609
rect -177 575 -165 609
rect -131 575 797 609
rect 831 575 1759 609
rect 1793 575 1805 609
rect -319 569 -273 575
rect -171 569 -125 575
rect 791 569 837 575
rect 1753 569 1799 575
rect -475 47 4027 62
rect -475 13 -389 47
rect -355 13 -317 47
rect -283 13 -239 47
rect -205 13 -161 47
rect -127 13 -89 47
rect -55 13 55 47
rect 89 13 127 47
rect 161 13 205 47
rect 239 13 283 47
rect 317 13 355 47
rect 389 13 499 47
rect 533 13 571 47
rect 605 13 643 47
rect 677 13 715 47
rect 749 13 805 47
rect 839 13 877 47
rect 911 13 949 47
rect 983 13 1021 47
rect 1055 13 1165 47
rect 1199 13 1237 47
rect 1271 13 1315 47
rect 1349 13 1393 47
rect 1427 13 1465 47
rect 1499 13 1609 47
rect 1643 13 1681 47
rect 1715 13 1753 47
rect 1787 13 1825 47
rect 1859 13 1915 47
rect 1949 13 1987 47
rect 2021 13 2059 47
rect 2093 13 2131 47
rect 2165 13 2275 47
rect 2309 13 2347 47
rect 2381 13 2425 47
rect 2459 13 2503 47
rect 2537 13 2575 47
rect 2609 13 2719 47
rect 2753 13 2791 47
rect 2825 13 2863 47
rect 2897 13 2935 47
rect 2969 13 3025 47
rect 3059 13 3097 47
rect 3131 13 3169 47
rect 3203 13 3241 47
rect 3275 13 3385 47
rect 3419 13 3457 47
rect 3491 13 3529 47
rect 3563 13 3601 47
rect 3635 13 3691 47
rect 3725 13 3763 47
rect 3797 13 3835 47
rect 3869 13 3907 47
rect 3941 13 4027 47
rect -475 0 4027 13
<< labels >>
rlabel metal1 3165 649 3199 683 1 Q
port 1 n
rlabel metal1 131 797 165 831 1 D
port 2 n
rlabel metal1 -313 575 -279 609 1 GATE_N
port 3 n
rlabel metal1 55 1505 89 1539 1 VDD
port 4 n
rlabel metal1 55 13 89 47 1 VSS
port 5 n
<< end >>
