* SPICE3 file created from AND3X1.ext - technology: sky130A

.subckt AND3X1 Y A B C VDD GND
M1000 VDD.t7 a_277_1050.t7 Y.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 VDD.t3 A.t0 a_277_1050.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 GND A.t1 a_91_103.t0 nshort w=-1.605u l=1.765u
+  ad=1.3199p pd=9.67u as=0p ps=0u
M1003 VDD.t2 B.t0 a_277_1050.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y a_277_1050.t9 GND.t1 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
M1005 VDD.t1 C.t1 a_277_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y.t2 a_277_1050.t8 VDD.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_277_1050.t6 A.t2 VDD.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_277_1050.t0 B.t2 VDD.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_277_1050.t5 C.t2 VDD.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 C B 0.18fF
C1 VDD B 0.05fF
C2 A B 0.18fF
C3 C VDD 0.06fF
C4 C A 0.02fF
C5 VDD Y 0.76fF
C6 VDD A 0.08fF
R0 a_277_1050.n5 a_277_1050.t7 512.525
R1 a_277_1050.n5 a_277_1050.t8 371.139
R2 a_277_1050.n6 a_277_1050.t9 210.434
R3 a_277_1050.n7 a_277_1050.n4 197.352
R4 a_277_1050.n9 a_277_1050.n7 193.073
R5 a_277_1050.n6 a_277_1050.n5 173.2
R6 a_277_1050.n7 a_277_1050.n6 153.043
R7 a_277_1050.n3 a_277_1050.n2 79.232
R8 a_277_1050.n4 a_277_1050.n3 63.152
R9 a_277_1050.n4 a_277_1050.n0 16.08
R10 a_277_1050.n3 a_277_1050.n1 16.08
R11 a_277_1050.n9 a_277_1050.n8 15.218
R12 a_277_1050.n0 a_277_1050.t1 14.282
R13 a_277_1050.n0 a_277_1050.t5 14.282
R14 a_277_1050.n1 a_277_1050.t2 14.282
R15 a_277_1050.n1 a_277_1050.t0 14.282
R16 a_277_1050.n2 a_277_1050.t4 14.282
R17 a_277_1050.n2 a_277_1050.t6 14.282
R18 a_277_1050.n10 a_277_1050.n9 12.014
R19 Y.n5 Y.n0 184.007
R20 Y.n5 Y.n4 179.015
R21 Y Y.n5 76
R22 Y.n4 Y.n3 30
R23 Y.n2 Y.n1 24.383
R24 Y.n4 Y.n2 23.684
R25 Y.n0 Y.t1 14.282
R26 Y.n0 Y.t2 14.282
R27 VDD.n68 VDD.n66 144.705
R28 VDD.n26 VDD.n25 77.792
R29 VDD.n35 VDD.n34 77.792
R30 VDD.n29 VDD.n23 76.145
R31 VDD.n29 VDD.n28 76
R32 VDD.n33 VDD.n32 76
R33 VDD.n39 VDD.n38 76
R34 VDD.n43 VDD.n42 76
R35 VDD.n70 VDD.n69 76
R36 VDD.n74 VDD.n73 76
R37 VDD.n78 VDD.n77 76
R38 VDD.n144 VDD.n143 76
R39 VDD.n139 VDD.n138 76
R40 VDD.n132 VDD.n131 76
R41 VDD.n127 VDD.n126 76
R42 VDD.n122 VDD.n121 76
R43 VDD.n115 VDD.n114 76
R44 VDD.n110 VDD.n109 76
R45 VDD.n105 VDD.n104 76
R46 VDD.n101 VDD.n100 76
R47 VDD.n141 VDD.n140 64.064
R48 VDD.n112 VDD.n111 59.488
R49 VDD.n106 VDD.t5 55.106
R50 VDD.n37 VDD.t6 55.106
R51 VDD.n24 VDD.t7 55.106
R52 VDD.n77 VDD.t1 55.106
R53 VDD.n117 VDD.n116 40.824
R54 VDD.n137 VDD.n136 40.824
R55 VDD.n59 VDD.n58 36.774
R56 VDD.n134 VDD.n133 27.456
R57 VDD.n119 VDD.n118 22.88
R58 VDD.n100 VDD.n97 21.841
R59 VDD.n23 VDD.n20 21.841
R60 VDD.n116 VDD.t0 14.282
R61 VDD.n116 VDD.t3 14.282
R62 VDD.n136 VDD.t4 14.282
R63 VDD.n136 VDD.t2 14.282
R64 VDD.n97 VDD.n80 14.167
R65 VDD.n80 VDD.n79 14.167
R66 VDD.n64 VDD.n45 14.167
R67 VDD.n45 VDD.n44 14.167
R68 VDD.n20 VDD.n19 14.167
R69 VDD.n19 VDD.n17 14.167
R70 VDD.n69 VDD.n65 14.167
R71 VDD.n124 VDD.n123 13.728
R72 VDD.n23 VDD.n22 13.653
R73 VDD.n22 VDD.n21 13.653
R74 VDD.n28 VDD.n27 13.653
R75 VDD.n27 VDD.n26 13.653
R76 VDD.n32 VDD.n31 13.653
R77 VDD.n31 VDD.n30 13.653
R78 VDD.n38 VDD.n36 13.653
R79 VDD.n36 VDD.n35 13.653
R80 VDD.n42 VDD.n41 13.653
R81 VDD.n41 VDD.n40 13.653
R82 VDD.n69 VDD.n68 13.653
R83 VDD.n68 VDD.n67 13.653
R84 VDD.n73 VDD.n72 13.653
R85 VDD.n72 VDD.n71 13.653
R86 VDD.n77 VDD.n76 13.653
R87 VDD.n76 VDD.n75 13.653
R88 VDD.n143 VDD.n142 13.653
R89 VDD.n142 VDD.n141 13.653
R90 VDD.n138 VDD.n135 13.653
R91 VDD.n135 VDD.n134 13.653
R92 VDD.n131 VDD.n130 13.653
R93 VDD.n130 VDD.n129 13.653
R94 VDD.n126 VDD.n125 13.653
R95 VDD.n125 VDD.n124 13.653
R96 VDD.n121 VDD.n120 13.653
R97 VDD.n120 VDD.n119 13.653
R98 VDD.n114 VDD.n113 13.653
R99 VDD.n113 VDD.n112 13.653
R100 VDD.n109 VDD.n108 13.653
R101 VDD.n108 VDD.n107 13.653
R102 VDD.n104 VDD.n103 13.653
R103 VDD.n103 VDD.n102 13.653
R104 VDD.n100 VDD.n99 13.653
R105 VDD.n99 VDD.n98 13.653
R106 VDD.n4 VDD.n2 12.915
R107 VDD.n4 VDD.n3 12.66
R108 VDD.n12 VDD.n11 12.343
R109 VDD.n10 VDD.n9 12.343
R110 VDD.n7 VDD.n6 12.343
R111 VDD.n129 VDD.n128 9.152
R112 VDD.n65 VDD.n64 7.674
R113 VDD.n49 VDD.n48 7.5
R114 VDD.n52 VDD.n51 7.5
R115 VDD.n54 VDD.n53 7.5
R116 VDD.n57 VDD.n56 7.5
R117 VDD.n64 VDD.n63 7.5
R118 VDD.n92 VDD.n91 7.5
R119 VDD.n86 VDD.n85 7.5
R120 VDD.n88 VDD.n87 7.5
R121 VDD.n94 VDD.n84 7.5
R122 VDD.n94 VDD.n82 7.5
R123 VDD.n97 VDD.n96 7.5
R124 VDD.n20 VDD.n16 7.5
R125 VDD.n2 VDD.n1 7.5
R126 VDD.n6 VDD.n5 7.5
R127 VDD.n9 VDD.n8 7.5
R128 VDD.n19 VDD.n18 7.5
R129 VDD.n14 VDD.n0 7.5
R130 VDD.n95 VDD.n81 6.772
R131 VDD.n93 VDD.n90 6.772
R132 VDD.n89 VDD.n86 6.772
R133 VDD.n89 VDD.n88 6.772
R134 VDD.n93 VDD.n92 6.772
R135 VDD.n96 VDD.n95 6.772
R136 VDD.n63 VDD.n62 6.772
R137 VDD.n50 VDD.n47 6.772
R138 VDD.n55 VDD.n52 6.772
R139 VDD.n60 VDD.n57 6.772
R140 VDD.n60 VDD.n59 6.772
R141 VDD.n55 VDD.n54 6.772
R142 VDD.n50 VDD.n49 6.772
R143 VDD.n62 VDD.n46 6.772
R144 VDD.n121 VDD.n117 6.69
R145 VDD.n16 VDD.n15 6.458
R146 VDD.n138 VDD.n137 6.296
R147 VDD.n84 VDD.n83 6.202
R148 VDD.n28 VDD.n24 1.967
R149 VDD.n38 VDD.n37 1.967
R150 VDD.n14 VDD.n7 1.329
R151 VDD.n14 VDD.n10 1.329
R152 VDD.n14 VDD.n12 1.329
R153 VDD.n14 VDD.n13 1.329
R154 VDD.n15 VDD.n14 0.696
R155 VDD.n14 VDD.n4 0.696
R156 VDD.n109 VDD.n106 0.393
R157 VDD.n94 VDD.n93 0.365
R158 VDD.n94 VDD.n89 0.365
R159 VDD.n95 VDD.n94 0.365
R160 VDD.n61 VDD.n60 0.365
R161 VDD.n61 VDD.n55 0.365
R162 VDD.n61 VDD.n50 0.365
R163 VDD.n62 VDD.n61 0.365
R164 VDD.n70 VDD.n43 0.29
R165 VDD.n101 VDD 0.207
R166 VDD.n132 VDD.n127 0.197
R167 VDD.n33 VDD.n29 0.157
R168 VDD.n39 VDD.n33 0.157
R169 VDD.n43 VDD.n39 0.145
R170 VDD.n74 VDD.n70 0.145
R171 VDD.n78 VDD.n74 0.145
R172 VDD.n144 VDD.n139 0.145
R173 VDD.n139 VDD.n132 0.145
R174 VDD.n127 VDD.n122 0.145
R175 VDD.n122 VDD.n115 0.145
R176 VDD.n115 VDD.n110 0.145
R177 VDD.n110 VDD.n105 0.145
R178 VDD.n105 VDD.n101 0.145
R179 VDD VDD.n78 0.086
R180 VDD VDD.n144 0.058
R181 A.n0 A.t0 512.525
R182 A.n0 A.t2 371.139
R183 A.n1 A.t1 314.221
R184 A.n1 A.n0 136.16
R185 A A.n1 76
R186 C.n0 C.t2 454.685
R187 C.n0 C.t1 428.979
R188 C.n1 C.t0 211.406
R189 C.n1 C.n0 125
R190 C C.n1 76
R191 a_372_210.n10 a_372_210.n8 82.852
R192 a_372_210.n11 a_372_210.n0 49.6
R193 a_372_210.n7 a_372_210.n6 32.833
R194 a_372_210.n8 a_372_210.t1 32.416
R195 a_372_210.n10 a_372_210.n9 27.2
R196 a_372_210.n3 a_372_210.n2 23.284
R197 a_372_210.n11 a_372_210.n10 22.4
R198 a_372_210.n7 a_372_210.n4 19.017
R199 a_372_210.n6 a_372_210.n5 13.494
R200 a_372_210.t1 a_372_210.n1 7.04
R201 a_372_210.t1 a_372_210.n3 5.727
R202 a_372_210.n8 a_372_210.n7 1.435
R203 B.n0 B.t0 479.223
R204 B.n0 B.t2 375.52
R205 B.n1 B.t1 241.707
R206 B.n1 B.n0 95.77
R207 B B.n1 76
R208 a_91_103.t0 a_91_103.n0 117.777
R209 a_91_103.n2 a_91_103.n1 55.228
R210 a_91_103.n4 a_91_103.n3 9.111
R211 a_91_103.t0 a_91_103.n2 4.04
R212 a_91_103.n8 a_91_103.n7 2.455
R213 a_91_103.n6 a_91_103.n4 1.964
R214 a_91_103.n6 a_91_103.n5 1.964
R215 a_91_103.n8 a_91_103.n6 0.636
R216 a_91_103.t0 a_91_103.n8 0.246
R217 GND.n30 GND.n29 219.745
R218 GND.n49 GND.n48 85.559
R219 GND.n30 GND.n28 85.529
R220 GND.n9 GND.n1 76.145
R221 GND.n43 GND.n42 76
R222 GND.n9 GND.n8 76
R223 GND.n17 GND.n16 76
R224 GND.n24 GND.n23 76
R225 GND.n27 GND.n26 76
R226 GND.n34 GND.n33 76
R227 GND.n37 GND.n36 76
R228 GND.n40 GND.n39 76
R229 GND.n69 GND.n68 76
R230 GND.n66 GND.n65 76
R231 GND.n63 GND.n62 76
R232 GND.n60 GND.n59 76
R233 GND.n57 GND.n56 76
R234 GND.n54 GND.n53 76
R235 GND.n51 GND.n50 76
R236 GND.n46 GND.n45 76
R237 GND.n5 GND.n4 35.01
R238 GND.n3 GND.n2 29.127
R239 GND.n12 GND.t1 20.794
R240 GND.n6 GND.n5 19.735
R241 GND.n14 GND.n13 19.735
R242 GND.n22 GND.n21 19.735
R243 GND.n5 GND.n3 19.017
R244 GND.n33 GND.n31 14.167
R245 GND.n45 GND.n44 13.653
R246 GND.n50 GND.n47 13.653
R247 GND.n53 GND.n52 13.653
R248 GND.n56 GND.n55 13.653
R249 GND.n59 GND.n58 13.653
R250 GND.n62 GND.n61 13.653
R251 GND.n65 GND.n64 13.653
R252 GND.n68 GND.n67 13.653
R253 GND.n39 GND.n38 13.653
R254 GND.n36 GND.n35 13.653
R255 GND.n33 GND.n32 13.653
R256 GND.n26 GND.n25 13.653
R257 GND.n23 GND.n18 13.653
R258 GND.n16 GND.n15 13.653
R259 GND.n8 GND.n7 13.653
R260 GND.n21 GND.n20 12.837
R261 GND.n20 GND.n19 7.566
R262 GND.n31 GND.n30 7.312
R263 GND.n11 GND.n10 4.551
R264 GND.n8 GND.n6 3.935
R265 GND.n23 GND.n22 3.541
R266 GND.t1 GND.n11 2.238
R267 GND.n1 GND.n0 0.596
R268 GND.n42 GND.n41 0.596
R269 GND.n13 GND.n12 0.358
R270 GND.n34 GND.n27 0.29
R271 GND.n43 GND 0.207
R272 GND.n63 GND.n60 0.197
R273 GND.n16 GND.n14 0.196
R274 GND.n50 GND.n49 0.196
R275 GND.n17 GND.n9 0.157
R276 GND.n24 GND.n17 0.157
R277 GND.n27 GND.n24 0.145
R278 GND.n37 GND.n34 0.145
R279 GND.n40 GND.n37 0.145
R280 GND.n69 GND.n66 0.145
R281 GND.n66 GND.n63 0.145
R282 GND.n60 GND.n57 0.145
R283 GND.n57 GND.n54 0.145
R284 GND.n54 GND.n51 0.145
R285 GND.n51 GND.n46 0.145
R286 GND.n46 GND.n43 0.145
R287 GND GND.n40 0.086
R288 GND GND.n69 0.058
C7 VDD GND 5.95fF
C8 a_91_103.n0 GND 0.03fF
C9 a_91_103.n1 GND 0.10fF
C10 a_91_103.n2 GND 0.10fF
C11 a_91_103.n3 GND 0.04fF
C12 a_91_103.n4 GND 0.03fF
C13 a_91_103.n5 GND 0.03fF
C14 a_91_103.n6 GND 0.03fF
C15 a_91_103.n7 GND 0.04fF
C16 a_372_210.n0 GND 0.02fF
C17 a_372_210.n1 GND 0.09fF
C18 a_372_210.n2 GND 0.13fF
C19 a_372_210.n3 GND 0.11fF
C20 a_372_210.t1 GND 0.30fF
C21 a_372_210.n4 GND 0.09fF
C22 a_372_210.n5 GND 0.06fF
C23 a_372_210.n6 GND 0.01fF
C24 a_372_210.n7 GND 0.03fF
C25 a_372_210.n8 GND 0.11fF
C26 a_372_210.n9 GND 0.02fF
C27 a_372_210.n10 GND 0.05fF
C28 a_372_210.n11 GND 0.02fF
C29 VDD.n0 GND 0.11fF
C30 VDD.n1 GND 0.02fF
C31 VDD.n2 GND 0.02fF
C32 VDD.n3 GND 0.04fF
C33 VDD.n4 GND 0.01fF
C34 VDD.n5 GND 0.02fF
C35 VDD.n6 GND 0.02fF
C36 VDD.n8 GND 0.02fF
C37 VDD.n9 GND 0.02fF
C38 VDD.n11 GND 0.02fF
C39 VDD.n14 GND 0.41fF
C40 VDD.n16 GND 0.03fF
C41 VDD.n17 GND 0.02fF
C42 VDD.n18 GND 0.02fF
C43 VDD.n19 GND 0.02fF
C44 VDD.n20 GND 0.03fF
C45 VDD.n21 GND 0.24fF
C46 VDD.n22 GND 0.02fF
C47 VDD.n23 GND 0.03fF
C48 VDD.n24 GND 0.05fF
C49 VDD.n25 GND 0.13fF
C50 VDD.n26 GND 0.18fF
C51 VDD.n27 GND 0.01fF
C52 VDD.n28 GND 0.01fF
C53 VDD.n29 GND 0.06fF
C54 VDD.n30 GND 0.15fF
C55 VDD.n31 GND 0.01fF
C56 VDD.n32 GND 0.02fF
C57 VDD.n33 GND 0.02fF
C58 VDD.n34 GND 0.13fF
C59 VDD.n35 GND 0.18fF
C60 VDD.n36 GND 0.01fF
C61 VDD.n37 GND 0.05fF
C62 VDD.n38 GND 0.01fF
C63 VDD.n39 GND 0.02fF
C64 VDD.n40 GND 0.24fF
C65 VDD.n41 GND 0.01fF
C66 VDD.n42 GND 0.02fF
C67 VDD.n43 GND 0.03fF
C68 VDD.n44 GND 0.02fF
C69 VDD.n45 GND 0.02fF
C70 VDD.n46 GND 0.02fF
C71 VDD.n47 GND 0.02fF
C72 VDD.n48 GND 0.02fF
C73 VDD.n49 GND 0.02fF
C74 VDD.n51 GND 0.02fF
C75 VDD.n52 GND 0.02fF
C76 VDD.n53 GND 0.02fF
C77 VDD.n54 GND 0.02fF
C78 VDD.n56 GND 0.03fF
C79 VDD.n57 GND 0.02fF
C80 VDD.n58 GND 0.21fF
C81 VDD.n59 GND 0.03fF
C82 VDD.n61 GND 0.24fF
C83 VDD.n63 GND 0.02fF
C84 VDD.n64 GND 0.02fF
C85 VDD.n65 GND 0.03fF
C86 VDD.n66 GND 0.02fF
C87 VDD.n67 GND 0.24fF
C88 VDD.n68 GND 0.01fF
C89 VDD.n69 GND 0.02fF
C90 VDD.n70 GND 0.03fF
C91 VDD.n71 GND 0.24fF
C92 VDD.n72 GND 0.01fF
C93 VDD.n73 GND 0.02fF
C94 VDD.n74 GND 0.02fF
C95 VDD.n75 GND 0.20fF
C96 VDD.n76 GND 0.01fF
C97 VDD.n77 GND 0.06fF
C98 VDD.n78 GND 0.02fF
C99 VDD.n79 GND 0.02fF
C100 VDD.n80 GND 0.02fF
C101 VDD.n81 GND 0.02fF
C102 VDD.n82 GND 0.18fF
C103 VDD.n83 GND 0.03fF
C104 VDD.n84 GND 0.02fF
C105 VDD.n85 GND 0.02fF
C106 VDD.n86 GND 0.02fF
C107 VDD.n87 GND 0.02fF
C108 VDD.n88 GND 0.02fF
C109 VDD.n90 GND 0.02fF
C110 VDD.n91 GND 0.02fF
C111 VDD.n92 GND 0.02fF
C112 VDD.n94 GND 0.41fF
C113 VDD.n96 GND 0.03fF
C114 VDD.n97 GND 0.03fF
C115 VDD.n98 GND 0.24fF
C116 VDD.n99 GND 0.02fF
C117 VDD.n100 GND 0.03fF
C118 VDD.n101 GND 0.02fF
C119 VDD.n102 GND 0.24fF
C120 VDD.n103 GND 0.01fF
C121 VDD.n104 GND 0.02fF
C122 VDD.n105 GND 0.02fF
C123 VDD.n106 GND 0.05fF
C124 VDD.n107 GND 0.20fF
C125 VDD.n108 GND 0.01fF
C126 VDD.n109 GND 0.01fF
C127 VDD.n110 GND 0.02fF
C128 VDD.n111 GND 0.12fF
C129 VDD.n112 GND 0.15fF
C130 VDD.n113 GND 0.01fF
C131 VDD.n114 GND 0.02fF
C132 VDD.n115 GND 0.02fF
C133 VDD.n116 GND 0.09fF
C134 VDD.n117 GND 0.02fF
C135 VDD.n118 GND 0.12fF
C136 VDD.n119 GND 0.14fF
C137 VDD.n120 GND 0.01fF
C138 VDD.n121 GND 0.01fF
C139 VDD.n122 GND 0.02fF
C140 VDD.n123 GND 0.16fF
C141 VDD.n124 GND 0.13fF
C142 VDD.n125 GND 0.01fF
C143 VDD.n126 GND 0.02fF
C144 VDD.n127 GND 0.02fF
C145 VDD.n128 GND 0.16fF
C146 VDD.n129 GND 0.13fF
C147 VDD.n130 GND 0.01fF
C148 VDD.n131 GND 0.02fF
C149 VDD.n132 GND 0.02fF
C150 VDD.n133 GND 0.12fF
C151 VDD.n134 GND 0.14fF
C152 VDD.n135 GND 0.01fF
C153 VDD.n136 GND 0.09fF
C154 VDD.n137 GND 0.02fF
C155 VDD.n138 GND 0.01fF
C156 VDD.n139 GND 0.02fF
C157 VDD.n140 GND 0.12fF
C158 VDD.n141 GND 0.15fF
C159 VDD.n142 GND 0.01fF
C160 VDD.n143 GND 0.02fF
C161 VDD.n144 GND 0.01fF
C162 Y.n0 GND 0.80fF
C163 Y.n1 GND 0.04fF
C164 Y.n2 GND 0.06fF
C165 Y.n3 GND 0.04fF
C166 Y.n4 GND 0.27fF
C167 Y.n5 GND 0.47fF
C168 a_277_1050.n0 GND 0.39fF
C169 a_277_1050.n1 GND 0.39fF
C170 a_277_1050.n2 GND 0.46fF
C171 a_277_1050.n3 GND 0.14fF
C172 a_277_1050.n4 GND 0.25fF
C173 a_277_1050.n5 GND 0.27fF
C174 a_277_1050.n6 GND 0.42fF
C175 a_277_1050.n7 GND 0.44fF
C176 a_277_1050.n8 GND 0.06fF
C177 a_277_1050.n9 GND 0.19fF
C178 a_277_1050.n10 GND 0.03fF
.ends
