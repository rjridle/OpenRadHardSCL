magic
tech sky130A
magscale 1 2
timestamp 1642373950
<< error_p >>
rect 261 322 262 323
rect 262 321 263 322
rect 277 291 278 292
rect 312 291 313 292
rect 277 188 278 189
rect 312 188 313 189
<< nwell >>
rect -36 591 619 1353
<< nmos >>
rect 232 322 262 375
rect 232 292 328 322
tri 328 292 358 322 sw
rect 232 188 262 292
tri 262 276 278 292 nw
tri 312 276 328 292 ne
tri 262 188 278 204 sw
tri 312 188 328 204 se
rect 328 188 358 292
tri 232 158 262 188 ne
rect 262 158 328 188
tri 328 158 358 188 nw
<< pmos >>
rect 56 629 86 1229
rect 144 629 174 1229
rect 232 629 262 1229
rect 320 629 350 1229
rect 408 629 438 1229
rect 497 629 527 1229
<< ndiff >>
rect 176 298 232 375
rect 262 322 412 375
rect 176 264 186 298
rect 220 264 232 298
tri 328 292 358 322 ne
rect 358 298 412 322
rect 176 215 232 264
rect 176 181 186 215
rect 220 181 232 215
tri 262 276 278 292 se
rect 278 276 312 292
tri 312 276 328 292 sw
rect 262 244 328 276
rect 262 210 274 244
rect 308 210 328 244
rect 262 204 328 210
tri 262 188 278 204 ne
rect 278 188 312 204
tri 312 188 328 204 nw
rect 358 264 370 298
rect 404 264 412 298
rect 358 215 412 264
rect 176 158 232 181
tri 232 158 262 188 sw
tri 328 158 358 188 se
rect 358 181 370 215
rect 404 181 412 215
rect 358 158 412 181
rect 176 147 412 158
rect 176 113 186 147
rect 220 113 274 147
rect 308 113 370 147
rect 404 113 412 147
rect 176 101 412 113
<< pdiff >>
rect 2 1213 56 1229
rect 2 1179 10 1213
rect 44 1179 56 1213
rect 2 1145 56 1179
rect 2 1111 10 1145
rect 44 1111 56 1145
rect 2 1077 56 1111
rect 2 1043 10 1077
rect 44 1043 56 1077
rect 2 1009 56 1043
rect 2 975 10 1009
rect 44 975 56 1009
rect 2 941 56 975
rect 2 907 10 941
rect 44 907 56 941
rect 2 873 56 907
rect 2 839 10 873
rect 44 839 56 873
rect 2 805 56 839
rect 2 771 10 805
rect 44 771 56 805
rect 2 737 56 771
rect 2 703 10 737
rect 44 703 56 737
rect 2 629 56 703
rect 86 1213 144 1229
rect 86 1179 98 1213
rect 132 1179 144 1213
rect 86 1145 144 1179
rect 86 1111 98 1145
rect 132 1111 144 1145
rect 86 1077 144 1111
rect 86 1043 98 1077
rect 132 1043 144 1077
rect 86 1009 144 1043
rect 86 975 98 1009
rect 132 975 144 1009
rect 86 941 144 975
rect 86 907 98 941
rect 132 907 144 941
rect 86 873 144 907
rect 86 839 98 873
rect 132 839 144 873
rect 86 805 144 839
rect 86 771 98 805
rect 132 771 144 805
rect 86 737 144 771
rect 86 703 98 737
rect 132 703 144 737
rect 86 629 144 703
rect 174 1213 232 1229
rect 174 1179 186 1213
rect 220 1179 232 1213
rect 174 1145 232 1179
rect 174 1111 186 1145
rect 220 1111 232 1145
rect 174 1077 232 1111
rect 174 1043 186 1077
rect 220 1043 232 1077
rect 174 1009 232 1043
rect 174 975 186 1009
rect 220 975 232 1009
rect 174 941 232 975
rect 174 907 186 941
rect 220 907 232 941
rect 174 873 232 907
rect 174 839 186 873
rect 220 839 232 873
rect 174 805 232 839
rect 174 771 186 805
rect 220 771 232 805
rect 174 737 232 771
rect 174 703 186 737
rect 220 703 232 737
rect 174 629 232 703
rect 262 1213 320 1229
rect 262 1179 274 1213
rect 308 1179 320 1213
rect 262 1145 320 1179
rect 262 1111 274 1145
rect 308 1111 320 1145
rect 262 1077 320 1111
rect 262 1043 274 1077
rect 308 1043 320 1077
rect 262 1009 320 1043
rect 262 975 274 1009
rect 308 975 320 1009
rect 262 941 320 975
rect 262 907 274 941
rect 308 907 320 941
rect 262 873 320 907
rect 262 839 274 873
rect 308 839 320 873
rect 262 805 320 839
rect 262 771 274 805
rect 308 771 320 805
rect 262 737 320 771
rect 262 703 274 737
rect 308 703 320 737
rect 262 629 320 703
rect 350 1213 408 1229
rect 350 1179 362 1213
rect 396 1179 408 1213
rect 350 1145 408 1179
rect 350 1111 362 1145
rect 396 1111 408 1145
rect 350 1077 408 1111
rect 350 1043 362 1077
rect 396 1043 408 1077
rect 350 1009 408 1043
rect 350 975 362 1009
rect 396 975 408 1009
rect 350 941 408 975
rect 350 907 362 941
rect 396 907 408 941
rect 350 873 408 907
rect 350 839 362 873
rect 396 839 408 873
rect 350 805 408 839
rect 350 771 362 805
rect 396 771 408 805
rect 350 737 408 771
rect 350 703 362 737
rect 396 703 408 737
rect 350 629 408 703
rect 438 1213 497 1229
rect 438 1179 450 1213
rect 484 1179 497 1213
rect 438 1145 497 1179
rect 438 1111 450 1145
rect 484 1111 497 1145
rect 438 1077 497 1111
rect 438 1043 450 1077
rect 484 1043 497 1077
rect 438 1009 497 1043
rect 438 975 450 1009
rect 484 975 497 1009
rect 438 941 497 975
rect 438 907 450 941
rect 484 907 497 941
rect 438 873 497 907
rect 438 839 450 873
rect 484 839 497 873
rect 438 805 497 839
rect 438 771 450 805
rect 484 771 497 805
rect 438 737 497 771
rect 438 703 450 737
rect 484 703 497 737
rect 438 629 497 703
rect 527 1213 581 1229
rect 527 1179 539 1213
rect 573 1179 581 1213
rect 527 1145 581 1179
rect 527 1111 539 1145
rect 573 1111 581 1145
rect 527 1077 581 1111
rect 527 1043 539 1077
rect 573 1043 581 1077
rect 527 1009 581 1043
rect 527 975 539 1009
rect 573 975 581 1009
rect 527 941 581 975
rect 527 907 539 941
rect 573 907 581 941
rect 527 873 581 907
rect 527 839 539 873
rect 573 839 581 873
rect 527 805 581 839
rect 527 771 539 805
rect 573 771 581 805
rect 527 737 581 771
rect 527 703 539 737
rect 573 703 581 737
rect 527 629 581 703
<< ndiffc >>
rect 186 264 220 298
rect 186 181 220 215
rect 274 210 308 244
rect 370 264 404 298
rect 370 181 404 215
rect 186 113 220 147
rect 274 113 308 147
rect 370 113 404 147
<< pdiffc >>
rect 10 1179 44 1213
rect 10 1111 44 1145
rect 10 1043 44 1077
rect 10 975 44 1009
rect 10 907 44 941
rect 10 839 44 873
rect 10 771 44 805
rect 10 703 44 737
rect 98 1179 132 1213
rect 98 1111 132 1145
rect 98 1043 132 1077
rect 98 975 132 1009
rect 98 907 132 941
rect 98 839 132 873
rect 98 771 132 805
rect 98 703 132 737
rect 186 1179 220 1213
rect 186 1111 220 1145
rect 186 1043 220 1077
rect 186 975 220 1009
rect 186 907 220 941
rect 186 839 220 873
rect 186 771 220 805
rect 186 703 220 737
rect 274 1179 308 1213
rect 274 1111 308 1145
rect 274 1043 308 1077
rect 274 975 308 1009
rect 274 907 308 941
rect 274 839 308 873
rect 274 771 308 805
rect 274 703 308 737
rect 362 1179 396 1213
rect 362 1111 396 1145
rect 362 1043 396 1077
rect 362 975 396 1009
rect 362 907 396 941
rect 362 839 396 873
rect 362 771 396 805
rect 362 703 396 737
rect 450 1179 484 1213
rect 450 1111 484 1145
rect 450 1043 484 1077
rect 450 975 484 1009
rect 450 907 484 941
rect 450 839 484 873
rect 450 771 484 805
rect 450 703 484 737
rect 539 1179 573 1213
rect 539 1111 573 1145
rect 539 1043 573 1077
rect 539 975 573 1009
rect 539 907 573 941
rect 539 839 573 873
rect 539 771 573 805
rect 539 703 573 737
<< psubdiff >>
rect 0 13 24 47
rect 58 13 93 47
rect 127 13 169 47
rect 203 13 237 47
rect 271 13 305 47
rect 339 13 374 47
rect 408 13 450 47
rect 484 13 518 47
rect 552 13 600 47
<< nsubdiff >>
rect 0 1283 24 1317
rect 58 1283 92 1317
rect 126 1283 160 1317
rect 195 1283 229 1317
rect 263 1283 297 1317
rect 331 1283 365 1317
rect 399 1283 433 1317
rect 468 1283 502 1317
rect 536 1283 580 1317
<< psubdiffcont >>
rect 24 13 58 47
rect 93 13 127 47
rect 169 13 203 47
rect 237 13 271 47
rect 305 13 339 47
rect 374 13 408 47
rect 450 13 484 47
rect 518 13 552 47
<< nsubdiffcont >>
rect 24 1283 58 1317
rect 92 1283 126 1317
rect 160 1283 195 1317
rect 229 1283 263 1317
rect 297 1283 331 1317
rect 365 1283 399 1317
rect 433 1283 468 1317
rect 502 1283 536 1317
<< poly >>
rect 56 1229 86 1255
rect 144 1229 174 1255
rect 232 1229 262 1255
rect 320 1229 350 1255
rect 408 1229 438 1255
rect 497 1229 527 1255
rect 56 612 86 629
rect 144 612 174 629
rect 232 612 262 629
rect 320 612 350 629
rect 408 612 438 629
rect 497 612 527 629
rect 56 582 527 612
rect 232 494 262 582
rect 196 478 262 494
rect 196 444 206 478
rect 240 444 262 478
rect 196 428 262 444
rect 232 375 262 428
<< polycont >>
rect 206 444 240 478
<< locali >>
rect 0 1317 580 1332
rect 0 1283 24 1317
rect 58 1283 92 1317
rect 126 1283 160 1317
rect 195 1283 229 1317
rect 263 1283 297 1317
rect 331 1283 365 1317
rect 399 1283 433 1317
rect 468 1283 502 1317
rect 536 1283 580 1317
rect 0 1270 580 1283
rect 10 1213 44 1270
rect 10 1145 44 1179
rect 10 1077 44 1111
rect 10 1009 44 1043
rect 10 941 44 975
rect 10 873 44 907
rect 10 805 44 839
rect 10 737 44 771
rect 10 627 44 703
rect 98 1213 132 1229
rect 98 1145 132 1179
rect 98 1077 132 1111
rect 98 1009 132 1043
rect 98 941 132 975
rect 98 873 132 907
rect 98 805 132 839
rect 98 737 132 771
rect 98 672 132 703
rect 186 1213 220 1270
rect 186 1145 220 1179
rect 186 1077 220 1111
rect 186 1009 220 1043
rect 186 941 220 975
rect 186 873 220 907
rect 186 805 220 839
rect 186 737 220 771
rect 186 627 220 703
rect 274 1213 308 1229
rect 274 1145 308 1179
rect 274 1077 308 1111
rect 274 1009 308 1043
rect 274 941 308 975
rect 274 873 308 907
rect 274 805 308 839
rect 274 737 308 771
rect 274 673 308 703
rect 206 478 240 494
rect 206 428 240 444
rect 186 298 220 343
rect 186 215 220 264
rect 274 244 308 638
rect 362 1213 396 1270
rect 362 1145 396 1179
rect 362 1077 396 1111
rect 362 1009 396 1043
rect 362 941 396 975
rect 362 873 396 907
rect 362 805 396 839
rect 362 737 396 771
rect 362 627 396 703
rect 450 1213 484 1229
rect 450 1145 484 1179
rect 450 1077 484 1111
rect 450 1009 484 1043
rect 450 941 484 975
rect 450 873 484 907
rect 450 805 484 839
rect 450 737 484 771
rect 450 673 484 703
rect 539 1213 573 1270
rect 539 1145 573 1179
rect 539 1077 573 1111
rect 539 1009 573 1043
rect 539 941 573 975
rect 539 873 573 907
rect 539 805 573 839
rect 539 737 573 771
rect 539 629 573 703
rect 274 194 308 210
rect 370 298 404 343
rect 370 215 404 264
rect 186 147 220 181
rect 370 147 404 181
rect 220 113 274 147
rect 308 113 370 147
rect 186 62 220 113
rect 370 62 404 113
rect 0 47 600 62
rect 0 13 24 47
rect 58 13 93 47
rect 127 13 169 47
rect 203 13 237 47
rect 271 13 305 47
rect 339 13 374 47
rect 408 13 450 47
rect 484 13 518 47
rect 552 13 600 47
rect 0 0 600 13
<< viali >>
rect 24 1283 58 1317
rect 92 1283 126 1317
rect 160 1283 195 1317
rect 229 1283 263 1317
rect 297 1283 331 1317
rect 365 1283 399 1317
rect 433 1283 468 1317
rect 502 1283 536 1317
rect 98 638 132 672
rect 274 638 308 673
rect 206 444 240 478
rect 450 639 484 673
rect 24 13 58 47
rect 93 13 127 47
rect 169 13 203 47
rect 237 13 271 47
rect 305 13 339 47
rect 374 13 408 47
rect 450 13 484 47
rect 518 13 552 47
<< metal1 >>
rect 0 1317 580 1332
rect 0 1283 24 1317
rect 58 1283 92 1317
rect 126 1283 160 1317
rect 195 1283 229 1317
rect 263 1283 297 1317
rect 331 1283 365 1317
rect 399 1283 433 1317
rect 468 1283 502 1317
rect 536 1283 580 1317
rect 0 1270 580 1283
rect 86 672 143 678
rect 262 673 320 679
rect 262 672 274 673
rect 86 638 98 672
rect 132 638 274 672
rect 308 672 320 673
rect 438 673 497 679
rect 438 672 450 673
rect 308 639 450 672
rect 484 639 497 673
rect 308 638 497 639
rect 86 632 143 638
rect 262 632 320 638
rect 438 632 497 638
rect 274 629 308 632
rect 206 485 240 502
rect 200 478 246 485
rect 200 444 206 478
rect 240 444 246 478
rect 200 437 246 444
rect 206 421 240 437
rect 0 47 600 62
rect 0 13 24 47
rect 58 13 93 47
rect 127 13 169 47
rect 203 13 237 47
rect 271 13 305 47
rect 339 13 374 47
rect 408 13 450 47
rect 484 13 518 47
rect 552 13 600 47
rect 0 0 600 13
<< labels >>
rlabel metal1 206 444 240 478 1 A
rlabel metal1 281 1301 281 1301 1 VDD
rlabel metal1 287 26 287 26 1 VSS
rlabel metal1 274 638 308 673 1 Y
<< end >>
