magic
tech sky130A
magscale 1 2
timestamp 1646004885
<< locali >>
rect -17 17 17 33
rect -17 -33 17 -17
<< viali >>
rect -17 -17 17 17
<< metal1 >>
rect -23 17 23 23
rect -53 -17 -17 17
rect 17 -17 29 17
rect -23 -23 23 -17
<< end >>
