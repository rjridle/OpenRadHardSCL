magic
tech sky130A
magscale 1 2
timestamp 1645648650
<< nmos >>
tri 145 222 161 238 se
rect 161 222 191 276
tri 55 192 85 222 se
rect 85 192 191 222
rect 55 92 85 192
tri 85 176 101 192 nw
tri 145 176 161 192 ne
tri 85 92 101 108 sw
tri 145 92 161 108 se
rect 161 92 191 192
tri 55 62 85 92 ne
rect 85 62 161 92
tri 161 62 191 92 nw
<< ndiff >>
rect -1 260 161 276
rect -1 226 9 260
rect 43 238 161 260
rect 43 226 145 238
rect -1 222 145 226
tri 145 222 161 238 nw
rect 191 260 247 276
rect 191 226 203 260
rect 237 226 247 260
rect -1 189 55 222
tri 55 192 85 222 nw
rect -1 155 9 189
rect 43 155 55 189
rect -1 121 55 155
rect -1 87 9 121
rect 43 87 55 121
tri 85 176 101 192 se
rect 101 176 145 192
tri 145 176 161 192 sw
rect 85 144 161 176
rect 85 110 106 144
rect 140 110 161 144
rect 85 108 161 110
tri 85 92 101 108 ne
rect 101 92 145 108
tri 145 92 161 108 nw
rect 191 189 247 226
rect 191 155 203 189
rect 237 155 247 189
rect 191 121 247 155
rect -1 62 55 87
tri 55 62 85 92 sw
tri 161 62 191 92 se
rect 191 87 203 121
rect 237 87 247 121
rect 191 62 247 87
rect -1 50 247 62
rect -1 16 9 50
rect 43 16 106 50
rect 140 16 203 50
rect 237 16 247 50
rect -1 0 247 16
<< ndiffc >>
rect 9 226 43 260
rect 203 226 237 260
rect 9 155 43 189
rect 9 87 43 121
rect 106 110 140 144
rect 203 155 237 189
rect 203 87 237 121
rect 9 16 43 50
rect 106 16 140 50
rect 203 16 237 50
<< poly >>
rect 161 276 191 309
<< locali >>
rect 9 260 43 276
rect 9 189 43 226
rect 203 260 237 276
rect 203 189 237 226
rect 9 121 43 155
rect 106 144 140 160
rect 106 94 140 110
rect 203 121 237 155
rect 9 50 43 87
rect 203 50 237 87
rect 43 16 106 50
rect 140 16 203 50
rect 9 0 43 16
rect 203 0 237 16
<< end >>
