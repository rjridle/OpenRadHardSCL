magic
tech sky130A
magscale 1 2
timestamp 1649546437
<< nwell >>
rect -84 832 5264 1575
<< nmos >>
rect 147 318 177 379
tri 177 318 193 334 sw
rect 447 318 477 379
rect 147 288 253 318
tri 253 288 283 318 sw
rect 147 187 177 288
tri 177 272 193 288 nw
tri 237 272 253 288 ne
tri 177 187 193 203 sw
tri 237 187 253 203 se
rect 253 187 283 288
tri 342 288 372 318 se
rect 372 288 477 318
rect 342 194 372 288
tri 372 272 388 288 nw
tri 431 272 447 288 ne
tri 372 194 388 210 sw
tri 431 194 447 210 se
rect 447 194 477 288
tri 147 157 177 187 ne
rect 177 157 253 187
tri 253 157 283 187 nw
tri 342 164 372 194 ne
rect 372 164 447 194
tri 447 164 477 194 nw
rect 649 326 679 379
tri 679 326 695 342 sw
rect 649 296 755 326
tri 755 296 785 326 sw
rect 649 195 679 296
tri 679 280 695 296 nw
tri 739 280 755 296 ne
tri 679 195 695 211 sw
tri 739 195 755 211 se
rect 755 195 785 296
tri 649 165 679 195 ne
rect 679 165 755 195
tri 755 165 785 195 nw
rect 1109 318 1139 379
tri 1139 318 1155 334 sw
rect 1409 318 1439 379
rect 1109 288 1215 318
tri 1215 288 1245 318 sw
rect 1109 187 1139 288
tri 1139 272 1155 288 nw
tri 1199 272 1215 288 ne
tri 1139 187 1155 203 sw
tri 1199 187 1215 203 se
rect 1215 187 1245 288
tri 1304 288 1334 318 se
rect 1334 288 1439 318
rect 1304 194 1334 288
tri 1334 272 1350 288 nw
tri 1393 272 1409 288 ne
tri 1334 194 1350 210 sw
tri 1393 194 1409 210 se
rect 1409 194 1439 288
tri 1109 157 1139 187 ne
rect 1139 157 1215 187
tri 1215 157 1245 187 nw
tri 1304 164 1334 194 ne
rect 1334 164 1409 194
tri 1409 164 1439 194 nw
rect 1611 326 1641 379
tri 1641 326 1657 342 sw
rect 1611 296 1717 326
tri 1717 296 1747 326 sw
rect 1611 195 1641 296
tri 1641 280 1657 296 nw
tri 1701 280 1717 296 ne
tri 1641 195 1657 211 sw
tri 1701 195 1717 211 se
rect 1717 195 1747 296
tri 1611 165 1641 195 ne
rect 1641 165 1717 195
tri 1717 165 1747 195 nw
rect 2092 316 2122 377
tri 2122 316 2138 332 sw
rect 2286 324 2316 377
tri 2316 324 2332 340 sw
rect 2092 286 2198 316
tri 2198 286 2228 316 sw
rect 2286 294 2392 324
tri 2392 294 2422 324 sw
rect 2092 185 2122 286
tri 2122 270 2138 286 nw
tri 2182 270 2198 286 ne
tri 2122 185 2138 201 sw
tri 2182 185 2198 201 se
rect 2198 185 2228 286
rect 2286 193 2316 294
tri 2316 278 2332 294 nw
tri 2376 278 2392 294 ne
tri 2316 193 2332 209 sw
tri 2376 193 2392 209 se
rect 2392 193 2422 294
tri 2092 155 2122 185 ne
rect 2122 155 2198 185
tri 2198 155 2228 185 nw
tri 2286 163 2316 193 ne
rect 2316 163 2392 193
tri 2392 163 2422 193 nw
rect 2737 318 2767 379
tri 2767 318 2783 334 sw
rect 3037 318 3067 379
rect 2737 288 2843 318
tri 2843 288 2873 318 sw
rect 2737 187 2767 288
tri 2767 272 2783 288 nw
tri 2827 272 2843 288 ne
tri 2767 187 2783 203 sw
tri 2827 187 2843 203 se
rect 2843 187 2873 288
tri 2932 288 2962 318 se
rect 2962 288 3067 318
rect 2932 194 2962 288
tri 2962 272 2978 288 nw
tri 3021 272 3037 288 ne
tri 2962 194 2978 210 sw
tri 3021 194 3037 210 se
rect 3037 194 3067 288
tri 2737 157 2767 187 ne
rect 2767 157 2843 187
tri 2843 157 2873 187 nw
tri 2932 164 2962 194 ne
rect 2962 164 3037 194
tri 3037 164 3067 194 nw
rect 3239 326 3269 379
tri 3269 326 3285 342 sw
rect 3239 296 3345 326
tri 3345 296 3375 326 sw
rect 3239 195 3269 296
tri 3269 280 3285 296 nw
tri 3329 280 3345 296 ne
tri 3269 195 3285 211 sw
tri 3329 195 3345 211 se
rect 3345 195 3375 296
tri 3239 165 3269 195 ne
rect 3269 165 3345 195
tri 3345 165 3375 195 nw
rect 3699 318 3729 379
tri 3729 318 3745 334 sw
rect 3999 318 4029 379
rect 3699 288 3805 318
tri 3805 288 3835 318 sw
rect 3699 187 3729 288
tri 3729 272 3745 288 nw
tri 3789 272 3805 288 ne
tri 3729 187 3745 203 sw
tri 3789 187 3805 203 se
rect 3805 187 3835 288
tri 3894 288 3924 318 se
rect 3924 288 4029 318
rect 3894 194 3924 288
tri 3924 272 3940 288 nw
tri 3983 272 3999 288 ne
tri 3924 194 3940 210 sw
tri 3983 194 3999 210 se
rect 3999 194 4029 288
tri 3699 157 3729 187 ne
rect 3729 157 3805 187
tri 3805 157 3835 187 nw
tri 3894 164 3924 194 ne
rect 3924 164 3999 194
tri 3999 164 4029 194 nw
rect 4201 326 4231 379
tri 4231 326 4247 342 sw
rect 4201 296 4307 326
tri 4307 296 4337 326 sw
rect 4201 195 4231 296
tri 4231 280 4247 296 nw
tri 4291 280 4307 296 ne
tri 4231 195 4247 211 sw
tri 4291 195 4307 211 se
rect 4307 195 4337 296
tri 4201 165 4231 195 ne
rect 4231 165 4307 195
tri 4307 165 4337 195 nw
rect 4682 316 4712 377
tri 4712 316 4728 332 sw
rect 4876 324 4906 377
tri 4906 324 4922 340 sw
rect 4682 286 4788 316
tri 4788 286 4818 316 sw
rect 4876 294 4982 324
tri 4982 294 5012 324 sw
rect 4682 185 4712 286
tri 4712 270 4728 286 nw
tri 4772 270 4788 286 ne
tri 4712 185 4728 201 sw
tri 4772 185 4788 201 se
rect 4788 185 4818 286
rect 4876 193 4906 294
tri 4906 278 4922 294 nw
tri 4966 278 4982 294 ne
tri 4906 193 4922 209 sw
tri 4966 193 4982 209 se
rect 4982 193 5012 294
tri 4682 155 4712 185 ne
rect 4712 155 4788 185
tri 4788 155 4818 185 nw
tri 4876 163 4906 193 ne
rect 4906 163 4982 193
tri 4982 163 5012 193 nw
<< pmos >>
rect 247 1050 277 1450
rect 335 1050 365 1450
rect 423 1050 453 1450
rect 511 1050 541 1450
rect 599 1050 629 1450
rect 687 1050 717 1450
rect 1209 1050 1239 1450
rect 1297 1050 1327 1450
rect 1385 1050 1415 1450
rect 1473 1050 1503 1450
rect 1561 1050 1591 1450
rect 1649 1050 1679 1450
rect 2111 1050 2141 1450
rect 2199 1050 2229 1450
rect 2287 1050 2317 1450
rect 2375 1050 2405 1450
rect 2837 1050 2867 1450
rect 2925 1050 2955 1450
rect 3013 1050 3043 1450
rect 3101 1050 3131 1450
rect 3189 1050 3219 1450
rect 3277 1050 3307 1450
rect 3799 1050 3829 1450
rect 3887 1050 3917 1450
rect 3975 1050 4005 1450
rect 4063 1050 4093 1450
rect 4151 1050 4181 1450
rect 4239 1050 4269 1450
rect 4701 1050 4731 1450
rect 4789 1050 4819 1450
rect 4877 1050 4907 1450
rect 4965 1050 4995 1450
<< ndiff >>
rect 91 363 147 379
rect 91 329 101 363
rect 135 329 147 363
rect 91 291 147 329
rect 177 363 447 379
rect 177 334 198 363
tri 177 318 193 334 ne
rect 193 329 198 334
rect 232 329 295 363
rect 329 329 392 363
rect 426 329 447 363
rect 193 318 447 329
rect 477 363 533 379
rect 477 329 489 363
rect 523 329 533 363
rect 91 257 101 291
rect 135 257 147 291
tri 253 288 283 318 ne
rect 283 291 342 318
rect 91 223 147 257
rect 91 189 101 223
rect 135 189 147 223
rect 91 157 147 189
tri 177 272 193 288 se
rect 193 272 237 288
tri 237 272 253 288 sw
rect 177 238 253 272
rect 177 204 198 238
rect 232 204 253 238
rect 177 203 253 204
tri 177 187 193 203 ne
rect 193 187 237 203
tri 237 187 253 203 nw
rect 283 257 295 291
rect 329 257 342 291
tri 342 288 372 318 nw
rect 283 223 342 257
rect 283 189 295 223
rect 329 189 342 223
tri 372 272 388 288 se
rect 388 272 431 288
tri 431 272 447 288 sw
rect 372 244 447 272
rect 372 210 393 244
rect 427 210 447 244
tri 372 194 388 210 ne
rect 388 194 431 210
tri 431 194 447 210 nw
tri 147 157 177 187 sw
tri 253 157 283 187 se
rect 283 164 342 189
tri 342 164 372 194 sw
tri 447 164 477 194 se
rect 477 164 533 329
rect 283 157 533 164
rect 91 153 533 157
rect 91 119 101 153
rect 135 119 295 153
rect 329 119 392 153
rect 426 119 489 153
rect 523 119 533 153
rect 91 103 533 119
rect 593 363 649 379
rect 593 329 603 363
rect 637 329 649 363
rect 593 291 649 329
rect 679 342 841 379
tri 679 326 695 342 ne
rect 695 326 841 342
tri 755 296 785 326 ne
rect 593 257 603 291
rect 637 257 649 291
rect 593 223 649 257
rect 593 189 603 223
rect 637 189 649 223
tri 679 280 695 296 se
rect 695 280 739 296
tri 739 280 755 296 sw
rect 679 247 755 280
rect 679 213 700 247
rect 734 213 755 247
rect 679 211 755 213
tri 679 195 695 211 ne
rect 695 195 739 211
tri 739 195 755 211 nw
rect 785 291 841 326
rect 785 257 797 291
rect 831 257 841 291
rect 785 223 841 257
rect 593 165 649 189
tri 649 165 679 195 sw
tri 755 165 785 195 se
rect 785 189 797 223
rect 831 189 841 223
rect 785 165 841 189
rect 593 153 841 165
rect 593 119 603 153
rect 637 119 700 153
rect 734 119 797 153
rect 831 119 841 153
rect 593 103 841 119
rect 1053 363 1109 379
rect 1053 329 1063 363
rect 1097 329 1109 363
rect 1053 291 1109 329
rect 1139 363 1409 379
rect 1139 334 1160 363
tri 1139 318 1155 334 ne
rect 1155 329 1160 334
rect 1194 329 1257 363
rect 1291 329 1354 363
rect 1388 329 1409 363
rect 1155 318 1409 329
rect 1439 363 1495 379
rect 1439 329 1451 363
rect 1485 329 1495 363
rect 1053 257 1063 291
rect 1097 257 1109 291
tri 1215 288 1245 318 ne
rect 1245 291 1304 318
rect 1053 223 1109 257
rect 1053 189 1063 223
rect 1097 189 1109 223
rect 1053 157 1109 189
tri 1139 272 1155 288 se
rect 1155 272 1199 288
tri 1199 272 1215 288 sw
rect 1139 238 1215 272
rect 1139 204 1160 238
rect 1194 204 1215 238
rect 1139 203 1215 204
tri 1139 187 1155 203 ne
rect 1155 187 1199 203
tri 1199 187 1215 203 nw
rect 1245 257 1257 291
rect 1291 257 1304 291
tri 1304 288 1334 318 nw
rect 1245 223 1304 257
rect 1245 189 1257 223
rect 1291 189 1304 223
tri 1334 272 1350 288 se
rect 1350 272 1393 288
tri 1393 272 1409 288 sw
rect 1334 244 1409 272
rect 1334 210 1355 244
rect 1389 210 1409 244
tri 1334 194 1350 210 ne
rect 1350 194 1393 210
tri 1393 194 1409 210 nw
tri 1109 157 1139 187 sw
tri 1215 157 1245 187 se
rect 1245 164 1304 189
tri 1304 164 1334 194 sw
tri 1409 164 1439 194 se
rect 1439 164 1495 329
rect 1245 157 1495 164
rect 1053 153 1495 157
rect 1053 119 1063 153
rect 1097 119 1257 153
rect 1291 119 1354 153
rect 1388 119 1451 153
rect 1485 119 1495 153
rect 1053 103 1495 119
rect 1555 363 1611 379
rect 1555 329 1565 363
rect 1599 329 1611 363
rect 1555 291 1611 329
rect 1641 342 1803 379
tri 1641 326 1657 342 ne
rect 1657 326 1803 342
tri 1717 296 1747 326 ne
rect 1555 257 1565 291
rect 1599 257 1611 291
rect 1555 223 1611 257
rect 1555 189 1565 223
rect 1599 189 1611 223
tri 1641 280 1657 296 se
rect 1657 280 1701 296
tri 1701 280 1717 296 sw
rect 1641 247 1717 280
rect 1641 213 1662 247
rect 1696 213 1717 247
rect 1641 211 1717 213
tri 1641 195 1657 211 ne
rect 1657 195 1701 211
tri 1701 195 1717 211 nw
rect 1747 291 1803 326
rect 1747 257 1759 291
rect 1793 257 1803 291
rect 1747 223 1803 257
rect 1555 165 1611 189
tri 1611 165 1641 195 sw
tri 1717 165 1747 195 se
rect 1747 189 1759 223
rect 1793 189 1803 223
rect 1747 165 1803 189
rect 1555 153 1803 165
rect 1555 119 1565 153
rect 1599 119 1662 153
rect 1696 119 1759 153
rect 1793 119 1803 153
rect 1555 103 1803 119
rect 2036 361 2092 377
rect 2036 327 2046 361
rect 2080 327 2092 361
rect 2036 289 2092 327
rect 2122 361 2286 377
rect 2122 332 2143 361
tri 2122 316 2138 332 ne
rect 2138 327 2143 332
rect 2177 327 2240 361
rect 2274 327 2286 361
rect 2138 316 2286 327
rect 2316 340 2478 377
tri 2316 324 2332 340 ne
rect 2332 324 2478 340
rect 2036 255 2046 289
rect 2080 255 2092 289
tri 2198 286 2228 316 ne
rect 2228 289 2286 316
tri 2392 294 2422 324 ne
rect 2036 221 2092 255
rect 2036 187 2046 221
rect 2080 187 2092 221
rect 2036 155 2092 187
tri 2122 270 2138 286 se
rect 2138 270 2182 286
tri 2182 270 2198 286 sw
rect 2122 236 2198 270
rect 2122 202 2143 236
rect 2177 202 2198 236
rect 2122 201 2198 202
tri 2122 185 2138 201 ne
rect 2138 185 2182 201
tri 2182 185 2198 201 nw
rect 2228 255 2240 289
rect 2274 255 2286 289
rect 2228 221 2286 255
rect 2228 187 2240 221
rect 2274 187 2286 221
tri 2316 278 2332 294 se
rect 2332 278 2376 294
tri 2376 278 2392 294 sw
rect 2316 245 2392 278
rect 2316 211 2337 245
rect 2371 211 2392 245
rect 2316 209 2392 211
tri 2316 193 2332 209 ne
rect 2332 193 2376 209
tri 2376 193 2392 209 nw
rect 2422 289 2478 324
rect 2422 255 2434 289
rect 2468 255 2478 289
rect 2422 221 2478 255
tri 2092 155 2122 185 sw
tri 2198 155 2228 185 se
rect 2228 163 2286 187
tri 2286 163 2316 193 sw
tri 2392 163 2422 193 se
rect 2422 187 2434 221
rect 2468 187 2478 221
rect 2422 163 2478 187
rect 2228 155 2478 163
rect 2036 151 2478 155
rect 2036 117 2046 151
rect 2080 117 2240 151
rect 2274 117 2337 151
rect 2371 117 2434 151
rect 2468 117 2478 151
rect 2036 101 2478 117
rect 2681 363 2737 379
rect 2681 329 2691 363
rect 2725 329 2737 363
rect 2681 291 2737 329
rect 2767 363 3037 379
rect 2767 334 2788 363
tri 2767 318 2783 334 ne
rect 2783 329 2788 334
rect 2822 329 2885 363
rect 2919 329 2982 363
rect 3016 329 3037 363
rect 2783 318 3037 329
rect 3067 363 3123 379
rect 3067 329 3079 363
rect 3113 329 3123 363
rect 2681 257 2691 291
rect 2725 257 2737 291
tri 2843 288 2873 318 ne
rect 2873 291 2932 318
rect 2681 223 2737 257
rect 2681 189 2691 223
rect 2725 189 2737 223
rect 2681 157 2737 189
tri 2767 272 2783 288 se
rect 2783 272 2827 288
tri 2827 272 2843 288 sw
rect 2767 238 2843 272
rect 2767 204 2788 238
rect 2822 204 2843 238
rect 2767 203 2843 204
tri 2767 187 2783 203 ne
rect 2783 187 2827 203
tri 2827 187 2843 203 nw
rect 2873 257 2885 291
rect 2919 257 2932 291
tri 2932 288 2962 318 nw
rect 2873 223 2932 257
rect 2873 189 2885 223
rect 2919 189 2932 223
tri 2962 272 2978 288 se
rect 2978 272 3021 288
tri 3021 272 3037 288 sw
rect 2962 244 3037 272
rect 2962 210 2983 244
rect 3017 210 3037 244
tri 2962 194 2978 210 ne
rect 2978 194 3021 210
tri 3021 194 3037 210 nw
tri 2737 157 2767 187 sw
tri 2843 157 2873 187 se
rect 2873 164 2932 189
tri 2932 164 2962 194 sw
tri 3037 164 3067 194 se
rect 3067 164 3123 329
rect 2873 157 3123 164
rect 2681 153 3123 157
rect 2681 119 2691 153
rect 2725 119 2885 153
rect 2919 119 2982 153
rect 3016 119 3079 153
rect 3113 119 3123 153
rect 2681 103 3123 119
rect 3183 363 3239 379
rect 3183 329 3193 363
rect 3227 329 3239 363
rect 3183 291 3239 329
rect 3269 342 3431 379
tri 3269 326 3285 342 ne
rect 3285 326 3431 342
tri 3345 296 3375 326 ne
rect 3183 257 3193 291
rect 3227 257 3239 291
rect 3183 223 3239 257
rect 3183 189 3193 223
rect 3227 189 3239 223
tri 3269 280 3285 296 se
rect 3285 280 3329 296
tri 3329 280 3345 296 sw
rect 3269 247 3345 280
rect 3269 213 3290 247
rect 3324 213 3345 247
rect 3269 211 3345 213
tri 3269 195 3285 211 ne
rect 3285 195 3329 211
tri 3329 195 3345 211 nw
rect 3375 291 3431 326
rect 3375 257 3387 291
rect 3421 257 3431 291
rect 3375 223 3431 257
rect 3183 165 3239 189
tri 3239 165 3269 195 sw
tri 3345 165 3375 195 se
rect 3375 189 3387 223
rect 3421 189 3431 223
rect 3375 165 3431 189
rect 3183 153 3431 165
rect 3183 119 3193 153
rect 3227 119 3290 153
rect 3324 119 3387 153
rect 3421 119 3431 153
rect 3183 103 3431 119
rect 3643 363 3699 379
rect 3643 329 3653 363
rect 3687 329 3699 363
rect 3643 291 3699 329
rect 3729 363 3999 379
rect 3729 334 3750 363
tri 3729 318 3745 334 ne
rect 3745 329 3750 334
rect 3784 329 3847 363
rect 3881 329 3944 363
rect 3978 329 3999 363
rect 3745 318 3999 329
rect 4029 363 4085 379
rect 4029 329 4041 363
rect 4075 329 4085 363
rect 3643 257 3653 291
rect 3687 257 3699 291
tri 3805 288 3835 318 ne
rect 3835 291 3894 318
rect 3643 223 3699 257
rect 3643 189 3653 223
rect 3687 189 3699 223
rect 3643 157 3699 189
tri 3729 272 3745 288 se
rect 3745 272 3789 288
tri 3789 272 3805 288 sw
rect 3729 238 3805 272
rect 3729 204 3750 238
rect 3784 204 3805 238
rect 3729 203 3805 204
tri 3729 187 3745 203 ne
rect 3745 187 3789 203
tri 3789 187 3805 203 nw
rect 3835 257 3847 291
rect 3881 257 3894 291
tri 3894 288 3924 318 nw
rect 3835 223 3894 257
rect 3835 189 3847 223
rect 3881 189 3894 223
tri 3924 272 3940 288 se
rect 3940 272 3983 288
tri 3983 272 3999 288 sw
rect 3924 244 3999 272
rect 3924 210 3945 244
rect 3979 210 3999 244
tri 3924 194 3940 210 ne
rect 3940 194 3983 210
tri 3983 194 3999 210 nw
tri 3699 157 3729 187 sw
tri 3805 157 3835 187 se
rect 3835 164 3894 189
tri 3894 164 3924 194 sw
tri 3999 164 4029 194 se
rect 4029 164 4085 329
rect 3835 157 4085 164
rect 3643 153 4085 157
rect 3643 119 3653 153
rect 3687 119 3847 153
rect 3881 119 3944 153
rect 3978 119 4041 153
rect 4075 119 4085 153
rect 3643 103 4085 119
rect 4145 363 4201 379
rect 4145 329 4155 363
rect 4189 329 4201 363
rect 4145 291 4201 329
rect 4231 342 4393 379
tri 4231 326 4247 342 ne
rect 4247 326 4393 342
tri 4307 296 4337 326 ne
rect 4145 257 4155 291
rect 4189 257 4201 291
rect 4145 223 4201 257
rect 4145 189 4155 223
rect 4189 189 4201 223
tri 4231 280 4247 296 se
rect 4247 280 4291 296
tri 4291 280 4307 296 sw
rect 4231 247 4307 280
rect 4231 213 4252 247
rect 4286 213 4307 247
rect 4231 211 4307 213
tri 4231 195 4247 211 ne
rect 4247 195 4291 211
tri 4291 195 4307 211 nw
rect 4337 291 4393 326
rect 4337 257 4349 291
rect 4383 257 4393 291
rect 4337 223 4393 257
rect 4145 165 4201 189
tri 4201 165 4231 195 sw
tri 4307 165 4337 195 se
rect 4337 189 4349 223
rect 4383 189 4393 223
rect 4337 165 4393 189
rect 4145 153 4393 165
rect 4145 119 4155 153
rect 4189 119 4252 153
rect 4286 119 4349 153
rect 4383 119 4393 153
rect 4145 103 4393 119
rect 4626 361 4682 377
rect 4626 327 4636 361
rect 4670 327 4682 361
rect 4626 289 4682 327
rect 4712 361 4876 377
rect 4712 332 4733 361
tri 4712 316 4728 332 ne
rect 4728 327 4733 332
rect 4767 327 4830 361
rect 4864 327 4876 361
rect 4728 316 4876 327
rect 4906 340 5068 377
tri 4906 324 4922 340 ne
rect 4922 324 5068 340
rect 4626 255 4636 289
rect 4670 255 4682 289
tri 4788 286 4818 316 ne
rect 4818 289 4876 316
tri 4982 294 5012 324 ne
rect 4626 221 4682 255
rect 4626 187 4636 221
rect 4670 187 4682 221
rect 4626 155 4682 187
tri 4712 270 4728 286 se
rect 4728 270 4772 286
tri 4772 270 4788 286 sw
rect 4712 236 4788 270
rect 4712 202 4733 236
rect 4767 202 4788 236
rect 4712 201 4788 202
tri 4712 185 4728 201 ne
rect 4728 185 4772 201
tri 4772 185 4788 201 nw
rect 4818 255 4830 289
rect 4864 255 4876 289
rect 4818 221 4876 255
rect 4818 187 4830 221
rect 4864 187 4876 221
tri 4906 278 4922 294 se
rect 4922 278 4966 294
tri 4966 278 4982 294 sw
rect 4906 245 4982 278
rect 4906 211 4927 245
rect 4961 211 4982 245
rect 4906 209 4982 211
tri 4906 193 4922 209 ne
rect 4922 193 4966 209
tri 4966 193 4982 209 nw
rect 5012 289 5068 324
rect 5012 255 5024 289
rect 5058 255 5068 289
rect 5012 221 5068 255
tri 4682 155 4712 185 sw
tri 4788 155 4818 185 se
rect 4818 163 4876 187
tri 4876 163 4906 193 sw
tri 4982 163 5012 193 se
rect 5012 187 5024 221
rect 5058 187 5068 221
rect 5012 163 5068 187
rect 4818 155 5068 163
rect 4626 151 5068 155
rect 4626 117 4636 151
rect 4670 117 4830 151
rect 4864 117 4927 151
rect 4961 117 5024 151
rect 5058 117 5068 151
rect 4626 101 5068 117
<< pdiff >>
rect 191 1412 247 1450
rect 191 1378 201 1412
rect 235 1378 247 1412
rect 191 1344 247 1378
rect 191 1310 201 1344
rect 235 1310 247 1344
rect 191 1276 247 1310
rect 191 1242 201 1276
rect 235 1242 247 1276
rect 191 1208 247 1242
rect 191 1174 201 1208
rect 235 1174 247 1208
rect 191 1139 247 1174
rect 191 1105 201 1139
rect 235 1105 247 1139
rect 191 1050 247 1105
rect 277 1412 335 1450
rect 277 1378 289 1412
rect 323 1378 335 1412
rect 277 1344 335 1378
rect 277 1310 289 1344
rect 323 1310 335 1344
rect 277 1276 335 1310
rect 277 1242 289 1276
rect 323 1242 335 1276
rect 277 1208 335 1242
rect 277 1174 289 1208
rect 323 1174 335 1208
rect 277 1139 335 1174
rect 277 1105 289 1139
rect 323 1105 335 1139
rect 277 1050 335 1105
rect 365 1412 423 1450
rect 365 1378 377 1412
rect 411 1378 423 1412
rect 365 1344 423 1378
rect 365 1310 377 1344
rect 411 1310 423 1344
rect 365 1276 423 1310
rect 365 1242 377 1276
rect 411 1242 423 1276
rect 365 1208 423 1242
rect 365 1174 377 1208
rect 411 1174 423 1208
rect 365 1050 423 1174
rect 453 1412 511 1450
rect 453 1378 465 1412
rect 499 1378 511 1412
rect 453 1344 511 1378
rect 453 1310 465 1344
rect 499 1310 511 1344
rect 453 1276 511 1310
rect 453 1242 465 1276
rect 499 1242 511 1276
rect 453 1208 511 1242
rect 453 1174 465 1208
rect 499 1174 511 1208
rect 453 1139 511 1174
rect 453 1105 465 1139
rect 499 1105 511 1139
rect 453 1050 511 1105
rect 541 1412 599 1450
rect 541 1378 553 1412
rect 587 1378 599 1412
rect 541 1344 599 1378
rect 541 1310 553 1344
rect 587 1310 599 1344
rect 541 1276 599 1310
rect 541 1242 553 1276
rect 587 1242 599 1276
rect 541 1208 599 1242
rect 541 1174 553 1208
rect 587 1174 599 1208
rect 541 1050 599 1174
rect 629 1412 687 1450
rect 629 1378 641 1412
rect 675 1378 687 1412
rect 629 1344 687 1378
rect 629 1310 641 1344
rect 675 1310 687 1344
rect 629 1276 687 1310
rect 629 1242 641 1276
rect 675 1242 687 1276
rect 629 1208 687 1242
rect 629 1174 641 1208
rect 675 1174 687 1208
rect 629 1139 687 1174
rect 629 1105 641 1139
rect 675 1105 687 1139
rect 629 1050 687 1105
rect 717 1412 771 1450
rect 717 1378 729 1412
rect 763 1378 771 1412
rect 717 1344 771 1378
rect 717 1310 729 1344
rect 763 1310 771 1344
rect 717 1276 771 1310
rect 717 1242 729 1276
rect 763 1242 771 1276
rect 717 1208 771 1242
rect 717 1174 729 1208
rect 763 1174 771 1208
rect 717 1050 771 1174
rect 1153 1412 1209 1450
rect 1153 1378 1163 1412
rect 1197 1378 1209 1412
rect 1153 1344 1209 1378
rect 1153 1310 1163 1344
rect 1197 1310 1209 1344
rect 1153 1276 1209 1310
rect 1153 1242 1163 1276
rect 1197 1242 1209 1276
rect 1153 1208 1209 1242
rect 1153 1174 1163 1208
rect 1197 1174 1209 1208
rect 1153 1139 1209 1174
rect 1153 1105 1163 1139
rect 1197 1105 1209 1139
rect 1153 1050 1209 1105
rect 1239 1412 1297 1450
rect 1239 1378 1251 1412
rect 1285 1378 1297 1412
rect 1239 1344 1297 1378
rect 1239 1310 1251 1344
rect 1285 1310 1297 1344
rect 1239 1276 1297 1310
rect 1239 1242 1251 1276
rect 1285 1242 1297 1276
rect 1239 1208 1297 1242
rect 1239 1174 1251 1208
rect 1285 1174 1297 1208
rect 1239 1139 1297 1174
rect 1239 1105 1251 1139
rect 1285 1105 1297 1139
rect 1239 1050 1297 1105
rect 1327 1412 1385 1450
rect 1327 1378 1339 1412
rect 1373 1378 1385 1412
rect 1327 1344 1385 1378
rect 1327 1310 1339 1344
rect 1373 1310 1385 1344
rect 1327 1276 1385 1310
rect 1327 1242 1339 1276
rect 1373 1242 1385 1276
rect 1327 1208 1385 1242
rect 1327 1174 1339 1208
rect 1373 1174 1385 1208
rect 1327 1050 1385 1174
rect 1415 1412 1473 1450
rect 1415 1378 1427 1412
rect 1461 1378 1473 1412
rect 1415 1344 1473 1378
rect 1415 1310 1427 1344
rect 1461 1310 1473 1344
rect 1415 1276 1473 1310
rect 1415 1242 1427 1276
rect 1461 1242 1473 1276
rect 1415 1208 1473 1242
rect 1415 1174 1427 1208
rect 1461 1174 1473 1208
rect 1415 1139 1473 1174
rect 1415 1105 1427 1139
rect 1461 1105 1473 1139
rect 1415 1050 1473 1105
rect 1503 1412 1561 1450
rect 1503 1378 1515 1412
rect 1549 1378 1561 1412
rect 1503 1344 1561 1378
rect 1503 1310 1515 1344
rect 1549 1310 1561 1344
rect 1503 1276 1561 1310
rect 1503 1242 1515 1276
rect 1549 1242 1561 1276
rect 1503 1208 1561 1242
rect 1503 1174 1515 1208
rect 1549 1174 1561 1208
rect 1503 1050 1561 1174
rect 1591 1412 1649 1450
rect 1591 1378 1603 1412
rect 1637 1378 1649 1412
rect 1591 1344 1649 1378
rect 1591 1310 1603 1344
rect 1637 1310 1649 1344
rect 1591 1276 1649 1310
rect 1591 1242 1603 1276
rect 1637 1242 1649 1276
rect 1591 1208 1649 1242
rect 1591 1174 1603 1208
rect 1637 1174 1649 1208
rect 1591 1139 1649 1174
rect 1591 1105 1603 1139
rect 1637 1105 1649 1139
rect 1591 1050 1649 1105
rect 1679 1412 1733 1450
rect 1679 1378 1691 1412
rect 1725 1378 1733 1412
rect 1679 1344 1733 1378
rect 1679 1310 1691 1344
rect 1725 1310 1733 1344
rect 1679 1276 1733 1310
rect 1679 1242 1691 1276
rect 1725 1242 1733 1276
rect 1679 1208 1733 1242
rect 1679 1174 1691 1208
rect 1725 1174 1733 1208
rect 1679 1050 1733 1174
rect 2055 1412 2111 1450
rect 2055 1378 2065 1412
rect 2099 1378 2111 1412
rect 2055 1344 2111 1378
rect 2055 1310 2065 1344
rect 2099 1310 2111 1344
rect 2055 1276 2111 1310
rect 2055 1242 2065 1276
rect 2099 1242 2111 1276
rect 2055 1208 2111 1242
rect 2055 1174 2065 1208
rect 2099 1174 2111 1208
rect 2055 1139 2111 1174
rect 2055 1105 2065 1139
rect 2099 1105 2111 1139
rect 2055 1050 2111 1105
rect 2141 1412 2199 1450
rect 2141 1378 2153 1412
rect 2187 1378 2199 1412
rect 2141 1344 2199 1378
rect 2141 1310 2153 1344
rect 2187 1310 2199 1344
rect 2141 1276 2199 1310
rect 2141 1242 2153 1276
rect 2187 1242 2199 1276
rect 2141 1208 2199 1242
rect 2141 1174 2153 1208
rect 2187 1174 2199 1208
rect 2141 1139 2199 1174
rect 2141 1105 2153 1139
rect 2187 1105 2199 1139
rect 2141 1050 2199 1105
rect 2229 1412 2287 1450
rect 2229 1378 2241 1412
rect 2275 1378 2287 1412
rect 2229 1344 2287 1378
rect 2229 1310 2241 1344
rect 2275 1310 2287 1344
rect 2229 1276 2287 1310
rect 2229 1242 2241 1276
rect 2275 1242 2287 1276
rect 2229 1208 2287 1242
rect 2229 1174 2241 1208
rect 2275 1174 2287 1208
rect 2229 1050 2287 1174
rect 2317 1412 2375 1450
rect 2317 1378 2329 1412
rect 2363 1378 2375 1412
rect 2317 1344 2375 1378
rect 2317 1310 2329 1344
rect 2363 1310 2375 1344
rect 2317 1276 2375 1310
rect 2317 1242 2329 1276
rect 2363 1242 2375 1276
rect 2317 1208 2375 1242
rect 2317 1174 2329 1208
rect 2363 1174 2375 1208
rect 2317 1139 2375 1174
rect 2317 1105 2329 1139
rect 2363 1105 2375 1139
rect 2317 1050 2375 1105
rect 2405 1412 2459 1450
rect 2405 1378 2417 1412
rect 2451 1378 2459 1412
rect 2405 1344 2459 1378
rect 2405 1310 2417 1344
rect 2451 1310 2459 1344
rect 2405 1276 2459 1310
rect 2405 1242 2417 1276
rect 2451 1242 2459 1276
rect 2405 1208 2459 1242
rect 2405 1174 2417 1208
rect 2451 1174 2459 1208
rect 2405 1050 2459 1174
rect 2781 1412 2837 1450
rect 2781 1378 2791 1412
rect 2825 1378 2837 1412
rect 2781 1344 2837 1378
rect 2781 1310 2791 1344
rect 2825 1310 2837 1344
rect 2781 1276 2837 1310
rect 2781 1242 2791 1276
rect 2825 1242 2837 1276
rect 2781 1208 2837 1242
rect 2781 1174 2791 1208
rect 2825 1174 2837 1208
rect 2781 1139 2837 1174
rect 2781 1105 2791 1139
rect 2825 1105 2837 1139
rect 2781 1050 2837 1105
rect 2867 1412 2925 1450
rect 2867 1378 2879 1412
rect 2913 1378 2925 1412
rect 2867 1344 2925 1378
rect 2867 1310 2879 1344
rect 2913 1310 2925 1344
rect 2867 1276 2925 1310
rect 2867 1242 2879 1276
rect 2913 1242 2925 1276
rect 2867 1208 2925 1242
rect 2867 1174 2879 1208
rect 2913 1174 2925 1208
rect 2867 1139 2925 1174
rect 2867 1105 2879 1139
rect 2913 1105 2925 1139
rect 2867 1050 2925 1105
rect 2955 1412 3013 1450
rect 2955 1378 2967 1412
rect 3001 1378 3013 1412
rect 2955 1344 3013 1378
rect 2955 1310 2967 1344
rect 3001 1310 3013 1344
rect 2955 1276 3013 1310
rect 2955 1242 2967 1276
rect 3001 1242 3013 1276
rect 2955 1208 3013 1242
rect 2955 1174 2967 1208
rect 3001 1174 3013 1208
rect 2955 1050 3013 1174
rect 3043 1412 3101 1450
rect 3043 1378 3055 1412
rect 3089 1378 3101 1412
rect 3043 1344 3101 1378
rect 3043 1310 3055 1344
rect 3089 1310 3101 1344
rect 3043 1276 3101 1310
rect 3043 1242 3055 1276
rect 3089 1242 3101 1276
rect 3043 1208 3101 1242
rect 3043 1174 3055 1208
rect 3089 1174 3101 1208
rect 3043 1139 3101 1174
rect 3043 1105 3055 1139
rect 3089 1105 3101 1139
rect 3043 1050 3101 1105
rect 3131 1412 3189 1450
rect 3131 1378 3143 1412
rect 3177 1378 3189 1412
rect 3131 1344 3189 1378
rect 3131 1310 3143 1344
rect 3177 1310 3189 1344
rect 3131 1276 3189 1310
rect 3131 1242 3143 1276
rect 3177 1242 3189 1276
rect 3131 1208 3189 1242
rect 3131 1174 3143 1208
rect 3177 1174 3189 1208
rect 3131 1050 3189 1174
rect 3219 1412 3277 1450
rect 3219 1378 3231 1412
rect 3265 1378 3277 1412
rect 3219 1344 3277 1378
rect 3219 1310 3231 1344
rect 3265 1310 3277 1344
rect 3219 1276 3277 1310
rect 3219 1242 3231 1276
rect 3265 1242 3277 1276
rect 3219 1208 3277 1242
rect 3219 1174 3231 1208
rect 3265 1174 3277 1208
rect 3219 1139 3277 1174
rect 3219 1105 3231 1139
rect 3265 1105 3277 1139
rect 3219 1050 3277 1105
rect 3307 1412 3361 1450
rect 3307 1378 3319 1412
rect 3353 1378 3361 1412
rect 3307 1344 3361 1378
rect 3307 1310 3319 1344
rect 3353 1310 3361 1344
rect 3307 1276 3361 1310
rect 3307 1242 3319 1276
rect 3353 1242 3361 1276
rect 3307 1208 3361 1242
rect 3307 1174 3319 1208
rect 3353 1174 3361 1208
rect 3307 1050 3361 1174
rect 3743 1412 3799 1450
rect 3743 1378 3753 1412
rect 3787 1378 3799 1412
rect 3743 1344 3799 1378
rect 3743 1310 3753 1344
rect 3787 1310 3799 1344
rect 3743 1276 3799 1310
rect 3743 1242 3753 1276
rect 3787 1242 3799 1276
rect 3743 1208 3799 1242
rect 3743 1174 3753 1208
rect 3787 1174 3799 1208
rect 3743 1139 3799 1174
rect 3743 1105 3753 1139
rect 3787 1105 3799 1139
rect 3743 1050 3799 1105
rect 3829 1412 3887 1450
rect 3829 1378 3841 1412
rect 3875 1378 3887 1412
rect 3829 1344 3887 1378
rect 3829 1310 3841 1344
rect 3875 1310 3887 1344
rect 3829 1276 3887 1310
rect 3829 1242 3841 1276
rect 3875 1242 3887 1276
rect 3829 1208 3887 1242
rect 3829 1174 3841 1208
rect 3875 1174 3887 1208
rect 3829 1139 3887 1174
rect 3829 1105 3841 1139
rect 3875 1105 3887 1139
rect 3829 1050 3887 1105
rect 3917 1412 3975 1450
rect 3917 1378 3929 1412
rect 3963 1378 3975 1412
rect 3917 1344 3975 1378
rect 3917 1310 3929 1344
rect 3963 1310 3975 1344
rect 3917 1276 3975 1310
rect 3917 1242 3929 1276
rect 3963 1242 3975 1276
rect 3917 1208 3975 1242
rect 3917 1174 3929 1208
rect 3963 1174 3975 1208
rect 3917 1050 3975 1174
rect 4005 1412 4063 1450
rect 4005 1378 4017 1412
rect 4051 1378 4063 1412
rect 4005 1344 4063 1378
rect 4005 1310 4017 1344
rect 4051 1310 4063 1344
rect 4005 1276 4063 1310
rect 4005 1242 4017 1276
rect 4051 1242 4063 1276
rect 4005 1208 4063 1242
rect 4005 1174 4017 1208
rect 4051 1174 4063 1208
rect 4005 1139 4063 1174
rect 4005 1105 4017 1139
rect 4051 1105 4063 1139
rect 4005 1050 4063 1105
rect 4093 1412 4151 1450
rect 4093 1378 4105 1412
rect 4139 1378 4151 1412
rect 4093 1344 4151 1378
rect 4093 1310 4105 1344
rect 4139 1310 4151 1344
rect 4093 1276 4151 1310
rect 4093 1242 4105 1276
rect 4139 1242 4151 1276
rect 4093 1208 4151 1242
rect 4093 1174 4105 1208
rect 4139 1174 4151 1208
rect 4093 1050 4151 1174
rect 4181 1412 4239 1450
rect 4181 1378 4193 1412
rect 4227 1378 4239 1412
rect 4181 1344 4239 1378
rect 4181 1310 4193 1344
rect 4227 1310 4239 1344
rect 4181 1276 4239 1310
rect 4181 1242 4193 1276
rect 4227 1242 4239 1276
rect 4181 1208 4239 1242
rect 4181 1174 4193 1208
rect 4227 1174 4239 1208
rect 4181 1139 4239 1174
rect 4181 1105 4193 1139
rect 4227 1105 4239 1139
rect 4181 1050 4239 1105
rect 4269 1412 4323 1450
rect 4269 1378 4281 1412
rect 4315 1378 4323 1412
rect 4269 1344 4323 1378
rect 4269 1310 4281 1344
rect 4315 1310 4323 1344
rect 4269 1276 4323 1310
rect 4269 1242 4281 1276
rect 4315 1242 4323 1276
rect 4269 1208 4323 1242
rect 4269 1174 4281 1208
rect 4315 1174 4323 1208
rect 4269 1050 4323 1174
rect 4645 1412 4701 1450
rect 4645 1378 4655 1412
rect 4689 1378 4701 1412
rect 4645 1344 4701 1378
rect 4645 1310 4655 1344
rect 4689 1310 4701 1344
rect 4645 1276 4701 1310
rect 4645 1242 4655 1276
rect 4689 1242 4701 1276
rect 4645 1208 4701 1242
rect 4645 1174 4655 1208
rect 4689 1174 4701 1208
rect 4645 1139 4701 1174
rect 4645 1105 4655 1139
rect 4689 1105 4701 1139
rect 4645 1050 4701 1105
rect 4731 1412 4789 1450
rect 4731 1378 4743 1412
rect 4777 1378 4789 1412
rect 4731 1344 4789 1378
rect 4731 1310 4743 1344
rect 4777 1310 4789 1344
rect 4731 1276 4789 1310
rect 4731 1242 4743 1276
rect 4777 1242 4789 1276
rect 4731 1208 4789 1242
rect 4731 1174 4743 1208
rect 4777 1174 4789 1208
rect 4731 1139 4789 1174
rect 4731 1105 4743 1139
rect 4777 1105 4789 1139
rect 4731 1050 4789 1105
rect 4819 1412 4877 1450
rect 4819 1378 4831 1412
rect 4865 1378 4877 1412
rect 4819 1344 4877 1378
rect 4819 1310 4831 1344
rect 4865 1310 4877 1344
rect 4819 1276 4877 1310
rect 4819 1242 4831 1276
rect 4865 1242 4877 1276
rect 4819 1208 4877 1242
rect 4819 1174 4831 1208
rect 4865 1174 4877 1208
rect 4819 1050 4877 1174
rect 4907 1412 4965 1450
rect 4907 1378 4919 1412
rect 4953 1378 4965 1412
rect 4907 1344 4965 1378
rect 4907 1310 4919 1344
rect 4953 1310 4965 1344
rect 4907 1276 4965 1310
rect 4907 1242 4919 1276
rect 4953 1242 4965 1276
rect 4907 1208 4965 1242
rect 4907 1174 4919 1208
rect 4953 1174 4965 1208
rect 4907 1139 4965 1174
rect 4907 1105 4919 1139
rect 4953 1105 4965 1139
rect 4907 1050 4965 1105
rect 4995 1412 5049 1450
rect 4995 1378 5007 1412
rect 5041 1378 5049 1412
rect 4995 1344 5049 1378
rect 4995 1310 5007 1344
rect 5041 1310 5049 1344
rect 4995 1276 5049 1310
rect 4995 1242 5007 1276
rect 5041 1242 5049 1276
rect 4995 1208 5049 1242
rect 4995 1174 5007 1208
rect 5041 1174 5049 1208
rect 4995 1050 5049 1174
<< ndiffc >>
rect 101 329 135 363
rect 198 329 232 363
rect 295 329 329 363
rect 392 329 426 363
rect 489 329 523 363
rect 101 257 135 291
rect 101 189 135 223
rect 198 204 232 238
rect 295 257 329 291
rect 295 189 329 223
rect 393 210 427 244
rect 101 119 135 153
rect 295 119 329 153
rect 392 119 426 153
rect 489 119 523 153
rect 603 329 637 363
rect 603 257 637 291
rect 603 189 637 223
rect 700 213 734 247
rect 797 257 831 291
rect 797 189 831 223
rect 603 119 637 153
rect 700 119 734 153
rect 797 119 831 153
rect 1063 329 1097 363
rect 1160 329 1194 363
rect 1257 329 1291 363
rect 1354 329 1388 363
rect 1451 329 1485 363
rect 1063 257 1097 291
rect 1063 189 1097 223
rect 1160 204 1194 238
rect 1257 257 1291 291
rect 1257 189 1291 223
rect 1355 210 1389 244
rect 1063 119 1097 153
rect 1257 119 1291 153
rect 1354 119 1388 153
rect 1451 119 1485 153
rect 1565 329 1599 363
rect 1565 257 1599 291
rect 1565 189 1599 223
rect 1662 213 1696 247
rect 1759 257 1793 291
rect 1759 189 1793 223
rect 1565 119 1599 153
rect 1662 119 1696 153
rect 1759 119 1793 153
rect 2046 327 2080 361
rect 2143 327 2177 361
rect 2240 327 2274 361
rect 2046 255 2080 289
rect 2046 187 2080 221
rect 2143 202 2177 236
rect 2240 255 2274 289
rect 2240 187 2274 221
rect 2337 211 2371 245
rect 2434 255 2468 289
rect 2434 187 2468 221
rect 2046 117 2080 151
rect 2240 117 2274 151
rect 2337 117 2371 151
rect 2434 117 2468 151
rect 2691 329 2725 363
rect 2788 329 2822 363
rect 2885 329 2919 363
rect 2982 329 3016 363
rect 3079 329 3113 363
rect 2691 257 2725 291
rect 2691 189 2725 223
rect 2788 204 2822 238
rect 2885 257 2919 291
rect 2885 189 2919 223
rect 2983 210 3017 244
rect 2691 119 2725 153
rect 2885 119 2919 153
rect 2982 119 3016 153
rect 3079 119 3113 153
rect 3193 329 3227 363
rect 3193 257 3227 291
rect 3193 189 3227 223
rect 3290 213 3324 247
rect 3387 257 3421 291
rect 3387 189 3421 223
rect 3193 119 3227 153
rect 3290 119 3324 153
rect 3387 119 3421 153
rect 3653 329 3687 363
rect 3750 329 3784 363
rect 3847 329 3881 363
rect 3944 329 3978 363
rect 4041 329 4075 363
rect 3653 257 3687 291
rect 3653 189 3687 223
rect 3750 204 3784 238
rect 3847 257 3881 291
rect 3847 189 3881 223
rect 3945 210 3979 244
rect 3653 119 3687 153
rect 3847 119 3881 153
rect 3944 119 3978 153
rect 4041 119 4075 153
rect 4155 329 4189 363
rect 4155 257 4189 291
rect 4155 189 4189 223
rect 4252 213 4286 247
rect 4349 257 4383 291
rect 4349 189 4383 223
rect 4155 119 4189 153
rect 4252 119 4286 153
rect 4349 119 4383 153
rect 4636 327 4670 361
rect 4733 327 4767 361
rect 4830 327 4864 361
rect 4636 255 4670 289
rect 4636 187 4670 221
rect 4733 202 4767 236
rect 4830 255 4864 289
rect 4830 187 4864 221
rect 4927 211 4961 245
rect 5024 255 5058 289
rect 5024 187 5058 221
rect 4636 117 4670 151
rect 4830 117 4864 151
rect 4927 117 4961 151
rect 5024 117 5058 151
<< pdiffc >>
rect 201 1378 235 1412
rect 201 1310 235 1344
rect 201 1242 235 1276
rect 201 1174 235 1208
rect 201 1105 235 1139
rect 289 1378 323 1412
rect 289 1310 323 1344
rect 289 1242 323 1276
rect 289 1174 323 1208
rect 289 1105 323 1139
rect 377 1378 411 1412
rect 377 1310 411 1344
rect 377 1242 411 1276
rect 377 1174 411 1208
rect 465 1378 499 1412
rect 465 1310 499 1344
rect 465 1242 499 1276
rect 465 1174 499 1208
rect 465 1105 499 1139
rect 553 1378 587 1412
rect 553 1310 587 1344
rect 553 1242 587 1276
rect 553 1174 587 1208
rect 641 1378 675 1412
rect 641 1310 675 1344
rect 641 1242 675 1276
rect 641 1174 675 1208
rect 641 1105 675 1139
rect 729 1378 763 1412
rect 729 1310 763 1344
rect 729 1242 763 1276
rect 729 1174 763 1208
rect 1163 1378 1197 1412
rect 1163 1310 1197 1344
rect 1163 1242 1197 1276
rect 1163 1174 1197 1208
rect 1163 1105 1197 1139
rect 1251 1378 1285 1412
rect 1251 1310 1285 1344
rect 1251 1242 1285 1276
rect 1251 1174 1285 1208
rect 1251 1105 1285 1139
rect 1339 1378 1373 1412
rect 1339 1310 1373 1344
rect 1339 1242 1373 1276
rect 1339 1174 1373 1208
rect 1427 1378 1461 1412
rect 1427 1310 1461 1344
rect 1427 1242 1461 1276
rect 1427 1174 1461 1208
rect 1427 1105 1461 1139
rect 1515 1378 1549 1412
rect 1515 1310 1549 1344
rect 1515 1242 1549 1276
rect 1515 1174 1549 1208
rect 1603 1378 1637 1412
rect 1603 1310 1637 1344
rect 1603 1242 1637 1276
rect 1603 1174 1637 1208
rect 1603 1105 1637 1139
rect 1691 1378 1725 1412
rect 1691 1310 1725 1344
rect 1691 1242 1725 1276
rect 1691 1174 1725 1208
rect 2065 1378 2099 1412
rect 2065 1310 2099 1344
rect 2065 1242 2099 1276
rect 2065 1174 2099 1208
rect 2065 1105 2099 1139
rect 2153 1378 2187 1412
rect 2153 1310 2187 1344
rect 2153 1242 2187 1276
rect 2153 1174 2187 1208
rect 2153 1105 2187 1139
rect 2241 1378 2275 1412
rect 2241 1310 2275 1344
rect 2241 1242 2275 1276
rect 2241 1174 2275 1208
rect 2329 1378 2363 1412
rect 2329 1310 2363 1344
rect 2329 1242 2363 1276
rect 2329 1174 2363 1208
rect 2329 1105 2363 1139
rect 2417 1378 2451 1412
rect 2417 1310 2451 1344
rect 2417 1242 2451 1276
rect 2417 1174 2451 1208
rect 2791 1378 2825 1412
rect 2791 1310 2825 1344
rect 2791 1242 2825 1276
rect 2791 1174 2825 1208
rect 2791 1105 2825 1139
rect 2879 1378 2913 1412
rect 2879 1310 2913 1344
rect 2879 1242 2913 1276
rect 2879 1174 2913 1208
rect 2879 1105 2913 1139
rect 2967 1378 3001 1412
rect 2967 1310 3001 1344
rect 2967 1242 3001 1276
rect 2967 1174 3001 1208
rect 3055 1378 3089 1412
rect 3055 1310 3089 1344
rect 3055 1242 3089 1276
rect 3055 1174 3089 1208
rect 3055 1105 3089 1139
rect 3143 1378 3177 1412
rect 3143 1310 3177 1344
rect 3143 1242 3177 1276
rect 3143 1174 3177 1208
rect 3231 1378 3265 1412
rect 3231 1310 3265 1344
rect 3231 1242 3265 1276
rect 3231 1174 3265 1208
rect 3231 1105 3265 1139
rect 3319 1378 3353 1412
rect 3319 1310 3353 1344
rect 3319 1242 3353 1276
rect 3319 1174 3353 1208
rect 3753 1378 3787 1412
rect 3753 1310 3787 1344
rect 3753 1242 3787 1276
rect 3753 1174 3787 1208
rect 3753 1105 3787 1139
rect 3841 1378 3875 1412
rect 3841 1310 3875 1344
rect 3841 1242 3875 1276
rect 3841 1174 3875 1208
rect 3841 1105 3875 1139
rect 3929 1378 3963 1412
rect 3929 1310 3963 1344
rect 3929 1242 3963 1276
rect 3929 1174 3963 1208
rect 4017 1378 4051 1412
rect 4017 1310 4051 1344
rect 4017 1242 4051 1276
rect 4017 1174 4051 1208
rect 4017 1105 4051 1139
rect 4105 1378 4139 1412
rect 4105 1310 4139 1344
rect 4105 1242 4139 1276
rect 4105 1174 4139 1208
rect 4193 1378 4227 1412
rect 4193 1310 4227 1344
rect 4193 1242 4227 1276
rect 4193 1174 4227 1208
rect 4193 1105 4227 1139
rect 4281 1378 4315 1412
rect 4281 1310 4315 1344
rect 4281 1242 4315 1276
rect 4281 1174 4315 1208
rect 4655 1378 4689 1412
rect 4655 1310 4689 1344
rect 4655 1242 4689 1276
rect 4655 1174 4689 1208
rect 4655 1105 4689 1139
rect 4743 1378 4777 1412
rect 4743 1310 4777 1344
rect 4743 1242 4777 1276
rect 4743 1174 4777 1208
rect 4743 1105 4777 1139
rect 4831 1378 4865 1412
rect 4831 1310 4865 1344
rect 4831 1242 4865 1276
rect 4831 1174 4865 1208
rect 4919 1378 4953 1412
rect 4919 1310 4953 1344
rect 4919 1242 4953 1276
rect 4919 1174 4953 1208
rect 4919 1105 4953 1139
rect 5007 1378 5041 1412
rect 5007 1310 5041 1344
rect 5007 1242 5041 1276
rect 5007 1174 5041 1208
<< psubdiff >>
rect -31 546 5211 572
rect -31 512 -17 546
rect 17 512 945 546
rect 979 512 1907 546
rect 1941 512 2573 546
rect 2607 512 3535 546
rect 3569 512 4497 546
rect 4531 512 5163 546
rect 5197 512 5211 546
rect -31 510 5211 512
rect -31 474 31 510
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect -31 368 -17 402
rect 17 368 31 402
rect 931 474 993 510
rect 931 440 945 474
rect 979 440 993 474
rect 931 402 993 440
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect 931 368 945 402
rect 979 368 993 402
rect 1893 474 1955 510
rect 1893 440 1907 474
rect 1941 440 1955 474
rect 1893 402 1955 440
rect 931 330 993 368
rect 931 296 945 330
rect 979 296 993 330
rect 931 258 993 296
rect 931 224 945 258
rect 979 224 993 258
rect 931 186 993 224
rect 931 152 945 186
rect 979 152 993 186
rect 931 114 993 152
rect -31 47 31 80
rect 931 80 945 114
rect 979 80 993 114
rect 1893 368 1907 402
rect 1941 368 1955 402
rect 2559 474 2621 510
rect 2559 440 2573 474
rect 2607 440 2621 474
rect 2559 402 2621 440
rect 1893 330 1955 368
rect 1893 296 1907 330
rect 1941 296 1955 330
rect 1893 258 1955 296
rect 1893 224 1907 258
rect 1941 224 1955 258
rect 1893 186 1955 224
rect 1893 152 1907 186
rect 1941 152 1955 186
rect 1893 114 1955 152
rect 931 47 993 80
rect 1893 80 1907 114
rect 1941 80 1955 114
rect 2559 368 2573 402
rect 2607 368 2621 402
rect 3521 474 3583 510
rect 3521 440 3535 474
rect 3569 440 3583 474
rect 3521 402 3583 440
rect 2559 330 2621 368
rect 2559 296 2573 330
rect 2607 296 2621 330
rect 2559 258 2621 296
rect 2559 224 2573 258
rect 2607 224 2621 258
rect 2559 186 2621 224
rect 2559 152 2573 186
rect 2607 152 2621 186
rect 2559 114 2621 152
rect 1893 47 1955 80
rect 2559 80 2573 114
rect 2607 80 2621 114
rect 3521 368 3535 402
rect 3569 368 3583 402
rect 4483 474 4545 510
rect 4483 440 4497 474
rect 4531 440 4545 474
rect 4483 402 4545 440
rect 3521 330 3583 368
rect 3521 296 3535 330
rect 3569 296 3583 330
rect 3521 258 3583 296
rect 3521 224 3535 258
rect 3569 224 3583 258
rect 3521 186 3583 224
rect 3521 152 3535 186
rect 3569 152 3583 186
rect 3521 114 3583 152
rect 2559 47 2621 80
rect 3521 80 3535 114
rect 3569 80 3583 114
rect 4483 368 4497 402
rect 4531 368 4545 402
rect 5149 474 5211 510
rect 5149 440 5163 474
rect 5197 440 5211 474
rect 5149 402 5211 440
rect 4483 330 4545 368
rect 4483 296 4497 330
rect 4531 296 4545 330
rect 4483 258 4545 296
rect 4483 224 4497 258
rect 4531 224 4545 258
rect 4483 186 4545 224
rect 4483 152 4497 186
rect 4531 152 4545 186
rect 4483 114 4545 152
rect 3521 47 3583 80
rect 4483 80 4497 114
rect 4531 80 4545 114
rect 5149 368 5163 402
rect 5197 368 5211 402
rect 5149 330 5211 368
rect 5149 296 5163 330
rect 5197 296 5211 330
rect 5149 258 5211 296
rect 5149 224 5163 258
rect 5197 224 5211 258
rect 5149 186 5211 224
rect 5149 152 5163 186
rect 5197 152 5211 186
rect 5149 114 5211 152
rect 4483 47 4545 80
rect 5149 80 5163 114
rect 5197 80 5211 114
rect 5149 47 5211 80
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 343 47
rect 377 13 415 47
rect 449 13 513 47
rect 547 13 585 47
rect 619 13 657 47
rect 691 13 729 47
rect 763 13 801 47
rect 835 13 873 47
rect 907 13 1017 47
rect 1051 13 1089 47
rect 1123 13 1161 47
rect 1195 13 1233 47
rect 1267 13 1305 47
rect 1339 13 1377 47
rect 1411 13 1475 47
rect 1509 13 1547 47
rect 1581 13 1619 47
rect 1653 13 1691 47
rect 1725 13 1763 47
rect 1797 13 1835 47
rect 1869 13 1979 47
rect 2013 13 2051 47
rect 2085 13 2123 47
rect 2157 13 2195 47
rect 2229 13 2285 47
rect 2319 13 2357 47
rect 2391 13 2429 47
rect 2463 13 2501 47
rect 2535 13 2645 47
rect 2679 13 2717 47
rect 2751 13 2789 47
rect 2823 13 2861 47
rect 2895 13 2933 47
rect 2967 13 3005 47
rect 3039 13 3103 47
rect 3137 13 3175 47
rect 3209 13 3247 47
rect 3281 13 3319 47
rect 3353 13 3391 47
rect 3425 13 3463 47
rect 3497 13 3607 47
rect 3641 13 3679 47
rect 3713 13 3751 47
rect 3785 13 3823 47
rect 3857 13 3895 47
rect 3929 13 3967 47
rect 4001 13 4065 47
rect 4099 13 4137 47
rect 4171 13 4209 47
rect 4243 13 4281 47
rect 4315 13 4353 47
rect 4387 13 4425 47
rect 4459 13 4569 47
rect 4603 13 4641 47
rect 4675 13 4713 47
rect 4747 13 4785 47
rect 4819 13 4875 47
rect 4909 13 4947 47
rect 4981 13 5019 47
rect 5053 13 5091 47
rect 5125 13 5211 47
rect -31 11 31 13
rect 931 11 993 13
rect 1893 11 1955 13
rect 2559 11 2621 13
rect 3521 11 3583 13
rect 4483 11 4545 13
rect 5149 11 5211 13
<< nsubdiff >>
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 343 1539
rect 377 1505 415 1539
rect 449 1505 513 1539
rect 547 1505 585 1539
rect 619 1505 657 1539
rect 691 1505 729 1539
rect 763 1505 801 1539
rect 835 1505 873 1539
rect 907 1505 1017 1539
rect 1051 1505 1089 1539
rect 1123 1505 1161 1539
rect 1195 1505 1233 1539
rect 1267 1505 1305 1539
rect 1339 1505 1377 1539
rect 1411 1505 1475 1539
rect 1509 1505 1547 1539
rect 1581 1505 1619 1539
rect 1653 1505 1691 1539
rect 1725 1505 1763 1539
rect 1797 1505 1835 1539
rect 1869 1505 1979 1539
rect 2013 1505 2051 1539
rect 2085 1505 2123 1539
rect 2157 1505 2195 1539
rect 2229 1505 2285 1539
rect 2319 1505 2357 1539
rect 2391 1505 2429 1539
rect 2463 1505 2501 1539
rect 2535 1505 2645 1539
rect 2679 1505 2717 1539
rect 2751 1505 2789 1539
rect 2823 1505 2861 1539
rect 2895 1505 2933 1539
rect 2967 1505 3005 1539
rect 3039 1505 3103 1539
rect 3137 1505 3175 1539
rect 3209 1505 3247 1539
rect 3281 1505 3319 1539
rect 3353 1505 3391 1539
rect 3425 1505 3463 1539
rect 3497 1505 3607 1539
rect 3641 1505 3679 1539
rect 3713 1505 3751 1539
rect 3785 1505 3823 1539
rect 3857 1505 3895 1539
rect 3929 1505 3967 1539
rect 4001 1505 4065 1539
rect 4099 1505 4137 1539
rect 4171 1505 4209 1539
rect 4243 1505 4281 1539
rect 4315 1505 4353 1539
rect 4387 1505 4425 1539
rect 4459 1505 4569 1539
rect 4603 1505 4641 1539
rect 4675 1505 4713 1539
rect 4747 1505 4785 1539
rect 4819 1505 4875 1539
rect 4909 1505 4947 1539
rect 4981 1505 5019 1539
rect 5053 1505 5091 1539
rect 5125 1505 5211 1539
rect -31 1470 31 1505
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect 931 1470 993 1505
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect -31 1038 31 1076
rect 931 1436 945 1470
rect 979 1436 993 1470
rect 1893 1470 1955 1505
rect 931 1398 993 1436
rect 931 1364 945 1398
rect 979 1364 993 1398
rect 931 1326 993 1364
rect 931 1292 945 1326
rect 979 1292 993 1326
rect 931 1254 993 1292
rect 931 1220 945 1254
rect 979 1220 993 1254
rect 931 1182 993 1220
rect 931 1148 945 1182
rect 979 1148 993 1182
rect 931 1110 993 1148
rect 931 1076 945 1110
rect 979 1076 993 1110
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect 931 1038 993 1076
rect 1893 1436 1907 1470
rect 1941 1436 1955 1470
rect 2559 1470 2621 1505
rect 1893 1398 1955 1436
rect 1893 1364 1907 1398
rect 1941 1364 1955 1398
rect 1893 1326 1955 1364
rect 1893 1292 1907 1326
rect 1941 1292 1955 1326
rect 1893 1254 1955 1292
rect 1893 1220 1907 1254
rect 1941 1220 1955 1254
rect 1893 1182 1955 1220
rect 1893 1148 1907 1182
rect 1941 1148 1955 1182
rect 1893 1110 1955 1148
rect 1893 1076 1907 1110
rect 1941 1076 1955 1110
rect 931 1004 945 1038
rect 979 1004 993 1038
rect 931 966 993 1004
rect -31 930 31 932
rect 931 932 945 966
rect 979 932 993 966
rect 1893 1038 1955 1076
rect 2559 1436 2573 1470
rect 2607 1436 2621 1470
rect 3521 1470 3583 1505
rect 2559 1398 2621 1436
rect 2559 1364 2573 1398
rect 2607 1364 2621 1398
rect 2559 1326 2621 1364
rect 2559 1292 2573 1326
rect 2607 1292 2621 1326
rect 2559 1254 2621 1292
rect 2559 1220 2573 1254
rect 2607 1220 2621 1254
rect 2559 1182 2621 1220
rect 2559 1148 2573 1182
rect 2607 1148 2621 1182
rect 2559 1110 2621 1148
rect 2559 1076 2573 1110
rect 2607 1076 2621 1110
rect 1893 1004 1907 1038
rect 1941 1004 1955 1038
rect 1893 966 1955 1004
rect 931 930 993 932
rect 1893 932 1907 966
rect 1941 932 1955 966
rect 2559 1038 2621 1076
rect 3521 1436 3535 1470
rect 3569 1436 3583 1470
rect 4483 1470 4545 1505
rect 3521 1398 3583 1436
rect 3521 1364 3535 1398
rect 3569 1364 3583 1398
rect 3521 1326 3583 1364
rect 3521 1292 3535 1326
rect 3569 1292 3583 1326
rect 3521 1254 3583 1292
rect 3521 1220 3535 1254
rect 3569 1220 3583 1254
rect 3521 1182 3583 1220
rect 3521 1148 3535 1182
rect 3569 1148 3583 1182
rect 3521 1110 3583 1148
rect 3521 1076 3535 1110
rect 3569 1076 3583 1110
rect 2559 1004 2573 1038
rect 2607 1004 2621 1038
rect 2559 966 2621 1004
rect 1893 930 1955 932
rect 2559 932 2573 966
rect 2607 932 2621 966
rect 3521 1038 3583 1076
rect 4483 1436 4497 1470
rect 4531 1436 4545 1470
rect 5149 1470 5211 1505
rect 4483 1398 4545 1436
rect 4483 1364 4497 1398
rect 4531 1364 4545 1398
rect 4483 1326 4545 1364
rect 4483 1292 4497 1326
rect 4531 1292 4545 1326
rect 4483 1254 4545 1292
rect 4483 1220 4497 1254
rect 4531 1220 4545 1254
rect 4483 1182 4545 1220
rect 4483 1148 4497 1182
rect 4531 1148 4545 1182
rect 4483 1110 4545 1148
rect 4483 1076 4497 1110
rect 4531 1076 4545 1110
rect 3521 1004 3535 1038
rect 3569 1004 3583 1038
rect 3521 966 3583 1004
rect 2559 930 2621 932
rect 3521 932 3535 966
rect 3569 932 3583 966
rect 4483 1038 4545 1076
rect 5149 1436 5163 1470
rect 5197 1436 5211 1470
rect 5149 1398 5211 1436
rect 5149 1364 5163 1398
rect 5197 1364 5211 1398
rect 5149 1326 5211 1364
rect 5149 1292 5163 1326
rect 5197 1292 5211 1326
rect 5149 1254 5211 1292
rect 5149 1220 5163 1254
rect 5197 1220 5211 1254
rect 5149 1182 5211 1220
rect 5149 1148 5163 1182
rect 5197 1148 5211 1182
rect 5149 1110 5211 1148
rect 5149 1076 5163 1110
rect 5197 1076 5211 1110
rect 4483 1004 4497 1038
rect 4531 1004 4545 1038
rect 4483 966 4545 1004
rect 3521 930 3583 932
rect 4483 932 4497 966
rect 4531 932 4545 966
rect 5149 1038 5211 1076
rect 5149 1004 5163 1038
rect 5197 1004 5211 1038
rect 5149 966 5211 1004
rect 4483 930 4545 932
rect 5149 932 5163 966
rect 5197 932 5211 966
rect 5149 930 5211 932
rect -31 868 5211 930
<< psubdiffcont >>
rect -17 512 17 546
rect 945 512 979 546
rect 1907 512 1941 546
rect 2573 512 2607 546
rect 3535 512 3569 546
rect 4497 512 4531 546
rect 5163 512 5197 546
rect -17 440 17 474
rect -17 368 17 402
rect 945 440 979 474
rect -17 296 17 330
rect -17 224 17 258
rect -17 152 17 186
rect -17 80 17 114
rect 945 368 979 402
rect 1907 440 1941 474
rect 945 296 979 330
rect 945 224 979 258
rect 945 152 979 186
rect 945 80 979 114
rect 1907 368 1941 402
rect 2573 440 2607 474
rect 1907 296 1941 330
rect 1907 224 1941 258
rect 1907 152 1941 186
rect 1907 80 1941 114
rect 2573 368 2607 402
rect 3535 440 3569 474
rect 2573 296 2607 330
rect 2573 224 2607 258
rect 2573 152 2607 186
rect 2573 80 2607 114
rect 3535 368 3569 402
rect 4497 440 4531 474
rect 3535 296 3569 330
rect 3535 224 3569 258
rect 3535 152 3569 186
rect 3535 80 3569 114
rect 4497 368 4531 402
rect 5163 440 5197 474
rect 4497 296 4531 330
rect 4497 224 4531 258
rect 4497 152 4531 186
rect 4497 80 4531 114
rect 5163 368 5197 402
rect 5163 296 5197 330
rect 5163 224 5197 258
rect 5163 152 5197 186
rect 5163 80 5197 114
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 343 13 377 47
rect 415 13 449 47
rect 513 13 547 47
rect 585 13 619 47
rect 657 13 691 47
rect 729 13 763 47
rect 801 13 835 47
rect 873 13 907 47
rect 1017 13 1051 47
rect 1089 13 1123 47
rect 1161 13 1195 47
rect 1233 13 1267 47
rect 1305 13 1339 47
rect 1377 13 1411 47
rect 1475 13 1509 47
rect 1547 13 1581 47
rect 1619 13 1653 47
rect 1691 13 1725 47
rect 1763 13 1797 47
rect 1835 13 1869 47
rect 1979 13 2013 47
rect 2051 13 2085 47
rect 2123 13 2157 47
rect 2195 13 2229 47
rect 2285 13 2319 47
rect 2357 13 2391 47
rect 2429 13 2463 47
rect 2501 13 2535 47
rect 2645 13 2679 47
rect 2717 13 2751 47
rect 2789 13 2823 47
rect 2861 13 2895 47
rect 2933 13 2967 47
rect 3005 13 3039 47
rect 3103 13 3137 47
rect 3175 13 3209 47
rect 3247 13 3281 47
rect 3319 13 3353 47
rect 3391 13 3425 47
rect 3463 13 3497 47
rect 3607 13 3641 47
rect 3679 13 3713 47
rect 3751 13 3785 47
rect 3823 13 3857 47
rect 3895 13 3929 47
rect 3967 13 4001 47
rect 4065 13 4099 47
rect 4137 13 4171 47
rect 4209 13 4243 47
rect 4281 13 4315 47
rect 4353 13 4387 47
rect 4425 13 4459 47
rect 4569 13 4603 47
rect 4641 13 4675 47
rect 4713 13 4747 47
rect 4785 13 4819 47
rect 4875 13 4909 47
rect 4947 13 4981 47
rect 5019 13 5053 47
rect 5091 13 5125 47
<< nsubdiffcont >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 343 1505 377 1539
rect 415 1505 449 1539
rect 513 1505 547 1539
rect 585 1505 619 1539
rect 657 1505 691 1539
rect 729 1505 763 1539
rect 801 1505 835 1539
rect 873 1505 907 1539
rect 1017 1505 1051 1539
rect 1089 1505 1123 1539
rect 1161 1505 1195 1539
rect 1233 1505 1267 1539
rect 1305 1505 1339 1539
rect 1377 1505 1411 1539
rect 1475 1505 1509 1539
rect 1547 1505 1581 1539
rect 1619 1505 1653 1539
rect 1691 1505 1725 1539
rect 1763 1505 1797 1539
rect 1835 1505 1869 1539
rect 1979 1505 2013 1539
rect 2051 1505 2085 1539
rect 2123 1505 2157 1539
rect 2195 1505 2229 1539
rect 2285 1505 2319 1539
rect 2357 1505 2391 1539
rect 2429 1505 2463 1539
rect 2501 1505 2535 1539
rect 2645 1505 2679 1539
rect 2717 1505 2751 1539
rect 2789 1505 2823 1539
rect 2861 1505 2895 1539
rect 2933 1505 2967 1539
rect 3005 1505 3039 1539
rect 3103 1505 3137 1539
rect 3175 1505 3209 1539
rect 3247 1505 3281 1539
rect 3319 1505 3353 1539
rect 3391 1505 3425 1539
rect 3463 1505 3497 1539
rect 3607 1505 3641 1539
rect 3679 1505 3713 1539
rect 3751 1505 3785 1539
rect 3823 1505 3857 1539
rect 3895 1505 3929 1539
rect 3967 1505 4001 1539
rect 4065 1505 4099 1539
rect 4137 1505 4171 1539
rect 4209 1505 4243 1539
rect 4281 1505 4315 1539
rect 4353 1505 4387 1539
rect 4425 1505 4459 1539
rect 4569 1505 4603 1539
rect 4641 1505 4675 1539
rect 4713 1505 4747 1539
rect 4785 1505 4819 1539
rect 4875 1505 4909 1539
rect 4947 1505 4981 1539
rect 5019 1505 5053 1539
rect 5091 1505 5125 1539
rect -17 1436 17 1470
rect -17 1364 17 1398
rect -17 1292 17 1326
rect -17 1220 17 1254
rect -17 1148 17 1182
rect -17 1076 17 1110
rect 945 1436 979 1470
rect 945 1364 979 1398
rect 945 1292 979 1326
rect 945 1220 979 1254
rect 945 1148 979 1182
rect 945 1076 979 1110
rect -17 1004 17 1038
rect -17 932 17 966
rect 1907 1436 1941 1470
rect 1907 1364 1941 1398
rect 1907 1292 1941 1326
rect 1907 1220 1941 1254
rect 1907 1148 1941 1182
rect 1907 1076 1941 1110
rect 945 1004 979 1038
rect 945 932 979 966
rect 2573 1436 2607 1470
rect 2573 1364 2607 1398
rect 2573 1292 2607 1326
rect 2573 1220 2607 1254
rect 2573 1148 2607 1182
rect 2573 1076 2607 1110
rect 1907 1004 1941 1038
rect 1907 932 1941 966
rect 3535 1436 3569 1470
rect 3535 1364 3569 1398
rect 3535 1292 3569 1326
rect 3535 1220 3569 1254
rect 3535 1148 3569 1182
rect 3535 1076 3569 1110
rect 2573 1004 2607 1038
rect 2573 932 2607 966
rect 4497 1436 4531 1470
rect 4497 1364 4531 1398
rect 4497 1292 4531 1326
rect 4497 1220 4531 1254
rect 4497 1148 4531 1182
rect 4497 1076 4531 1110
rect 3535 1004 3569 1038
rect 3535 932 3569 966
rect 5163 1436 5197 1470
rect 5163 1364 5197 1398
rect 5163 1292 5197 1326
rect 5163 1220 5197 1254
rect 5163 1148 5197 1182
rect 5163 1076 5197 1110
rect 4497 1004 4531 1038
rect 4497 932 4531 966
rect 5163 1004 5197 1038
rect 5163 932 5197 966
<< poly >>
rect 247 1450 277 1476
rect 335 1450 365 1476
rect 423 1450 453 1476
rect 511 1450 541 1476
rect 599 1450 629 1476
rect 687 1450 717 1476
rect 1209 1450 1239 1476
rect 1297 1450 1327 1476
rect 1385 1450 1415 1476
rect 1473 1450 1503 1476
rect 1561 1450 1591 1476
rect 1649 1450 1679 1476
rect 247 1019 277 1050
rect 335 1019 365 1050
rect 423 1019 453 1050
rect 511 1019 541 1050
rect 195 1003 365 1019
rect 195 969 205 1003
rect 239 989 365 1003
rect 417 1003 541 1019
rect 239 969 249 989
rect 195 953 249 969
rect 417 969 427 1003
rect 461 989 541 1003
rect 599 1019 629 1050
rect 687 1019 717 1050
rect 599 1003 717 1019
rect 599 989 649 1003
rect 461 969 471 989
rect 417 953 471 969
rect 639 969 649 989
rect 683 989 717 1003
rect 2111 1450 2141 1476
rect 2199 1450 2229 1476
rect 2287 1450 2317 1476
rect 2375 1450 2405 1476
rect 1209 1019 1239 1050
rect 1297 1019 1327 1050
rect 1385 1019 1415 1050
rect 1473 1019 1503 1050
rect 683 969 693 989
rect 639 953 693 969
rect 1157 1003 1327 1019
rect 1157 969 1167 1003
rect 1201 989 1327 1003
rect 1379 1003 1503 1019
rect 1201 969 1211 989
rect 1157 953 1211 969
rect 1379 969 1389 1003
rect 1423 989 1503 1003
rect 1561 1019 1591 1050
rect 1649 1019 1679 1050
rect 1561 1003 1679 1019
rect 1561 989 1611 1003
rect 1423 969 1433 989
rect 1379 953 1433 969
rect 1601 969 1611 989
rect 1645 989 1679 1003
rect 2837 1450 2867 1476
rect 2925 1450 2955 1476
rect 3013 1450 3043 1476
rect 3101 1450 3131 1476
rect 3189 1450 3219 1476
rect 3277 1450 3307 1476
rect 1645 969 1655 989
rect 1601 953 1655 969
rect 2111 1019 2141 1050
rect 2199 1019 2229 1050
rect 2287 1019 2317 1050
rect 2375 1019 2405 1050
rect 2111 1003 2229 1019
rect 2111 989 2129 1003
rect 2119 969 2129 989
rect 2163 989 2229 1003
rect 2273 1003 2405 1019
rect 2163 969 2173 989
rect 2119 953 2173 969
rect 2273 969 2283 1003
rect 2317 989 2405 1003
rect 3799 1450 3829 1476
rect 3887 1450 3917 1476
rect 3975 1450 4005 1476
rect 4063 1450 4093 1476
rect 4151 1450 4181 1476
rect 4239 1450 4269 1476
rect 2837 1019 2867 1050
rect 2925 1019 2955 1050
rect 3013 1019 3043 1050
rect 3101 1019 3131 1050
rect 2317 969 2327 989
rect 2273 953 2327 969
rect 2785 1003 2955 1019
rect 2785 969 2795 1003
rect 2829 989 2955 1003
rect 3007 1003 3131 1019
rect 2829 969 2839 989
rect 2785 953 2839 969
rect 3007 969 3017 1003
rect 3051 989 3131 1003
rect 3189 1019 3219 1050
rect 3277 1019 3307 1050
rect 3189 1003 3307 1019
rect 3189 989 3239 1003
rect 3051 969 3061 989
rect 3007 953 3061 969
rect 3229 969 3239 989
rect 3273 989 3307 1003
rect 4701 1450 4731 1476
rect 4789 1450 4819 1476
rect 4877 1450 4907 1476
rect 4965 1450 4995 1476
rect 3799 1019 3829 1050
rect 3887 1019 3917 1050
rect 3975 1019 4005 1050
rect 4063 1019 4093 1050
rect 3273 969 3283 989
rect 3229 953 3283 969
rect 3747 1003 3917 1019
rect 3747 969 3757 1003
rect 3791 989 3917 1003
rect 3969 1003 4093 1019
rect 3791 969 3801 989
rect 3747 953 3801 969
rect 3969 969 3979 1003
rect 4013 989 4093 1003
rect 4151 1019 4181 1050
rect 4239 1019 4269 1050
rect 4151 1003 4269 1019
rect 4151 989 4201 1003
rect 4013 969 4023 989
rect 3969 953 4023 969
rect 4191 969 4201 989
rect 4235 989 4269 1003
rect 4235 969 4245 989
rect 4191 953 4245 969
rect 4701 1019 4731 1050
rect 4789 1019 4819 1050
rect 4877 1019 4907 1050
rect 4965 1019 4995 1050
rect 4701 1003 4819 1019
rect 4701 989 4719 1003
rect 4709 969 4719 989
rect 4753 989 4819 1003
rect 4863 1003 4995 1019
rect 4753 969 4763 989
rect 4709 953 4763 969
rect 4863 969 4873 1003
rect 4907 989 4995 1003
rect 4907 969 4917 989
rect 4863 953 4917 969
rect 195 461 249 477
rect 195 441 205 461
rect 147 427 205 441
rect 239 427 249 461
rect 147 411 249 427
rect 417 461 471 477
rect 417 427 427 461
rect 461 441 471 461
rect 639 461 693 477
rect 461 427 477 441
rect 417 411 477 427
rect 639 427 649 461
rect 683 427 693 461
rect 639 411 693 427
rect 1157 461 1211 477
rect 1157 441 1167 461
rect 147 379 177 411
rect 447 379 477 411
rect 649 379 679 411
rect 1109 427 1167 441
rect 1201 427 1211 461
rect 1109 411 1211 427
rect 1379 461 1433 477
rect 1379 427 1389 461
rect 1423 441 1433 461
rect 1601 461 1655 477
rect 1423 427 1439 441
rect 1379 411 1439 427
rect 1601 427 1611 461
rect 1645 427 1655 461
rect 1601 411 1655 427
rect 2119 461 2173 477
rect 2119 441 2129 461
rect 1109 379 1139 411
rect 1409 379 1439 411
rect 1611 379 1641 411
rect 2092 427 2129 441
rect 2163 427 2173 461
rect 2092 411 2173 427
rect 2267 461 2321 477
rect 2267 427 2277 461
rect 2311 427 2321 461
rect 2267 411 2321 427
rect 2785 461 2839 477
rect 2785 441 2795 461
rect 2092 377 2122 411
rect 2286 377 2316 411
rect 2737 427 2795 441
rect 2829 427 2839 461
rect 2737 411 2839 427
rect 3007 461 3061 477
rect 3007 427 3017 461
rect 3051 441 3061 461
rect 3229 461 3283 477
rect 3051 427 3067 441
rect 3007 411 3067 427
rect 3229 427 3239 461
rect 3273 427 3283 461
rect 3229 411 3283 427
rect 3747 461 3801 477
rect 3747 441 3757 461
rect 2737 379 2767 411
rect 3037 379 3067 411
rect 3239 379 3269 411
rect 3699 427 3757 441
rect 3791 427 3801 461
rect 3699 411 3801 427
rect 3969 461 4023 477
rect 3969 427 3979 461
rect 4013 441 4023 461
rect 4191 461 4245 477
rect 4013 427 4029 441
rect 3969 411 4029 427
rect 4191 427 4201 461
rect 4235 427 4245 461
rect 4191 411 4245 427
rect 4709 461 4763 477
rect 4709 441 4719 461
rect 3699 379 3729 411
rect 3999 379 4029 411
rect 4201 379 4231 411
rect 4682 427 4719 441
rect 4753 427 4763 461
rect 4682 411 4763 427
rect 4857 461 4911 477
rect 4857 427 4867 461
rect 4901 427 4911 461
rect 4857 411 4911 427
rect 4682 377 4712 411
rect 4876 377 4906 411
<< polycont >>
rect 205 969 239 1003
rect 427 969 461 1003
rect 649 969 683 1003
rect 1167 969 1201 1003
rect 1389 969 1423 1003
rect 1611 969 1645 1003
rect 2129 969 2163 1003
rect 2283 969 2317 1003
rect 2795 969 2829 1003
rect 3017 969 3051 1003
rect 3239 969 3273 1003
rect 3757 969 3791 1003
rect 3979 969 4013 1003
rect 4201 969 4235 1003
rect 4719 969 4753 1003
rect 4873 969 4907 1003
rect 205 427 239 461
rect 427 427 461 461
rect 649 427 683 461
rect 1167 427 1201 461
rect 1389 427 1423 461
rect 1611 427 1645 461
rect 2129 427 2163 461
rect 2277 427 2311 461
rect 2795 427 2829 461
rect 3017 427 3051 461
rect 3239 427 3273 461
rect 3757 427 3791 461
rect 3979 427 4013 461
rect 4201 427 4235 461
rect 4719 427 4753 461
rect 4867 427 4901 461
<< locali >>
rect -31 1539 5211 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 343 1539
rect 377 1505 415 1539
rect 449 1505 513 1539
rect 547 1505 585 1539
rect 619 1505 657 1539
rect 691 1505 729 1539
rect 763 1505 801 1539
rect 835 1505 873 1539
rect 907 1505 1017 1539
rect 1051 1505 1089 1539
rect 1123 1505 1161 1539
rect 1195 1505 1233 1539
rect 1267 1505 1305 1539
rect 1339 1505 1377 1539
rect 1411 1505 1475 1539
rect 1509 1505 1547 1539
rect 1581 1505 1619 1539
rect 1653 1505 1691 1539
rect 1725 1505 1763 1539
rect 1797 1505 1835 1539
rect 1869 1505 1979 1539
rect 2013 1505 2051 1539
rect 2085 1505 2123 1539
rect 2157 1505 2195 1539
rect 2229 1505 2285 1539
rect 2319 1505 2357 1539
rect 2391 1505 2429 1539
rect 2463 1505 2501 1539
rect 2535 1505 2645 1539
rect 2679 1505 2717 1539
rect 2751 1505 2789 1539
rect 2823 1505 2861 1539
rect 2895 1505 2933 1539
rect 2967 1505 3005 1539
rect 3039 1505 3103 1539
rect 3137 1505 3175 1539
rect 3209 1505 3247 1539
rect 3281 1505 3319 1539
rect 3353 1505 3391 1539
rect 3425 1505 3463 1539
rect 3497 1505 3607 1539
rect 3641 1505 3679 1539
rect 3713 1505 3751 1539
rect 3785 1505 3823 1539
rect 3857 1505 3895 1539
rect 3929 1505 3967 1539
rect 4001 1505 4065 1539
rect 4099 1505 4137 1539
rect 4171 1505 4209 1539
rect 4243 1505 4281 1539
rect 4315 1505 4353 1539
rect 4387 1505 4425 1539
rect 4459 1505 4569 1539
rect 4603 1505 4641 1539
rect 4675 1505 4713 1539
rect 4747 1505 4785 1539
rect 4819 1505 4875 1539
rect 4909 1505 4947 1539
rect 4981 1505 5019 1539
rect 5053 1505 5091 1539
rect 5125 1505 5211 1539
rect -31 1492 5211 1505
rect -31 1470 31 1492
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect 201 1412 235 1492
rect 201 1344 235 1378
rect 201 1276 235 1310
rect 201 1208 235 1242
rect 201 1139 235 1174
rect 201 1089 235 1105
rect 289 1412 323 1450
rect 289 1344 323 1378
rect 289 1276 323 1310
rect 289 1208 323 1242
rect 289 1139 323 1174
rect 377 1412 411 1492
rect 377 1344 411 1378
rect 377 1276 411 1310
rect 377 1208 411 1242
rect 377 1157 411 1174
rect 465 1412 499 1450
rect 465 1344 499 1378
rect 465 1276 499 1310
rect 465 1208 499 1242
rect 289 1094 323 1105
rect 465 1139 499 1174
rect 553 1412 587 1492
rect 553 1344 587 1378
rect 553 1276 587 1310
rect 553 1208 587 1242
rect 553 1157 587 1174
rect 641 1412 675 1450
rect 641 1344 675 1378
rect 641 1276 675 1310
rect 641 1208 675 1242
rect 465 1094 499 1105
rect 641 1139 675 1174
rect 729 1412 763 1492
rect 729 1344 763 1378
rect 729 1276 763 1310
rect 729 1208 763 1242
rect 729 1157 763 1174
rect 931 1470 993 1492
rect 931 1436 945 1470
rect 979 1436 993 1470
rect 931 1398 993 1436
rect 931 1364 945 1398
rect 979 1364 993 1398
rect 931 1326 993 1364
rect 931 1292 945 1326
rect 979 1292 993 1326
rect 931 1254 993 1292
rect 931 1220 945 1254
rect 979 1220 993 1254
rect 931 1182 993 1220
rect 641 1094 675 1105
rect 931 1148 945 1182
rect 979 1148 993 1182
rect 931 1110 993 1148
rect -31 1038 31 1076
rect 289 1060 831 1094
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect -31 868 31 932
rect 205 1003 239 1019
rect 205 905 239 969
rect -31 546 31 572
rect -31 512 -17 546
rect 17 512 31 546
rect -31 474 31 512
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect 205 461 239 871
rect 205 411 239 427
rect 427 1003 461 1019
rect 427 461 461 945
rect 427 411 461 427
rect 649 1003 683 1019
rect 649 757 683 969
rect 649 461 683 723
rect 649 411 683 427
rect 797 831 831 1060
rect 931 1076 945 1110
rect 979 1076 993 1110
rect 1163 1412 1197 1492
rect 1163 1344 1197 1378
rect 1163 1276 1197 1310
rect 1163 1208 1197 1242
rect 1163 1139 1197 1174
rect 1163 1089 1197 1105
rect 1251 1412 1285 1450
rect 1251 1344 1285 1378
rect 1251 1276 1285 1310
rect 1251 1208 1285 1242
rect 1251 1139 1285 1174
rect 1339 1412 1373 1492
rect 1339 1344 1373 1378
rect 1339 1276 1373 1310
rect 1339 1208 1373 1242
rect 1339 1157 1373 1174
rect 1427 1412 1461 1450
rect 1427 1344 1461 1378
rect 1427 1276 1461 1310
rect 1427 1208 1461 1242
rect 1251 1094 1285 1105
rect 1427 1139 1461 1174
rect 1515 1412 1549 1492
rect 1515 1344 1549 1378
rect 1515 1276 1549 1310
rect 1515 1208 1549 1242
rect 1515 1157 1549 1174
rect 1603 1412 1637 1450
rect 1603 1344 1637 1378
rect 1603 1276 1637 1310
rect 1603 1208 1637 1242
rect 1427 1094 1461 1105
rect 1603 1139 1637 1174
rect 1691 1412 1725 1492
rect 1691 1344 1725 1378
rect 1691 1276 1725 1310
rect 1691 1208 1725 1242
rect 1691 1157 1725 1174
rect 1893 1470 1955 1492
rect 1893 1436 1907 1470
rect 1941 1436 1955 1470
rect 1893 1398 1955 1436
rect 1893 1364 1907 1398
rect 1941 1364 1955 1398
rect 1893 1326 1955 1364
rect 1893 1292 1907 1326
rect 1941 1292 1955 1326
rect 1893 1254 1955 1292
rect 1893 1220 1907 1254
rect 1941 1220 1955 1254
rect 1893 1182 1955 1220
rect 1603 1094 1637 1105
rect 1893 1148 1907 1182
rect 1941 1148 1955 1182
rect 1893 1110 1955 1148
rect 931 1038 993 1076
rect 1251 1060 1793 1094
rect 931 1004 945 1038
rect 979 1004 993 1038
rect 931 966 993 1004
rect 931 932 945 966
rect 979 932 993 966
rect 931 868 993 932
rect 1167 1003 1201 1019
rect -31 368 -17 402
rect 17 368 31 402
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect 101 363 135 379
rect 295 363 329 379
rect 489 363 523 379
rect 135 329 198 363
rect 232 329 295 363
rect 329 329 392 363
rect 426 329 489 363
rect 101 291 135 329
rect 101 223 135 257
rect 295 291 329 329
rect 489 313 523 329
rect 603 363 637 379
rect 797 378 831 797
rect 1167 831 1201 969
rect 603 291 637 329
rect 101 153 135 189
rect 101 103 135 119
rect 198 238 232 254
rect -31 62 31 80
rect 198 62 232 204
rect 295 223 329 257
rect 393 244 427 260
rect 603 244 637 257
rect 427 223 637 244
rect 427 210 603 223
rect 393 194 427 210
rect 295 153 329 189
rect 700 344 831 378
rect 931 546 993 572
rect 931 512 945 546
rect 979 512 993 546
rect 931 474 993 512
rect 931 440 945 474
rect 979 440 993 474
rect 931 402 993 440
rect 1167 461 1201 797
rect 1167 411 1201 427
rect 1389 1003 1423 1019
rect 1389 683 1423 969
rect 1389 461 1423 649
rect 1389 411 1423 427
rect 1611 1003 1645 1019
rect 1611 535 1645 969
rect 1611 461 1645 501
rect 1611 411 1645 427
rect 1759 757 1793 1060
rect 1893 1076 1907 1110
rect 1941 1076 1955 1110
rect 1893 1038 1955 1076
rect 2065 1412 2099 1492
rect 2065 1344 2099 1378
rect 2065 1276 2099 1310
rect 2065 1208 2099 1242
rect 2065 1139 2099 1174
rect 2065 1073 2099 1105
rect 2153 1412 2187 1450
rect 2153 1344 2187 1378
rect 2153 1276 2187 1310
rect 2153 1208 2187 1242
rect 2153 1139 2187 1174
rect 2241 1412 2275 1492
rect 2241 1344 2275 1378
rect 2241 1276 2275 1310
rect 2241 1208 2275 1242
rect 2241 1157 2275 1174
rect 2329 1412 2363 1450
rect 2329 1344 2363 1378
rect 2329 1276 2363 1310
rect 2329 1208 2363 1242
rect 2153 1103 2187 1105
rect 2329 1139 2363 1174
rect 2417 1412 2451 1492
rect 2417 1344 2451 1378
rect 2417 1276 2451 1310
rect 2417 1208 2451 1242
rect 2417 1157 2451 1174
rect 2559 1470 2621 1492
rect 2559 1436 2573 1470
rect 2607 1436 2621 1470
rect 2559 1398 2621 1436
rect 2559 1364 2573 1398
rect 2607 1364 2621 1398
rect 2559 1326 2621 1364
rect 2559 1292 2573 1326
rect 2607 1292 2621 1326
rect 2559 1254 2621 1292
rect 2559 1220 2573 1254
rect 2607 1220 2621 1254
rect 2559 1182 2621 1220
rect 2329 1103 2363 1105
rect 2559 1148 2573 1182
rect 2607 1148 2621 1182
rect 2559 1110 2621 1148
rect 2153 1069 2459 1103
rect 1893 1004 1907 1038
rect 1941 1004 1955 1038
rect 1893 966 1955 1004
rect 1893 932 1907 966
rect 1941 932 1955 966
rect 1893 868 1955 932
rect 2129 1003 2163 1019
rect 2283 1003 2317 1019
rect 931 368 945 402
rect 979 368 993 402
rect 700 247 734 344
rect 931 330 993 368
rect 700 197 734 213
rect 797 291 831 307
rect 797 223 831 257
rect 489 153 523 169
rect 329 119 392 153
rect 426 119 489 153
rect 295 103 329 119
rect 489 103 523 119
rect 603 153 637 189
rect 797 153 831 189
rect 637 119 700 153
rect 734 119 797 153
rect 603 103 637 119
rect 797 103 831 119
rect 931 296 945 330
rect 979 296 993 330
rect 931 258 993 296
rect 931 224 945 258
rect 979 224 993 258
rect 931 186 993 224
rect 931 152 945 186
rect 979 152 993 186
rect 931 114 993 152
rect 931 80 945 114
rect 979 80 993 114
rect 1063 363 1097 379
rect 1257 363 1291 379
rect 1451 363 1485 379
rect 1097 329 1160 363
rect 1194 329 1257 363
rect 1291 329 1354 363
rect 1388 329 1451 363
rect 1063 291 1097 329
rect 1063 223 1097 257
rect 1257 291 1291 329
rect 1451 313 1485 329
rect 1565 363 1599 379
rect 1759 378 1793 723
rect 2129 757 2163 969
rect 1565 291 1599 329
rect 1063 153 1097 189
rect 1063 103 1097 119
rect 1160 238 1194 254
rect 931 62 993 80
rect 1160 62 1194 204
rect 1257 223 1291 257
rect 1355 244 1389 260
rect 1565 244 1599 257
rect 1389 223 1599 244
rect 1389 210 1565 223
rect 1355 194 1389 210
rect 1257 153 1291 189
rect 1662 344 1793 378
rect 1893 546 1955 572
rect 1893 512 1907 546
rect 1941 512 1955 546
rect 1893 474 1955 512
rect 1893 440 1907 474
rect 1941 440 1955 474
rect 1893 402 1955 440
rect 2129 461 2163 723
rect 2129 411 2163 427
rect 2277 969 2283 988
rect 2277 953 2317 969
rect 2277 905 2311 953
rect 2277 461 2311 871
rect 2277 411 2311 427
rect 2425 757 2459 1069
rect 2559 1076 2573 1110
rect 2607 1076 2621 1110
rect 2791 1412 2825 1492
rect 2791 1344 2825 1378
rect 2791 1276 2825 1310
rect 2791 1208 2825 1242
rect 2791 1139 2825 1174
rect 2791 1089 2825 1105
rect 2879 1412 2913 1450
rect 2879 1344 2913 1378
rect 2879 1276 2913 1310
rect 2879 1208 2913 1242
rect 2879 1139 2913 1174
rect 2967 1412 3001 1492
rect 2967 1344 3001 1378
rect 2967 1276 3001 1310
rect 2967 1208 3001 1242
rect 2967 1157 3001 1174
rect 3055 1412 3089 1450
rect 3055 1344 3089 1378
rect 3055 1276 3089 1310
rect 3055 1208 3089 1242
rect 2879 1094 2913 1105
rect 3055 1139 3089 1174
rect 3143 1412 3177 1492
rect 3143 1344 3177 1378
rect 3143 1276 3177 1310
rect 3143 1208 3177 1242
rect 3143 1157 3177 1174
rect 3231 1412 3265 1450
rect 3231 1344 3265 1378
rect 3231 1276 3265 1310
rect 3231 1208 3265 1242
rect 3055 1094 3089 1105
rect 3231 1139 3265 1174
rect 3319 1412 3353 1492
rect 3319 1344 3353 1378
rect 3319 1276 3353 1310
rect 3319 1208 3353 1242
rect 3319 1157 3353 1174
rect 3521 1470 3583 1492
rect 3521 1436 3535 1470
rect 3569 1436 3583 1470
rect 3521 1398 3583 1436
rect 3521 1364 3535 1398
rect 3569 1364 3583 1398
rect 3521 1326 3583 1364
rect 3521 1292 3535 1326
rect 3569 1292 3583 1326
rect 3521 1254 3583 1292
rect 3521 1220 3535 1254
rect 3569 1220 3583 1254
rect 3521 1182 3583 1220
rect 3231 1094 3265 1105
rect 3521 1148 3535 1182
rect 3569 1148 3583 1182
rect 3521 1110 3583 1148
rect 2559 1038 2621 1076
rect 2879 1060 3421 1094
rect 2559 1004 2573 1038
rect 2607 1004 2621 1038
rect 2559 966 2621 1004
rect 2559 932 2573 966
rect 2607 932 2621 966
rect 2559 868 2621 932
rect 2795 1003 2829 1019
rect 1893 368 1907 402
rect 1941 368 1955 402
rect 1662 247 1696 344
rect 1893 330 1955 368
rect 1662 197 1696 213
rect 1759 291 1793 307
rect 1759 223 1793 257
rect 1451 153 1485 169
rect 1291 119 1354 153
rect 1388 119 1451 153
rect 1257 103 1291 119
rect 1451 103 1485 119
rect 1565 153 1599 189
rect 1759 153 1793 189
rect 1599 119 1662 153
rect 1696 119 1759 153
rect 1565 103 1599 119
rect 1759 103 1793 119
rect 1893 296 1907 330
rect 1941 296 1955 330
rect 1893 258 1955 296
rect 1893 224 1907 258
rect 1941 224 1955 258
rect 1893 186 1955 224
rect 1893 152 1907 186
rect 1941 152 1955 186
rect 1893 114 1955 152
rect 1893 80 1907 114
rect 1941 80 1955 114
rect 2046 361 2080 377
rect 2240 361 2274 377
rect 2425 376 2459 723
rect 2795 757 2829 969
rect 2080 327 2143 361
rect 2177 327 2240 361
rect 2046 289 2080 327
rect 2046 221 2080 255
rect 2240 289 2274 327
rect 2046 151 2080 187
rect 2046 101 2080 117
rect 2143 236 2177 252
rect 1893 62 1955 80
rect 2143 62 2177 202
rect 2240 221 2274 255
rect 2337 342 2459 376
rect 2559 546 2621 572
rect 2559 512 2573 546
rect 2607 512 2621 546
rect 2559 474 2621 512
rect 2559 440 2573 474
rect 2607 440 2621 474
rect 2559 402 2621 440
rect 2795 461 2829 723
rect 2795 411 2829 427
rect 3017 1003 3051 1019
rect 3017 461 3051 945
rect 3017 411 3051 427
rect 3239 1003 3273 1019
rect 3239 535 3273 969
rect 3239 461 3273 501
rect 3239 411 3273 427
rect 3387 905 3421 1060
rect 2559 368 2573 402
rect 2607 368 2621 402
rect 2337 245 2371 342
rect 2559 330 2621 368
rect 2337 195 2371 211
rect 2434 289 2468 305
rect 2434 221 2468 255
rect 2240 151 2274 187
rect 2434 151 2468 187
rect 2274 117 2337 151
rect 2371 117 2434 151
rect 2240 101 2274 117
rect 2434 101 2468 117
rect 2559 296 2573 330
rect 2607 296 2621 330
rect 2559 258 2621 296
rect 2559 224 2573 258
rect 2607 224 2621 258
rect 2559 186 2621 224
rect 2559 152 2573 186
rect 2607 152 2621 186
rect 2559 114 2621 152
rect 2559 80 2573 114
rect 2607 80 2621 114
rect 2691 363 2725 379
rect 2885 363 2919 379
rect 3079 363 3113 379
rect 2725 329 2788 363
rect 2822 329 2885 363
rect 2919 329 2982 363
rect 3016 329 3079 363
rect 2691 291 2725 329
rect 2691 223 2725 257
rect 2885 291 2919 329
rect 3079 313 3113 329
rect 3193 363 3227 379
rect 3387 378 3421 871
rect 3521 1076 3535 1110
rect 3569 1076 3583 1110
rect 3753 1412 3787 1492
rect 3753 1344 3787 1378
rect 3753 1276 3787 1310
rect 3753 1208 3787 1242
rect 3753 1139 3787 1174
rect 3753 1089 3787 1105
rect 3841 1412 3875 1450
rect 3841 1344 3875 1378
rect 3841 1276 3875 1310
rect 3841 1208 3875 1242
rect 3841 1139 3875 1174
rect 3929 1412 3963 1492
rect 3929 1344 3963 1378
rect 3929 1276 3963 1310
rect 3929 1208 3963 1242
rect 3929 1157 3963 1174
rect 4017 1412 4051 1450
rect 4017 1344 4051 1378
rect 4017 1276 4051 1310
rect 4017 1208 4051 1242
rect 3841 1094 3875 1105
rect 4017 1139 4051 1174
rect 4105 1412 4139 1492
rect 4105 1344 4139 1378
rect 4105 1276 4139 1310
rect 4105 1208 4139 1242
rect 4105 1157 4139 1174
rect 4193 1412 4227 1450
rect 4193 1344 4227 1378
rect 4193 1276 4227 1310
rect 4193 1208 4227 1242
rect 4017 1094 4051 1105
rect 4193 1139 4227 1174
rect 4281 1412 4315 1492
rect 4281 1344 4315 1378
rect 4281 1276 4315 1310
rect 4281 1208 4315 1242
rect 4281 1157 4315 1174
rect 4483 1470 4545 1492
rect 4483 1436 4497 1470
rect 4531 1436 4545 1470
rect 4483 1398 4545 1436
rect 4483 1364 4497 1398
rect 4531 1364 4545 1398
rect 4483 1326 4545 1364
rect 4483 1292 4497 1326
rect 4531 1292 4545 1326
rect 4483 1254 4545 1292
rect 4483 1220 4497 1254
rect 4531 1220 4545 1254
rect 4483 1182 4545 1220
rect 4193 1094 4227 1105
rect 4483 1148 4497 1182
rect 4531 1148 4545 1182
rect 4483 1110 4545 1148
rect 3521 1038 3583 1076
rect 3841 1060 4383 1094
rect 3521 1004 3535 1038
rect 3569 1004 3583 1038
rect 3521 966 3583 1004
rect 3521 932 3535 966
rect 3569 932 3583 966
rect 3521 868 3583 932
rect 3757 1003 3791 1019
rect 3757 831 3791 969
rect 3193 291 3227 329
rect 2691 153 2725 189
rect 2691 103 2725 119
rect 2788 238 2822 254
rect 2559 62 2621 80
rect 2788 62 2822 204
rect 2885 223 2919 257
rect 2983 244 3017 260
rect 3193 244 3227 257
rect 3017 223 3227 244
rect 3017 210 3193 223
rect 2983 194 3017 210
rect 2885 153 2919 189
rect 3290 344 3421 378
rect 3521 546 3583 572
rect 3521 512 3535 546
rect 3569 512 3583 546
rect 3521 474 3583 512
rect 3521 440 3535 474
rect 3569 440 3583 474
rect 3521 402 3583 440
rect 3757 461 3791 797
rect 3757 411 3791 427
rect 3979 1003 4013 1019
rect 3979 535 4013 969
rect 3979 461 4013 501
rect 3979 411 4013 427
rect 4201 1003 4235 1019
rect 4201 831 4235 969
rect 4201 461 4235 797
rect 4201 411 4235 427
rect 4349 757 4383 1060
rect 4483 1076 4497 1110
rect 4531 1076 4545 1110
rect 4483 1038 4545 1076
rect 4655 1412 4689 1492
rect 4655 1344 4689 1378
rect 4655 1276 4689 1310
rect 4655 1208 4689 1242
rect 4655 1139 4689 1174
rect 4655 1073 4689 1105
rect 4743 1412 4777 1450
rect 4743 1344 4777 1378
rect 4743 1276 4777 1310
rect 4743 1208 4777 1242
rect 4743 1139 4777 1174
rect 4831 1412 4865 1492
rect 4831 1344 4865 1378
rect 4831 1276 4865 1310
rect 4831 1208 4865 1242
rect 4831 1157 4865 1174
rect 4919 1412 4953 1450
rect 4919 1344 4953 1378
rect 4919 1276 4953 1310
rect 4919 1208 4953 1242
rect 4743 1103 4777 1105
rect 4919 1139 4953 1174
rect 5007 1412 5041 1492
rect 5007 1344 5041 1378
rect 5007 1276 5041 1310
rect 5007 1208 5041 1242
rect 5007 1157 5041 1174
rect 5149 1470 5211 1492
rect 5149 1436 5163 1470
rect 5197 1436 5211 1470
rect 5149 1398 5211 1436
rect 5149 1364 5163 1398
rect 5197 1364 5211 1398
rect 5149 1326 5211 1364
rect 5149 1292 5163 1326
rect 5197 1292 5211 1326
rect 5149 1254 5211 1292
rect 5149 1220 5163 1254
rect 5197 1220 5211 1254
rect 5149 1182 5211 1220
rect 4919 1103 4953 1105
rect 5149 1148 5163 1182
rect 5197 1148 5211 1182
rect 5149 1110 5211 1148
rect 4743 1069 5049 1103
rect 4483 1004 4497 1038
rect 4531 1004 4545 1038
rect 4483 966 4545 1004
rect 4483 932 4497 966
rect 4531 932 4545 966
rect 4483 868 4545 932
rect 4719 1003 4753 1019
rect 4873 1003 4907 1019
rect 3521 368 3535 402
rect 3569 368 3583 402
rect 3290 247 3324 344
rect 3521 330 3583 368
rect 3290 197 3324 213
rect 3387 291 3421 307
rect 3387 223 3421 257
rect 3079 153 3113 169
rect 2919 119 2982 153
rect 3016 119 3079 153
rect 2885 103 2919 119
rect 3079 103 3113 119
rect 3193 153 3227 189
rect 3387 153 3421 189
rect 3227 119 3290 153
rect 3324 119 3387 153
rect 3193 103 3227 119
rect 3387 103 3421 119
rect 3521 296 3535 330
rect 3569 296 3583 330
rect 3521 258 3583 296
rect 3521 224 3535 258
rect 3569 224 3583 258
rect 3521 186 3583 224
rect 3521 152 3535 186
rect 3569 152 3583 186
rect 3521 114 3583 152
rect 3521 80 3535 114
rect 3569 80 3583 114
rect 3653 363 3687 379
rect 3847 363 3881 379
rect 4041 363 4075 379
rect 3687 329 3750 363
rect 3784 329 3847 363
rect 3881 329 3944 363
rect 3978 329 4041 363
rect 3653 291 3687 329
rect 3653 223 3687 257
rect 3847 291 3881 329
rect 4041 313 4075 329
rect 4155 363 4189 379
rect 4349 378 4383 723
rect 4719 757 4753 969
rect 4155 291 4189 329
rect 3653 153 3687 189
rect 3653 103 3687 119
rect 3750 238 3784 254
rect 3521 62 3583 80
rect 3750 62 3784 204
rect 3847 223 3881 257
rect 3945 244 3979 260
rect 4155 244 4189 257
rect 3979 223 4189 244
rect 3979 210 4155 223
rect 3945 194 3979 210
rect 3847 153 3881 189
rect 4252 344 4383 378
rect 4483 546 4545 572
rect 4483 512 4497 546
rect 4531 512 4545 546
rect 4483 474 4545 512
rect 4483 440 4497 474
rect 4531 440 4545 474
rect 4483 402 4545 440
rect 4719 461 4753 723
rect 4719 411 4753 427
rect 4867 969 4873 988
rect 4867 953 4907 969
rect 4867 905 4901 953
rect 4867 461 4901 871
rect 4867 411 4901 427
rect 5015 831 5049 1069
rect 5149 1076 5163 1110
rect 5197 1076 5211 1110
rect 5149 1038 5211 1076
rect 5149 1004 5163 1038
rect 5197 1004 5211 1038
rect 5149 966 5211 1004
rect 5149 932 5163 966
rect 5197 932 5211 966
rect 5149 868 5211 932
rect 4483 368 4497 402
rect 4531 368 4545 402
rect 4252 247 4286 344
rect 4483 330 4545 368
rect 4252 197 4286 213
rect 4349 291 4383 307
rect 4349 223 4383 257
rect 4041 153 4075 169
rect 3881 119 3944 153
rect 3978 119 4041 153
rect 3847 103 3881 119
rect 4041 103 4075 119
rect 4155 153 4189 189
rect 4349 153 4383 189
rect 4189 119 4252 153
rect 4286 119 4349 153
rect 4155 103 4189 119
rect 4349 103 4383 119
rect 4483 296 4497 330
rect 4531 296 4545 330
rect 4483 258 4545 296
rect 4483 224 4497 258
rect 4531 224 4545 258
rect 4483 186 4545 224
rect 4483 152 4497 186
rect 4531 152 4545 186
rect 4483 114 4545 152
rect 4483 80 4497 114
rect 4531 80 4545 114
rect 4636 361 4670 377
rect 4830 361 4864 377
rect 5015 376 5049 797
rect 4670 327 4733 361
rect 4767 327 4830 361
rect 4636 289 4670 327
rect 4636 221 4670 255
rect 4830 289 4864 327
rect 4636 151 4670 187
rect 4636 101 4670 117
rect 4733 236 4767 252
rect 4483 62 4545 80
rect 4733 62 4767 202
rect 4830 221 4864 255
rect 4927 342 5049 376
rect 5149 546 5211 572
rect 5149 512 5163 546
rect 5197 512 5211 546
rect 5149 474 5211 512
rect 5149 440 5163 474
rect 5197 440 5211 474
rect 5149 402 5211 440
rect 5149 368 5163 402
rect 5197 368 5211 402
rect 4927 245 4961 342
rect 5149 330 5211 368
rect 4927 195 4961 211
rect 5024 289 5058 305
rect 5024 221 5058 255
rect 4830 151 4864 187
rect 5024 151 5058 187
rect 4864 117 4927 151
rect 4961 117 5024 151
rect 4830 101 4864 117
rect 5024 101 5058 117
rect 5149 296 5163 330
rect 5197 296 5211 330
rect 5149 258 5211 296
rect 5149 224 5163 258
rect 5197 224 5211 258
rect 5149 186 5211 224
rect 5149 152 5163 186
rect 5197 152 5211 186
rect 5149 114 5211 152
rect 5149 80 5163 114
rect 5197 80 5211 114
rect 5149 62 5211 80
rect -31 47 5211 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 343 47
rect 377 13 415 47
rect 449 13 513 47
rect 547 13 585 47
rect 619 13 657 47
rect 691 13 729 47
rect 763 13 801 47
rect 835 13 873 47
rect 907 13 1017 47
rect 1051 13 1089 47
rect 1123 13 1161 47
rect 1195 13 1233 47
rect 1267 13 1305 47
rect 1339 13 1377 47
rect 1411 13 1475 47
rect 1509 13 1547 47
rect 1581 13 1619 47
rect 1653 13 1691 47
rect 1725 13 1763 47
rect 1797 13 1835 47
rect 1869 13 1979 47
rect 2013 13 2051 47
rect 2085 13 2123 47
rect 2157 13 2195 47
rect 2229 13 2285 47
rect 2319 13 2357 47
rect 2391 13 2429 47
rect 2463 13 2501 47
rect 2535 13 2645 47
rect 2679 13 2717 47
rect 2751 13 2789 47
rect 2823 13 2861 47
rect 2895 13 2933 47
rect 2967 13 3005 47
rect 3039 13 3103 47
rect 3137 13 3175 47
rect 3209 13 3247 47
rect 3281 13 3319 47
rect 3353 13 3391 47
rect 3425 13 3463 47
rect 3497 13 3607 47
rect 3641 13 3679 47
rect 3713 13 3751 47
rect 3785 13 3823 47
rect 3857 13 3895 47
rect 3929 13 3967 47
rect 4001 13 4065 47
rect 4099 13 4137 47
rect 4171 13 4209 47
rect 4243 13 4281 47
rect 4315 13 4353 47
rect 4387 13 4425 47
rect 4459 13 4569 47
rect 4603 13 4641 47
rect 4675 13 4713 47
rect 4747 13 4785 47
rect 4819 13 4875 47
rect 4909 13 4947 47
rect 4981 13 5019 47
rect 5053 13 5091 47
rect 5125 13 5211 47
rect -31 0 5211 13
<< viali >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 343 1505 377 1539
rect 415 1505 449 1539
rect 513 1505 547 1539
rect 585 1505 619 1539
rect 657 1505 691 1539
rect 729 1505 763 1539
rect 801 1505 835 1539
rect 873 1505 907 1539
rect 1017 1505 1051 1539
rect 1089 1505 1123 1539
rect 1161 1505 1195 1539
rect 1233 1505 1267 1539
rect 1305 1505 1339 1539
rect 1377 1505 1411 1539
rect 1475 1505 1509 1539
rect 1547 1505 1581 1539
rect 1619 1505 1653 1539
rect 1691 1505 1725 1539
rect 1763 1505 1797 1539
rect 1835 1505 1869 1539
rect 1979 1505 2013 1539
rect 2051 1505 2085 1539
rect 2123 1505 2157 1539
rect 2195 1505 2229 1539
rect 2285 1505 2319 1539
rect 2357 1505 2391 1539
rect 2429 1505 2463 1539
rect 2501 1505 2535 1539
rect 2645 1505 2679 1539
rect 2717 1505 2751 1539
rect 2789 1505 2823 1539
rect 2861 1505 2895 1539
rect 2933 1505 2967 1539
rect 3005 1505 3039 1539
rect 3103 1505 3137 1539
rect 3175 1505 3209 1539
rect 3247 1505 3281 1539
rect 3319 1505 3353 1539
rect 3391 1505 3425 1539
rect 3463 1505 3497 1539
rect 3607 1505 3641 1539
rect 3679 1505 3713 1539
rect 3751 1505 3785 1539
rect 3823 1505 3857 1539
rect 3895 1505 3929 1539
rect 3967 1505 4001 1539
rect 4065 1505 4099 1539
rect 4137 1505 4171 1539
rect 4209 1505 4243 1539
rect 4281 1505 4315 1539
rect 4353 1505 4387 1539
rect 4425 1505 4459 1539
rect 4569 1505 4603 1539
rect 4641 1505 4675 1539
rect 4713 1505 4747 1539
rect 4785 1505 4819 1539
rect 4875 1505 4909 1539
rect 4947 1505 4981 1539
rect 5019 1505 5053 1539
rect 5091 1505 5125 1539
rect 205 871 239 905
rect 427 969 461 979
rect 427 945 461 969
rect 649 723 683 757
rect 797 797 831 831
rect 1167 797 1201 831
rect 1389 649 1423 683
rect 1611 501 1645 535
rect 1759 723 1793 757
rect 2129 723 2163 757
rect 2277 871 2311 905
rect 2425 723 2459 757
rect 2795 723 2829 757
rect 3017 969 3051 979
rect 3017 945 3051 969
rect 3239 501 3273 535
rect 3387 871 3421 905
rect 3757 797 3791 831
rect 3979 501 4013 535
rect 4201 797 4235 831
rect 4349 723 4383 757
rect 4719 723 4753 757
rect 4867 871 4901 905
rect 5015 797 5049 831
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 343 13 377 47
rect 415 13 449 47
rect 513 13 547 47
rect 585 13 619 47
rect 657 13 691 47
rect 729 13 763 47
rect 801 13 835 47
rect 873 13 907 47
rect 1017 13 1051 47
rect 1089 13 1123 47
rect 1161 13 1195 47
rect 1233 13 1267 47
rect 1305 13 1339 47
rect 1377 13 1411 47
rect 1475 13 1509 47
rect 1547 13 1581 47
rect 1619 13 1653 47
rect 1691 13 1725 47
rect 1763 13 1797 47
rect 1835 13 1869 47
rect 1979 13 2013 47
rect 2051 13 2085 47
rect 2123 13 2157 47
rect 2195 13 2229 47
rect 2285 13 2319 47
rect 2357 13 2391 47
rect 2429 13 2463 47
rect 2501 13 2535 47
rect 2645 13 2679 47
rect 2717 13 2751 47
rect 2789 13 2823 47
rect 2861 13 2895 47
rect 2933 13 2967 47
rect 3005 13 3039 47
rect 3103 13 3137 47
rect 3175 13 3209 47
rect 3247 13 3281 47
rect 3319 13 3353 47
rect 3391 13 3425 47
rect 3463 13 3497 47
rect 3607 13 3641 47
rect 3679 13 3713 47
rect 3751 13 3785 47
rect 3823 13 3857 47
rect 3895 13 3929 47
rect 3967 13 4001 47
rect 4065 13 4099 47
rect 4137 13 4171 47
rect 4209 13 4243 47
rect 4281 13 4315 47
rect 4353 13 4387 47
rect 4425 13 4459 47
rect 4569 13 4603 47
rect 4641 13 4675 47
rect 4713 13 4747 47
rect 4785 13 4819 47
rect 4875 13 4909 47
rect 4947 13 4981 47
rect 5019 13 5053 47
rect 5091 13 5125 47
<< metal1 >>
rect -31 1539 5211 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 343 1539
rect 377 1505 415 1539
rect 449 1505 513 1539
rect 547 1505 585 1539
rect 619 1505 657 1539
rect 691 1505 729 1539
rect 763 1505 801 1539
rect 835 1505 873 1539
rect 907 1505 1017 1539
rect 1051 1505 1089 1539
rect 1123 1505 1161 1539
rect 1195 1505 1233 1539
rect 1267 1505 1305 1539
rect 1339 1505 1377 1539
rect 1411 1505 1475 1539
rect 1509 1505 1547 1539
rect 1581 1505 1619 1539
rect 1653 1505 1691 1539
rect 1725 1505 1763 1539
rect 1797 1505 1835 1539
rect 1869 1505 1979 1539
rect 2013 1505 2051 1539
rect 2085 1505 2123 1539
rect 2157 1505 2195 1539
rect 2229 1505 2285 1539
rect 2319 1505 2357 1539
rect 2391 1505 2429 1539
rect 2463 1505 2501 1539
rect 2535 1505 2645 1539
rect 2679 1505 2717 1539
rect 2751 1505 2789 1539
rect 2823 1505 2861 1539
rect 2895 1505 2933 1539
rect 2967 1505 3005 1539
rect 3039 1505 3103 1539
rect 3137 1505 3175 1539
rect 3209 1505 3247 1539
rect 3281 1505 3319 1539
rect 3353 1505 3391 1539
rect 3425 1505 3463 1539
rect 3497 1505 3607 1539
rect 3641 1505 3679 1539
rect 3713 1505 3751 1539
rect 3785 1505 3823 1539
rect 3857 1505 3895 1539
rect 3929 1505 3967 1539
rect 4001 1505 4065 1539
rect 4099 1505 4137 1539
rect 4171 1505 4209 1539
rect 4243 1505 4281 1539
rect 4315 1505 4353 1539
rect 4387 1505 4425 1539
rect 4459 1505 4569 1539
rect 4603 1505 4641 1539
rect 4675 1505 4713 1539
rect 4747 1505 4785 1539
rect 4819 1505 4875 1539
rect 4909 1505 4947 1539
rect 4981 1505 5019 1539
rect 5053 1505 5091 1539
rect 5125 1505 5211 1539
rect -31 1492 5211 1505
rect 421 979 467 985
rect 3011 979 3057 985
rect 415 945 427 979
rect 461 945 3017 979
rect 3051 945 3063 979
rect 421 939 467 945
rect 3011 939 3057 945
rect 199 905 245 911
rect 2271 905 2317 911
rect 3381 905 3427 911
rect 4861 905 4907 911
rect 193 871 205 905
rect 239 871 2277 905
rect 2311 871 3387 905
rect 3421 871 4867 905
rect 4901 871 4913 905
rect 199 865 245 871
rect 2271 865 2317 871
rect 3381 865 3427 871
rect 4861 865 4907 871
rect 791 831 837 837
rect 1161 831 1207 837
rect 3751 831 3797 837
rect 4195 831 4241 837
rect 5009 831 5055 837
rect 785 797 797 831
rect 831 797 1167 831
rect 1201 797 3757 831
rect 3791 797 3803 831
rect 4189 797 4201 831
rect 4235 797 5015 831
rect 5049 797 5061 831
rect 791 791 837 797
rect 1161 791 1207 797
rect 3751 791 3797 797
rect 4195 791 4241 797
rect 5009 791 5055 797
rect 643 757 689 763
rect 1753 757 1799 763
rect 2123 757 2169 763
rect 2419 757 2465 763
rect 2789 757 2835 763
rect 4343 757 4389 763
rect 4713 757 4759 763
rect 637 723 649 757
rect 683 723 1759 757
rect 1793 723 2129 757
rect 2163 723 2175 757
rect 2413 723 2425 757
rect 2459 723 2795 757
rect 2829 723 2841 757
rect 4337 723 4349 757
rect 4383 723 4719 757
rect 4753 723 4765 757
rect 643 717 689 723
rect 1753 717 1799 723
rect 2123 717 2169 723
rect 2419 717 2465 723
rect 2789 717 2835 723
rect 4343 717 4389 723
rect 4713 717 4759 723
rect 1383 683 1429 689
rect 1353 649 1389 683
rect 1423 649 1435 683
rect 1383 643 1429 649
rect 1605 535 1651 541
rect 3233 535 3279 541
rect 3973 535 4019 541
rect 1599 501 1611 535
rect 1645 501 3239 535
rect 3273 501 3979 535
rect 4013 501 4025 535
rect 1605 495 1651 501
rect 3233 495 3279 501
rect 3973 495 4019 501
rect -31 47 5211 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 343 47
rect 377 13 415 47
rect 449 13 513 47
rect 547 13 585 47
rect 619 13 657 47
rect 691 13 729 47
rect 763 13 801 47
rect 835 13 873 47
rect 907 13 1017 47
rect 1051 13 1089 47
rect 1123 13 1161 47
rect 1195 13 1233 47
rect 1267 13 1305 47
rect 1339 13 1377 47
rect 1411 13 1475 47
rect 1509 13 1547 47
rect 1581 13 1619 47
rect 1653 13 1691 47
rect 1725 13 1763 47
rect 1797 13 1835 47
rect 1869 13 1979 47
rect 2013 13 2051 47
rect 2085 13 2123 47
rect 2157 13 2195 47
rect 2229 13 2285 47
rect 2319 13 2357 47
rect 2391 13 2429 47
rect 2463 13 2501 47
rect 2535 13 2645 47
rect 2679 13 2717 47
rect 2751 13 2789 47
rect 2823 13 2861 47
rect 2895 13 2933 47
rect 2967 13 3005 47
rect 3039 13 3103 47
rect 3137 13 3175 47
rect 3209 13 3247 47
rect 3281 13 3319 47
rect 3353 13 3391 47
rect 3425 13 3463 47
rect 3497 13 3607 47
rect 3641 13 3679 47
rect 3713 13 3751 47
rect 3785 13 3823 47
rect 3857 13 3895 47
rect 3929 13 3967 47
rect 4001 13 4065 47
rect 4099 13 4137 47
rect 4171 13 4209 47
rect 4243 13 4281 47
rect 4315 13 4353 47
rect 4387 13 4425 47
rect 4459 13 4569 47
rect 4603 13 4641 47
rect 4675 13 4713 47
rect 4747 13 4785 47
rect 4819 13 4875 47
rect 4909 13 4947 47
rect 4981 13 5019 47
rect 5053 13 5091 47
rect 5125 13 5211 47
rect -31 0 5211 13
<< labels >>
rlabel metal1 5015 797 5049 831 1 Q
port 1 n
rlabel metal1 4349 723 4383 757 1 QN
port 2 n
rlabel metal1 1389 649 1423 683 1 D
port 3 n
rlabel metal1 427 945 461 979 1 CLK
port 4 n
rlabel metal1 1611 501 1645 535 1 RN
port 5 n
rlabel metal1 55 1505 89 1539 1 VDD
port 6 n
rlabel metal1 55 13 89 47 1 VSS
port 7 n
<< end >>
