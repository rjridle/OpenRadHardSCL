magic
tech sky130A
magscale 1 2
timestamp 1643666983
<< nwell >>
rect -36 1337 470 1353
rect -36 1334 484 1337
rect -52 1267 484 1334
rect -36 1261 484 1267
rect -36 1061 470 1261
rect -36 956 472 1061
rect -36 950 -7 956
rect -36 893 470 950
rect 4 758 429 893
<< psubdiff >>
rect -49 501 482 552
rect -49 13 24 47
rect 58 13 93 47
rect 127 13 169 47
rect 203 13 237 47
rect 271 13 306 47
rect 340 13 374 47
rect 408 13 482 47
<< nsubdiff >>
rect -49 1283 24 1317
rect 58 1283 92 1317
rect 126 1283 160 1317
rect 195 1283 229 1317
rect 263 1283 297 1317
rect 331 1283 482 1317
rect -111 795 482 846
<< psubdiffcont >>
rect 24 13 58 47
rect 93 13 127 47
rect 169 13 203 47
rect 237 13 271 47
rect 306 13 340 47
rect 374 13 408 47
<< nsubdiffcont >>
rect 24 1283 58 1317
rect 92 1283 126 1317
rect 160 1283 195 1317
rect 229 1283 263 1317
rect 297 1283 331 1317
<< poly >>
rect 60 403 92 469
<< locali >>
rect -49 1317 482 1332
rect -49 1283 24 1317
rect 58 1283 92 1317
rect 126 1283 160 1317
rect 195 1283 229 1317
rect 263 1283 297 1317
rect 331 1283 482 1317
rect -49 1270 482 1283
rect 194 1230 228 1270
rect 18 1019 52 1029
rect 18 977 52 985
rect 370 1019 404 1029
rect 370 977 404 985
rect 108 290 142 657
rect 292 290 326 296
rect 292 250 326 256
rect 16 62 50 109
rect 108 62 142 117
rect 200 62 234 107
rect 292 62 326 117
rect 384 62 418 101
rect -49 47 482 62
rect -49 13 24 47
rect 58 13 93 47
rect 127 13 169 47
rect 203 13 237 47
rect 271 13 306 47
rect 340 13 374 47
rect 408 13 482 47
rect -49 0 482 13
<< viali >>
rect 24 1283 58 1317
rect 92 1283 126 1317
rect 160 1283 195 1317
rect 229 1283 263 1317
rect 297 1283 331 1317
rect 18 985 52 1019
rect 370 985 404 1019
rect 108 256 142 290
rect 292 256 326 290
rect 24 13 58 47
rect 93 13 127 47
rect 169 13 203 47
rect 237 13 271 47
rect 306 13 340 47
rect 374 13 408 47
<< metal1 >>
rect -49 1317 482 1332
rect -49 1283 24 1317
rect 58 1283 92 1317
rect 126 1283 160 1317
rect 195 1283 229 1317
rect 263 1283 297 1317
rect 331 1283 482 1317
rect -49 1270 482 1283
rect 12 1019 58 1025
rect 364 1019 410 1025
rect 6 985 18 1019
rect 52 985 370 1019
rect 404 985 416 1019
rect 12 979 58 985
rect 108 750 142 985
rect 364 979 410 985
rect 102 290 148 296
rect 286 290 332 296
rect 96 256 108 290
rect 142 256 292 290
rect 326 256 338 290
rect 102 255 332 256
rect 102 250 148 255
rect 286 250 332 255
rect -49 47 482 62
rect -49 13 24 47
rect 58 13 93 47
rect 127 13 169 47
rect 203 13 237 47
rect 271 13 306 47
rect 340 13 374 47
rect 408 13 482 47
rect -49 0 482 13
use M1_M2_contact  M1_M2_contact_0 ./pcells
timestamp 1643652910
transform 1 0 -64 0 1 4
box 64 391 130 473
use diff_ring_side  diff_ring_side_1 pcells
timestamp 1643181737
transform 1 0 588 0 1 0
box -159 0 9 1353
use diff_ring_side  diff_ring_side_0
timestamp 1643181737
transform 1 0 -5 0 1 0
box -159 0 9 1353
use pmos  pmos_1 pcells
timestamp 1643179034
transform 1 0 184 0 1 1228
box -36 -312 264 42
use pmos  pmos_0
timestamp 1643179034
transform 1 0 8 0 1 1228
box -36 -312 264 42
use nmos_top_left  nmos_top_left_1 pcells
timestamp 1643656170
transform 1 0 235 0 1 165
box -45 -64 193 238
use nmos_top_left  nmos_top_left_0
timestamp 1643656170
transform 1 0 51 0 1 165
box -45 -64 193 238
<< labels >>
rlabel metal1 161 1325 161 1325 1 VDD
port 1 n
rlabel metal1 148 31 148 31 1 VSS
port 2 n
rlabel metal1 370 985 404 1019 1 YN
port 5 n
<< end >>
