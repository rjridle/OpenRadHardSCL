* HSPICE file created from tmp.ext - technology: sky130A

.option scale=5000u

.subckt tmp A Y VDD VSS
X0 Y A VDD VDD sky130_fd_pr__pfet_01v8 ad=11600 pd=458 as=22000 ps=910 w=400 l=30 M=2
X1 Y A VSS VSS sky130_fd_pr__nfet_01v8 ad=7088 pd=312 as=46290 ps=1624 w=598 l=30
.ends

** hspice subcircuit dictionary
