magic
tech sky130A
magscale 1 2
timestamp 1651077592
<< metal1 >>
rect -31 1492 2251 1554
rect 131 871 165 905
rect 2055 871 2089 905
rect 1611 723 1645 757
rect -31 0 2251 62
use xor2X1_pcell  xor2X1_pcell_0 pcells
timestamp 1648314317
transform 1 0 0 0 1 0
box -84 0 2304 1575
<< labels >>
rlabel metal1 1611 723 1645 757 1 Y
port 1 n
rlabel metal1 131 871 165 905 1 A
port 2 n
rlabel metal1 2055 871 2089 905 1 B
port 3 n
rlabel metal1 -31 1492 2251 1554 1 VDD
rlabel metal1 -31 0 2251 62 1 GND
<< end >>
