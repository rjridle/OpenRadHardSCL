magic
tech sky130A
magscale 1 2
timestamp 1648324032
<< nwell >>
rect -84 832 1490 1575
<< nmos >>
rect 164 316 194 377
tri 194 316 210 332 sw
rect 358 324 388 377
tri 388 324 404 340 sw
rect 164 286 270 316
tri 270 286 300 316 sw
rect 358 294 464 324
tri 464 294 494 324 sw
rect 164 185 194 286
tri 194 270 210 286 nw
tri 254 270 270 286 ne
tri 194 185 210 201 sw
tri 254 185 270 201 se
rect 270 185 300 286
rect 358 193 388 294
tri 388 278 404 294 nw
tri 448 278 464 294 ne
tri 388 193 404 209 sw
tri 448 193 464 209 se
rect 464 193 494 294
tri 164 155 194 185 ne
rect 194 155 270 185
tri 270 155 300 185 nw
tri 358 163 388 193 ne
rect 388 163 464 193
tri 464 163 494 193 nw
tri 752 316 768 332 se
rect 768 316 798 377
tri 662 286 692 316 se
rect 692 286 798 316
rect 662 185 692 286
tri 692 270 708 286 nw
tri 752 270 768 286 ne
tri 692 185 708 201 sw
tri 752 185 768 201 se
rect 768 185 798 286
tri 662 155 692 185 ne
rect 692 155 768 185
tri 768 155 798 185 nw
rect 1117 324 1147 377
tri 1147 324 1163 340 sw
rect 1117 294 1223 324
tri 1223 294 1253 324 sw
rect 1117 193 1147 294
tri 1147 278 1163 294 nw
tri 1207 278 1223 294 ne
tri 1147 193 1163 209 sw
tri 1207 193 1223 209 se
rect 1223 193 1253 294
tri 1117 163 1147 193 ne
rect 1147 163 1223 193
tri 1223 163 1253 193 nw
<< pmos >>
rect 193 1051 223 1451
rect 281 1051 311 1451
rect 369 1051 399 1451
rect 457 1051 487 1451
rect 653 1051 683 1451
rect 741 1051 771 1451
rect 1125 1050 1155 1450
rect 1213 1050 1243 1450
<< ndiff >>
rect 108 361 164 377
rect 108 327 118 361
rect 152 327 164 361
rect 108 289 164 327
rect 194 361 358 377
rect 194 332 215 361
tri 194 316 210 332 ne
rect 210 327 215 332
rect 249 327 312 361
rect 346 327 358 361
rect 210 316 358 327
rect 388 340 550 377
tri 388 324 404 340 ne
rect 404 324 550 340
rect 108 255 118 289
rect 152 255 164 289
tri 270 286 300 316 ne
rect 300 289 358 316
tri 464 294 494 324 ne
rect 108 221 164 255
rect 108 187 118 221
rect 152 187 164 221
rect 108 155 164 187
tri 194 270 210 286 se
rect 210 270 254 286
tri 254 270 270 286 sw
rect 194 236 270 270
rect 194 202 215 236
rect 249 202 270 236
rect 194 201 270 202
tri 194 185 210 201 ne
rect 210 185 254 201
tri 254 185 270 201 nw
rect 300 255 312 289
rect 346 255 358 289
rect 300 221 358 255
rect 300 187 312 221
rect 346 187 358 221
tri 388 278 404 294 se
rect 404 278 448 294
tri 448 278 464 294 sw
rect 388 245 464 278
rect 388 211 409 245
rect 443 211 464 245
rect 388 209 464 211
tri 388 193 404 209 ne
rect 404 193 448 209
tri 448 193 464 209 nw
rect 494 289 550 324
rect 494 255 506 289
rect 540 255 550 289
rect 494 221 550 255
tri 164 155 194 185 sw
tri 270 155 300 185 se
rect 300 163 358 187
tri 358 163 388 193 sw
tri 464 163 494 193 se
rect 494 187 506 221
rect 540 187 550 221
rect 494 163 550 187
rect 300 155 550 163
rect 108 151 550 155
rect 108 117 118 151
rect 152 117 312 151
rect 346 117 409 151
rect 443 117 506 151
rect 540 117 550 151
rect 108 101 550 117
rect 606 361 768 377
rect 606 327 616 361
rect 650 327 713 361
rect 747 332 768 361
rect 747 327 752 332
rect 606 316 752 327
tri 752 316 768 332 nw
rect 798 361 854 377
rect 798 327 810 361
rect 844 327 854 361
rect 606 289 662 316
rect 606 255 616 289
rect 650 255 662 289
tri 662 286 692 316 nw
rect 798 289 854 327
rect 606 221 662 255
rect 606 187 616 221
rect 650 187 662 221
rect 606 155 662 187
tri 692 270 708 286 se
rect 708 270 752 286
tri 752 270 768 286 sw
rect 692 236 768 270
rect 692 202 713 236
rect 747 202 768 236
rect 692 201 768 202
tri 692 185 708 201 ne
rect 708 185 752 201
tri 752 185 768 201 nw
rect 798 255 810 289
rect 844 255 854 289
rect 798 221 854 255
rect 798 187 810 221
rect 844 187 854 221
tri 662 155 692 185 sw
tri 768 155 798 185 se
rect 798 155 854 187
rect 606 151 854 155
rect 606 117 616 151
rect 650 117 810 151
rect 844 117 854 151
rect 606 101 854 117
rect 1061 361 1117 377
rect 1061 327 1071 361
rect 1105 327 1117 361
rect 1061 289 1117 327
rect 1147 361 1307 377
rect 1147 340 1265 361
tri 1147 324 1163 340 ne
rect 1163 327 1265 340
rect 1299 327 1307 361
rect 1163 324 1307 327
tri 1223 294 1253 324 ne
rect 1061 255 1071 289
rect 1105 255 1117 289
rect 1061 221 1117 255
rect 1061 187 1071 221
rect 1105 187 1117 221
tri 1147 278 1163 294 se
rect 1163 278 1207 294
tri 1207 278 1223 294 sw
rect 1147 245 1223 278
rect 1147 211 1167 245
rect 1201 211 1223 245
rect 1147 209 1223 211
tri 1147 193 1163 209 ne
rect 1163 193 1207 209
tri 1207 193 1223 209 nw
rect 1253 289 1307 324
rect 1253 255 1265 289
rect 1299 255 1307 289
rect 1253 221 1307 255
rect 1061 163 1117 187
tri 1117 163 1147 193 sw
tri 1223 163 1253 193 se
rect 1253 187 1265 221
rect 1299 187 1307 221
rect 1253 163 1307 187
rect 1061 151 1307 163
rect 1061 117 1071 151
rect 1105 117 1167 151
rect 1201 117 1265 151
rect 1299 117 1307 151
rect 1061 101 1307 117
<< pdiff >>
rect 137 1411 193 1451
rect 137 1377 147 1411
rect 181 1377 193 1411
rect 137 1343 193 1377
rect 137 1309 147 1343
rect 181 1309 193 1343
rect 137 1275 193 1309
rect 137 1241 147 1275
rect 181 1241 193 1275
rect 137 1207 193 1241
rect 137 1173 147 1207
rect 181 1173 193 1207
rect 137 1051 193 1173
rect 223 1411 281 1451
rect 223 1377 235 1411
rect 269 1377 281 1411
rect 223 1343 281 1377
rect 223 1309 235 1343
rect 269 1309 281 1343
rect 223 1275 281 1309
rect 223 1241 235 1275
rect 269 1241 281 1275
rect 223 1207 281 1241
rect 223 1173 235 1207
rect 269 1173 281 1207
rect 223 1139 281 1173
rect 223 1105 235 1139
rect 269 1105 281 1139
rect 223 1051 281 1105
rect 311 1411 369 1451
rect 311 1377 323 1411
rect 357 1377 369 1411
rect 311 1343 369 1377
rect 311 1309 323 1343
rect 357 1309 369 1343
rect 311 1275 369 1309
rect 311 1241 323 1275
rect 357 1241 369 1275
rect 311 1207 369 1241
rect 311 1173 323 1207
rect 357 1173 369 1207
rect 311 1051 369 1173
rect 399 1413 457 1451
rect 399 1377 411 1413
rect 445 1377 457 1413
rect 399 1343 457 1377
rect 399 1309 411 1343
rect 445 1309 457 1343
rect 399 1275 457 1309
rect 399 1241 411 1275
rect 445 1241 457 1275
rect 399 1207 457 1241
rect 399 1173 411 1207
rect 445 1173 457 1207
rect 399 1139 457 1173
rect 399 1105 411 1139
rect 445 1105 457 1139
rect 399 1051 457 1105
rect 487 1411 541 1451
rect 487 1377 499 1411
rect 533 1377 541 1411
rect 487 1343 541 1377
rect 487 1309 499 1343
rect 533 1309 541 1343
rect 487 1275 541 1309
rect 487 1241 499 1275
rect 533 1241 541 1275
rect 487 1207 541 1241
rect 487 1173 499 1207
rect 533 1173 541 1207
rect 487 1051 541 1173
rect 597 1343 653 1451
rect 597 1309 607 1343
rect 641 1309 653 1343
rect 597 1275 653 1309
rect 597 1241 607 1275
rect 641 1241 653 1275
rect 597 1207 653 1241
rect 597 1173 607 1207
rect 641 1173 653 1207
rect 597 1051 653 1173
rect 683 1343 741 1451
rect 683 1309 695 1343
rect 729 1309 741 1343
rect 683 1275 741 1309
rect 683 1241 695 1275
rect 729 1241 741 1275
rect 683 1207 741 1241
rect 683 1173 695 1207
rect 729 1173 741 1207
rect 683 1051 741 1173
rect 771 1343 825 1451
rect 771 1309 783 1343
rect 817 1309 825 1343
rect 771 1275 825 1309
rect 771 1241 783 1275
rect 817 1241 825 1275
rect 771 1207 825 1241
rect 771 1173 783 1207
rect 817 1173 825 1207
rect 771 1051 825 1173
rect 1069 1412 1125 1450
rect 1069 1378 1079 1412
rect 1113 1378 1125 1412
rect 1069 1344 1125 1378
rect 1069 1310 1079 1344
rect 1113 1310 1125 1344
rect 1069 1276 1125 1310
rect 1069 1242 1079 1276
rect 1113 1242 1125 1276
rect 1069 1208 1125 1242
rect 1069 1174 1079 1208
rect 1113 1174 1125 1208
rect 1069 1139 1125 1174
rect 1069 1105 1079 1139
rect 1113 1105 1125 1139
rect 1069 1050 1125 1105
rect 1155 1412 1213 1450
rect 1155 1378 1167 1412
rect 1201 1378 1213 1412
rect 1155 1344 1213 1378
rect 1155 1310 1167 1344
rect 1201 1310 1213 1344
rect 1155 1276 1213 1310
rect 1155 1242 1167 1276
rect 1201 1242 1213 1276
rect 1155 1208 1213 1242
rect 1155 1174 1167 1208
rect 1201 1174 1213 1208
rect 1155 1139 1213 1174
rect 1155 1105 1167 1139
rect 1201 1105 1213 1139
rect 1155 1050 1213 1105
rect 1243 1412 1297 1450
rect 1243 1378 1255 1412
rect 1289 1378 1297 1412
rect 1243 1344 1297 1378
rect 1243 1310 1255 1344
rect 1289 1310 1297 1344
rect 1243 1276 1297 1310
rect 1243 1242 1255 1276
rect 1289 1242 1297 1276
rect 1243 1208 1297 1242
rect 1243 1174 1255 1208
rect 1289 1174 1297 1208
rect 1243 1139 1297 1174
rect 1243 1105 1255 1139
rect 1289 1105 1297 1139
rect 1243 1050 1297 1105
<< ndiffc >>
rect 118 327 152 361
rect 215 327 249 361
rect 312 327 346 361
rect 118 255 152 289
rect 118 187 152 221
rect 215 202 249 236
rect 312 255 346 289
rect 312 187 346 221
rect 409 211 443 245
rect 506 255 540 289
rect 506 187 540 221
rect 118 117 152 151
rect 312 117 346 151
rect 409 117 443 151
rect 506 117 540 151
rect 616 327 650 361
rect 713 327 747 361
rect 810 327 844 361
rect 616 255 650 289
rect 616 187 650 221
rect 713 202 747 236
rect 810 255 844 289
rect 810 187 844 221
rect 616 117 650 151
rect 810 117 844 151
rect 1071 327 1105 361
rect 1265 327 1299 361
rect 1071 255 1105 289
rect 1071 187 1105 221
rect 1167 211 1201 245
rect 1265 255 1299 289
rect 1265 187 1299 221
rect 1071 117 1105 151
rect 1167 117 1201 151
rect 1265 117 1299 151
<< pdiffc >>
rect 147 1377 181 1411
rect 147 1309 181 1343
rect 147 1241 181 1275
rect 147 1173 181 1207
rect 235 1377 269 1411
rect 235 1309 269 1343
rect 235 1241 269 1275
rect 235 1173 269 1207
rect 235 1105 269 1139
rect 323 1377 357 1411
rect 323 1309 357 1343
rect 323 1241 357 1275
rect 323 1173 357 1207
rect 411 1377 445 1413
rect 411 1309 445 1343
rect 411 1241 445 1275
rect 411 1173 445 1207
rect 411 1105 445 1139
rect 499 1377 533 1411
rect 499 1309 533 1343
rect 499 1241 533 1275
rect 499 1173 533 1207
rect 607 1309 641 1343
rect 607 1241 641 1275
rect 607 1173 641 1207
rect 695 1309 729 1343
rect 695 1241 729 1275
rect 695 1173 729 1207
rect 783 1309 817 1343
rect 783 1241 817 1275
rect 783 1173 817 1207
rect 1079 1378 1113 1412
rect 1079 1310 1113 1344
rect 1079 1242 1113 1276
rect 1079 1174 1113 1208
rect 1079 1105 1113 1139
rect 1167 1378 1201 1412
rect 1167 1310 1201 1344
rect 1167 1242 1201 1276
rect 1167 1174 1201 1208
rect 1167 1105 1201 1139
rect 1255 1378 1289 1412
rect 1255 1310 1289 1344
rect 1255 1242 1289 1276
rect 1255 1174 1289 1208
rect 1255 1105 1289 1139
<< psubdiff >>
rect -31 571 635 572
rect 931 571 1437 572
rect -31 546 1437 571
rect -31 512 -17 546
rect 17 512 945 546
rect 979 512 1389 546
rect 1423 512 1437 546
rect -31 510 1437 512
rect -31 474 31 510
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect -31 368 -17 402
rect 17 368 31 402
rect 931 474 993 510
rect 931 440 945 474
rect 979 440 993 474
rect 931 402 993 440
rect 1375 474 1437 510
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect 931 368 945 402
rect 979 368 993 402
rect 1375 440 1389 474
rect 1423 440 1437 474
rect 1375 402 1437 440
rect 931 330 993 368
rect 931 296 945 330
rect 979 296 993 330
rect 931 258 993 296
rect 931 224 945 258
rect 979 224 993 258
rect 931 186 993 224
rect 931 152 945 186
rect 979 152 993 186
rect 931 114 993 152
rect -31 47 31 80
rect 931 80 945 114
rect 979 80 993 114
rect 1375 368 1389 402
rect 1423 368 1437 402
rect 1375 330 1437 368
rect 1375 296 1389 330
rect 1423 296 1437 330
rect 1375 258 1437 296
rect 1375 224 1389 258
rect 1423 224 1437 258
rect 1375 186 1437 224
rect 1375 152 1389 186
rect 1423 152 1437 186
rect 1375 114 1437 152
rect 931 47 993 80
rect 1375 80 1389 114
rect 1423 80 1437 114
rect 1375 47 1437 80
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 343 47
rect 377 13 415 47
rect 449 13 513 47
rect 547 13 585 47
rect 619 13 657 47
rect 691 13 729 47
rect 763 13 801 47
rect 835 13 873 47
rect 907 13 1017 47
rect 1051 13 1089 47
rect 1123 13 1167 47
rect 1201 13 1245 47
rect 1279 13 1317 47
rect 1351 13 1437 47
rect -31 11 31 13
rect 931 11 993 13
rect 1375 11 1437 13
<< nsubdiff >>
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 343 1539
rect 377 1505 415 1539
rect 449 1505 513 1539
rect 547 1505 585 1539
rect 619 1505 657 1539
rect 691 1505 729 1539
rect 763 1505 801 1539
rect 835 1505 873 1539
rect 907 1505 1017 1539
rect 1051 1505 1089 1539
rect 1123 1505 1167 1539
rect 1201 1505 1245 1539
rect 1279 1505 1317 1539
rect 1351 1505 1437 1539
rect -31 1470 31 1505
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect 931 1470 993 1505
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect -31 1038 31 1076
rect 931 1436 945 1470
rect 979 1436 993 1470
rect 1375 1470 1437 1505
rect 931 1398 993 1436
rect 931 1364 945 1398
rect 979 1364 993 1398
rect 931 1326 993 1364
rect 931 1292 945 1326
rect 979 1292 993 1326
rect 931 1254 993 1292
rect 931 1220 945 1254
rect 979 1220 993 1254
rect 931 1182 993 1220
rect 931 1148 945 1182
rect 979 1148 993 1182
rect 931 1110 993 1148
rect 931 1076 945 1110
rect 979 1076 993 1110
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect 931 1038 993 1076
rect 1375 1436 1389 1470
rect 1423 1436 1437 1470
rect 1375 1398 1437 1436
rect 1375 1364 1389 1398
rect 1423 1364 1437 1398
rect 1375 1326 1437 1364
rect 1375 1292 1389 1326
rect 1423 1292 1437 1326
rect 1375 1254 1437 1292
rect 1375 1220 1389 1254
rect 1423 1220 1437 1254
rect 1375 1182 1437 1220
rect 1375 1148 1389 1182
rect 1423 1148 1437 1182
rect 1375 1110 1437 1148
rect 1375 1076 1389 1110
rect 1423 1076 1437 1110
rect 931 1004 945 1038
rect 979 1004 993 1038
rect 931 966 993 1004
rect -31 930 31 932
rect 931 932 945 966
rect 979 932 993 966
rect 1375 1038 1437 1076
rect 1375 1004 1389 1038
rect 1423 1004 1437 1038
rect 1375 966 1437 1004
rect 931 930 993 932
rect 1375 932 1389 966
rect 1423 932 1437 966
rect 1375 930 1437 932
rect -31 868 1437 930
<< psubdiffcont >>
rect -17 512 17 546
rect 945 512 979 546
rect 1389 512 1423 546
rect -17 440 17 474
rect -17 368 17 402
rect 945 440 979 474
rect -17 296 17 330
rect -17 224 17 258
rect -17 152 17 186
rect -17 80 17 114
rect 945 368 979 402
rect 1389 440 1423 474
rect 945 296 979 330
rect 945 224 979 258
rect 945 152 979 186
rect 945 80 979 114
rect 1389 368 1423 402
rect 1389 296 1423 330
rect 1389 224 1423 258
rect 1389 152 1423 186
rect 1389 80 1423 114
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 343 13 377 47
rect 415 13 449 47
rect 513 13 547 47
rect 585 13 619 47
rect 657 13 691 47
rect 729 13 763 47
rect 801 13 835 47
rect 873 13 907 47
rect 1017 13 1051 47
rect 1089 13 1123 47
rect 1167 13 1201 47
rect 1245 13 1279 47
rect 1317 13 1351 47
<< nsubdiffcont >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 343 1505 377 1539
rect 415 1505 449 1539
rect 513 1505 547 1539
rect 585 1505 619 1539
rect 657 1505 691 1539
rect 729 1505 763 1539
rect 801 1505 835 1539
rect 873 1505 907 1539
rect 1017 1505 1051 1539
rect 1089 1505 1123 1539
rect 1167 1505 1201 1539
rect 1245 1505 1279 1539
rect 1317 1505 1351 1539
rect -17 1436 17 1470
rect -17 1364 17 1398
rect -17 1292 17 1326
rect -17 1220 17 1254
rect -17 1148 17 1182
rect -17 1076 17 1110
rect 945 1436 979 1470
rect 945 1364 979 1398
rect 945 1292 979 1326
rect 945 1220 979 1254
rect 945 1148 979 1182
rect 945 1076 979 1110
rect -17 1004 17 1038
rect -17 932 17 966
rect 1389 1436 1423 1470
rect 1389 1364 1423 1398
rect 1389 1292 1423 1326
rect 1389 1220 1423 1254
rect 1389 1148 1423 1182
rect 1389 1076 1423 1110
rect 945 1004 979 1038
rect 945 932 979 966
rect 1389 1004 1423 1038
rect 1389 932 1423 966
<< poly >>
rect 193 1451 223 1477
rect 281 1451 311 1477
rect 369 1451 399 1477
rect 457 1451 487 1477
rect 653 1451 683 1477
rect 741 1451 771 1477
rect 1125 1450 1155 1476
rect 1213 1450 1243 1476
rect 193 1020 223 1051
rect 281 1020 311 1051
rect 369 1020 399 1051
rect 457 1020 487 1051
rect 193 1004 311 1020
rect 193 990 205 1004
rect 195 970 205 990
rect 239 990 311 1004
rect 359 1004 487 1020
rect 239 970 249 990
rect 195 954 249 970
rect 359 970 369 1004
rect 403 990 487 1004
rect 653 1020 683 1051
rect 741 1020 771 1051
rect 653 1004 841 1020
rect 653 990 797 1004
rect 403 970 413 990
rect 359 954 413 970
rect 787 970 797 990
rect 831 970 841 1004
rect 787 954 841 970
rect 1125 1019 1155 1050
rect 1213 1019 1243 1050
rect 1083 1003 1243 1019
rect 1083 969 1093 1003
rect 1127 989 1243 1003
rect 1127 969 1137 989
rect 1083 953 1137 969
rect 195 461 249 477
rect 195 441 205 461
rect 164 427 205 441
rect 239 427 249 461
rect 164 411 249 427
rect 343 461 397 477
rect 343 427 353 461
rect 387 427 397 461
rect 787 461 841 477
rect 787 441 797 461
rect 343 411 397 427
rect 768 427 797 441
rect 831 427 841 461
rect 768 411 841 427
rect 164 377 194 411
rect 358 377 388 411
rect 768 377 798 411
rect 1083 461 1137 477
rect 1083 427 1093 461
rect 1127 441 1137 461
rect 1127 427 1147 441
rect 1083 411 1147 427
rect 1117 377 1147 411
<< polycont >>
rect 205 970 239 1004
rect 369 970 403 1004
rect 797 970 831 1004
rect 1093 969 1127 1003
rect 205 427 239 461
rect 353 427 387 461
rect 797 427 831 461
rect 1093 427 1127 461
<< locali >>
rect -31 1539 1437 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 343 1539
rect 377 1505 415 1539
rect 449 1505 513 1539
rect 547 1505 585 1539
rect 619 1505 657 1539
rect 691 1505 729 1539
rect 763 1505 801 1539
rect 835 1505 873 1539
rect 907 1505 1017 1539
rect 1051 1505 1089 1539
rect 1123 1505 1167 1539
rect 1201 1505 1245 1539
rect 1279 1505 1317 1539
rect 1351 1505 1437 1539
rect -31 1492 1437 1505
rect -31 1470 31 1492
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect 147 1411 181 1492
rect 147 1343 181 1377
rect 147 1275 181 1309
rect 147 1207 181 1241
rect 147 1157 181 1173
rect 235 1411 269 1445
rect 235 1343 269 1377
rect 235 1275 269 1309
rect 235 1207 269 1241
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect -31 1038 31 1076
rect 235 1139 269 1173
rect 323 1411 357 1492
rect 323 1343 357 1377
rect 323 1275 357 1309
rect 323 1207 357 1241
rect 323 1157 357 1173
rect 411 1413 445 1429
rect 411 1343 445 1377
rect 411 1275 445 1309
rect 411 1207 445 1241
rect 411 1139 445 1173
rect 499 1411 533 1492
rect 931 1470 993 1492
rect 499 1343 533 1377
rect 499 1275 533 1309
rect 499 1207 533 1241
rect 499 1157 533 1173
rect 607 1411 817 1445
rect 607 1343 641 1411
rect 607 1275 641 1309
rect 607 1207 641 1241
rect 607 1105 641 1173
rect 235 1071 641 1105
rect 695 1343 729 1359
rect 695 1275 729 1309
rect 695 1207 729 1241
rect 695 1105 729 1173
rect 783 1343 817 1411
rect 783 1275 817 1309
rect 783 1207 817 1241
rect 783 1157 817 1173
rect 931 1436 945 1470
rect 979 1436 993 1470
rect 931 1398 993 1436
rect 931 1364 945 1398
rect 979 1364 993 1398
rect 931 1326 993 1364
rect 931 1292 945 1326
rect 979 1292 993 1326
rect 931 1254 993 1292
rect 931 1220 945 1254
rect 979 1220 993 1254
rect 931 1182 993 1220
rect 931 1148 945 1182
rect 979 1148 993 1182
rect 931 1110 993 1148
rect 695 1071 757 1105
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect -31 868 31 932
rect 205 1004 239 1020
rect 369 1004 403 1020
rect 205 609 239 970
rect -31 546 31 572
rect -31 512 -17 546
rect 17 512 31 546
rect -31 474 31 512
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect 205 461 239 575
rect 205 411 239 427
rect 353 970 369 988
rect 353 954 403 970
rect 353 683 387 954
rect 353 461 387 649
rect 353 411 387 427
rect 723 905 757 1071
rect 931 1076 945 1110
rect 979 1076 993 1110
rect 1079 1412 1113 1492
rect 1079 1344 1113 1378
rect 1079 1276 1113 1310
rect 1079 1208 1113 1242
rect 1079 1139 1113 1174
rect 1079 1083 1113 1105
rect 1167 1412 1201 1450
rect 1167 1344 1201 1378
rect 1167 1276 1201 1310
rect 1167 1208 1201 1242
rect 1167 1139 1201 1174
rect 931 1038 993 1076
rect 723 757 757 871
rect -31 368 -17 402
rect 17 368 31 402
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect 118 361 152 377
rect 312 361 346 377
rect 616 373 650 377
rect 152 327 215 361
rect 249 327 312 361
rect 118 289 152 327
rect 118 221 152 255
rect 312 289 346 327
rect 118 151 152 187
rect 118 101 152 117
rect 215 236 249 252
rect -31 62 31 80
rect 215 62 249 202
rect 312 221 346 255
rect 409 361 650 373
rect 723 361 757 723
rect 797 1004 831 1020
rect 797 461 831 970
rect 931 1004 945 1038
rect 979 1004 993 1038
rect 931 966 993 1004
rect 931 932 945 966
rect 979 932 993 966
rect 931 868 993 932
rect 1093 1003 1127 1019
rect 1093 905 1127 969
rect 1167 979 1201 1105
rect 1255 1412 1289 1492
rect 1255 1344 1289 1378
rect 1255 1276 1289 1310
rect 1255 1208 1289 1242
rect 1255 1139 1289 1174
rect 1255 1083 1289 1105
rect 1375 1470 1437 1492
rect 1375 1436 1389 1470
rect 1423 1436 1437 1470
rect 1375 1398 1437 1436
rect 1375 1364 1389 1398
rect 1423 1364 1437 1398
rect 1375 1326 1437 1364
rect 1375 1292 1389 1326
rect 1423 1292 1437 1326
rect 1375 1254 1437 1292
rect 1375 1220 1389 1254
rect 1423 1220 1437 1254
rect 1375 1182 1437 1220
rect 1375 1148 1389 1182
rect 1423 1148 1437 1182
rect 1375 1110 1437 1148
rect 1375 1076 1389 1110
rect 1423 1076 1437 1110
rect 1375 1038 1437 1076
rect 1375 1004 1389 1038
rect 1423 1004 1437 1038
rect 1167 945 1275 979
rect 797 411 831 427
rect 931 546 993 572
rect 931 512 945 546
rect 979 512 993 546
rect 931 474 993 512
rect 931 440 945 474
rect 979 440 993 474
rect 931 402 993 440
rect 1093 461 1127 871
rect 1241 757 1275 945
rect 1375 966 1437 1004
rect 1375 932 1389 966
rect 1423 932 1437 966
rect 1375 868 1437 932
rect 1241 461 1275 723
rect 1093 411 1127 427
rect 1167 427 1275 461
rect 1375 546 1437 572
rect 1375 512 1389 546
rect 1423 512 1437 546
rect 1375 474 1437 512
rect 1375 440 1389 474
rect 1423 440 1437 474
rect 810 361 844 377
rect 409 339 616 361
rect 409 245 443 339
rect 650 327 713 361
rect 747 327 810 361
rect 409 195 443 211
rect 506 289 540 305
rect 506 221 540 255
rect 312 151 346 187
rect 506 151 540 187
rect 346 117 409 151
rect 443 117 506 151
rect 312 101 346 117
rect 506 101 540 117
rect 616 289 650 327
rect 616 221 650 255
rect 810 289 844 327
rect 616 151 650 187
rect 616 101 650 117
rect 713 236 747 252
rect 713 62 747 202
rect 810 221 844 255
rect 810 151 844 187
rect 810 101 844 117
rect 931 368 945 402
rect 979 368 993 402
rect 931 330 993 368
rect 931 296 945 330
rect 979 296 993 330
rect 931 258 993 296
rect 931 224 945 258
rect 979 224 993 258
rect 931 186 993 224
rect 931 152 945 186
rect 979 152 993 186
rect 931 114 993 152
rect 931 80 945 114
rect 979 80 993 114
rect 931 62 993 80
rect 1071 361 1105 377
rect 1071 289 1105 327
rect 1071 221 1105 255
rect 1167 245 1201 427
rect 1375 402 1437 440
rect 1167 195 1201 211
rect 1265 361 1299 377
rect 1265 289 1299 327
rect 1265 221 1299 255
rect 1071 151 1105 187
rect 1265 151 1299 187
rect 1105 117 1167 151
rect 1201 117 1265 151
rect 1071 62 1105 117
rect 1168 62 1202 117
rect 1265 62 1299 117
rect 1375 368 1389 402
rect 1423 368 1437 402
rect 1375 330 1437 368
rect 1375 296 1389 330
rect 1423 296 1437 330
rect 1375 258 1437 296
rect 1375 224 1389 258
rect 1423 224 1437 258
rect 1375 186 1437 224
rect 1375 152 1389 186
rect 1423 152 1437 186
rect 1375 114 1437 152
rect 1375 80 1389 114
rect 1423 80 1437 114
rect 1375 62 1437 80
rect -31 47 1437 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 343 47
rect 377 13 415 47
rect 449 13 513 47
rect 547 13 585 47
rect 619 13 657 47
rect 691 13 729 47
rect 763 13 801 47
rect 835 13 873 47
rect 907 13 1017 47
rect 1051 13 1089 47
rect 1123 13 1167 47
rect 1201 13 1245 47
rect 1279 13 1317 47
rect 1351 13 1437 47
rect -31 0 1437 13
<< viali >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 343 1505 377 1539
rect 415 1505 449 1539
rect 513 1505 547 1539
rect 585 1505 619 1539
rect 657 1505 691 1539
rect 729 1505 763 1539
rect 801 1505 835 1539
rect 873 1505 907 1539
rect 1017 1505 1051 1539
rect 1089 1505 1123 1539
rect 1167 1505 1201 1539
rect 1245 1505 1279 1539
rect 1317 1505 1351 1539
rect 205 575 239 609
rect 353 649 387 683
rect 723 871 757 905
rect 723 723 757 757
rect 1093 871 1127 905
rect 1241 723 1275 757
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 343 13 377 47
rect 415 13 449 47
rect 513 13 547 47
rect 585 13 619 47
rect 657 13 691 47
rect 729 13 763 47
rect 801 13 835 47
rect 873 13 907 47
rect 1017 13 1051 47
rect 1089 13 1123 47
rect 1167 13 1201 47
rect 1245 13 1279 47
rect 1317 13 1351 47
<< metal1 >>
rect -31 1539 1437 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 343 1539
rect 377 1505 415 1539
rect 449 1505 513 1539
rect 547 1505 585 1539
rect 619 1505 657 1539
rect 691 1505 729 1539
rect 763 1505 801 1539
rect 835 1505 873 1539
rect 907 1505 1017 1539
rect 1051 1505 1089 1539
rect 1123 1505 1167 1539
rect 1201 1505 1245 1539
rect 1279 1505 1317 1539
rect 1351 1505 1437 1539
rect -31 1492 1437 1505
rect 717 905 763 911
rect 1087 905 1133 911
rect 711 871 723 905
rect 757 871 1093 905
rect 1127 871 1139 905
rect 717 865 763 871
rect 1087 865 1133 871
rect 717 757 763 763
rect 1235 757 1281 763
rect 687 723 723 757
rect 757 723 769 757
rect 1229 723 1241 757
rect 1275 723 1311 757
rect 717 717 763 723
rect 1235 717 1281 723
rect 347 683 393 689
rect 317 649 353 683
rect 387 649 399 683
rect 347 643 393 649
rect 199 609 245 615
rect 169 575 205 609
rect 239 575 251 609
rect 199 569 245 575
rect -31 47 1437 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 343 47
rect 377 13 415 47
rect 449 13 513 47
rect 547 13 585 47
rect 619 13 657 47
rect 691 13 729 47
rect 763 13 801 47
rect 835 13 873 47
rect 907 13 1017 47
rect 1051 13 1089 47
rect 1123 13 1167 47
rect 1201 13 1245 47
rect 1279 13 1317 47
rect 1351 13 1437 47
rect -31 0 1437 13
<< labels >>
rlabel metal1 1241 723 1275 757 1 Y
port 1 n
rlabel metal1 205 575 239 609 1 A
port 2 n
rlabel metal1 353 649 387 683 1 B
port 3 n
rlabel metal1 723 723 757 757 1 C
port 4 n
rlabel metal1 55 1505 89 1539 1 VDD
port 5 n
rlabel metal1 55 13 89 47 1 VSS
port 6 n
<< end >>
