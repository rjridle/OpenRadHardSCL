* NGSPICE file created from 21T_ms_rhbd.ext - technology: sky130A

