* SPICE3 file created from DFFQNX1.ext - technology: sky130A

.subckt DFFQNX1 QN D CLK VDD GND
X0 VDD.t51 a_1845_1050.t5 a_147_187.t4 `��<*V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X1 QN.t3 a_277_1050.t7 VDD.t1 0�<*V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X2 VDD.t11 CLK.t0 a_277_1050.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X3 QN.t4 a_3303_411.t5 VDD.t33 VDD.t32 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X4 GND a_1845_1050.t6 a_2406_101.t0 GND sky130_fd_pr__nfet_01v8 ad=1.0746p pd=9.42u as=0p ps=0u w=0u l=0u
X5 VDD.t39 CLK.t1 a_147_187.t1 �ɨ� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X6 VDD.t19 a_599_989.t5 a_277_1050.t2 �ɨ� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X7 a_3303_411.t4 QN.t5 VDD.t9 �ɨ� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X8 QN a_3303_411.t6 a_3072_101.t0 GND sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=0p ps=0u w=0u l=0u
X9 VDD.t13 a_277_1050.t9 a_599_989.t2  �ɨ� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X10 VDD.t31 a_147_187.t6 a_3303_411.t2 VDD.t30 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X11 a_1845_1050.t1 a_147_187.t7 VDD.t29  �ɨ� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X12 GND a_147_187.t10 a_91_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X13 a_3303_411.t1 a_147_187.t8 VDD.t27 VDD.t26 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X14 VDD.t7 D.t1 a_599_989.t0  �ɨ� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X15 a_277_1050.t4 a_147_187.t9 VDD.t25 �ɨ� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X16 GND a_599_989.t8 a_1740_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X17 VDD.t47 a_599_989.t7 a_1845_1050.t3  �ɨ� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X18 a_277_1050.t5 CLK.t2 VDD.t37 �ɨ� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X19 a_147_187.t2 CLK.t3 VDD.t41  �ɨ� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X20 VDD.t15 a_277_1050.t10 QN.t2 �ɨ� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X21 GND QN.t6 a_3738_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X22 a_277_1050.t1 a_599_989.t9 VDD.t17  �ɨ� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X23 a_599_989.t1 a_277_1050.t11 VDD.t5 �ɨ� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X24 a_147_187.t3 a_1845_1050.t7 VDD.t49  �ɨ� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X25 GND a_277_1050.t12 a_1074_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X26 VDD.t3 a_3303_411.t7 QN.t1 �ɨ� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X27 VDD.t43 QN.t7 a_3303_411.t3  �ɨ� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X28 a_599_989.t3 D.t2 VDD.t35 �ɨ� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X29 GND a_277_1050.t8 a_3072_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X30 a_1845_1050.t2 a_599_989.t10 VDD.t45  �ɨ� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X31 VDD.t23 a_147_187.t11 a_1845_1050.t0 �ɨ� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X32 VDD.t21 a_147_187.t13 a_277_1050.t3  �ɨ� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
C0 VDD D 0.32fF
C1 CLK D 0.07fF
C2 QN VDD 2.20fF
C3 VDD CLK 1.85fF
R0 a_1845_1050.n3 a_1845_1050.t5 480.392
R1 a_1845_1050.n3 a_1845_1050.t7 403.272
R2 a_1845_1050.n4 a_1845_1050.t6 357.204
R3 a_1845_1050.n7 a_1845_1050.n5 312.103
R4 a_1845_1050.n4 a_1845_1050.n3 171.288
R5 a_1845_1050.n5 a_1845_1050.n2 159.999
R6 a_1845_1050.n2 a_1845_1050.n1 157.964
R7 a_1845_1050.n2 a_1845_1050.n0 91.706
R8 a_1845_1050.n7 a_1845_1050.n6 15.218
R9 a_1845_1050.n0 a_1845_1050.t0 14.282
R10 a_1845_1050.n0 a_1845_1050.t1 14.282
R11 a_1845_1050.n1 a_1845_1050.t3 14.282
R12 a_1845_1050.n1 a_1845_1050.t2 14.282
R13 a_1845_1050.n8 a_1845_1050.n7 12.014
R14 a_1845_1050.n5 a_1845_1050.n4 10.615
R15 a_147_187.n7 a_147_187.t13 512.525
R16 a_147_187.n5 a_147_187.t11 472.359
R17 a_147_187.n3 a_147_187.t6 472.359
R18 a_147_187.n8 a_147_187.t10 417.109
R19 a_147_187.n5 a_147_187.t7 384.527
R20 a_147_187.n3 a_147_187.t8 384.527
R21 a_147_187.n7 a_147_187.t9 371.139
R22 a_147_187.n6 a_147_187.t12 370.613
R23 a_147_187.n4 a_147_187.t5 370.613
R24 a_147_187.n13 a_147_187.n11 367.82
R25 a_147_187.n8 a_147_187.n7 179.837
R26 a_147_187.n2 a_147_187.n1 157.964
R27 a_147_187.n6 a_147_187.n5 127.096
R28 a_147_187.n4 a_147_187.n3 127.096
R29 a_147_187.n11 a_147_187.n2 104.282
R30 a_147_187.n2 a_147_187.n0 91.706
R31 a_147_187.n13 a_147_187.n12 15.218
R32 a_147_187.n0 a_147_187.t1 14.282
R33 a_147_187.n0 a_147_187.t2 14.282
R34 a_147_187.n1 a_147_187.t4 14.282
R35 a_147_187.n1 a_147_187.t3 14.282
R36 a_147_187.n14 a_147_187.n13 12.014
R37 a_147_187.n9 a_147_187.n8 11.134
R38 a_147_187.n10 a_147_187.n4 8.957
R39 a_147_187.n9 a_147_187.n6 4.65
R40 a_147_187.n11 a_147_187.n10 4.65
R41 a_147_187.n10 a_147_187.n9 2.947
R42 VDD.n297 VDD.n286 144.705
R43 VDD.n193 VDD.n186 144.705
R44 VDD.n354 VDD.n347 144.705
R45 VDD.n136 VDD.n129 144.705
R46 VDD.n79 VDD.n68 144.705
R47 VDD.n263 VDD.t19 143.754
R48 VDD.n322 VDD.t7 143.754
R49 VDD.n196 VDD.t23 143.754
R50 VDD.n139 VDD.t39 143.754
R51 VDD.n82 VDD.t3 143.754
R52 VDD.n24 VDD.t31 143.754
R53 VDD.n228 VDD.t25 135.17
R54 VDD.n300 VDD.t5 135.17
R55 VDD.n357 VDD.t45 135.17
R56 VDD.n161 VDD.t49 135.17
R57 VDD.n104 VDD.t1 135.17
R58 VDD.n46 VDD.t9 135.17
R59 VDD.n238 VDD.n237 129.472
R60 VDD.n254 VDD.n253 129.472
R61 VDD.n314 VDD.n313 129.472
R62 VDD.n371 VDD.n370 129.472
R63 VDD.n149 VDD.n148 129.472
R64 VDD.n92 VDD.n91 129.472
R65 VDD.n34 VDD.n33 129.472
R66 VDD.n64 VDD.n63 92.5
R67 VDD.n62 VDD.n61 92.5
R68 VDD.n60 VDD.n59 92.5
R69 VDD.n58 VDD.n57 92.5
R70 VDD.n66 VDD.n65 92.5
R71 VDD.n125 VDD.n124 92.5
R72 VDD.n123 VDD.n122 92.5
R73 VDD.n121 VDD.n120 92.5
R74 VDD.n119 VDD.n118 92.5
R75 VDD.n127 VDD.n126 92.5
R76 VDD.n182 VDD.n181 92.5
R77 VDD.n180 VDD.n179 92.5
R78 VDD.n178 VDD.n177 92.5
R79 VDD.n176 VDD.n175 92.5
R80 VDD.n184 VDD.n183 92.5
R81 VDD.n343 VDD.n342 92.5
R82 VDD.n341 VDD.n340 92.5
R83 VDD.n339 VDD.n338 92.5
R84 VDD.n337 VDD.n336 92.5
R85 VDD.n345 VDD.n344 92.5
R86 VDD.n282 VDD.n281 92.5
R87 VDD.n280 VDD.n279 92.5
R88 VDD.n278 VDD.n277 92.5
R89 VDD.n276 VDD.n275 92.5
R90 VDD.n284 VDD.n283 92.5
R91 VDD.n212 VDD.n211 92.5
R92 VDD.n210 VDD.n209 92.5
R93 VDD.n208 VDD.n207 92.5
R94 VDD.n206 VDD.n205 92.5
R95 VDD.n214 VDD.n213 92.5
R96 VDD.n14 VDD.n1 92.5
R97 VDD.n5 VDD.n4 92.5
R98 VDD.n7 VDD.n6 92.5
R99 VDD.n9 VDD.n8 92.5
R100 VDD.n11 VDD.n10 92.5
R101 VDD.n13 VDD.n12 92.5
R102 VDD.n21 VDD.n20 92.059
R103 VDD.n78 VDD.n77 92.059
R104 VDD.n135 VDD.n134 92.059
R105 VDD.n192 VDD.n191 92.059
R106 VDD.n353 VDD.n352 92.059
R107 VDD.n296 VDD.n295 92.059
R108 VDD.n220 VDD.n219 92.059
R109 VDD.n20 VDD.n16 67.194
R110 VDD.n20 VDD.n17 67.194
R111 VDD.n20 VDD.n18 67.194
R112 VDD.n20 VDD.n19 67.194
R113 VDD.n204 VDD.n203 44.141
R114 VDD.n335 VDD.n334 44.141
R115 VDD.n174 VDD.n173 44.141
R116 VDD.n117 VDD.n116 44.141
R117 VDD.n5 VDD.n3 44.141
R118 VDD.n334 VDD.n332 44.107
R119 VDD.n173 VDD.n171 44.107
R120 VDD.n116 VDD.n114 44.107
R121 VDD.n203 VDD.n201 44.107
R122 VDD.n3 VDD.n2 44.107
R123 VDD.n20 VDD.n15 41.052
R124 VDD.n72 VDD.n70 39.742
R125 VDD.n72 VDD.n71 39.742
R126 VDD.n74 VDD.n73 39.742
R127 VDD.n131 VDD.n130 39.742
R128 VDD.n188 VDD.n187 39.742
R129 VDD.n349 VDD.n348 39.742
R130 VDD.n216 VDD.n215 39.742
R131 VDD.n294 VDD.n291 39.742
R132 VDD.n294 VDD.n293 39.742
R133 VDD.n290 VDD.n289 39.742
R134 VDD.n116 VDD.n115 38
R135 VDD.n173 VDD.n172 38
R136 VDD.n334 VDD.n333 38
R137 VDD.n203 VDD.n202 38
R138 VDD.n332 VDD.n331 36.774
R139 VDD.n171 VDD.n170 36.774
R140 VDD.n114 VDD.n113 36.774
R141 VDD.n70 VDD.n69 36.774
R142 VDD.n293 VDD.n292 36.774
R143 VDD.n257 �ɨ� 35.8
R144 VDD.n233 �ɨ� 33.243
R145 VDD.n1 VDD.n0 30.923
R146 VDD.n77 VDD.n75 26.38
R147 VDD.n77 VDD.n74 26.38
R148 VDD.n77 VDD.n72 26.38
R149 VDD.n77 VDD.n76 26.38
R150 VDD.n134 VDD.n132 26.38
R151 VDD.n134 VDD.n131 26.38
R152 VDD.n134 VDD.n133 26.38
R153 VDD.n191 VDD.n189 26.38
R154 VDD.n191 VDD.n188 26.38
R155 VDD.n191 VDD.n190 26.38
R156 VDD.n352 VDD.n350 26.38
R157 VDD.n352 VDD.n349 26.38
R158 VDD.n352 VDD.n351 26.38
R159 VDD.n219 VDD.n217 26.38
R160 VDD.n219 VDD.n216 26.38
R161 VDD.n219 VDD.n218 26.38
R162 VDD.n295 VDD.n294 26.38
R163 VDD.n295 VDD.n290 26.38
R164 VDD.n295 VDD.n288 26.38
R165 VDD.n295 VDD.n287 26.38
R166 VDD.n222 VDD.n214 22.915
R167 VDD.n23 VDD.n14 22.915
R168 VDD.n29 VDD.t30 20.457
R169 VDD.n87 �ɨ� 20.457
R170 VDD.n144 �ɨ� 20.457
R171 VDD.n375 �ɨ� 20.457
R172 VDD.n318  �ɨ� 20.457
R173 VDD.n42 �ɨ� 17.9
R174 VDD.n100 0�<*V 17.9
R175 VDD.n157  �ɨ� 17.9
R176 VDD.n362  �ɨ� 17.9
R177 VDD.n305 �ɨ� 17.9
R178 VDD.n251  �ɨ� 15.343
R179 VDD.n214 VDD.n212 14.864
R180 VDD.n212 VDD.n210 14.864
R181 VDD.n210 VDD.n208 14.864
R182 VDD.n208 VDD.n206 14.864
R183 VDD.n206 VDD.n204 14.864
R184 VDD.n345 VDD.n343 14.864
R185 VDD.n343 VDD.n341 14.864
R186 VDD.n341 VDD.n339 14.864
R187 VDD.n339 VDD.n337 14.864
R188 VDD.n337 VDD.n335 14.864
R189 VDD.n184 VDD.n182 14.864
R190 VDD.n182 VDD.n180 14.864
R191 VDD.n180 VDD.n178 14.864
R192 VDD.n178 VDD.n176 14.864
R193 VDD.n176 VDD.n174 14.864
R194 VDD.n127 VDD.n125 14.864
R195 VDD.n125 VDD.n123 14.864
R196 VDD.n123 VDD.n121 14.864
R197 VDD.n121 VDD.n119 14.864
R198 VDD.n119 VDD.n117 14.864
R199 VDD.n66 VDD.n64 14.864
R200 VDD.n64 VDD.n62 14.864
R201 VDD.n62 VDD.n60 14.864
R202 VDD.n60 VDD.n58 14.864
R203 VDD.n58 VDD.n56 14.864
R204 VDD.n56 VDD.n55 14.864
R205 VDD.n284 VDD.n282 14.864
R206 VDD.n282 VDD.n280 14.864
R207 VDD.n280 VDD.n278 14.864
R208 VDD.n278 VDD.n276 14.864
R209 VDD.n276 VDD.n274 14.864
R210 VDD.n274 VDD.n273 14.864
R211 VDD.n14 VDD.n13 14.864
R212 VDD.n13 VDD.n11 14.864
R213 VDD.n11 VDD.n9 14.864
R214 VDD.n9 VDD.n7 14.864
R215 VDD.n7 VDD.n5 14.864
R216 VDD.n80 VDD.n67 14.864
R217 VDD.n137 VDD.n128 14.864
R218 VDD.n194 VDD.n185 14.864
R219 VDD.n355 VDD.n346 14.864
R220 VDD.n298 VDD.n285 14.864
R221 VDD.n237 VDD.t37 14.282
R222 VDD.n237 VDD.t21 14.282
R223 VDD.n253 VDD.t17 14.282
R224 VDD.n253 VDD.t11 14.282
R225 VDD.n313 VDD.t35 14.282
R226 VDD.n313 VDD.t13 14.282
R227 VDD.n370 VDD.t29 14.282
R228 VDD.n370 VDD.t47 14.282
R229 VDD.n148 VDD.t41 14.282
R230 VDD.n148 VDD.t51 14.282
R231 VDD.n91 VDD.t33 14.282
R232 VDD.n91 VDD.t15 14.282
R233 VDD.n33 VDD.t27 14.282
R234 VDD.n33 VDD.t43 14.282
R235 VDD.n239  �ɨ� 12.786
R236 VDD.n36 VDD.n34 9.083
R237 VDD.n94 VDD.n92 9.083
R238 VDD.n151 VDD.n149 9.083
R239 VDD.n373 VDD.n371 9.083
R240 VDD.n316 VDD.n314 9.083
R241 VDD.n23 VDD.n22 8.855
R242 VDD.n22 VDD.n21 8.855
R243 VDD.n27 VDD.n26 8.855
R244 VDD.n26 VDD.n25 8.855
R245 VDD.n31 VDD.n30 8.855
R246 VDD.n30 VDD.n29 8.855
R247 VDD.n36 VDD.n35 8.855
R248 VDD.n35 VDD.t26 8.855
R249 VDD.n40 VDD.n39 8.855
R250 VDD.n39 VDD.n38 8.855
R251 VDD.n44 VDD.n43 8.855
R252 VDD.n43 VDD.n42 8.855
R253 VDD.n49 VDD.n48 8.855
R254 VDD.n48 VDD.n47 8.855
R255 VDD.n53 VDD.n52 8.855
R256 VDD.n52 VDD.n51 8.855
R257 VDD.n80 VDD.n79 8.855
R258 VDD.n79 VDD.n78 8.855
R259 VDD.n85 VDD.n84 8.855
R260 VDD.n84 VDD.n83 8.855
R261 VDD.n89 VDD.n88 8.855
R262 VDD.n88 VDD.n87 8.855
R263 VDD.n94 VDD.n93 8.855
R264 VDD.n93 VDD.t32 8.855
R265 VDD.n98 VDD.n97 8.855
R266 VDD.n97 VDD.n96 8.855
R267 VDD.n102 VDD.n101 8.855
R268 VDD.n101 VDD.n100 8.855
R269 VDD.n107 VDD.n106 8.855
R270 VDD.n106 VDD.n105 8.855
R271 VDD.n111 VDD.n110 8.855
R272 VDD.n110 VDD.n109 8.855
R273 VDD.n137 VDD.n136 8.855
R274 VDD.n136 VDD.n135 8.855
R275 VDD.n142 VDD.n141 8.855
R276 VDD.n141 VDD.n140 8.855
R277 VDD.n146 VDD.n145 8.855
R278 VDD.n145 VDD.n144 8.855
R279 VDD.n151 VDD.n150 8.855
R280 VDD.n150  �ɨ� 8.855
R281 VDD.n155 VDD.n154 8.855
R282 VDD.n154 VDD.n153 8.855
R283 VDD.n159 VDD.n158 8.855
R284 VDD.n158 VDD.n157 8.855
R285 VDD.n164 VDD.n163 8.855
R286 VDD.n163 VDD.n162 8.855
R287 VDD.n168 VDD.n167 8.855
R288 VDD.n167 VDD.n166 8.855
R289 VDD.n194 VDD.n193 8.855
R290 VDD.n193 VDD.n192 8.855
R291 VDD.n199 VDD.n198 8.855
R292 VDD.n198 VDD.n197 8.855
R293 VDD.n377 VDD.n376 8.855
R294 VDD.n376 VDD.n375 8.855
R295 VDD.n373 VDD.n372 8.855
R296 VDD.n372  �ɨ� 8.855
R297 VDD.n368 VDD.n367 8.855
R298 VDD.n367 VDD.n366 8.855
R299 VDD.n364 VDD.n363 8.855
R300 VDD.n363 VDD.n362 8.855
R301 VDD.n360 VDD.n359 8.855
R302 VDD.n359 VDD.n358 8.855
R303 VDD.n355 VDD.n354 8.855
R304 VDD.n354 VDD.n353 8.855
R305 VDD.n329 VDD.n328 8.855
R306 VDD.n328 VDD.n327 8.855
R307 VDD.n325 VDD.n324 8.855
R308 VDD.n324 VDD.n323 8.855
R309 VDD.n320 VDD.n319 8.855
R310 VDD.n319 VDD.n318 8.855
R311 VDD.n316 VDD.n315 8.855
R312 VDD.n315 �ɨ� 8.855
R313 VDD.n311 VDD.n310 8.855
R314 VDD.n310 VDD.n309 8.855
R315 VDD.n307 VDD.n306 8.855
R316 VDD.n306 VDD.n305 8.855
R317 VDD.n303 VDD.n302 8.855
R318 VDD.n302 VDD.n301 8.855
R319 VDD.n298 VDD.n297 8.855
R320 VDD.n297 VDD.n296 8.855
R321 VDD.n271 VDD.n270 8.855
R322 VDD.n270 VDD.n269 8.855
R323 VDD.n267 VDD.n266 8.855
R324 VDD.n266 VDD.n265 8.855
R325 VDD.n263 VDD.n262 8.855
R326 VDD.n262 VDD.n261 8.855
R327 VDD.n259 VDD.n258 8.855
R328 VDD.n258 VDD.n257 8.855
R329 VDD.n255 VDD.n252 8.855
R330 VDD.n252 VDD.n251 8.855
R331 VDD.n249 VDD.n248 8.855
R332 VDD.n248 VDD.n247 8.855
R333 VDD.n245 VDD.n244 8.855
R334 VDD.n244 VDD.n243 8.855
R335 VDD.n241 VDD.n240 8.855
R336 VDD.n240 VDD.n239 8.855
R337 VDD.n235 VDD.n234 8.855
R338 VDD.n234 VDD.n233 8.855
R339 VDD.n231 VDD.n230 8.855
R340 VDD.n230 VDD.n229 8.855
R341 VDD.n226 VDD.n225 8.855
R342 VDD.n225 VDD.n224 8.855
R343 VDD.n222 VDD.n221 8.855
R344 VDD.n221 VDD.n220 8.855
R345 VDD.n346 VDD.n345 8.051
R346 VDD.n185 VDD.n184 8.051
R347 VDD.n128 VDD.n127 8.051
R348 VDD.n67 VDD.n66 8.051
R349 VDD.n285 VDD.n284 8.051
R350 VDD.n243 �ɨ� 7.671
R351 VDD.n241 VDD.n238 7.019
R352 VDD.n255 VDD.n254 6.606
R353 VDD.n247 �0=*V 5.114
R354 VDD.n32 VDD.n31 4.65
R355 VDD.n37 VDD.n36 4.65
R356 VDD.n41 VDD.n40 4.65
R357 VDD.n45 VDD.n44 4.65
R358 VDD.n50 VDD.n49 4.65
R359 VDD.n54 VDD.n53 4.65
R360 VDD.n81 VDD.n80 4.65
R361 VDD.n86 VDD.n85 4.65
R362 VDD.n90 VDD.n89 4.65
R363 VDD.n95 VDD.n94 4.65
R364 VDD.n99 VDD.n98 4.65
R365 VDD.n103 VDD.n102 4.65
R366 VDD.n108 VDD.n107 4.65
R367 VDD.n112 VDD.n111 4.65
R368 VDD.n138 VDD.n137 4.65
R369 VDD.n143 VDD.n142 4.65
R370 VDD.n147 VDD.n146 4.65
R371 VDD.n152 VDD.n151 4.65
R372 VDD.n156 VDD.n155 4.65
R373 VDD.n160 VDD.n159 4.65
R374 VDD.n165 VDD.n164 4.65
R375 VDD.n169 VDD.n168 4.65
R376 VDD.n195 VDD.n194 4.65
R377 VDD.n200 VDD.n199 4.65
R378 VDD.n378 VDD.n377 4.65
R379 VDD.n374 VDD.n373 4.65
R380 VDD.n369 VDD.n368 4.65
R381 VDD.n365 VDD.n364 4.65
R382 VDD.n361 VDD.n360 4.65
R383 VDD.n356 VDD.n355 4.65
R384 VDD.n330 VDD.n329 4.65
R385 VDD.n326 VDD.n325 4.65
R386 VDD.n321 VDD.n320 4.65
R387 VDD.n317 VDD.n316 4.65
R388 VDD.n312 VDD.n311 4.65
R389 VDD.n308 VDD.n307 4.65
R390 VDD.n304 VDD.n303 4.65
R391 VDD.n299 VDD.n298 4.65
R392 VDD.n272 VDD.n271 4.65
R393 VDD.n268 VDD.n267 4.65
R394 VDD.n264 VDD.n263 4.65
R395 VDD.n260 VDD.n259 4.65
R396 VDD.n256 VDD.n255 4.65
R397 VDD.n250 VDD.n249 4.65
R398 VDD.n246 VDD.n245 4.65
R399 VDD.n242 VDD.n241 4.65
R400 VDD.n236 VDD.n235 4.65
R401 VDD.n232 VDD.n231 4.65
R402 VDD.n227 VDD.n226 4.65
R403 VDD.n223 VDD.n222 4.65
R404 VDD.n28 VDD.n23 2.933
R405 VDD.n49 VDD.n46 2.89
R406 VDD.n107 VDD.n104 2.89
R407 VDD.n164 VDD.n161 2.89
R408 VDD.n360 VDD.n357 2.89
R409 VDD.n303 VDD.n300 2.89
R410 VDD.n28 VDD.n27 2.844
R411 VDD.n38  �ɨ� 2.557
R412 VDD.n96 �ɨ� 2.557
R413 VDD.n153 `��<*V 2.557
R414 VDD.n366  �ɨ� 2.557
R415 VDD.n309  �ɨ� 2.557
R416 VDD.n27 VDD.n24 2.477
R417 VDD.n85 VDD.n82 2.477
R418 VDD.n142 VDD.n139 2.477
R419 VDD.n199 VDD.n196 2.477
R420 VDD.n325 VDD.n322 2.477
R421 VDD.n32 VDD.n28 1.063
R422 VDD.n231 VDD.n228 0.412
R423 VDD.n81 VDD.n54 0.29
R424 VDD.n138 VDD.n112 0.29
R425 VDD.n195 VDD.n169 0.29
R426 VDD.n356 VDD.n330 0.29
R427 VDD.n299 VDD.n272 0.29
R428 VDD.n223 VDD 0.207
R429 VDD.n250 VDD.n246 0.197
R430 VDD.n41 VDD.n37 0.181
R431 VDD.n99 VDD.n95 0.181
R432 VDD.n156 VDD.n152 0.181
R433 VDD.n374 VDD.n369 0.181
R434 VDD.n317 VDD.n312 0.181
R435 VDD.n37 VDD.n32 0.145
R436 VDD.n45 VDD.n41 0.145
R437 VDD.n50 VDD.n45 0.145
R438 VDD.n54 VDD.n50 0.145
R439 VDD.n86 VDD.n81 0.145
R440 VDD.n90 VDD.n86 0.145
R441 VDD.n95 VDD.n90 0.145
R442 VDD.n103 VDD.n99 0.145
R443 VDD.n108 VDD.n103 0.145
R444 VDD.n112 VDD.n108 0.145
R445 VDD.n143 VDD.n138 0.145
R446 VDD.n147 VDD.n143 0.145
R447 VDD.n152 VDD.n147 0.145
R448 VDD.n160 VDD.n156 0.145
R449 VDD.n165 VDD.n160 0.145
R450 VDD.n169 VDD.n165 0.145
R451 VDD.n200 VDD.n195 0.145
R452 VDD.n378 VDD.n374 0.145
R453 VDD.n369 VDD.n365 0.145
R454 VDD.n365 VDD.n361 0.145
R455 VDD.n361 VDD.n356 0.145
R456 VDD.n330 VDD.n326 0.145
R457 VDD.n326 VDD.n321 0.145
R458 VDD.n321 VDD.n317 0.145
R459 VDD.n312 VDD.n308 0.145
R460 VDD.n308 VDD.n304 0.145
R461 VDD.n304 VDD.n299 0.145
R462 VDD.n272 VDD.n268 0.145
R463 VDD.n268 VDD.n264 0.145
R464 VDD.n264 VDD.n260 0.145
R465 VDD.n260 VDD.n256 0.145
R466 VDD.n256 VDD.n250 0.145
R467 VDD.n246 VDD.n242 0.145
R468 VDD.n242 VDD.n236 0.145
R469 VDD.n236 VDD.n232 0.145
R470 VDD.n232 VDD.n227 0.145
R471 VDD.n227 VDD.n223 0.145
R472 VDD VDD.n378 0.137
R473 VDD VDD.n200 0.008
R474 a_277_1050.n4 a_277_1050.t9 480.392
R475 a_277_1050.n2 a_277_1050.t10 480.392
R476 a_277_1050.n4 a_277_1050.t11 403.272
R477 a_277_1050.n2 a_277_1050.t7 403.272
R478 a_277_1050.n5 a_277_1050.t12 385.063
R479 a_277_1050.n3 a_277_1050.t8 385.063
R480 a_277_1050.n8 a_277_1050.n7 357.814
R481 a_277_1050.n11 a_277_1050.n10 161.352
R482 a_277_1050.n9 a_277_1050.n8 151.34
R483 a_277_1050.n5 a_277_1050.n4 143.429
R484 a_277_1050.n3 a_277_1050.n2 143.429
R485 a_277_1050.n9 a_277_1050.n1 95.095
R486 a_277_1050.n10 a_277_1050.n0 95.095
R487 a_277_1050.n10 a_277_1050.n9 66.258
R488 a_277_1050.n1 a_277_1050.t2 14.282
R489 a_277_1050.n1 a_277_1050.t1 14.282
R490 a_277_1050.n0 a_277_1050.t0 14.282
R491 a_277_1050.n0 a_277_1050.t5 14.282
R492 a_277_1050.n11 a_277_1050.t3 14.282
R493 a_277_1050.t4 a_277_1050.n11 14.282
R494 a_277_1050.n6 a_277_1050.n3 11.95
R495 a_277_1050.n8 a_277_1050.n6 5.965
R496 a_277_1050.n6 a_277_1050.n5 4.65
R497 QN.n0 QN.t7 480.392
R498 QN.n0 QN.t5 403.272
R499 QN.n1 QN.t6 357.204
R500 QN.n9 QN.n8 305.581
R501 QN.n1 QN.n0 171.288
R502 QN.n9 QN.n4 159.999
R503 QN.n4 QN.n3 157.964
R504 QN.n4 QN.n2 91.706
R505 QN.n8 QN.n7 30
R506 QN.n6 QN.n5 24.383
R507 QN.n8 QN.n6 23.684
R508 QN.n2 QN.t1 14.282
R509 QN.n2 QN.t4 14.282
R510 QN.n3 QN.t2 14.282
R511 QN.n3 QN.t3 14.282
R512 QN QN.n9 5.919
R513 QN.n10 QN.n1 4.65
R514 QN.n10 QN 0.046
R515 a_3072_101.t0 a_3072_101.n1 93.333
R516 a_3072_101.n4 a_3072_101.n2 79.092
R517 a_3072_101.t0 a_3072_101.n0 8.137
R518 a_3072_101.n4 a_3072_101.n3 4.614
R519 a_3072_101.t0 a_3072_101.n4 0.111
R520 GND.n144 GND.n143 237.558
R521 GND.n96 GND.n95 237.558
R522 GND.n177 GND.n176 237.558
R523 GND.n63 GND.n62 237.558
R524 GND.n31 GND.n30 237.558
R525 GND.n28 GND.n27 210.82
R526 GND.n146 GND.n145 210.82
R527 GND.n179 GND.n178 210.82
R528 GND.n93 GND.n92 210.82
R529 GND.n60 GND.n59 210.82
R530 GND.n49 GND.n48 166.605
R531 GND.n189 GND.n188 166.605
R532 GND.n113 GND.n112 152.358
R533 GND.n17 GND.n16 151.605
R534 GND.n82 GND.n81 151.605
R535 GND.n157 GND.n156 151.605
R536 GND.n16 GND.n15 28.421
R537 GND.n81 GND.n80 28.421
R538 GND.n156 GND.n155 28.421
R539 GND.n112 GND.n111 28.421
R540 GND.n16 GND.n14 25.263
R541 GND.n81 GND.n79 25.263
R542 GND.n156 GND.n154 25.263
R543 GND.n112 GND.n110 25.263
R544 GND.n14 GND.n13 24.383
R545 GND.n79 GND.n78 24.383
R546 GND.n154 GND.n153 24.383
R547 GND.n110 GND.n109 24.383
R548 GND.n48 GND.n46 23.03
R549 GND.n188 GND.n186 23.03
R550 GND.n29 GND.n28 18.953
R551 GND.n147 GND.n146 18.953
R552 GND.n180 GND.n179 18.953
R553 GND.n94 GND.n93 18.953
R554 GND.n61 GND.n60 18.953
R555 GND.n32 GND.n29 14.864
R556 GND.n64 GND.n61 14.864
R557 GND.n97 GND.n94 14.864
R558 GND.n181 GND.n180 14.864
R559 GND.n148 GND.n147 14.864
R560 GND.n106 GND.n105 9.154
R561 GND.n114 GND.n108 9.154
R562 GND.n117 GND.n116 9.154
R563 GND.n120 GND.n119 9.154
R564 GND.n123 GND.n122 9.154
R565 GND.n126 GND.n125 9.154
R566 GND.n129 GND.n128 9.154
R567 GND.n132 GND.n131 9.154
R568 GND.n135 GND.n134 9.154
R569 GND.n138 GND.n137 9.154
R570 GND.n141 GND.n140 9.154
R571 GND.n148 GND.n144 9.154
R572 GND.n151 GND.n150 9.154
R573 GND.n159 GND.n158 9.154
R574 GND.n162 GND.n161 9.154
R575 GND.n165 GND.n164 9.154
R576 GND.n168 GND.n167 9.154
R577 GND.n171 GND.n170 9.154
R578 GND.n174 GND.n173 9.154
R579 GND.n181 GND.n177 9.154
R580 GND.n184 GND.n183 9.154
R581 GND.n191 GND.n190 9.154
R582 GND.n194 GND.n193 9.154
R583 GND.n197 GND.n196 9.154
R584 GND.n200 GND.n199 9.154
R585 GND.n100 GND.n99 9.154
R586 GND.n97 GND.n96 9.154
R587 GND.n90 GND.n89 9.154
R588 GND.n87 GND.n86 9.154
R589 GND.n84 GND.n83 9.154
R590 GND.n76 GND.n75 9.154
R591 GND.n73 GND.n72 9.154
R592 GND.n70 GND.n69 9.154
R593 GND.n67 GND.n66 9.154
R594 GND.n64 GND.n63 9.154
R595 GND.n57 GND.n56 9.154
R596 GND.n54 GND.n53 9.154
R597 GND.n51 GND.n50 9.154
R598 GND.n44 GND.n43 9.154
R599 GND.n41 GND.n40 9.154
R600 GND.n38 GND.n37 9.154
R601 GND.n35 GND.n34 9.154
R602 GND.n32 GND.n31 9.154
R603 GND.n25 GND.n24 9.154
R604 GND.n22 GND.n21 9.154
R605 GND.n19 GND.n18 9.154
R606 GND.n11 GND.n10 9.154
R607 GND.n8 GND.n7 9.154
R608 GND.n5 GND.n4 9.154
R609 GND.n2 GND.n1 9.154
R610 GND.n48 GND.n47 8.128
R611 GND.n188 GND.n187 8.128
R612 GND.n104 GND.n103 4.65
R613 GND.n6 GND.n5 4.65
R614 GND.n9 GND.n8 4.65
R615 GND.n12 GND.n11 4.65
R616 GND.n20 GND.n19 4.65
R617 GND.n23 GND.n22 4.65
R618 GND.n26 GND.n25 4.65
R619 GND.n33 GND.n32 4.65
R620 GND.n36 GND.n35 4.65
R621 GND.n39 GND.n38 4.65
R622 GND.n42 GND.n41 4.65
R623 GND.n45 GND.n44 4.65
R624 GND.n52 GND.n51 4.65
R625 GND.n55 GND.n54 4.65
R626 GND.n58 GND.n57 4.65
R627 GND.n65 GND.n64 4.65
R628 GND.n68 GND.n67 4.65
R629 GND.n71 GND.n70 4.65
R630 GND.n74 GND.n73 4.65
R631 GND.n77 GND.n76 4.65
R632 GND.n85 GND.n84 4.65
R633 GND.n88 GND.n87 4.65
R634 GND.n91 GND.n90 4.65
R635 GND.n98 GND.n97 4.65
R636 GND.n101 GND.n100 4.65
R637 GND.n201 GND.n200 4.65
R638 GND.n198 GND.n197 4.65
R639 GND.n195 GND.n194 4.65
R640 GND.n192 GND.n191 4.65
R641 GND.n185 GND.n184 4.65
R642 GND.n182 GND.n181 4.65
R643 GND.n175 GND.n174 4.65
R644 GND.n172 GND.n171 4.65
R645 GND.n169 GND.n168 4.65
R646 GND.n166 GND.n165 4.65
R647 GND.n163 GND.n162 4.65
R648 GND.n160 GND.n159 4.65
R649 GND.n152 GND.n151 4.65
R650 GND.n149 GND.n148 4.65
R651 GND.n142 GND.n141 4.65
R652 GND.n139 GND.n138 4.65
R653 GND.n136 GND.n135 4.65
R654 GND.n133 GND.n132 4.65
R655 GND.n130 GND.n129 4.65
R656 GND.n127 GND.n126 4.65
R657 GND.n124 GND.n123 4.65
R658 GND.n121 GND.n120 4.65
R659 GND.n118 GND.n117 4.65
R660 GND.n115 GND.n114 4.65
R661 GND.n107 GND.n106 4.65
R662 GND.n19 GND.n17 4.129
R663 GND.n51 GND.n49 4.129
R664 GND.n84 GND.n82 4.129
R665 GND.n191 GND.n189 4.129
R666 GND.n159 GND.n157 4.129
R667 GND.n3 GND.n0 3.407
R668 GND.n3 GND.n2 2.844
R669 GND.n6 GND.n3 1.063
R670 GND.n103 GND.n102 0.474
R671 GND.n33 GND.n26 0.29
R672 GND.n65 GND.n58 0.29
R673 GND.n98 GND.n91 0.29
R674 GND.n182 GND.n175 0.29
R675 GND.n149 GND.n142 0.29
R676 GND.n104 GND 0.207
R677 GND.n114 GND.n113 0.206
R678 GND.n127 GND.n124 0.197
R679 GND.n12 GND.n9 0.181
R680 GND.n45 GND.n42 0.181
R681 GND.n77 GND.n74 0.181
R682 GND.n198 GND.n195 0.181
R683 GND.n166 GND.n163 0.181
R684 GND.n9 GND.n6 0.145
R685 GND.n20 GND.n12 0.145
R686 GND.n23 GND.n20 0.145
R687 GND.n26 GND.n23 0.145
R688 GND.n36 GND.n33 0.145
R689 GND.n39 GND.n36 0.145
R690 GND.n42 GND.n39 0.145
R691 GND.n52 GND.n45 0.145
R692 GND.n55 GND.n52 0.145
R693 GND.n58 GND.n55 0.145
R694 GND.n68 GND.n65 0.145
R695 GND.n71 GND.n68 0.145
R696 GND.n74 GND.n71 0.145
R697 GND.n85 GND.n77 0.145
R698 GND.n88 GND.n85 0.145
R699 GND.n91 GND.n88 0.145
R700 GND.n101 GND.n98 0.145
R701 GND.n201 GND.n198 0.145
R702 GND.n195 GND.n192 0.145
R703 GND.n192 GND.n185 0.145
R704 GND.n185 GND.n182 0.145
R705 GND.n175 GND.n172 0.145
R706 GND.n172 GND.n169 0.145
R707 GND.n169 GND.n166 0.145
R708 GND.n163 GND.n160 0.145
R709 GND.n160 GND.n152 0.145
R710 GND.n152 GND.n149 0.145
R711 GND.n142 GND.n139 0.145
R712 GND.n139 GND.n136 0.145
R713 GND.n136 GND.n133 0.145
R714 GND.n133 GND.n130 0.145
R715 GND.n130 GND.n127 0.145
R716 GND.n124 GND.n121 0.145
R717 GND.n121 GND.n118 0.145
R718 GND.n118 GND.n115 0.145
R719 GND.n115 GND.n107 0.145
R720 GND.n107 GND.n104 0.145
R721 GND GND.n201 0.137
R722 GND GND.n101 0.008
R723 CLK.n0 CLK.t1 472.359
R724 CLK.n2 CLK.t0 459.505
R725 CLK.n3 CLK.t4 399.181
R726 CLK.n1 CLK.t5 398.558
R727 CLK.n2 CLK.t2 384.527
R728 CLK.n0 CLK.t3 384.527
R729 CLK.n3 CLK.n2 33.832
R730 CLK.n1 CLK.n0 32.394
R731 CLK.n4 CLK.n1 9.575
R732 CLK.n4 CLK.n3 2.079
R733 CLK.n4 CLK 0.046
R734 a_3303_411.n0 a_3303_411.t7 472.359
R735 a_3303_411.n0 a_3303_411.t5 384.527
R736 a_3303_411.n1 a_3303_411.t6 342.755
R737 a_3303_411.n6 a_3303_411.n5 333.44
R738 a_3303_411.n8 a_3303_411.n7 157.964
R739 a_3303_411.n1 a_3303_411.n0 154.955
R740 a_3303_411.n8 a_3303_411.n6 132.141
R741 a_3303_411.n9 a_3303_411.n8 91.705
R742 a_3303_411.n5 a_3303_411.n4 30
R743 a_3303_411.n3 a_3303_411.n2 24.383
R744 a_3303_411.n5 a_3303_411.n3 23.684
R745 a_3303_411.n7 a_3303_411.t3 14.282
R746 a_3303_411.n7 a_3303_411.t4 14.282
R747 a_3303_411.t2 a_3303_411.n9 14.282
R748 a_3303_411.n9 a_3303_411.t1 14.282
R749 a_3303_411.n6 a_3303_411.n1 12.247
R750 a_3738_101.n3 a_3738_101.n1 42.788
R751 a_3738_101.t0 a_3738_101.n0 8.137
R752 a_3738_101.n3 a_3738_101.n2 4.665
R753 a_3738_101.t0 a_3738_101.n3 0.06
R754 a_599_989.n1 a_599_989.t7 480.392
R755 a_599_989.n3 a_599_989.t9 454.685
R756 a_599_989.n3 a_599_989.t5 428.979
R757 a_599_989.n1 a_599_989.t10 403.272
R758 a_599_989.n2 a_599_989.t8 357.204
R759 a_599_989.n7 a_599_989.n6 327.32
R760 a_599_989.n4 a_599_989.t6 311.683
R761 a_599_989.n4 a_599_989.n3 171.288
R762 a_599_989.n2 a_599_989.n1 171.288
R763 a_599_989.n8 a_599_989.n7 159.999
R764 a_599_989.n9 a_599_989.n8 157.963
R765 a_599_989.n8 a_599_989.n0 91.706
R766 a_599_989.n0 a_599_989.t0 14.282
R767 a_599_989.n0 a_599_989.t3 14.282
R768 a_599_989.t2 a_599_989.n9 14.282
R769 a_599_989.n9 a_599_989.t1 14.282
R770 a_599_989.n5 a_599_989.n4 7.597
R771 a_599_989.n5 a_599_989.n2 5.965
R772 a_599_989.n7 a_599_989.n5 4.65
R773 D.n0 D.t1 472.359
R774 D.n0 D.t2 384.527
R775 D.n1 D.t0 219.801
R776 D.n1 D.n0 210.673
R777 D.n2 D.n1 4.65
R778 D.n2 D 0.046
R779 a_1074_101.n11 a_1074_101.n10 68.43
R780 a_1074_101.n3 a_1074_101.n2 62.817
R781 a_1074_101.n7 a_1074_101.n6 38.626
R782 a_1074_101.n6 a_1074_101.n5 35.955
R783 a_1074_101.n3 a_1074_101.n1 26.202
R784 a_1074_101.t0 a_1074_101.n3 19.737
R785 a_1074_101.t1 a_1074_101.n8 8.137
R786 a_1074_101.t0 a_1074_101.n4 7.273
R787 a_1074_101.t0 a_1074_101.n0 6.109
R788 a_1074_101.t1 a_1074_101.n7 4.864
R789 a_1074_101.t0 a_1074_101.n12 2.074
R790 a_1074_101.n12 a_1074_101.t1 0.937
R791 a_1074_101.t1 a_1074_101.n11 0.763
R792 a_1074_101.n11 a_1074_101.n9 0.185
R793 a_372_210.n9 a_372_210.n7 171.558
R794 a_372_210.t0 a_372_210.n9 75.765
R795 a_372_210.n3 a_372_210.n1 74.827
R796 a_372_210.n3 a_372_210.n2 27.476
R797 a_372_210.n7 a_372_210.n6 27.2
R798 a_372_210.n5 a_372_210.n4 23.498
R799 a_372_210.n7 a_372_210.n5 22.4
R800 a_372_210.t0 a_372_210.n11 20.241
R801 a_372_210.t0 a_372_210.n3 13.984
R802 a_372_210.n11 a_372_210.n10 13.494
R803 a_372_210.t0 a_372_210.n0 8.137
R804 a_372_210.n9 a_372_210.n8 1.505
R805 a_2406_101.n3 a_2406_101.n1 42.788
R806 a_2406_101.t0 a_2406_101.n0 8.137
R807 a_2406_101.n3 a_2406_101.n2 4.665
R808 a_2406_101.t0 a_2406_101.n3 0.06
R809 a_91_103.t0 a_91_103.n7 59.616
R810 a_91_103.n4 a_91_103.n2 54.496
R811 a_91_103.n4 a_91_103.n3 54.496
R812 a_91_103.n1 a_91_103.n0 24.679
R813 a_91_103.t0 a_91_103.n1 7.505
R814 a_91_103.n6 a_91_103.n5 2.455
R815 a_91_103.n6 a_91_103.n4 0.636
R816 a_91_103.t0 a_91_103.n6 0.246
R817 a_1740_101.n11 a_1740_101.n10 68.43
R818 a_1740_101.n3 a_1740_101.n2 62.817
R819 a_1740_101.n7 a_1740_101.n6 38.626
R820 a_1740_101.n6 a_1740_101.n5 35.955
R821 a_1740_101.n3 a_1740_101.n1 26.202
R822 a_1740_101.t0 a_1740_101.n3 19.737
R823 a_1740_101.t1 a_1740_101.n8 8.137
R824 a_1740_101.t0 a_1740_101.n4 7.273
R825 a_1740_101.t0 a_1740_101.n0 6.109
R826 a_1740_101.t1 a_1740_101.n7 4.864
R827 a_1740_101.t0 a_1740_101.n12 2.074
R828 a_1740_101.n12 a_1740_101.t1 0.937
R829 a_1740_101.t1 a_1740_101.n11 0.763
R830 a_1740_101.n11 a_1740_101.n9 0.185
C4 VDD GND 6.94fF
C5 a_1740_101.n0 GND 0.02fF
C6 a_1740_101.n1 GND 0.09fF
C7 a_1740_101.n2 GND 0.08fF
C8 a_1740_101.n3 GND 0.03fF
C9 a_1740_101.n4 GND 0.01fF
C10 a_1740_101.n5 GND 0.04fF
C11 a_1740_101.n6 GND 0.04fF
C12 a_1740_101.n7 GND 0.02fF
C13 a_1740_101.n8 GND 0.05fF
C14 a_1740_101.n9 GND 0.15fF
C15 a_1740_101.n10 GND 0.08fF
C16 a_1740_101.n11 GND 0.08fF
C17 a_1740_101.t1 GND 0.23fF
C18 a_1740_101.n12 GND 0.01fF
C19 a_91_103.n0 GND 0.08fF
C20 a_91_103.n1 GND 0.07fF
C21 a_91_103.n2 GND 0.04fF
C22 a_91_103.n3 GND 0.06fF
C23 a_91_103.n4 GND 0.03fF
C24 a_91_103.n5 GND 0.03fF
C25 a_91_103.n7 GND 0.08fF
C26 a_2406_101.n0 GND 0.05fF
C27 a_2406_101.n1 GND 0.12fF
C28 a_2406_101.n2 GND 0.04fF
C29 a_2406_101.n3 GND 0.17fF
C30 a_372_210.n0 GND 0.07fF
C31 a_372_210.n1 GND 0.09fF
C32 a_372_210.n2 GND 0.12fF
C33 a_372_210.n3 GND 0.08fF
C34 a_372_210.n4 GND 0.02fF
C35 a_372_210.n5 GND 0.03fF
C36 a_372_210.n6 GND 0.02fF
C37 a_372_210.n7 GND 0.03fF
C38 a_372_210.n8 GND 0.02fF
C39 a_372_210.n9 GND 0.13fF
C40 a_372_210.n10 GND 0.08fF
C41 a_372_210.n11 GND 0.02fF
C42 a_372_210.t0 GND 0.31fF
C43 a_1074_101.n0 GND 0.02fF
C44 a_1074_101.n1 GND 0.09fF
C45 a_1074_101.n2 GND 0.08fF
C46 a_1074_101.n3 GND 0.03fF
C47 a_1074_101.n4 GND 0.01fF
C48 a_1074_101.n5 GND 0.04fF
C49 a_1074_101.n6 GND 0.04fF
C50 a_1074_101.n7 GND 0.02fF
C51 a_1074_101.n8 GND 0.05fF
C52 a_1074_101.n9 GND 0.15fF
C53 a_1074_101.n10 GND 0.08fF
C54 a_1074_101.n11 GND 0.08fF
C55 a_1074_101.t1 GND 0.23fF
C56 a_1074_101.n12 GND 0.01fF
C57 a_599_989.n0 GND 0.40fF
C58 a_599_989.n1 GND 0.34fF
C59 a_599_989.n2 GND 0.49fF
C60 a_599_989.n3 GND 0.34fF
C61 a_599_989.t6 GND 0.54fF
C62 a_599_989.n4 GND 0.57fF
C63 a_599_989.n5 GND 0.88fF
C64 a_599_989.n6 GND 0.34fF
C65 a_599_989.n7 GND 0.53fF
C66 a_599_989.n8 GND 0.60fF
C67 a_599_989.n9 GND 0.51fF
C68 a_3738_101.n0 GND 0.05fF
C69 a_3738_101.n1 GND 0.12fF
C70 a_3738_101.n2 GND 0.04fF
C71 a_3738_101.n3 GND 0.16fF
C72 a_3303_411.n0 GND 0.30fF
C73 a_3303_411.n1 GND 0.77fF
C74 a_3303_411.n2 GND 0.04fF
C75 a_3303_411.n3 GND 0.05fF
C76 a_3303_411.n4 GND 0.03fF
C77 a_3303_411.n5 GND 0.26fF
C78 a_3303_411.n6 GND 0.87fF
C79 a_3303_411.n7 GND 0.50fF
C80 a_3303_411.n8 GND 0.56fF
C81 a_3303_411.n9 GND 0.39fF
C82 a_3072_101.n0 GND 0.05fF
C83 a_3072_101.n1 GND 0.02fF
C84 a_3072_101.n2 GND 0.12fF
C85 a_3072_101.n3 GND 0.04fF
C86 a_3072_101.n4 GND 0.17fF
C87 QN.n0 GND 0.30fF
C88 QN.n1 GND 0.39fF
C89 QN.n2 GND 0.35fF
C90 QN.n3 GND 0.45fF
C91 QN.n4 GND 0.53fF
C92 QN.n5 GND 0.04fF
C93 QN.n6 GND 0.05fF
C94 QN.n7 GND 0.03fF
C95 QN.n8 GND 0.20fF
C96 QN.n9 GND 0.49fF
C97 QN.n10 GND 0.03fF
C98 a_277_1050.n0 GND 0.49fF
C99 a_277_1050.n1 GND 0.49fF
C100 a_277_1050.n2 GND 0.38fF
C101 a_277_1050.n3 GND 1.20fF
C102 a_277_1050.n4 GND 0.38fF
C103 a_277_1050.n5 GND 0.55fF
C104 a_277_1050.n6 GND 1.82fF
C105 a_277_1050.n7 GND 0.46fF
C106 a_277_1050.n8 GND 0.73fF
C107 a_277_1050.n9 GND 0.53fF
C108 a_277_1050.n10 GND 0.60fF
C109 a_277_1050.n11 GND 0.63fF
C110 VDD.n1 GND 0.03fF
C111 VDD.n2 GND 0.13fF
C112 VDD.n3 GND 0.03fF
C113 VDD.n4 GND 0.02fF
C114 VDD.n5 GND 0.06fF
C115 VDD.n6 GND 0.02fF
C116 VDD.n7 GND 0.02fF
C117 VDD.n8 GND 0.02fF
C118 VDD.n9 GND 0.02fF
C119 VDD.n10 GND 0.02fF
C120 VDD.n11 GND 0.02fF
C121 VDD.n12 GND 0.02fF
C122 VDD.n13 GND 0.02fF
C123 VDD.n14 GND 0.04fF
C124 VDD.n15 GND 0.01fF
C125 VDD.n20 GND 0.45fF
C126 VDD.n21 GND 0.27fF
C127 VDD.n22 GND 0.02fF
C128 VDD.n23 GND 0.03fF
C129 VDD.n24 GND 0.06fF
C130 VDD.n25 GND 0.24fF
C131 VDD.n26 GND 0.01fF
C132 VDD.n27 GND 0.01fF
C133 VDD.n28 GND 0.01fF
C134 VDD.n29 GND 0.17fF
C135 VDD.n30 GND 0.01fF
C136 VDD.n31 GND 0.02fF
C137 VDD.n32 GND 0.08fF
C138 VDD.n33 GND 0.08fF
C139 VDD.n34 GND 0.05fF
C140 VDD.n35 GND 0.01fF
C141 VDD.n36 GND 0.02fF
C142 VDD.n37 GND 0.03fF
C143 VDD.n38 GND 0.14fF
C144 VDD.n39 GND 0.01fF
C145 VDD.n40 GND 0.02fF
C146 VDD.n41 GND 0.03fF
C147 VDD.n42 GND 0.16fF
C148 VDD.n43 GND 0.01fF
C149 VDD.n44 GND 0.02fF
C150 VDD.n45 GND 0.02fF
C151 VDD.n46 GND 0.06fF
C152 VDD.n47 GND 0.25fF
C153 VDD.n48 GND 0.01fF
C154 VDD.n49 GND 0.01fF
C155 VDD.n50 GND 0.02fF
C156 VDD.n51 GND 0.27fF
C157 VDD.n52 GND 0.01fF
C158 VDD.n53 GND 0.02fF
C159 VDD.n54 GND 0.03fF
C160 VDD.n55 GND 0.05fF
C161 VDD.n56 GND 0.02fF
C162 VDD.n57 GND 0.02fF
C163 VDD.n58 GND 0.02fF
C164 VDD.n59 GND 0.02fF
C165 VDD.n60 GND 0.02fF
C166 VDD.n61 GND 0.02fF
C167 VDD.n62 GND 0.02fF
C168 VDD.n63 GND 0.02fF
C169 VDD.n64 GND 0.02fF
C170 VDD.n65 GND 0.02fF
C171 VDD.n66 GND 0.02fF
C172 VDD.n67 GND 0.03fF
C173 VDD.n68 GND 0.02fF
C174 VDD.n69 GND 0.22fF
C175 VDD.n70 GND 0.02fF
C176 VDD.n71 GND 0.02fF
C177 VDD.n73 GND 0.02fF
C178 VDD.n77 GND 0.27fF
C179 VDD.n78 GND 0.27fF
C180 VDD.n79 GND 0.01fF
C181 VDD.n80 GND 0.02fF
C182 VDD.n81 GND 0.03fF
C183 VDD.n82 GND 0.06fF
C184 VDD.n83 GND 0.24fF
C185 VDD.n84 GND 0.01fF
C186 VDD.n85 GND 0.01fF
C187 VDD.n86 GND 0.02fF
C188 VDD.n87 GND 0.17fF
C189 VDD.n88 GND 0.01fF
C190 VDD.n89 GND 0.02fF
C191 VDD.n90 GND 0.02fF
C192 VDD.n91 GND 0.08fF
C193 VDD.n92 GND 0.05fF
C194 VDD.n93 GND 0.01fF
C195 VDD.n94 GND 0.02fF
C196 VDD.n95 GND 0.03fF
C197 VDD.n96 GND 0.14fF
C198 VDD.n97 GND 0.01fF
C199 VDD.n98 GND 0.02fF
C200 VDD.n99 GND 0.03fF
C201 VDD.n100 GND 0.16fF
C202 VDD.n101 GND 0.01fF
C203 VDD.n102 GND 0.02fF
C204 VDD.n103 GND 0.02fF
C205 VDD.n104 GND 0.06fF
C206 VDD.n105 GND 0.25fF
C207 VDD.n106 GND 0.01fF
C208 VDD.n107 GND 0.01fF
C209 VDD.n108 GND 0.02fF
C210 VDD.n109 GND 0.27fF
C211 VDD.n110 GND 0.01fF
C212 VDD.n111 GND 0.02fF
C213 VDD.n112 GND 0.03fF
C214 VDD.n113 GND 0.21fF
C215 VDD.n114 GND 0.02fF
C216 VDD.n115 GND 0.02fF
C217 VDD.n116 GND 0.02fF
C218 VDD.n117 GND 0.06fF
C219 VDD.n118 GND 0.02fF
C220 VDD.n119 GND 0.02fF
C221 VDD.n120 GND 0.02fF
C222 VDD.n121 GND 0.02fF
C223 VDD.n122 GND 0.02fF
C224 VDD.n123 GND 0.02fF
C225 VDD.n124 GND 0.02fF
C226 VDD.n125 GND 0.02fF
C227 VDD.n126 GND 0.02fF
C228 VDD.n127 GND 0.02fF
C229 VDD.n128 GND 0.03fF
C230 VDD.n129 GND 0.02fF
C231 VDD.n130 GND 0.02fF
C232 VDD.n134 GND 0.27fF
C233 VDD.n135 GND 0.27fF
C234 VDD.n136 GND 0.01fF
C235 VDD.n137 GND 0.02fF
C236 VDD.n138 GND 0.03fF
C237 VDD.n139 GND 0.06fF
C238 VDD.n140 GND 0.24fF
C239 VDD.n141 GND 0.01fF
C240 VDD.n142 GND 0.01fF
C241 VDD.n143 GND 0.02fF
C242 VDD.n144 GND 0.17fF
C243 VDD.n145 GND 0.01fF
C244 VDD.n146 GND 0.02fF
C245 VDD.n147 GND 0.02fF
C246 VDD.n148 GND 0.08fF
C247 VDD.n149 GND 0.05fF
C248 VDD.n150 GND 0.01fF
C249 VDD.n151 GND 0.02fF
C250 VDD.n152 GND 0.03fF
C251 VDD.n153 GND 0.14fF
C252 VDD.n154 GND 0.01fF
C253 VDD.n155 GND 0.02fF
C254 VDD.n156 GND 0.03fF
C255 VDD.n157 GND 0.16fF
C256 VDD.n158 GND 0.01fF
C257 VDD.n159 GND 0.02fF
C258 VDD.n160 GND 0.02fF
C259 VDD.n161 GND 0.06fF
C260 VDD.n162 GND 0.25fF
C261 VDD.n163 GND 0.01fF
C262 VDD.n164 GND 0.01fF
C263 VDD.n165 GND 0.02fF
C264 VDD.n166 GND 0.27fF
C265 VDD.n167 GND 0.01fF
C266 VDD.n168 GND 0.02fF
C267 VDD.n169 GND 0.03fF
C268 VDD.n170 GND 0.21fF
C269 VDD.n171 GND 0.02fF
C270 VDD.n172 GND 0.02fF
C271 VDD.n173 GND 0.02fF
C272 VDD.n174 GND 0.06fF
C273 VDD.n175 GND 0.02fF
C274 VDD.n176 GND 0.02fF
C275 VDD.n177 GND 0.02fF
C276 VDD.n178 GND 0.02fF
C277 VDD.n179 GND 0.02fF
C278 VDD.n180 GND 0.02fF
C279 VDD.n181 GND 0.02fF
C280 VDD.n182 GND 0.02fF
C281 VDD.n183 GND 0.02fF
C282 VDD.n184 GND 0.02fF
C283 VDD.n185 GND 0.03fF
C284 VDD.n186 GND 0.02fF
C285 VDD.n187 GND 0.02fF
C286 VDD.n191 GND 0.27fF
C287 VDD.n192 GND 0.27fF
C288 VDD.n193 GND 0.01fF
C289 VDD.n194 GND 0.02fF
C290 VDD.n195 GND 0.03fF
C291 VDD.n196 GND 0.06fF
C292 VDD.n197 GND 0.24fF
C293 VDD.n198 GND 0.01fF
C294 VDD.n199 GND 0.01fF
C295 VDD.n200 GND 0.01fF
C296 VDD.n201 GND 0.18fF
C297 VDD.n202 GND 0.02fF
C298 VDD.n203 GND 0.02fF
C299 VDD.n204 GND 0.06fF
C300 VDD.n205 GND 0.02fF
C301 VDD.n206 GND 0.02fF
C302 VDD.n207 GND 0.02fF
C303 VDD.n208 GND 0.02fF
C304 VDD.n209 GND 0.02fF
C305 VDD.n210 GND 0.02fF
C306 VDD.n211 GND 0.02fF
C307 VDD.n212 GND 0.02fF
C308 VDD.n213 GND 0.03fF
C309 VDD.n214 GND 0.04fF
C310 VDD.n215 GND 0.02fF
C311 VDD.n219 GND 0.45fF
C312 VDD.n220 GND 0.27fF
C313 VDD.n221 GND 0.02fF
C314 VDD.n222 GND 0.03fF
C315 VDD.n223 GND 0.03fF
C316 VDD.n224 GND 0.27fF
C317 VDD.n225 GND 0.01fF
C318 VDD.n226 GND 0.02fF
C319 VDD.n227 GND 0.02fF
C320 VDD.n228 GND 0.06fF
C321 VDD.n229 GND 0.22fF
C322 VDD.n230 GND 0.01fF
C323 VDD.n231 GND 0.01fF
C324 VDD.n232 GND 0.02fF
C325 VDD.n233 GND 0.17fF
C326 VDD.n234 GND 0.01fF
C327 VDD.n235 GND 0.02fF
C328 VDD.n236 GND 0.02fF
C329 VDD.n237 GND 0.08fF
C330 VDD.n238 GND 0.05fF
C331 VDD.n239 GND 0.15fF
C332 VDD.n240 GND 0.01fF
C333 VDD.n241 GND 0.02fF
C334 VDD.n242 GND 0.02fF
C335 VDD.n243 GND 0.15fF
C336 VDD.n244 GND 0.01fF
C337 VDD.n245 GND 0.02fF
C338 VDD.n246 GND 0.03fF
C339 VDD.n247 GND 0.14fF
C340 VDD.n248 GND 0.01fF
C341 VDD.n249 GND 0.02fF
C342 VDD.n250 GND 0.03fF
C343 VDD.n251 GND 0.16fF
C344 VDD.n252 GND 0.01fF
C345 VDD.n253 GND 0.08fF
C346 VDD.n254 GND 0.05fF
C347 VDD.n255 GND 0.02fF
C348 VDD.n256 GND 0.02fF
C349 VDD.n257 GND 0.17fF
C350 VDD.n258 GND 0.01fF
C351 VDD.n259 GND 0.02fF
C352 VDD.n260 GND 0.02fF
C353 VDD.n261 GND 0.22fF
C354 VDD.n262 GND 0.01fF
C355 VDD.n263 GND 0.07fF
C356 VDD.n264 GND 0.02fF
C357 VDD.n265 GND 0.27fF
C358 VDD.n266 GND 0.01fF
C359 VDD.n267 GND 0.02fF
C360 VDD.n268 GND 0.02fF
C361 VDD.n269 GND 0.27fF
C362 VDD.n270 GND 0.01fF
C363 VDD.n271 GND 0.02fF
C364 VDD.n272 GND 0.03fF
C365 VDD.n273 GND 0.05fF
C366 VDD.n274 GND 0.02fF
C367 VDD.n275 GND 0.02fF
C368 VDD.n276 GND 0.02fF
C369 VDD.n277 GND 0.02fF
C370 VDD.n278 GND 0.02fF
C371 VDD.n279 GND 0.02fF
C372 VDD.n280 GND 0.02fF
C373 VDD.n281 GND 0.02fF
C374 VDD.n282 GND 0.02fF
C375 VDD.n283 GND 0.02fF
C376 VDD.n284 GND 0.02fF
C377 VDD.n285 GND 0.03fF
C378 VDD.n286 GND 0.02fF
C379 VDD.n289 GND 0.02fF
C380 VDD.n291 GND 0.02fF
C381 VDD.n292 GND 0.26fF
C382 VDD.n293 GND 0.02fF
C383 VDD.n295 GND 0.27fF
C384 VDD.n296 GND 0.27fF
C385 VDD.n297 GND 0.01fF
C386 VDD.n298 GND 0.02fF
C387 VDD.n299 GND 0.03fF
C388 VDD.n300 GND 0.06fF
C389 VDD.n301 GND 0.25fF
C390 VDD.n302 GND 0.01fF
C391 VDD.n303 GND 0.01fF
C392 VDD.n304 GND 0.02fF
C393 VDD.n305 GND 0.16fF
C394 VDD.n306 GND 0.01fF
C395 VDD.n307 GND 0.02fF
C396 VDD.n308 GND 0.02fF
C397 VDD.n309 GND 0.14fF
C398 VDD.n310 GND 0.01fF
C399 VDD.n311 GND 0.02fF
C400 VDD.n312 GND 0.03fF
C401 VDD.n313 GND 0.08fF
C402 VDD.n314 GND 0.05fF
C403 VDD.n315 GND 0.01fF
C404 VDD.n316 GND 0.02fF
C405 VDD.n317 GND 0.03fF
C406 VDD.n318 GND 0.17fF
C407 VDD.n319 GND 0.01fF
C408 VDD.n320 GND 0.02fF
C409 VDD.n321 GND 0.02fF
C410 VDD.n322 GND 0.06fF
C411 VDD.n323 GND 0.24fF
C412 VDD.n324 GND 0.01fF
C413 VDD.n325 GND 0.01fF
C414 VDD.n326 GND 0.02fF
C415 VDD.n327 GND 0.27fF
C416 VDD.n328 GND 0.01fF
C417 VDD.n329 GND 0.02fF
C418 VDD.n330 GND 0.03fF
C419 VDD.n331 GND 0.21fF
C420 VDD.n332 GND 0.02fF
C421 VDD.n333 GND 0.02fF
C422 VDD.n334 GND 0.02fF
C423 VDD.n335 GND 0.06fF
C424 VDD.n336 GND 0.02fF
C425 VDD.n337 GND 0.02fF
C426 VDD.n338 GND 0.02fF
C427 VDD.n339 GND 0.02fF
C428 VDD.n340 GND 0.02fF
C429 VDD.n341 GND 0.02fF
C430 VDD.n342 GND 0.02fF
C431 VDD.n343 GND 0.02fF
C432 VDD.n344 GND 0.02fF
C433 VDD.n345 GND 0.02fF
C434 VDD.n346 GND 0.03fF
C435 VDD.n347 GND 0.02fF
C436 VDD.n348 GND 0.02fF
C437 VDD.n352 GND 0.27fF
C438 VDD.n353 GND 0.27fF
C439 VDD.n354 GND 0.01fF
C440 VDD.n355 GND 0.02fF
C441 VDD.n356 GND 0.03fF
C442 VDD.n357 GND 0.06fF
C443 VDD.n358 GND 0.25fF
C444 VDD.n359 GND 0.01fF
C445 VDD.n360 GND 0.01fF
C446 VDD.n361 GND 0.02fF
C447 VDD.n362 GND 0.16fF
C448 VDD.n363 GND 0.01fF
C449 VDD.n364 GND 0.02fF
C450 VDD.n365 GND 0.02fF
C451 VDD.n366 GND 0.14fF
C452 VDD.n367 GND 0.01fF
C453 VDD.n368 GND 0.02fF
C454 VDD.n369 GND 0.03fF
C455 VDD.n370 GND 0.08fF
C456 VDD.n371 GND 0.05fF
C457 VDD.n372 GND 0.01fF
C458 VDD.n373 GND 0.02fF
C459 VDD.n374 GND 0.03fF
C460 VDD.n375 GND 0.17fF
C461 VDD.n376 GND 0.01fF
C462 VDD.n377 GND 0.02fF
C463 VDD.n378 GND 0.02fF
C464 a_147_187.n0 GND 0.56fF
C465 a_147_187.n1 GND 0.71fF
C466 a_147_187.n2 GND 0.75fF
C467 a_147_187.n3 GND 0.40fF
C468 a_147_187.t5 GND 0.83fF
C469 a_147_187.n4 GND 0.91fF
C470 a_147_187.n5 GND 0.40fF
C471 a_147_187.t12 GND 0.83fF
C472 a_147_187.n6 GND 0.56fF
C473 a_147_187.n7 GND 0.41fF
C474 a_147_187.n8 GND 1.32fF
C475 a_147_187.n9 GND 1.99fF
C476 a_147_187.n10 GND 1.57fF
C477 a_147_187.n11 GND 0.73fF
C478 a_147_187.n12 GND 0.12fF
C479 a_147_187.n13 GND 0.40fF
C480 a_147_187.n14 GND 0.07fF
C481 a_1845_1050.n0 GND 0.37fF
C482 a_1845_1050.n1 GND 0.47fF
C483 a_1845_1