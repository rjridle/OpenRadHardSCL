magic
tech sky130A
magscale 1 2
timestamp 1643177486
<< nmos >>
rect 11 150 41 212
rect 11 120 107 150
tri 107 120 137 150 sw
rect 11 28 41 120
tri 41 104 57 120 nw
tri 91 104 107 120 ne
tri 41 28 57 44 sw
tri 91 28 107 44 se
rect 107 28 137 120
tri 11 -2 41 28 ne
rect 41 -2 107 28
tri 107 -2 137 28 nw
<< ndiff >>
rect -45 196 11 212
rect -45 162 -35 196
rect -1 162 11 196
rect -45 125 11 162
rect 41 196 193 212
rect 41 162 149 196
rect 183 162 193 196
rect 41 150 193 162
rect -45 91 -35 125
rect -1 91 11 125
tri 107 120 137 150 ne
rect 137 125 193 150
rect -45 57 11 91
rect -45 23 -35 57
rect -1 23 11 57
tri 41 104 57 120 se
rect 57 104 91 120
tri 91 104 107 120 sw
rect 41 91 107 104
rect 41 57 57 91
rect 91 57 107 91
rect 41 44 107 57
tri 41 28 57 44 ne
rect 57 28 91 44
tri 91 28 107 44 nw
rect 137 91 149 125
rect 183 91 193 125
rect 137 57 193 91
rect -45 -2 11 23
tri 11 -2 41 28 sw
tri 107 -2 137 28 se
rect 137 23 149 57
rect 183 23 193 57
rect 137 -2 193 23
rect -45 -14 193 -2
rect -45 -48 -35 -14
rect -1 -48 57 -14
rect 91 -48 149 -14
rect 183 -48 193 -14
rect -45 -64 193 -48
<< ndiffc >>
rect -35 162 -1 196
rect 149 162 183 196
rect -35 91 -1 125
rect -35 23 -1 57
rect 57 57 91 91
rect 149 91 183 125
rect 149 23 183 57
rect -35 -48 -1 -14
rect 57 -48 91 -14
rect 149 -48 183 -14
<< poly >>
rect 11 212 41 238
<< locali >>
rect -35 196 -1 212
rect -35 125 -1 162
rect 149 196 183 212
rect 149 125 183 162
rect -35 57 -1 91
rect 57 91 91 107
rect 57 41 91 57
rect 149 57 183 91
rect -35 -14 -1 23
rect 149 -14 183 23
rect -1 -48 57 -14
rect 91 -48 149 -14
rect -35 -64 -1 -48
rect 149 -64 183 -48
<< end >>
