magic
tech sky130A
magscale 1 2
timestamp 1645636714
<< nmos >>
tri 144 222 160 238 se
rect 160 222 190 276
tri 54 192 84 222 se
rect 84 192 190 222
rect 54 92 84 192
tri 84 176 100 192 nw
tri 144 176 160 192 ne
tri 84 92 100 108 sw
tri 144 92 160 108 se
rect 160 92 190 192
tri 54 62 84 92 ne
rect 84 62 160 92
tri 160 62 190 92 nw
<< ndiff >>
rect -1 260 160 276
rect -1 226 9 260
rect 43 238 160 260
rect 43 226 144 238
rect -1 222 144 226
tri 144 222 160 238 nw
rect 190 260 246 276
rect 190 226 202 260
rect 236 226 246 260
rect -1 189 54 222
tri 54 192 84 222 nw
rect -1 155 9 189
rect 43 155 54 189
rect -1 121 54 155
rect -1 87 9 121
rect 43 87 54 121
tri 84 176 100 192 se
rect 100 176 144 192
tri 144 176 160 192 sw
rect 84 148 160 176
rect 84 114 105 148
rect 139 114 160 148
rect 84 108 160 114
tri 84 92 100 108 ne
rect 100 92 144 108
tri 144 92 160 108 nw
rect 190 189 246 226
rect 190 155 202 189
rect 236 155 246 189
rect 190 121 246 155
rect -1 62 54 87
tri 54 62 84 92 sw
tri 160 62 190 92 se
rect 190 87 202 121
rect 236 87 246 121
rect 190 62 246 87
rect -1 50 246 62
rect -1 16 9 50
rect 43 16 110 50
rect 144 16 202 50
rect 236 16 246 50
rect -1 0 246 16
<< ndiffc >>
rect 9 226 43 260
rect 202 226 236 260
rect 9 155 43 189
rect 9 87 43 121
rect 105 114 139 148
rect 202 155 236 189
rect 202 87 236 121
rect 9 16 43 50
rect 110 16 144 50
rect 202 16 236 50
<< poly >>
rect 160 276 190 309
<< locali >>
rect 9 260 43 276
rect 9 189 43 226
rect 202 260 236 276
rect 202 189 236 226
rect 9 121 43 155
rect 105 148 139 164
rect 105 98 139 114
rect 202 121 236 155
rect 9 50 43 87
rect 202 50 236 87
rect 43 16 110 50
rect 144 16 202 50
rect 9 0 43 16
rect 202 0 236 16
<< end >>
