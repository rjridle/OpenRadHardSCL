* NGSPICE file created from NAND2X1.ext - technology: sky130A

.subckt NAND2X1 VDD VSS Y A B
X0 VSS A nmos_bottom_0/a_0_0# VSS sky130_fd_pr__nfet_01v8 ad=1.772e+11p pd=1.56e+06u as=0p ps=0u w=3e+06u l=150000u
X1 Y B nmos_bottom_0/a_0_0# VSS sky130_fd_pr__nfet_01v8 ad=1.772e+11p pd=1.56e+06u as=0p ps=0u w=3e+06u l=150000u
X2 Y A VDD VDD sky130_fd_pr__pfet_01v8 ad=-8.675e+09p pd=9.165e+06u as=2.27525e+12p ps=1.3685e+07u w=2e+06u l=150000u M=2
X3 Y B VDD VDD sky130_fd_pr__pfet_01v8 ad=-0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
.ends
