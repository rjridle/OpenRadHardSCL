* SPICE3 file created from DFFSNRNQX1.ext - technology: sky130A

.subckt DFFSNRNQX1 Q D CLK SN RN VDD GND
X0 GND a_4125_1050.t7 a_4901_103.t0 GND sky130_fd_pr__nfet_01v8 ad=1.0746p pd=9.42u as=0p ps=0u w=0u l=0u
X1 a_599_989.t6 CLK.t0 VDD.t65 �H���U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X2 VDD.t55 a_277_1050.t7 a_2201_1050.t4  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X3 VDD.t63 CLK.t1 a_1561_989.t4 VDD.t62 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X4 VDD.t41 RN.t0 a_277_1050.t3  �Y�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X5 a_599_989.t1 a_1561_989.t7 VDD.t17 ��Y�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X6 VDD.t31 RN.t1 a_1561_989.t1  �Y�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X7 a_4125_1050.t6 a_599_989.t8 VDD.t67 ��Y�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X8 VDD.t71 SN.t1 a_2201_1050.t6  �Y�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X9 a_1561_989.t3 CLK.t4 VDD.t61 ��Y�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X10 a_4125_1050.t4 Q.t7 VDD.t49  �Y�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X11 VDD.t15 a_599_989.t9 a_277_1050.t6 ��Y�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X12 GND D.t1 a_91_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X13 VDD.t69 a_1561_989.t8 a_2201_1050.t5  �Y�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X14 a_1561_989.t6 a_2201_1050.t7 VDD.t47 ��Y�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X15 a_4125_1050.t2 RN.t2 VDD.t1  �Y�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X16 VDD.t9 a_4125_1050.t8 Q.t3 ��Y�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X17 a_277_1050.t1 D.t0 VDD.t5  �Y�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X18 VDD.t39 a_277_1050.t8 a_599_989.t3 ��Y�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X19 VDD.t13 a_1561_989.t9 a_599_989.t0  �Y�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X20 VDD.t57 SN.t2 Q.t1 ��Y�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X21 a_277_1050.t2 RN.t3 VDD.t7  �Y�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X22 VDD.t59 CLK.t5 a_599_989.t5 ��Y�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X23 a_2201_1050.t1 SN.t3 VDD.t33  �Y�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X24 a_1561_989.t0 RN.t4 VDD.t25 ��Y�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X25 VDD.t11 a_1561_989.t10 Q.t6  �Y�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X26 GND a_277_1050.t11 a_2015_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X27 Q a_1561_989.t15 a_5182_210.t1 GND sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=0p ps=0u w=0u l=0u
X28 a_599_989.t4 a_277_1050.t9 VDD.t53 ��Y�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X29 VDD.t51 RN.t5 a_4125_1050.t1  �Y�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X30 a_277_1050.t5 a_599_989.t11 VDD.t45 ��Y�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X31 a_2201_1050.t3 a_277_1050.t10 VDD.t37  �Y�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X32 GND a_2201_1050.t8 a_2977_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X33 a_2201_1050.t2 a_1561_989.t12 VDD.t35 ��Y�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X34 VDD.t43 a_599_989.t12 a_4125_1050.t5  �Y�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X35 VDD.t29 Q.t9 a_4125_1050.t3 ��Y�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X36 Q.t2 a_4125_1050.t9 VDD.t23  �Y�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X37 GND a_277_1050.t12 a_1053_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X38 Q.t5 a_1561_989.t14 VDD.t27 ��Y�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X39 GND a_599_989.t7 a_3939_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X40 VDD.t21 a_2201_1050.t9 a_1561_989.t5  �Y�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X41 Q.t0 SN.t4 VDD.t19 ��Y�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X42 VDD.t3 D.t2 a_277_1050.t0  �Y�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
C0 D VDD 0.35fF
C1 VDD RN 4.40fF
C2 VDD CLK 0.59fF
C3 D RN 0.18fF
C4 Q VDD 2.79fF
C5 SN VDD 0.59fF
C6 RN CLK 0.73fF
C7 Q RN 0.18fF
C8 SN RN 0.37fF
C9 SN CLK 0.48fF
C10 Q SN 0.39fF
R0 CLK.n2 CLK.t5 479.223
R1 CLK.n0 CLK.t1 479.223
R2 CLK.n2 CLK.t0 375.52
R3 CLK.n0 CLK.t4 375.52
R4 CLK.n3 CLK.t2 287.572
R5 CLK.n1 CLK.t3 287.572
R6 CLK.n3 CLK.n2 196.47
R7 CLK.n1 CLK.n0 196.47
R8 CLK.n4 CLK.n1 11.678
R9 CLK.n4 CLK.n3 4.65
R10 CLK.n4 CLK 0.046
R11 VDD.n336 VDD.n325 144.705
R12 VDD.n466 VDD.n459 144.705
R13 VDD.n411 VDD.n404 144.705
R14 VDD.n172 VDD.n165 144.705
R15 VDD.n97 VDD.n86 144.705
R16 VDD.n302 VDD.t15 143.754
R17 VDD.n378 VDD.t13 143.754
R18 VDD.n453 VDD.t69 143.754
R19 VDD.n181 VDD.t31 143.754
R20 VDD.n106 VDD.t29 143.754
R21 VDD.n30 VDD.t11 143.754
R22 VDD.n267 VDD.t5 135.17
R23 VDD.n343 VDD.t53 135.17
R24 VDD.n418 VDD.t37 135.17
R25 VDD.n211 VDD.t47 135.17
R26 VDD.n136 VDD.t67 135.17
R27 VDD.n60 VDD.t23 135.17
R28 VDD.n277 VDD.n276 129.472
R29 VDD.n293 VDD.n292 129.472
R30 VDD.n353 VDD.n352 129.472
R31 VDD.n369 VDD.n368 129.472
R32 VDD.n428 VDD.n427 129.472
R33 VDD.n444 VDD.n443 129.472
R34 VDD.n202 VDD.n201 129.472
R35 VDD.n190 VDD.n189 129.472
R36 VDD.n127 VDD.n126 129.472
R37 VDD.n115 VDD.n114 129.472
R38 VDD.n51 VDD.n50 129.472
R39 VDD.n39 VDD.n38 129.472
R40 VDD.n82 VDD.n81 92.5
R41 VDD.n80 VDD.n79 92.5
R42 VDD.n78 VDD.n77 92.5
R43 VDD.n76 VDD.n75 92.5
R44 VDD.n84 VDD.n83 92.5
R45 VDD.n161 VDD.n160 92.5
R46 VDD.n159 VDD.n158 92.5
R47 VDD.n157 VDD.n156 92.5
R48 VDD.n155 VDD.n154 92.5
R49 VDD.n163 VDD.n162 92.5
R50 VDD.n232 VDD.n231 92.5
R51 VDD.n230 VDD.n229 92.5
R52 VDD.n228 VDD.n227 92.5
R53 VDD.n226 VDD.n225 92.5
R54 VDD.n234 VDD.n233 92.5
R55 VDD.n400 VDD.n399 92.5
R56 VDD.n398 VDD.n397 92.5
R57 VDD.n396 VDD.n395 92.5
R58 VDD.n394 VDD.n393 92.5
R59 VDD.n402 VDD.n401 92.5
R60 VDD.n321 VDD.n320 92.5
R61 VDD.n319 VDD.n318 92.5
R62 VDD.n317 VDD.n316 92.5
R63 VDD.n315 VDD.n314 92.5
R64 VDD.n323 VDD.n322 92.5
R65 VDD.n251 VDD.n250 92.5
R66 VDD.n249 VDD.n248 92.5
R67 VDD.n247 VDD.n246 92.5
R68 VDD.n245 VDD.n244 92.5
R69 VDD.n253 VDD.n252 92.5
R70 VDD.n14 VDD.n1 92.5
R71 VDD.n5 VDD.n4 92.5
R72 VDD.n7 VDD.n6 92.5
R73 VDD.n9 VDD.n8 92.5
R74 VDD.n11 VDD.n10 92.5
R75 VDD.n13 VDD.n12 92.5
R76 VDD.n21 VDD.n20 92.059
R77 VDD.n96 VDD.n95 92.059
R78 VDD.n171 VDD.n170 92.059
R79 VDD.n465 VDD.n464 92.059
R80 VDD.n410 VDD.n409 92.059
R81 VDD.n335 VDD.n334 92.059
R82 VDD.n259 VDD.n258 92.059
R83 VDD.n20 VDD.n16 67.194
R84 VDD.n20 VDD.n17 67.194
R85 VDD.n20 VDD.n18 67.194
R86 VDD.n20 VDD.n19 67.194
R87 VDD.n243 VDD.n242 44.141
R88 VDD.n392 VDD.n391 44.141
R89 VDD.n224 VDD.n223 44.141
R90 VDD.n153 VDD.n152 44.141
R91 VDD.n5 VDD.n3 44.141
R92 VDD.n391 VDD.n389 44.107
R93 VDD.n223 VDD.n221 44.107
R94 VDD.n152 VDD.n150 44.107
R95 VDD.n242 VDD.n240 44.107
R96 VDD.n3 VDD.n2 44.107
R97 VDD.n20 VDD.n15 41.052
R98 VDD.n90 VDD.n88 39.742
R99 VDD.n90 VDD.n89 39.742
R100 VDD.n92 VDD.n91 39.742
R101 VDD.n167 VDD.n166 39.742
R102 VDD.n461 VDD.n460 39.742
R103 VDD.n406 VDD.n405 39.742
R104 VDD.n255 VDD.n254 39.742
R105 VDD.n333 VDD.n330 39.742
R106 VDD.n333 VDD.n332 39.742
R107 VDD.n329 VDD.n328 39.742
R108 VDD.n152 VDD.n151 38
R109 VDD.n223 VDD.n222 38
R110 VDD.n391 VDD.n390 38
R111 VDD.n242 VDD.n241 38
R112 VDD.n389 VDD.n388 36.774
R113 VDD.n221 VDD.n220 36.774
R114 VDD.n150 VDD.n149 36.774
R115 VDD.n88 VDD.n87 36.774
R116 VDD.n332 VDD.n331 36.774
R117 VDD.n32  �Y�� 35.8
R118 VDD.n108 ��Y�� 35.8
R119 VDD.n183  �Y�� 35.8
R120 VDD.n447  �Y�� 35.8
R121 VDD.n372  �Y�� 35.8
R122 VDD.n296 ��Y�� 35.8
R123 VDD.n56  �Y�� 33.243
R124 VDD.n132 ��Y�� 33.243
R125 VDD.n207 ��Y�� 33.243
R126 VDD.n423  �Y�� 33.243
R127 VDD.n348 ��Y�� 33.243
R128 VDD.n272  �Y�� 33.243
R129 VDD.n1 VDD.n0 30.923
R130 VDD.n95 VDD.n93 26.38
R131 VDD.n95 VDD.n92 26.38
R132 VDD.n95 VDD.n90 26.38
R133 VDD.n95 VDD.n94 26.38
R134 VDD.n170 VDD.n168 26.38
R135 VDD.n170 VDD.n167 26.38
R136 VDD.n170 VDD.n169 26.38
R137 VDD.n464 VDD.n462 26.38
R138 VDD.n464 VDD.n461 26.38
R139 VDD.n464 VDD.n463 26.38
R140 VDD.n409 VDD.n407 26.38
R141 VDD.n409 VDD.n406 26.38
R142 VDD.n409 VDD.n408 26.38
R143 VDD.n258 VDD.n256 26.38
R144 VDD.n258 VDD.n255 26.38
R145 VDD.n258 VDD.n257 26.38
R146 VDD.n334 VDD.n333 26.38
R147 VDD.n334 VDD.n329 26.38
R148 VDD.n334 VDD.n327 26.38
R149 VDD.n334 VDD.n326 26.38
R150 VDD.n261 VDD.n253 22.915
R151 VDD.n23 VDD.n14 22.915
R152 VDD.n36 ��Y�� 15.343
R153 VDD.n112  �Y�� 15.343
R154 VDD.n187 ��Y�� 15.343
R155 VDD.n441 ��Y�� 15.343
R156 VDD.n366 ��Y�� 15.343
R157 VDD.n290 ��Y�� 15.343
R158 VDD.n253 VDD.n251 14.864
R159 VDD.n251 VDD.n249 14.864
R160 VDD.n249 VDD.n247 14.864
R161 VDD.n247 VDD.n245 14.864
R162 VDD.n245 VDD.n243 14.864
R163 VDD.n402 VDD.n400 14.864
R164 VDD.n400 VDD.n398 14.864
R165 VDD.n398 VDD.n396 14.864
R166 VDD.n396 VDD.n394 14.864
R167 VDD.n394 VDD.n392 14.864
R168 VDD.n234 VDD.n232 14.864
R169 VDD.n232 VDD.n230 14.864
R170 VDD.n230 VDD.n228 14.864
R171 VDD.n228 VDD.n226 14.864
R172 VDD.n226 VDD.n224 14.864
R173 VDD.n163 VDD.n161 14.864
R174 VDD.n161 VDD.n159 14.864
R175 VDD.n159 VDD.n157 14.864
R176 VDD.n157 VDD.n155 14.864
R177 VDD.n155 VDD.n153 14.864
R178 VDD.n84 VDD.n82 14.864
R179 VDD.n82 VDD.n80 14.864
R180 VDD.n80 VDD.n78 14.864
R181 VDD.n78 VDD.n76 14.864
R182 VDD.n76 VDD.n74 14.864
R183 VDD.n74 VDD.n73 14.864
R184 VDD.n323 VDD.n321 14.864
R185 VDD.n321 VDD.n319 14.864
R186 VDD.n319 VDD.n317 14.864
R187 VDD.n317 VDD.n315 14.864
R188 VDD.n315 VDD.n313 14.864
R189 VDD.n313 VDD.n312 14.864
R190 VDD.n14 VDD.n13 14.864
R191 VDD.n13 VDD.n11 14.864
R192 VDD.n11 VDD.n9 14.864
R193 VDD.n9 VDD.n7 14.864
R194 VDD.n7 VDD.n5 14.864
R195 VDD.n98 VDD.n85 14.864
R196 VDD.n173 VDD.n164 14.864
R197 VDD.n238 VDD.n235 14.864
R198 VDD.n412 VDD.n403 14.864
R199 VDD.n337 VDD.n324 14.864
R200 VDD.n276 VDD.t7 14.282
R201 VDD.n276 VDD.t3 14.282
R202 VDD.n292 VDD.t45 14.282
R203 VDD.n292 VDD.t41 14.282
R204 VDD.n352 VDD.t65 14.282
R205 VDD.n352 VDD.t39 14.282
R206 VDD.n368 VDD.t17 14.282
R207 VDD.n368 VDD.t59 14.282
R208 VDD.n427 VDD.t33 14.282
R209 VDD.n427 VDD.t55 14.282
R210 VDD.n443 VDD.t35 14.282
R211 VDD.n443 VDD.t71 14.282
R212 VDD.n201 VDD.t61 14.282
R213 VDD.n201 VDD.t21 14.282
R214 VDD.n189 VDD.t25 14.282
R215 VDD.n189 VDD.t63 14.282
R216 VDD.n126 VDD.t1 14.282
R217 VDD.n126 VDD.t43 14.282
R218 VDD.n114 VDD.t49 14.282
R219 VDD.n114 VDD.t51 14.282
R220 VDD.n50 VDD.t19 14.282
R221 VDD.n50 VDD.t9 14.282
R222 VDD.n38 VDD.t27 14.282
R223 VDD.n38 VDD.t57 14.282
R224 VDD.n52 ��Y�� 12.786
R225 VDD.n128  �Y�� 12.786
R226 VDD.n203  �Y�� 12.786
R227 VDD.n429  M���U 12.786
R228 VDD.n354 ��Y�� 12.786
R229 VDD.n278  �Y�� 12.786
R230 VDD.n23 VDD.n22 8.855
R231 VDD.n22 VDD.n21 8.855
R232 VDD.n26 VDD.n25 8.855
R233 VDD.n25 VDD.n24 8.855
R234 VDD.n30 VDD.n29 8.855
R235 VDD.n29 VDD.n28 8.855
R236 VDD.n34 VDD.n33 8.855
R237 VDD.n33 VDD.n32 8.855
R238 VDD.n40 VDD.n37 8.855
R239 VDD.n37 VDD.n36 8.855
R240 VDD.n44 VDD.n43 8.855
R241 VDD.n43 VDD.n42 8.855
R242 VDD.n48 VDD.n47 8.855
R243 VDD.n47 VDD.n46 8.855
R244 VDD.n54 VDD.n53 8.855
R245 VDD.n53 VDD.n52 8.855
R246 VDD.n58 VDD.n57 8.855
R247 VDD.n57 VDD.n56 8.855
R248 VDD.n63 VDD.n62 8.855
R249 VDD.n62 VDD.n61 8.855
R250 VDD.n67 VDD.n66 8.855
R251 VDD.n66 VDD.n65 8.855
R252 VDD.n71 VDD.n70 8.855
R253 VDD.n70 VDD.n69 8.855
R254 VDD.n98 VDD.n97 8.855
R255 VDD.n97 VDD.n96 8.855
R256 VDD.n102 VDD.n101 8.855
R257 VDD.n101 VDD.n100 8.855
R258 VDD.n106 VDD.n105 8.855
R259 VDD.n105 VDD.n104 8.855
R260 VDD.n110 VDD.n109 8.855
R261 VDD.n109 VDD.n108 8.855
R262 VDD.n116 VDD.n113 8.855
R263 VDD.n113 VDD.n112 8.855
R264 VDD.n120 VDD.n119 8.855
R265 VDD.n119 VDD.n118 8.855
R266 VDD.n124 VDD.n123 8.855
R267 VDD.n123 VDD.n122 8.855
R268 VDD.n130 VDD.n129 8.855
R269 VDD.n129 VDD.n128 8.855
R270 VDD.n134 VDD.n133 8.855
R271 VDD.n133 VDD.n132 8.855
R272 VDD.n139 VDD.n138 8.855
R273 VDD.n138 VDD.n137 8.855
R274 VDD.n143 VDD.n142 8.855
R275 VDD.n142 VDD.n141 8.855
R276 VDD.n147 VDD.n146 8.855
R277 VDD.n146 VDD.n145 8.855
R278 VDD.n173 VDD.n172 8.855
R279 VDD.n172 VDD.n171 8.855
R280 VDD.n177 VDD.n176 8.855
R281 VDD.n176 VDD.n175 8.855
R282 VDD.n181 VDD.n180 8.855
R283 VDD.n180 VDD.n179 8.855
R284 VDD.n185 VDD.n184 8.855
R285 VDD.n184 VDD.n183 8.855
R286 VDD.n191 VDD.n188 8.855
R287 VDD.n188 VDD.n187 8.855
R288 VDD.n195 VDD.n194 8.855
R289 VDD.n194 VDD.n193 8.855
R290 VDD.n199 VDD.n198 8.855
R291 VDD.n198 VDD.n197 8.855
R292 VDD.n205 VDD.n204 8.855
R293 VDD.n204 VDD.n203 8.855
R294 VDD.n209 VDD.n208 8.855
R295 VDD.n208 VDD.n207 8.855
R296 VDD.n214 VDD.n213 8.855
R297 VDD.n213 VDD.n212 8.855
R298 VDD.n218 VDD.n217 8.855
R299 VDD.n217 VDD.n216 8.855
R300 VDD.n238 VDD.n237 8.855
R301 VDD.n237 VDD.n236 8.855
R302 VDD.n467 VDD.n466 8.855
R303 VDD.n466 VDD.n465 8.855
R304 VDD.n457 VDD.n456 8.855
R305 VDD.n456 VDD.n455 8.855
R306 VDD.n453 VDD.n452 8.855
R307 VDD.n452 VDD.n451 8.855
R308 VDD.n449 VDD.n448 8.855
R309 VDD.n448 VDD.n447 8.855
R310 VDD.n445 VDD.n442 8.855
R311 VDD.n442 VDD.n441 8.855
R312 VDD.n439 VDD.n438 8.855
R313 VDD.n438 VDD.n437 8.855
R314 VDD.n435 VDD.n434 8.855
R315 VDD.n434 VDD.n433 8.855
R316 VDD.n431 VDD.n430 8.855
R317 VDD.n430 VDD.n429 8.855
R318 VDD.n425 VDD.n424 8.855
R319 VDD.n424 VDD.n423 8.855
R320 VDD.n421 VDD.n420 8.855
R321 VDD.n420 VDD.n419 8.855
R322 VDD.n416 VDD.n415 8.855
R323 VDD.n415 VDD.n414 8.855
R324 VDD.n412 VDD.n411 8.855
R325 VDD.n411 VDD.n410 8.855
R326 VDD.n386 VDD.n385 8.855
R327 VDD.n385 VDD.n384 8.855
R328 VDD.n382 VDD.n381 8.855
R329 VDD.n381 VDD.n380 8.855
R330 VDD.n378 VDD.n377 8.855
R331 VDD.n377 VDD.n376 8.855
R332 VDD.n374 VDD.n373 8.855
R333 VDD.n373 VDD.n372 8.855
R334 VDD.n370 VDD.n367 8.855
R335 VDD.n367 VDD.n366 8.855
R336 VDD.n364 VDD.n363 8.855
R337 VDD.n363 VDD.n362 8.855
R338 VDD.n360 VDD.n359 8.855
R339 VDD.n359 VDD.n358 8.855
R340 VDD.n356 VDD.n355 8.855
R341 VDD.n355 VDD.n354 8.855
R342 VDD.n350 VDD.n349 8.855
R343 VDD.n349 VDD.n348 8.855
R344 VDD.n346 VDD.n345 8.855
R345 VDD.n345 VDD.n344 8.855
R346 VDD.n341 VDD.n340 8.855
R347 VDD.n340 VDD.n339 8.855
R348 VDD.n337 VDD.n336 8.855
R349 VDD.n336 VDD.n335 8.855
R350 VDD.n310 VDD.n309 8.855
R351 VDD.n309 VDD.n308 8.855
R352 VDD.n306 VDD.n305 8.855
R353 VDD.n305 VDD.n304 8.855
R354 VDD.n302 VDD.n301 8.855
R355 VDD.n301 VDD.n300 8.855
R356 VDD.n298 VDD.n297 8.855
R357 VDD.n297 VDD.n296 8.855
R358 VDD.n294 VDD.n291 8.855
R359 VDD.n291 VDD.n290 8.855
R360 VDD.n288 VDD.n287 8.855
R361 VDD.n287 VDD.n286 8.855
R362 VDD.n284 VDD.n283 8.855
R363 VDD.n283 VDD.n282 8.855
R364 VDD.n280 VDD.n279 8.855
R365 VDD.n279 VDD.n278 8.855
R366 VDD.n274 VDD.n273 8.855
R367 VDD.n273 VDD.n272 8.855
R368 VDD.n270 VDD.n269 8.855
R369 VDD.n269 VDD.n268 8.855
R370 VDD.n265 VDD.n264 8.855
R371 VDD.n264 VDD.n263 8.855
R372 VDD.n261 VDD.n260 8.855
R373 VDD.n260 VDD.n259 8.855
R374 VDD.n403 VDD.n402 8.051
R375 VDD.n235 VDD.n234 8.051
R376 VDD.n164 VDD.n163 8.051
R377 VDD.n85 VDD.n84 8.051
R378 VDD.n324 VDD.n323 8.051
R379 VDD.n46 ��Y�� 7.671
R380 VDD.n122  �Y�� 7.671
R381 VDD.n197 ��Y�� 7.671
R382 VDD.n433  �Y�� 7.671
R383 VDD.n358 �H���U 7.671
R384 VDD.n282  �Y�� 7.671
R385 VDD.n54 VDD.n51 7.019
R386 VDD.n130 VDD.n127 7.019
R387 VDD.n205 VDD.n202 7.019
R388 VDD.n431 VDD.n428 7.019
R389 VDD.n356 VDD.n353 7.019
R390 VDD.n280 VDD.n277 7.019
R391 VDD.n40 VDD.n39 6.606
R392 VDD.n116 VDD.n115 6.606
R393 VDD.n191 VDD.n190 6.606
R394 VDD.n445 VDD.n444 6.606
R395 VDD.n370 VDD.n369 6.606
R396 VDD.n294 VDD.n293 6.606
R397 VDD.n42 ��Y�� 5.114
R398 VDD.n118  �Y�� 5.114
R399 VDD.n193 VDD.t62 5.114
R400 VDD.n437  �Y�� 5.114
R401 VDD.n362 ��Y�� 5.114
R402 VDD.n286  �Y�� 5.114
R403 VDD.n31 VDD.n30 4.65
R404 VDD.n35 VDD.n34 4.65
R405 VDD.n41 VDD.n40 4.65
R406 VDD.n45 VDD.n44 4.65
R407 VDD.n49 VDD.n48 4.65
R408 VDD.n55 VDD.n54 4.65
R409 VDD.n59 VDD.n58 4.65
R410 VDD.n64 VDD.n63 4.65
R411 VDD.n68 VDD.n67 4.65
R412 VDD.n72 VDD.n71 4.65
R413 VDD.n99 VDD.n98 4.65
R414 VDD.n103 VDD.n102 4.65
R415 VDD.n107 VDD.n106 4.65
R416 VDD.n111 VDD.n110 4.65
R417 VDD.n117 VDD.n116 4.65
R418 VDD.n121 VDD.n120 4.65
R419 VDD.n125 VDD.n124 4.65
R420 VDD.n131 VDD.n130 4.65
R421 VDD.n135 VDD.n134 4.65
R422 VDD.n140 VDD.n139 4.65
R423 VDD.n144 VDD.n143 4.65
R424 VDD.n148 VDD.n147 4.65
R425 VDD.n174 VDD.n173 4.65
R426 VDD.n178 VDD.n177 4.65
R427 VDD.n182 VDD.n181 4.65
R428 VDD.n186 VDD.n185 4.65
R429 VDD.n192 VDD.n191 4.65
R430 VDD.n196 VDD.n195 4.65
R431 VDD.n200 VDD.n199 4.65
R432 VDD.n206 VDD.n205 4.65
R433 VDD.n210 VDD.n209 4.65
R434 VDD.n215 VDD.n214 4.65
R435 VDD.n219 VDD.n218 4.65
R436 VDD.n239 VDD.n238 4.65
R437 VDD.n468 VDD.n467 4.65
R438 VDD.n458 VDD.n457 4.65
R439 VDD.n454 VDD.n453 4.65
R440 VDD.n450 VDD.n449 4.65
R441 VDD.n446 VDD.n445 4.65
R442 VDD.n440 VDD.n439 4.65
R443 VDD.n436 VDD.n435 4.65
R444 VDD.n432 VDD.n431 4.65
R445 VDD.n426 VDD.n425 4.65
R446 VDD.n422 VDD.n421 4.65
R447 VDD.n417 VDD.n416 4.65
R448 VDD.n413 VDD.n412 4.65
R449 VDD.n387 VDD.n386 4.65
R450 VDD.n383 VDD.n382 4.65
R451 VDD.n379 VDD.n378 4.65
R452 VDD.n375 VDD.n374 4.65
R453 VDD.n371 VDD.n370 4.65
R454 VDD.n365 VDD.n364 4.65
R455 VDD.n361 VDD.n360 4.65
R456 VDD.n357 VDD.n356 4.65
R457 VDD.n351 VDD.n350 4.65
R458 VDD.n347 VDD.n346 4.65
R459 VDD.n342 VDD.n341 4.65
R460 VDD.n338 VDD.n337 4.65
R461 VDD.n311 VDD.n310 4.65
R462 VDD.n307 VDD.n306 4.65
R463 VDD.n303 VDD.n302 4.65
R464 VDD.n299 VDD.n298 4.65
R465 VDD.n295 VDD.n294 4.65
R466 VDD.n289 VDD.n288 4.65
R467 VDD.n285 VDD.n284 4.65
R468 VDD.n281 VDD.n280 4.65
R469 VDD.n275 VDD.n274 4.65
R470 VDD.n271 VDD.n270 4.65
R471 VDD.n266 VDD.n265 4.65
R472 VDD.n262 VDD.n261 4.65
R473 VDD.n27 VDD.n23 2.933
R474 VDD.n27 VDD.n26 2.844
R475 VDD.n31 VDD.n27 1.063
R476 VDD.n63 VDD.n60 0.412
R477 VDD.n139 VDD.n136 0.412
R478 VDD.n214 VDD.n211 0.412
R479 VDD.n421 VDD.n418 0.412
R480 VDD.n346 VDD.n343 0.412
R481 VDD.n270 VDD.n267 0.412
R482 VDD.n99 VDD.n72 0.29
R483 VDD.n174 VDD.n148 0.29
R484 VDD.n413 VDD.n387 0.29
R485 VDD.n338 VDD.n311 0.29
R486 VDD.n262 VDD 0.207
R487 VDD.n49 VDD.n45 0.197
R488 VDD.n125 VDD.n121 0.197
R489 VDD.n200 VDD.n196 0.197
R490 VDD.n440 VDD.n436 0.197
R491 VDD.n365 VDD.n361 0.197
R492 VDD.n289 VDD.n285 0.197
R493 VDD.n35 VDD.n31 0.145
R494 VDD.n41 VDD.n35 0.145
R495 VDD.n45 VDD.n41 0.145
R496 VDD.n55 VDD.n49 0.145
R497 VDD.n59 VDD.n55 0.145
R498 VDD.n64 VDD.n59 0.145
R499 VDD.n68 VDD.n64 0.145
R500 VDD.n72 VDD.n68 0.145
R501 VDD.n103 VDD.n99 0.145
R502 VDD.n107 VDD.n103 0.145
R503 VDD.n111 VDD.n107 0.145
R504 VDD.n117 VDD.n111 0.145
R505 VDD.n121 VDD.n117 0.145
R506 VDD.n131 VDD.n125 0.145
R507 VDD.n135 VDD.n131 0.145
R508 VDD.n140 VDD.n135 0.145
R509 VDD.n144 VDD.n140 0.145
R510 VDD.n148 VDD.n144 0.145
R511 VDD.n178 VDD.n174 0.145
R512 VDD.n182 VDD.n178 0.145
R513 VDD.n186 VDD.n182 0.145
R514 VDD.n192 VDD.n186 0.145
R515 VDD.n196 VDD.n192 0.145
R516 VDD.n206 VDD.n200 0.145
R517 VDD.n210 VDD.n206 0.145
R518 VDD.n215 VDD.n210 0.145
R519 VDD.n219 VDD.n215 0.145
R520 VDD.n239 VDD.n219 0.145
R521 VDD VDD.n239 0.145
R522 VDD VDD.n468 0.145
R523 VDD.n468 VDD.n458 0.145
R524 VDD.n458 VDD.n454 0.145
R525 VDD.n454 VDD.n450 0.145
R526 VDD.n450 VDD.n446 0.145
R527 VDD.n446 VDD.n440 0.145
R528 VDD.n436 VDD.n432 0.145
R529 VDD.n432 VDD.n426 0.145
R530 VDD.n426 VDD.n422 0.145
R531 VDD.n422 VDD.n417 0.145
R532 VDD.n417 VDD.n413 0.145
R533 VDD.n387 VDD.n383 0.145
R534 VDD.n383 VDD.n379 0.145
R535 VDD.n379 VDD.n375 0.145
R536 VDD.n375 VDD.n371 0.145
R537 VDD.n371 VDD.n365 0.145
R538 VDD.n361 VDD.n357 0.145
R539 VDD.n357 VDD.n351 0.145
R540 VDD.n351 VDD.n347 0.145
R541 VDD.n347 VDD.n342 0.145
R542 VDD.n342 VDD.n338 0.145
R543 VDD.n311 VDD.n307 0.145
R544 VDD.n307 VDD.n303 0.145
R545 VDD.n303 VDD.n299 0.145
R546 VDD.n299 VDD.n295 0.145
R547 VDD.n295 VDD.n289 0.145
R548 VDD.n285 VDD.n281 0.145
R549 VDD.n281 VDD.n275 0.145
R550 VDD.n275 VDD.n271 0.145
R551 VDD.n271 VDD.n266 0.145
R552 VDD.n266 VDD.n262 0.145
R553 a_599_989.n1 a_599_989.t12 512.525
R554 a_599_989.n3 a_599_989.t11 454.685
R555 a_599_989.n3 a_599_989.t9 428.979
R556 a_599_989.n1 a_599_989.t8 371.139
R557 a_599_989.n2 a_599_989.t7 361.392
R558 a_599_989.n7 a_599_989.n6 329.955
R559 a_599_989.n4 a_599_989.t10 311.683
R560 a_599_989.n2 a_599_989.n1 235.554
R561 a_599_989.n8 a_599_989.n7 179.199
R562 a_599_989.n4 a_599_989.n3 171.288
R563 a_599_989.n10 a_599_989.n9 161.352
R564 a_599_989.n8 a_599_989.n0 95.095
R565 a_599_989.n11 a_599_989.n10 95.094
R566 a_599_989.n10 a_599_989.n8 66.258
R567 a_599_989.n0 a_599_989.t0 14.282
R568 a_599_989.n0 a_599_989.t1 14.282
R569 a_599_989.n9 a_599_989.t3 14.282
R570 a_599_989.n9 a_599_989.t4 14.282
R571 a_599_989.n11 a_599_989.t5 14.282
R572 a_599_989.t6 a_599_989.n11 14.282
R573 a_599_989.n5 a_599_989.n2 13.038
R574 a_599_989.n5 a_599_989.n4 8.685
R575 a_599_989.n7 a_599_989.n5 4.65
R576 a_3939_103.t0 a_3939_103.n0 117.777
R577 a_3939_103.n2 a_3939_103.n1 66.629
R578 a_3939_103.t0 a_3939_103.n8 59.616
R579 a_3939_103.n5 a_3939_103.n3 54.496
R580 a_3939_103.n5 a_3939_103.n4 54.496
R581 a_3939_103.t0 a_3939_103.n2 20.262
R582 a_3939_103.n7 a_3939_103.n6 2.455
R583 a_3939_103.n7 a_3939_103.n5 0.636
R584 a_3939_103.t0 a_3939_103.n7 0.246
R585 GND.n164 GND.n163 237.558
R586 GND.n248 GND.n247 237.558
R587 GND.n206 GND.n205 237.558
R588 GND.n87 GND.n86 237.558
R589 GND.n43 GND.n42 237.558
R590 GND.n40 GND.n39 210.82
R591 GND.n166 GND.n165 210.82
R592 GND.n208 GND.n207 210.82
R593 GND.n245 GND.n244 210.82
R594 GND.n84 GND.n83 210.82
R595 GND.n116 GND.n115 173.365
R596 GND.n217 GND.n216 173.365
R597 GND.n175 GND.n174 173.365
R598 GND.n133 GND.n132 173.365
R599 GND.n74 GND.n73 167.358
R600 GND.n30 GND.n29 152.358
R601 GND.n29 GND.n28 28.421
R602 GND.n29 GND.n27 25.263
R603 GND.n27 GND.n26 24.383
R604 GND.n73 GND.n71 23.03
R605 GND.n41 GND.n40 18.953
R606 GND.n167 GND.n166 18.953
R607 GND.n209 GND.n208 18.953
R608 GND.n246 GND.n245 18.953
R609 GND.n85 GND.n84 18.953
R610 GND.n44 GND.n41 14.864
R611 GND.n88 GND.n85 14.864
R612 GND.n249 GND.n246 14.864
R613 GND.n210 GND.n209 14.864
R614 GND.n168 GND.n167 14.864
R615 GND.n129 GND.n128 9.154
R616 GND.n134 GND.n131 9.154
R617 GND.n137 GND.n136 9.154
R618 GND.n140 GND.n139 9.154
R619 GND.n143 GND.n142 9.154
R620 GND.n146 GND.n145 9.154
R621 GND.n149 GND.n148 9.154
R622 GND.n152 GND.n151 9.154
R623 GND.n155 GND.n154 9.154
R624 GND.n158 GND.n157 9.154
R625 GND.n161 GND.n160 9.154
R626 GND.n168 GND.n164 9.154
R627 GND.n171 GND.n170 9.154
R628 GND.n176 GND.n173 9.154
R629 GND.n179 GND.n178 9.154
R630 GND.n182 GND.n181 9.154
R631 GND.n185 GND.n184 9.154
R632 GND.n188 GND.n187 9.154
R633 GND.n191 GND.n190 9.154
R634 GND.n194 GND.n193 9.154
R635 GND.n197 GND.n196 9.154
R636 GND.n200 GND.n199 9.154
R637 GND.n203 GND.n202 9.154
R638 GND.n210 GND.n206 9.154
R639 GND.n213 GND.n212 9.154
R640 GND.n218 GND.n215 9.154
R641 GND.n221 GND.n220 9.154
R642 GND.n224 GND.n223 9.154
R643 GND.n227 GND.n226 9.154
R644 GND.n230 GND.n229 9.154
R645 GND.n233 GND.n232 9.154
R646 GND.n236 GND.n235 9.154
R647 GND.n239 GND.n238 9.154
R648 GND.n242 GND.n241 9.154
R649 GND.n249 GND.n248 9.154
R650 GND.n123 GND.n122 9.154
R651 GND.n120 GND.n119 9.154
R652 GND.n117 GND.n114 9.154
R653 GND.n112 GND.n111 9.154
R654 GND.n109 GND.n108 9.154
R655 GND.n106 GND.n105 9.154
R656 GND.n103 GND.n102 9.154
R657 GND.n100 GND.n99 9.154
R658 GND.n97 GND.n96 9.154
R659 GND.n94 GND.n93 9.154
R660 GND.n91 GND.n90 9.154
R661 GND.n88 GND.n87 9.154
R662 GND.n81 GND.n80 9.154
R663 GND.n78 GND.n77 9.154
R664 GND.n75 GND.n70 9.154
R665 GND.n68 GND.n67 9.154
R666 GND.n65 GND.n64 9.154
R667 GND.n62 GND.n61 9.154
R668 GND.n59 GND.n58 9.154
R669 GND.n56 GND.n55 9.154
R670 GND.n53 GND.n52 9.154
R671 GND.n50 GND.n49 9.154
R672 GND.n47 GND.n46 9.154
R673 GND.n44 GND.n43 9.154
R674 GND.n37 GND.n36 9.154
R675 GND.n34 GND.n33 9.154
R676 GND.n31 GND.n25 9.154
R677 GND.n23 GND.n22 9.154
R678 GND.n20 GND.n19 9.154
R679 GND.n17 GND.n16 9.154
R680 GND.n14 GND.n13 9.154
R681 GND.n11 GND.n10 9.154
R682 GND.n8 GND.n7 9.154
R683 GND.n5 GND.n4 9.154
R684 GND.n2 GND.n1 9.154
R685 GND.n73 GND.n72 8.128
R686 GND.n127 GND.n126 4.65
R687 GND.n6 GND.n5 4.65
R688 GND.n9 GND.n8 4.65
R689 GND.n12 GND.n11 4.65
R690 GND.n15 GND.n14 4.65
R691 GND.n18 GND.n17 4.65
R692 GND.n21 GND.n20 4.65
R693 GND.n24 GND.n23 4.65
R694 GND.n32 GND.n31 4.65
R695 GND.n35 GND.n34 4.65
R696 GND.n38 GND.n37 4.65
R697 GND.n45 GND.n44 4.65
R698 GND.n48 GND.n47 4.65
R699 GND.n51 GND.n50 4.65
R700 GND.n54 GND.n53 4.65
R701 GND.n57 GND.n56 4.65
R702 GND.n60 GND.n59 4.65
R703 GND.n63 GND.n62 4.65
R704 GND.n66 GND.n65 4.65
R705 GND.n69 GND.n68 4.65
R706 GND.n76 GND.n75 4.65
R707 GND.n79 GND.n78 4.65
R708 GND.n82 GND.n81 4.65
R709 GND.n89 GND.n88 4.65
R710 GND.n92 GND.n91 4.65
R711 GND.n95 GND.n94 4.65
R712 GND.n98 GND.n97 4.65
R713 GND.n101 GND.n100 4.65
R714 GND.n104 GND.n103 4.65
R715 GND.n107 GND.n106 4.65
R716 GND.n110 GND.n109 4.65
R717 GND.n113 GND.n112 4.65
R718 GND.n118 GND.n117 4.65
R719 GND.n121 GND.n120 4.65
R720 GND.n124 GND.n123 4.65
R721 GND.n250 GND.n249 4.65
R722 GND.n243 GND.n242 4.65
R723 GND.n240 GND.n239 4.65
R724 GND.n237 GND.n236 4.65
R725 GND.n234 GND.n233 4.65
R726 GND.n231 GND.n230 4.65
R727 GND.n228 GND.n227 4.65
R728 GND.n225 GND.n224 4.65
R729 GND.n222 GND.n221 4.65
R730 GND.n219 GND.n218 4.65
R731 GND.n214 GND.n213 4.65
R732 GND.n211 GND.n210 4.65
R733 GND.n204 GND.n203 4.65
R734 GND.n201 GND.n200 4.65
R735 GND.n198 GND.n197 4.65
R736 GND.n195 GND.n194 4.65
R737 GND.n192 GND.n191 4.65
R738 GND.n189 GND.n188 4.65
R739 GND.n186 GND.n185 4.65
R740 GND.n183 GND.n182 4.65
R741 GND.n180 GND.n179 4.65
R742 GND.n177 GND.n176 4.65
R743 GND.n172 GND.n171 4.65
R744 GND.n169 GND.n168 4.65
R745 GND.n162 GND.n161 4.65
R746 GND.n159 GND.n158 4.65
R747 GND.n156 GND.n155 4.65
R748 GND.n153 GND.n152 4.65
R749 GND.n150 GND.n149 4.65
R750 GND.n147 GND.n146 4.65
R751 GND.n144 GND.n143 4.65
R752 GND.n141 GND.n140 4.65
R753 GND.n138 GND.n137 4.65
R754 GND.n135 GND.n134 4.65
R755 GND.n130 GND.n129 4.65
R756 GND.n3 GND.n0 3.407
R757 GND.n3 GND.n2 2.844
R758 GND.n6 GND.n3 1.063
R759 GND.n126 GND.n125 0.474
R760 GND.n45 GND.n38 0.29
R761 GND.n89 GND.n82 0.29
R762 GND.n211 GND.n204 0.29
R763 GND.n169 GND.n162 0.29
R764 GND.n127 GND 0.207
R765 GND.n31 GND.n30 0.206
R766 GND.n75 GND.n74 0.206
R767 GND.n117 GND.n116 0.206
R768 GND.n218 GND.n217 0.206
R769 GND.n176 GND.n175 0.206
R770 GND.n134 GND.n133 0.206
R771 GND.n18 GND.n15 0.197
R772 GND.n63 GND.n60 0.197
R773 GND.n107 GND.n104 0.197
R774 GND.n231 GND.n228 0.197
R775 GND.n189 GND.n186 0.197
R776 GND.n147 GND.n144 0.197
R777 GND.n9 GND.n6 0.145
R778 GND.n12 GND.n9 0.145
R779 GND.n15 GND.n12 0.145
R780 GND.n21 GND.n18 0.145
R781 GND.n24 GND.n21 0.145
R782 GND.n32 GND.n24 0.145
R783 GND.n35 GND.n32 0.145
R784 GND.n38 GND.n35 0.145
R785 GND.n48 GND.n45 0.145
R786 GND.n51 GND.n48 0.145
R787 GND.n54 GND.n51 0.145
R788 GND.n57 GND.n54 0.145
R789 GND.n60 GND.n57 0.145
R790 GND.n66 GND.n63 0.145
R791 GND.n69 GND.n66 0.145
R792 GND.n76 GND.n69 0.145
R793 GND.n79 GND.n76 0.145
R794 GND.n82 GND.n79 0.145
R795 GND.n92 GND.n89 0.145
R796 GND.n95 GND.n92 0.145
R797 GND.n98 GND.n95 0.145
R798 GND.n101 GND.n98 0.145
R799 GND.n104 GND.n101 0.145
R800 GND.n110 GND.n107 0.145
R801 GND.n113 GND.n110 0.145
R802 GND.n118 GND.n113 0.145
R803 GND.n121 GND.n118 0.145
R804 GND.n124 GND.n121 0.145
R805 GND GND.n124 0.145
R806 GND GND.n250 0.145
R807 GND.n250 GND.n243 0.145
R808 GND.n243 GND.n240 0.145
R809 GND.n240 GND.n237 0.145
R810 GND.n237 GND.n234 0.145
R811 GND.n234 GND.n231 0.145
R812 GND.n228 GND.n225 0.145
R813 GND.n225 GND.n222 0.145
R814 GND.n222 GND.n219 0.145
R815 GND.n219 GND.n214 0.145
R816 GND.n214 GND.n211 0.145
R817 GND.n204 GND.n201 0.145
R818 GND.n201 GND.n198 0.145
R819 GND.n198 GND.n195 0.145
R820 GND.n195 GND.n192 0.145
R821 GND.n192 GND.n189 0.145
R822 GND.n186 GND.n183 0.145
R823 GND.n183 GND.n180 0.145
R824 GND.n180 GND.n177 0.145
R825 GND.n177 GND.n172 0.145
R826 GND.n172 GND.n169 0.145
R827 GND.n162 GND.n159 0.145
R828 GND.n159 GND.n156 0.145
R829 GND.n156 GND.n153 0.145
R830 GND.n153 GND.n150 0.145
R831 GND.n150 GND.n147 0.145
R832 GND.n144 GND.n141 0.145
R833 GND.n141 GND.n138 0.145
R834 GND.n138 GND.n135 0.145
R835 GND.n135 GND.n130 0.145
R836 GND.n130 GND.n127 0.145
R837 a_277_1050.n2 a_277_1050.t8 512.525
R838 a_277_1050.n0 a_277_1050.t7 512.525
R839 a_277_1050.n2 a_277_1050.t9 371.139
R840 a_277_1050.n0 a_277_1050.t10 371.139
R841 a_277_1050.n3 a_277_1050.t12 306.051
R842 a_277_1050.n1 a_277_1050.t11 306.051
R843 a_277_1050.n3 a_277_1050.n2 290.895
R844 a_277_1050.n1 a_277_1050.n0 290.895
R845 a_277_1050.n9 a_277_1050.n8 252.875
R846 a_277_1050.n13 a_277_1050.n9 234.54
R847 a_277_1050.n12 a_277_1050.n11 161.352
R848 a_277_1050.n12 a_277_1050.n10 95.095
R849 a_277_1050.n14 a_277_1050.n13 95.094
R850 a_277_1050.n13 a_277_1050.n12 66.258
R851 a_277_1050.n8 a_277_1050.n7 30
R852 a_277_1050.n6 a_277_1050.n5 24.383
R853 a_277_1050.n8 a_277_1050.n6 23.684
R854 a_277_1050.n10 a_277_1050.t3 14.282
R855 a_277_1050.n10 a_277_1050.t2 14.282
R856 a_277_1050.n11 a_277_1050.t0 14.282
R857 a_277_1050.n11 a_277_1050.t1 14.282
R858 a_277_1050.t6 a_277_1050.n14 14.282
R859 a_277_1050.n14 a_277_1050.t5 14.282
R860 a_277_1050.n4 a_277_1050.n1 8.141
R861 a_277_1050.n9 a_277_1050.n4 5.965
R862 a_277_1050.n4 a_277_1050.n3 4.65
R863 a_2201_1050.n2 a_2201_1050.t9 512.525
R864 a_2201_1050.n2 a_2201_1050.t7 371.139
R865 a_2201_1050.n3 a_2201_1050.t8 305.674
R866 a_2201_1050.n3 a_2201_1050.n2 291.272
R867 a_2201_1050.n5 a_2201_1050.n4 274.237
R868 a_2201_1050.n6 a_2201_1050.n5 234.917
R869 a_2201_1050.n8 a_2201_1050.n7 161.352
R870 a_2201_1050.n6 a_2201_1050.n1 95.095
R871 a_2201_1050.n7 a_2201_1050.n0 95.095
R872 a_2201_1050.n7 a_2201_1050.n6 66.258
R873 a_2201_1050.n1 a_2201_1050.t5 14.282
R874 a_2201_1050.n1 a_2201_1050.t2 14.282
R875 a_2201_1050.n0 a_2201_1050.t6 14.282
R876 a_2201_1050.n0 a_2201_1050.t1 14.282
R877 a_2201_1050.t4 a_2201_1050.n8 14.282
R878 a_2201_1050.n8 a_2201_1050.t3 14.282
R879 a_2201_1050.n5 a_2201_1050.n3 10.615
R880 a_1561_989.n3 a_1561_989.t12 454.685
R881 a_1561_989.n5 a_1561_989.t7 454.685
R882 a_1561_989.n1 a_1561_989.t14 454.685
R883 a_1561_989.n3 a_1561_989.t8 428.979
R884 a_1561_989.n5 a_1561_989.t9 428.979
R885 a_1561_989.n1 a_1561_989.t10 428.979
R886 a_1561_989.n10 a_1561_989.n9 357.814
R887 a_1561_989.n4 a_1561_989.t11 339.542
R888 a_1561_989.n2 a_1561_989.t15 339.542
R889 a_1561_989.n6 a_1561_989.t13 339.186
R890 a_1561_989.n13 a_1561_989.n12 161.352
R891 a_1561_989.n11 a_1561_989.n10 151.34
R892 a_1561_989.n4 a_1561_989.n3 143.429
R893 a_1561_989.n2 a_1561_989.n1 143.429
R894 a_1561_989.n6 a_1561_989.n5 143.074
R895 a_1561_989.n11 a_1561_989.n0 95.095
R896 a_1561_989.n14 a_1561_989.n13 95.094
R897 a_1561_989.n13 a_1561_989.n11 66.258
R898 a_1561_989.n0 a_1561_989.t1 14.282
R899 a_1561_989.n0 a_1561_989.t0 14.282
R900 a_1561_989.n12 a_1561_989.t5 14.282
R901 a_1561_989.n12 a_1561_989.t6 14.282
R902 a_1561_989.t4 a_1561_989.n14 14.282
R903 a_1561_989.n14 a_1561_989.t3 14.282
R904 a_1561_989.n8 a_1561_989.n2 11.134
R905 a_1561_989.n7 a_1561_989.n6 8.145
R906 a_1561_989.n7 a_1561_989.n4 4.65
R907 a_1561_989.n10 a_1561_989.n8 4.65
R908 a_1561_989.n8 a_1561_989.n7 4.035
R909 RN.n5 RN.t0 479.223
R910 RN.n0 RN.t5 479.223
R911 RN.n2 RN.t4 454.685
R912 RN.n2 RN.t1 428.979
R913 RN.n5 RN.t3 375.52
R914 RN.n0 RN.t2 375.52
R915 RN.n6 RN.t6 371.148
R916 RN.n1 RN.t8 371.148
R917 RN.n3 RN.t7 367.4
R918 RN.n3 RN.n2 115.571
R919 RN.n6 RN.n5 112.894
R920 RN.n1 RN.n0 112.894
R921 RN.n7 RN.n4 11.381
R922 RN.n4 RN.n1 7.325
R923 RN.n4 RN.n3 4.65
R924 RN.n7 RN.n6 4.65
R925 RN.n7 RN 0.046
R926 a_1053_103.n5 a_1053_103.n4 66.708
R927 a_1053_103.n2 a_1053_103.n0 32.662
R928 a_1053_103.n5 a_1053_103.n3 19.496
R929 a_1053_103.t0 a_1053_103.n5 13.756
R930 a_1053_103.t0 a_1053_103.n2 3.034
R931 a_1053_103.n2 a_1053_103.n1 0.443
R932 a_1334_210.n10 a_1334_210.n8 171.558
R933 a_1334_210.n8 a_1334_210.t1 75.764
R934 a_1334_210.n11 a_1334_210.n0 49.6
R935 a_1334_210.n3 a_1334_210.n2 27.476
R936 a_1334_210.n10 a_1334_210.n9 27.2
R937 a_1334_210.n11 a_1334_210.n10 22.4
R938 a_1334_210.t1 a_1334_210.n5 20.241
R939 a_1334_210.n7 a_1334_210.n6 19.952
R940 a_1334_210.t1 a_1334_210.n3 13.984
R941 a_1334_210.n5 a_1334_210.n4 13.494
R942 a_1334_210.t1 a_1334_210.n1 7.04
R943 a_1334_210.n8 a_1334_210.n7 1.505
R944 a_2977_103.t0 a_2977_103.n7 59.616
R945 a_2977_103.n4 a_2977_103.n2 54.496
R946 a_2977_103.n4 a_2977_103.n3 54.496
R947 a_2977_103.n1 a_2977_103.n0 24.679
R948 a_2977_103.n6 a_2977_103.n4 7.859
R949 a_2977_103.t0 a_2977_103.n1 7.505
R950 a_2977_103.t0 a_2977_103.n6 3.034
R951 a_2977_103.n6 a_2977_103.n5 0.443
R952 a_3258_210.n8 a_3258_210.n6 185.173
R953 a_3258_210.t0 a_3258_210.n8 75.765
R954 a_3258_210.n3 a_3258_210.n1 74.827
R955 a_3258_210.n3 a_3258_210.n2 27.476
R956 a_3258_210.n6 a_3258_210.n5 22.349
R957 a_3258_210.t0 a_3258_210.n10 20.241
R958 a_3258_210.t0 a_3258_210.n3 13.984
R959 a_3258_210.n10 a_3258_210.n9 13.494
R960 a_3258_210.n6 a_3258_210.n4 8.443
R961 a_3258_210.t0 a_3258_210.n0 8.137
R962 a_3258_210.n8 a_3258_210.n7 1.505
R963 SN.n2 SN.t1 479.223
R964 SN.n0 SN.t2 479.223
R965 SN.n2 SN.t3 375.52
R966 SN.n0 SN.t4 375.52
R967 SN.n1 SN.n0 252.188
R968 SN.n3 SN.n2 251.811
R969 SN.n3 SN.t5 232.231
R970 SN.n1 SN.t0 231.854
R971 SN.n4 SN.n1 15.211
R972 SN.n4 SN.n3 4.65
R973 SN.n4 SN 0.046
R974 a_4901_103.n5 a_4901_103.n4 66.708
R975 a_4901_103.n2 a_4901_103.n0 32.662
R976 a_4901_103.n5 a_4901_103.n3 19.496
R977 a_4901_103.t0 a_4901_103.n5 13.756
R978 a_4901_103.t0 a_4901_103.n2 3.034
R979 a_4901_103.n2 a_4901_103.n1 0.443
R980 a_5182_210.n12 a_5182_210.n10 171.558
R981 a_5182_210.n7 a_5182_210.n6 117.622
R982 a_5182_210.n5 a_5182_210.n4 92.5
R983 a_5182_210.n9 a_5182_210.n8 92.5
R984 a_5182_210.n10 a_5182_210.t1 75.764
R985 a_5182_210.n5 a_5182_210.n3 65.02
R986 a_5182_210.n13 a_5182_210.n0 49.6
R987 a_5182_210.n7 a_5182_210.n5 36.517
R988 a_5182_210.n3 a_5182_210.n2 35.865
R989 a_5182_210.n12 a_5182_210.n11 27.2
R990 a_5182_210.n13 a_5182_210.n12 22.4
R991 a_5182_210.n9 a_5182_210.n7 19.952
R992 a_5182_210.t1 a_5182_210.n1 7.04
R993 a_5182_210.n10 a_5182_210.n9 1.505
R994 a_4125_1050.n1 a_4125_1050.t8 512.525
R995 a_4125_1050.n1 a_4125_1050.t9 371.139
R996 a_4125_1050.n2 a_4125_1050.t7 333.533
R997 a_4125_1050.n4 a_4125_1050.n3 302.096
R998 a_4125_1050.n2 a_4125_1050.n1 263.413
R999 a_4125_1050.n5 a_4125_1050.n4 207.058
R1000 a_4125_1050.n7 a_4125_1050.n6 161.352
R1001 a_4125_1050.n5 a_4125_1050.n0 95.095
R1002 a_4125_1050.n8 a_4125_1050.n7 95.094
R1003 a_4125_1050.n7 a_4125_1050.n5 66.258
R1004 a_4125_1050.n0 a_4125_1050.t3 14.282
R1005 a_4125_1050.n0 a_4125_1050.t4 14.282
R1006 a_4125_1050.n6 a_4125_1050.t5 14.282
R1007 a_4125_1050.n6 a_4125_1050.t6 14.282
R1008 a_4125_1050.n8 a_4125_1050.t1 14.282
R1009 a_4125_1050.t2 a_4125_1050.n8 14.282
R1010 a_4125_1050.n4 a_4125_1050.n2 10.615
R1011 Q.n7 Q.t7 454.685
R1012 Q.n7 Q.t9 428.979
R1013 Q.n6 Q.n5 329.955
R1014 Q.n8 Q.t8 311.683
R1015 Q.n6 Q.n4 179.199
R1016 Q.n8 Q.n7 171.288
R1017 Q.n3 Q.n2 161.352
R1018 Q.n4 Q.n0 95.095
R1019 Q.n3 Q.n1 95.095
R1020 Q.n4 Q.n3 66.258
R1021 Q.n0 Q.t6 14.282
R1022 Q.n0 Q.t5 14.282
R1023 Q.n1 Q.t1 14.282
R1024 Q.n1 Q.t0 14.282
R1025 Q.n2 Q.t3 14.282
R1026 Q.n2 Q.t2 14.282
R1027 Q Q.n8 8.639
R1028 Q.n9 Q.n6 4.65
R1029 Q.n9 Q 0.046
R1030 a_372_210.n10 a_372_210.n8 171.558
R1031 a_372_210.n8 a_372_210.t1 75.764
R1032 a_372_210.n3 a_372_210.n2 27.476
R1033 a_372_210.n10 a_372_210.n9 27.2
R1034 a_372_210.n11 a_372_210.n0 23.498
R1035 a_372_210.n11 a_372_210.n10 22.4
R1036 a_372_210.t1 a_372_210.n5 20.241
R1037 a_372_210.n7 a_372_210.n6 19.952
R1038 a_372_210.t1 a_372_210.n3 13.984
R1039 a_372_210.n5 a_372_210.n4 13.494
R1040 a_372_210.t1 a_372_210.n1 7.04
R1041 a_372_210.n8 a_372_210.n7 1.505
R1042 D.n0 D.t2 512.525
R1043 D.n0 D.t0 371.139
R1044 D.n1 D.t1 305.674
R1045 D.n1 D.n0 291.272
R1046 D.n2 D.n1 4.65
R1047 D.n2 D 0.046
R1048 a_91_103.n5 a_91_103.n4 66.708
R1049 a_91_103.n2 a_91_103.n0 25.439
R1050 a_91_103.n5 a_91_103.n3 19.496
R1051 a_91_103.t0 a_91_103.n5 13.756
R1052 a_91_103.n2 a_91_103.n1 2.455
R1053 a_91_103.t0 a_91_103.n2 0.246
R1054 a_2296_210.n10 a_2296_210.n8 171.558
R1055 a_2296_210.n8 a_2296_210.t1 75.764
R1056 a_2296_210.n3 a_2296_210.n2 27.476
R1057 a_2296_210.n10 a_2296_210.n9 27.2
R1058 a_2296_210.n11 a_2296_210.n0 23.498
R1059 a_2296_210.n11 a_2296_210.n10 22.4
R1060 a_2296_210.t1 a_2296_210.n5 20.241
R1061 a_2296_210.n7 a_2296_210.n6 19.952
R1062 a_2296_210.t1 a_2296_210.n3 13.984
R1063 a_2296_210.n5 a_2296_210.n4 13.494
R1064 a_2296_210.t1 a_2296_210.n1 7.04
R1065 a_2296_210.n8 a_2296_210.n7 1.505
R1066 a_4220_210.n10 a_4220_210.n8 171.558
R1067 a_4220_210.n8 a_4220_210.t1 75.764
R1068 a_4220_210.n11 a_4220_210.n0 49.6
R1069 a_4220_210.n3 a_4220_210.n2 27.476
R1070 a_4220_210.n10 a_4220_210.n9 27.2
R1071 a_4220_210.n11 a_4220_210.n10 22.4
R1072 a_4220_210.t1 a_4220_210.n5 20.241
R1073 a_4220_210.n7 a_4220_210.n6 19.952
R1074 a_4220_210.t1 a_4220_210.n3 13.984
R1075 a_4220_210.n5 a_4220_210.n4 13.494
R1076 a_4220_210.t1 a_4220_210.n1 7.04
R1077 a_4220_210.n8 a_4220_210.n7 1.505
R1078 a_2015_103.t0 a_2015_103.n7 59.616
R1079 a_2015_103.n4 a_2015_103.n2 54.496
R1080 a_2015_103.n4 a_2015_103.n3 54.496
R1081 a_2015_103.n1 a_2015_103.n0 24.679
R1082 a_2015_103.t0 a_2015_103.n1 7.505
R1083 a_2015_103.n6 a_2015_103.n5 2.455
R1084 a_2015_103.n6 a_2015_103.n4 0.636
R1085 a_2015_103.t0 a_2015_103.n6 0.246
C11 SN GND 1.67fF
C12 VDD GND 9.61fF
C13 a_2015_103.n0 GND 0.08fF
C14 a_2015_103.n1 GND 0.07fF
C15 a_2015_103.n2 GND 0.04fF
C16 a_2015_103.n3 GND 0.06fF
C17 a_2015_103.n4 GND 0.03fF
C18 a_2015_103.n5 GND 0.04fF
C19 a_2015_103.n7 GND 0.08fF
C20 a_4220_210.n0 GND 0.02fF
C21 a_4220_210.n1 GND 0.09fF
C22 a_4220_210.n2 GND 0.12fF
C23 a_4220_210.n3 GND 0.08fF
C24 a_4220_210.n4 GND 0.08fF
C25 a_4220_210.n5 GND 0.02fF
C26 a_4220_210.t1 GND 0.29fF
C27 a_4220_210.n6 GND 0.09fF
C28 a_4220_210.n7 GND 0.02fF
C29 a_4220_210.n8 GND 0.13fF
C30 a_4220_210.n9 GND 0.02fF
C31 a_4220_210.n10 GND 0.03fF
C32 a_4220_210.n11 GND 0.02fF
C33 a_2296_210.n0 GND 0.02fF
C34 a_2296_210.n1 GND 0.09fF
C35 a_2296_210.n2 GND 0.12fF
C36 a_2296_210.n3 GND 0.08fF
C37 a_2296_210.n4 GND 0.08fF
C38 a_2296_210.n5 GND 0.02fF
C39 a_2296_210.t1 GND 0.29fF
C40 a_2296_210.n6 GND 0.09fF
C41 a_2296_210.n7 GND 0.02fF
C42 a_2296_210.n8 GND 0.13fF
C43 a_2296_210.n9 GND 0.02fF
C44 a_2296_210.n10 GND 0.03fF
C45 a_2296_210.n11 GND 0.03fF
C46 a_91_103.n0 GND 0.10fF
C47 a_91_103.n1 GND 0.03fF
C48 a_91_103.n2 GND 0.03fF
C49 a_91_103.n3 GND 0.07fF
C50 a_91_103.n4 GND 0.08fF
C51 a_91_103.n5 GND 0.03fF
C52 a_372_210.n0 GND 0.02fF
C53 a_372_210.n1 GND 0.09fF
C54 a_372_210.n2 GND 0.12fF
C55 a_372_210.n3 GND 0.08fF
C56 a_372_210.n4 GND 0.08fF
C57 a_372_210.n5 GND 0.02fF
C58 a_372_210.t1 GND 0.29fF
C59 a_372_210.n6 GND 0.09fF
C60 a_372_210.n7 GND 0.02fF
C61 a_372_210.n8 GND 0.13fF
C62 a_372_210.n9 GND 0.02fF
C63 a_372_210.n10 GND 0.03fF
C64 a_372_210.n11 GND 0.03fF
C65 Q.n0 GND 0.38fF
C66 Q.n1 GND 0.38fF
C67 Q.n2 GND 0.48fF
C68 Q.n3 GND 0.46fF
C69 Q.n4 GND 0.44fF
C70 Q.n5 GND 0.33fF
C71 Q.n6 GND 0.52fF
C72 Q.n7 GND 0.32fF
C73 Q.t8 GND 0.52fF
C74 Q.n8 GND 0.61fF
C75 Q.n9 GND 0.03fF
C76 a_4125_1050.n0 GND 0.33fF
C77 a_4125_1050.n1 GND 0.29fF
C78 a_4125_1050.n2 GND 0.54fF
C79 a_4125_1050.n3 GND 0.26fF
C80 a_4125_1050.n4 GND 0.60fF
C81 a_4125_1050.n5 GND 0.40fF
C82 a_4125_1050.n6 GND 0.41fF
C83 a_4125_1050.n7 GND 0.39fF
C84 a_4125_1050.n8 GND 0.33fF
C85 a_5182_210.n0 GND 0.02fF
C86 a_5182_210.n1 GND 0.09fF
C87 a_5182_210.n2 GND 0.09fF
C88 a_5182_210.n3 GND 0.07fF
C89 a_5182_210.n4 GND 0.04fF
C90 a_5182_210.n5 GND 0.08fF
C91 a_5182_210.n6 GND 0.09fF
C92 a_5182_210.n7 GND 0.04fF
C93 a_5182_210.n8 GND 0.02fF
C94 a_5182_210.n9 GND 0.01fF
C95 a_5182_210.n10 GND 0.13fF
C96 a_5182_210.n11 GND 0.02fF
C97 a_5182_210.n12 GND 0.03fF
C98 a_5182_210.n13 GND 0.02fF
C99 a_4901_103.n0 GND 0.13fF
C100 a_4901_103.n1 GND 0.04fF
C101 a_4901_103.n2 GND 0.09fF
C102 a_4901_103.n3 GND 0.07fF
C103 a_4901_103.n4 GND 0.08fF
C104 a_4901_103.n5 GND 0.03fF
C105 SN.n0 GND 0.47fF
C106 SN.t0 GND 0.51fF
C107 SN.n1 GND 1.35fF
C108 SN.n2 GND 0.47fF
C109 SN.t5 GND 0.51fF
C110 SN.n3 GND 0.43fF
C111 SN.n4 GND 1.72fF
C112 a_3258_210.n0 GND 0.07fF
C113 a_3258_210.n1 GND 0.09fF
C114 a_3258_210.n2 GND 0.12fF
C115 a_3258_210.n3 GND 0.08fF
C116 a_3258_210.n4 GND 0.02fF
C117 a_3258_210.n5 GND 0.03fF
C118 a_3258_210.n6 GND 0.05fF
C119 a_3258_210.n7 GND 0.02fF
C120 a_3258_210.n8 GND 0.14fF
C121 a_3258_210.n9 GND 0.08fF
C122 a_3258_210.n10 GND 0.02fF
C123 a_3258_210.t0 GND 0.31fF
C124 a_2977_103.n0 GND 0.08fF
C125 a_2977_103.n1 GND 0.07fF
C126 a_2977_103.n2 GND 0.04fF
C127 a_2977_103.n3 GND 0.06fF
C128 a_2977_103.n4 GND 0.11fF
C129 a_2977_103.n5 GND 0.04fF
C130 a_2977_103.n7 GND 0.08fF
C131 a_1334_210.n0 GND 0.02fF
C132 a_1334_210.n1 GND 0.09fF
C133 a_1334_210.n2 GND 0.12fF
C134 a_1334_210.n3 GND 0.08fF
C135 a_1334_210.n4 GND 0.08fF
C136 a_1334_210.n5 GND 0.02fF
C137 a_1334_210.t1 GND 0.29fF
C138 a_1334_210.n6 GND 0.09fF
C139 a_1334_210.n7 GND 0.02fF
C140 a_1334_210.n8 GND 0.13fF
C141 a_1334_210.n9 GND 0.02fF
C142 a_1334_210.n10 GND 0.03fF
C143 a_1334_210.n11 GND 0.02fF
C144 a_1053_103.n0 GND 0.13fF
C145 a_1053_103.n1 GND 0.04fF
C146 a_1053_103.n2 GND 0.09fF
C147 a_1053_103.n3 GND 0.07fF
C148 a_1053_103.n4 GND 0.08fF
C149 a_1053_103.n5 GND 0.03fF
C150 RN.n0 GND 0.43fF
C151 RN.t8 GND 0.83fF
C152 RN.n1 GND 0.78fF
C153 RN.n2 GND 0.41fF
C154 RN.t7 GND 0.84fF
C155 RN.n3 GND 0.60fF
C156 RN.n4 GND 2.61fF
C157 RN.n5 GND 0.43fF
C158 RN.t6 GND 0.83fF
C159 RN.n6 GND 0.61fF
C160 RN.n7 GND 1.87fF
C161 a_1561_989.n0 GND 0.54fF
C162 a_1561_989.n1 GND 0.42fF
C163 a_1561_989.n2 GND 1.18fF
C164 a_1561_989.n3 GND 0.42fF
C165 a_1561_989.t11 GND 0.77fF
C166 a_1561_989.n4 GND 0.57fF
C167 a_1561_989.n5 GND 0.42fF
C168 a_1561_989.t13 GND 0.77fF
C169 a_1561_989.n6 GND 0.83fF
C170 a_1561_989.n7 GND 1.52fF
C171 a_1561_989.n8 GND 2.08fF
C172 a_1561_989.n9 GND 0.51fF
C173 a_1561_989.n10 GND 0.75fF
C174 a_1561_989.n11 GND 0.58fF
C175 a_1561_989.n12 GND 0.69fF
C176 a_1561_989.n13 GND 0.65fF
C177 a_1561_989.n14 GND 0.54fF
C178 a_2201_1050.n0 GND 0.37fF
C179 a_2201_1050.n1 GND 0.37fF
C180 a_2201_1050.n2 GND 0.35fF
C181 a_2201_1050.n3 GND 0.61fF
C182 a_2201_1050.n4 GND 0.26fF
C183 a_2201_1050.n5 GND 0.67fF
C184 a_2201_1050.n6 GND 0.48fF
C185 a_2201_1050.n7 GND 0.44fF
C186 a_2201_1050.n8 GND 0.47fF
C187 a_277_1050.n0 GND 0.33fF
C188 a_277_1050.n1 GND 0.57fF
C189 a_277_1050.n2 GND 0.33fF
C190 a_277_1050.n3 GND 0.41fF
C191 a_277_1050.n4 GND 0.82fF
C192 a_277_1050.n5 GND 0.04fF
C193 a_277_1050.n6 GND 0.05fF
C194 a_277_1050.n7 GND 0.03fF
C195 a_277_1050.n8 GND 0.15fF
C196 a_277_1050.n9 GND 0.49fF
C197 a_277_1050.n10 GND 0.34fF
C198 a_277_1050.n11 GND 0.44fF
C199 a_277_1050.n12 GND 0.41fF
C200 a_277_1050.n13 GND 0.45fF
C201 a_277_1050.n14 GND 0.34fF
C202 a_3939_103.n0 GND 0.03fF
C203 a_3939_103.n1 GND 0.09fF
C204 a_3939_103.n2 GND 0.08fF
C205 a_3939_103.n3 GND 0.04fF
C206 a_3939_103.n4 GND 0.05fF
C207 a_3939_103.n5 GND 0.03fF
C208 a_3939_103.n6 GND 0.04fF
C209 a_3939_103.n8 GND 0.08fF
C210 a_599_989.n0 GND 0.56fF
C211 a_599_989.n1 GND 0.46fF
C212 a_599_989.n2 GND 1.56fF
C213 a_599_989.n3 GND 0.47fF
C214 a_599_989.t10 GND 0.75fF
C215 a_599_989.n4 GND 0.90fF
C216 a_599_989.n5 GND 2.84fF
C217 a_599_989.n6 GND 0.48fF
C218 a_599_989.n7 GND 0.77fF
C219 a_599_989.n8 GND 0.64fF
C220 a_599_989.n9 GND 0.71fF
C221 a_599_989.n10 GND 0.67fF
C222 a_599_989.n11 GND 0.56fF
C223 VDD.n1 GND 0.03fF
C224 VDD.n2 GND 0.17fF
C225 VDD.n3 GND 0.03fF
C226 VDD.n4 GND 0.02fF
C227 VDD.n5 GND 0.06fF
C228 VDD.n6 GND 0.02fF
C229 VDD.n7 GND 0.02fF
C230 VDD.n8 GND 0.02fF
C231 VDD.n9 GND 0.02fF
C232 VDD.n10 GND 0.02fF
C233 VDD.n11 GND 0.02fF
C234 VDD.n12 GND 0.02fF
C235 VDD.n13 GND 0.02fF
C236 VDD.n14 GND 0.03fF
C237 VDD.n15 GND 0.01fF
C238 VDD.n20 GND 0.43fF
C239 VDD.n21 GND 0.26fF
C240 VDD.n22 GND 0.02fF
C241 VDD.n23 GND 0.03fF
C242 VDD.n24 GND 0.26fF
C243 VDD.n25 GND 0.01fF
C244 VDD.n26 GND 0.02fF
C245 VDD.n27 GND 0.01fF
C246 VDD.n28 GND 0.21fF
C247 VDD.n29 GND 0.01fF
C248 VDD.n30 GND 0.07fF
C249 VDD.n31 GND 0.07fF
C250 VDD.n32 GND 0.16fF
C251 VDD.n33 GND 0.01fF
C252 VDD.n34 GND 0.02fF
C253 VDD.n35 GND 0.02fF
C254 VDD.n36 GND 0.15fF
C255 VDD.n37 GND 0.01fF
C256 VDD.n38 GND 0.08fF
C257 VDD.n39 GND 0.05fF
C258 VDD.n40 GND 0.02fF
C259 VDD.n41 GND 0.02fF
C260 VDD.n42 GND 0.14fF
C261 VDD.n43 GND 0.01fF
C262 VDD.n44 GND 0.02fF
C263 VDD.n45 GND 0.03fF
C264 VDD.n46 GND 0.14fF
C265 VDD.n47 GND 0.01fF
C266 VDD.n48 GND 0.02fF
C267 VDD.n49 GND 0.03fF
C268 VDD.n50 GND 0.08fF
C269 VDD.n51 GND 0.05fF
C270 VDD.n52 GND 0.15fF
C271 VDD.n53 GND 0.01fF
C272 VDD.n54 GND 0.02fF
C273 VDD.n55 GND 0.02fF
C274 VDD.n56 GND 0.16fF
C275 VDD.n57 GND 0.01fF
C276 VDD.n58 GND 0.02fF
C277 VDD.n59 GND 0.02fF
C278 VDD.n60 GND 0.06fF
C279 VDD.n61 GND 0.21fF
C280 VDD.n62 GND 0.01fF
C281 VDD.n63 GND 0.01fF
C282 VDD.n64 GND 0.02fF
C283 VDD.n65 GND 0.26fF
C284 VDD.n66 GND 0.01fF
C285 VDD.n67 GND 0.02fF
C286 VDD.n68 GND 0.02fF
C287 VDD.n69 GND 0.26fF
C288 VDD.n70 GND 0.01fF
C289 VDD.n71 GND 0.02fF
C290 VDD.n72 GND 0.03fF
C291 VDD.n73 GND 0.05fF
C292 VDD.n74 GND 0.02fF
C293 VDD.n75 GND 0.02fF
C294 VDD.n76 GND 0.02fF
C295 VDD.n77 GND 0.02fF
C296 VDD.n78 GND 0.02fF
C297 VDD.n79 GND 0.02fF
C298 VDD.n80 GND 0.02fF
C299 VDD.n81 GND 0.02fF
C300 VDD.n82 GND 0.02fF
C301 VDD.n83 GND 0.02fF
C302 VDD.n84 GND 0.02fF
C303 VDD.n85 GND 0.03fF
C304 VDD.n86 GND 0.02fF
C305 VDD.n87 GND 0.29fF
C306 VDD.n88 GND 0.02fF
C307 VDD.n89 GND 0.02fF
C308 VDD.n91 GND 0.02fF
C309 VDD.n95 GND 0.26fF
C310 VDD.n96 GND 0.26fF
C311 VDD.n97 GND 0.01fF
C312 VDD.n98 GND 0.02fF
C313 VDD.n99 GND 0.03fF
C314 VDD.n100 GND 0.26fF
C315 VDD.n101 GND 0.01fF
C316 VDD.n102 GND 0.02fF
C317 VDD.n103 GND 0.02fF
C318 VDD.n104 GND 0.21fF
C319 VDD.n105 GND 0.01fF
C320 VDD.n106 GND 0.07fF
C321 VDD.n107 GND 0.02fF
C322 VDD.n108 GND 0.16fF
C323 VDD.n109 GND 0.01fF
C324 VDD.n110 GND 0.02fF
C325 VDD.n111 GND 0.02fF
C326 VDD.n112 GND 0.15fF
C327 VDD.n113 GND 0.01fF
C328 VDD.n114 GND 0.08fF
C329 VDD.n115 GND 0.05fF
C330 VDD.n116 GND 0.02fF
C331 VDD.n117 GND 0.02fF
C332 VDD.n118 GND 0.14fF
C333 VDD.n119 GND 0.01fF
C334 VDD.n120 GND 0.02fF
C335 VDD.n121 GND 0.03fF
C336 VDD.n122 GND 0.14fF
C337 VDD.n123 GND 0.01fF
C338 VDD.n124 GND 0.02fF
C339 VDD.n125 GND 0.03fF
C340 VDD.n126 GND 0.08fF
C341 VDD.n127 GND 0.05fF
C342 VDD.n128 GND 0.15fF
C343 VDD.n129 GND 0.01fF
C344 VDD.n130 GND 0.02fF
C345 VDD.n131 GND 0.02fF
C346 VDD.n132 GND 0.16fF
C347 VDD.n133 GND 0.01fF
C348 VDD.n134 GND 0.02fF
C349 VDD.n135 GND 0.02fF
C350 VDD.n136 GND 0.06fF
C351 VDD.n137 GND 0.21fF
C352 VDD.n138 GND 0.01fF
C353 VDD.n139 GND 0.01fF
C354 VDD.n140 GND 0.02fF
C355 VDD.n141 GND 0.26fF
C356 VDD.n142 GND 0.01fF
C357 VDD.n143 GND 0.02fF
C358 VDD.n144 GND 0.02fF
C359 VDD.n145 GND 0.26fF
C360 VDD.n146 GND 0.01fF
C361 VDD.n147 GND 0.02fF
C362 VDD.n148 GND 0.03fF
C363 VDD.n149 GND 0.29fF
C364 VDD.n150 GND 0.02fF
C365 VDD.n151 GND 0.02fF
C366 VDD.n152 GND 0.02fF
C367 VDD.n153 GND 0.06fF
C368 VDD.n154 GND 0.02fF
C369 VDD.n155 GND 0.02fF
C370 VDD.n156 GND 0.02fF
C371 VDD.n157 GND 0.02fF
C372 VDD.n158 GND 0.02fF
C373 VDD.n159 GND 0.02fF
C374 VDD.n160 GND 0.02fF
C375 VDD.n161 GND 0.02fF
C376 VDD.n162 GND 0.02fF
C377 VDD.n163 GND 0.02fF
C378 VDD.n164 GND 0.03fF
C379 VDD.n165 GND 0.02fF
C380 VDD.n166 GND 0.02fF
C381 VDD.n170 GND 0.26fF
C382 VDD.n171 GND 0.26fF
C383 VDD.n172 GND 0.01fF
C384 VDD.n173 GND 0.02fF
C385 VDD.n174 GND 0.03fF
C386 VDD.n175 GND 0.26fF
C387 VDD.n176 GND 0.01fF
C388 VDD.n177 GND 0.02fF
C389 VDD.n178 GND 0.02fF
C390 VDD.n179 GND 0.21fF
C391 VDD.n180 GND 0.01fF
C392 VDD.n181 GND 0.07fF
C393 VDD.n182 GND 0.02fF
C394 VDD.n183 GND 0.16fF
C395 VDD.n184 GND 0.01fF
C396 VDD.n185 GND 0.02fF
C397 VDD.n186 GND 0.02fF
C398 VDD.n187 GND 0.15fF
C399 VDD.n188 GND 0.01fF
C400 VDD.n189 GND 0.08fF
C401 VDD.n190 GND 0.05fF
C402 VDD.n191 GND 0.02fF
C403 VDD.n192 GND 0.02fF
C404 VDD.n193 GND 0.14fF
C405 VDD.n194 GND 0.01fF
C406 VDD.n195 GND 0.02fF
C407 VDD.n196 GND 0.03fF
C408 VDD.n197 GND 0.14fF
C409 VDD.n198 GND 0.01fF
C410 VDD.n199 GND 0.02fF
C411 VDD.n200 GND 0.03fF
C412 VDD.n201 GND 0.08fF
C413 VDD.n202 GND 0.05fF
C414 VDD.n203 GND 0.15fF
C415 VDD.n204 GND 0.01fF
C416 VDD.n205 GND 0.02fF
C417 VDD.n206 GND 0.02fF
C418 VDD.n207 GND 0.16fF
C419 VDD.n208 GND 0.01fF
C420 VDD.n209 GND 0.02fF
C421 VDD.n210 GND 0.02fF
C422 VDD.n211 GND 0.06fF
C423 VDD.n212 GND 0.21fF
C424 VDD.n213 GND 0.01fF
C425 VDD.n214 GND 0.01fF
C426 VDD.n215 GND 0.02fF
C427 VDD.n216 GND 0.26fF
C428 VDD.n217 GND 0.01fF
C429 VDD.n218 GND 0.02fF
C430 VDD.n219 GND 0.02fF
C431 VDD.n220 GND 0.29fF
C432 VDD.n221 GND 0.02fF
C433 VDD.n222 GND 0.02fF
C434 VDD.n223 GND 0.02fF
C435 VDD.n224 GND 0.06fF
C436 VDD.n225 GND 0.02fF
C437 VDD.n226 GND 0.02fF
C438 VDD.n227 GND 0.02fF
C439 VDD.n228 GND 0.02fF
C440 VDD.n229 GND 0.02fF
C441 VDD.n230 GND 0.02fF
C442 VDD.n231 GND 0.02fF
C443 VDD.n232 GND 0.02fF
C444 VDD.n233 GND 0.02fF
C445 VDD.n234 GND 0.02fF
C446 VDD.n235 GND 0.03fF
C447 VDD.n236 GND 0.26fF
C448 VDD.n237 GND 0.01fF
C449 VDD.n238 GND 0.02fF
C450 VDD.n239 GND 0.02fF
C451 VDD.n240 GND 0.17fF
C452 VDD.n241 GND 0.02fF
C453 VDD.n242 GND 0.02fF
C454 VDD.n243 GND 0.06fF
C455 VDD.n244 GND 0.02fF
C456 VDD.n245 GND 0.02fF
C457 VDD.n246 GND 0.02fF
C458 VDD.n247 GND 0.02fF
C459 VDD.n248 GND 0.02fF
C460 VDD.n249 GND 0.02fF
C461 VDD.n250 GND 0.02fF
C462 VDD.n251 GND 0.02fF
C463 VDD.n252 GND 0.03fF
C464 VDD.n253 GND 0.03fF
C465 VDD.n254 GND 0.02fF
C466 VDD.n258 GND 0.43fF
C467 VDD.n259 GND 0.26fF
C468 VDD.n260 GND 0.02fF
C469 VDD.n261 GND 0.03fF
C470 VDD.n262 GND 0.03fF
C471 VDD.n263 GND 0.26fF
C472 VDD.n264 GND 0.01fF
C473 VDD.n265 GND 0.02fF
C474 VDD.n266 GND 0.02fF
C475 VDD.n267 GND 0.06fF
C476 VDD.n268 GND 0.21fF
C477 VDD.n269 GND 0.01fF
C478 VDD.n270 GND 0.01fF
C479 VDD.n271 GND 0.02fF
C480 VDD.n272 GND 0.16fF
C481 VDD.n273 GND 0.01fF
C482 VDD.n274 GND 0.02fF
C483 VDD.n275 GND 0.02fF
C484 VDD.n276 GND 0.08fF
C485 VDD.n277 GND 0.05fF
C486 VDD.n278 GND 0.15fF
C487 VDD.n279 GND 0.01fF
C488 VDD.n280 GND 0.02fF
C489 VDD.n281 GND 0.02fF
C490 VDD.n282 GND 0.14fF
C491 VDD.n283 GND 0.01fF
C492 VDD.n284 GND 0.02fF
C493 VDD.n285 GND 0.03fF
C494 VDD.n286 GND 0.14fF
C495 VDD.n287 GND 0.01fF
C496 VDD.n288 GND 0.02fF
C497 VDD.n289 GND 0.03fF
C498 VDD.n290 GND 0.15fF
C499 VDD.n291 GND 0.01fF
C500 VDD.n292 GND 0.08fF
C501 VDD.n293 GND 0.05fF
C502 VDD.n294 GND 0.02fF
C503 VDD.n295 GND 0.02fF
C504 VDD.n296 GND 0.16fF
C505 VDD.n297 GND 0.01fF
C506 VDD.n298 GND 0.02fF
C507 VDD.n299 GND 0.02fF
C508 VDD.n300 GND 0.21fF
C509 VDD.n301 GND 0.01fF
C510 VDD.n302 GND 0.07fF
C511 VDD.n303 GND 0.02fF
C512 VDD.n304 GND 0.26fF
C513 VDD.n305 GND 0.01fF
C514 VDD.n306 GND 0.02fF
C515 VDD.n307 GND 0.02fF
C516 VDD.n308 GND 0.26fF
C517 VDD.n309 GND 0.01fF
C518 VDD.n310 GND 0.02fF
C519 VDD.n311 GND 0.03fF
C520 VDD.n312 GND 0.05fF
C521 VDD.n313 GND 0.02fF
C522 VDD.n314 GND 0.02fF
C523 VDD.n315 GND 0.02fF
C524 VDD.n316 GND 0.02fF
C525 VDD.n317 GND 0.02fF
C526 VDD.n318 GND 0.02fF
C527 VDD.n319 GND 0.02fF
C528 VDD.n320 GND 0.02fF
C529 VDD.n321 GND 0.02fF
C530 VDD.n322 GND 0.02fF
C531 VDD.n323 GND 0.02fF
C532 VDD.n324 GND 0.03fF
C533 VDD.n325 GND 0.02fF
C534 VDD.n328 GND 0.02fF
C535 VDD.n330 GND 0.02fF
C536 VDD.n331 GND 0.29fF
C537 VDD.n332 GND 0.02fF
C538 VDD.n334 GND 0.26fF
C539 VDD.n335 GND 0.26fF
C540 VDD.n336 GND 0.01fF
C541 VDD.n337 GND 0.02fF
C542 VDD.n338 GND 0.03fF
C543 VDD.n339 GND 0.26fF
C544 VDD.n340 GND 0.01fF
C545 VDD.n341 GND 0.02fF
C546 VDD.n342 GND 0.02fF
C547 VDD.n343 GND 0.06fF
C548 VDD.n344 GND 0.21fF
C549 VDD.n345 GND 0.01fF
C550 VDD.n346 GND 0.01fF
C551 VDD.n347 GND 0.02fF
C552 VDD.n348 GND 0.16fF
C553 VDD.n349 GND 0.01fF
C554 VDD.n350 GND 0.02fF
C555 VDD.n351 GND 0.02fF
C556 VDD.n352 GND 0.08fF
C557 VDD.n353 GND 0.05fF
C558 VDD.n354 GND 0.15fF
C559 VDD.n355 GND 0.01fF
C560 VDD.n356 GND 0.02fF
C561 VDD.n357 GND 0.02fF
C562 VDD.n358 GND 0.14fF
C563 VDD.n359 GND 0.01fF
C564 VDD.n360 GND 0.02fF
C565 VDD.n361 GND 0.03fF
C566 VDD.n362 GND 0.14fF
C567 VDD.n363 GND 0.01fF
C568 VDD.n364 GND 0.02fF
C569 VDD.n365 GND 0.03fF
C570 VDD.n366 GND 0.15fF
C571 VDD.n367 GND 0.01fF
C572 VDD.n368 GND 0.08fF
C573 VDD.n369 GND 0.05fF
C574 VDD.n370 GND 0.02fF
C575 VDD.n371 GND 0.02fF
C576 VDD.n372 GND 0.16fF
C577 VDD.n373 GND 0.01fF
C578 VDD.n374 GND 0.02fF
C579 VDD.n375 GND 0.02fF
C580 VDD.n376 GND 0.21fF
C581 VDD.n377 GND 0.01fF
C582 VDD.n378 GND 0.07fF
C583 VDD.n379 GND 0.02fF
C584 VDD.n380 GND 0.26fF
C585 VDD.n381 GND 0.01fF
C586 VDD.n382 GND 0.02fF
C587 VDD.n383 GND 0.02fF
C588 VDD.n384 GND 0.26fF
C589 VDD.n385 GND 0.01fF
C590 VDD.n386 GND 0.02fF
C591 VDD.n387 GND 0.03fF
C592 VDD.n388 GND 0.29fF
C593 VDD.n389 GND 0.02fF
C594 VDD.n390 GND 0.02fF
C595 VDD.n391 GND 0.02fF
C596 VDD.n392 GND 0.06fF
C597 VDD.n393 GN