* SPICE3 file created from XOR2X1.ext - technology: sky130A

.subckt XOR2X1 Y A B VDD GND
X0 GND A.t1 a_556_101.t0 GND sky130_fd_pr__nfet_01v8 ad=2.6398p pd=1.934u as=0p ps=0u w=0u l=0u
X1 a_807_990.t2 B.t0 VDD.t13 ��+�
V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X2 a_185_209.t2 A.t0 VDD.t15 @R`�
V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X3 Y a_185_209.t3 a_1222_101.t0 GND sky130_fd_pr__nfet_01v8 ad=3.582p pd=3.14u as=0p ps=0u w=0u l=0u
X4 a_575_1051.t3 a_807_990.t3 Y.t4 ��ϕ
V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X5 a_1241_1051.t3 B.t1 VDD.t11  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X6 Y B.t3 a_556_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X7 Y.t3 a_807_990.t4 a_575_1051.t2 VDD.t1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X8 a_1241_1051.t1 a_185_209.t4 Y.t0  ̻Ӿ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X9 VDD.t19 A.t3 a_575_1051.t1 �˻Ӿ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X10 VDD.t5 A.t4 a_185_209.t1  ̻Ӿ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X11 VDD.t9 B.t4 a_1241_1051.t2 �˻Ӿ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X12 GND a_807_990.t5 a_1222_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X13 a_575_1051.t0 A.t5 VDD.t17  ̻Ӿ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X14 Y.t2 a_185_209.t5 a_1241_1051.t0 �˻Ӿ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X15 VDD.t7 B.t5 a_807_990.t1  ̻Ӿ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
C0 B VDD 1.45fF
C1 B Y 0.62fF
C2 A VDD 1.26fF
C3 Y A 0.08fF
C4 Y VDD 1.04fF
C5 B A 0.04fF
R0 B.n0 B.t0 512.525
R1 B.n3 B.t1 480.392
R2 B.n3 B.t4 403.272
R3 B.n0 B.t5 371.139
R4 B.n1 B.t3 299.455
R5 B.n1 B.t2 227.134
R6 B.n2 B.n0 163.771
R7 B.n2 B.n1 139.294
R8 B B.n3 123.226
R9 B.n4 B.n2 4.65
R10 B.n4 B 0.046
R11 VDD.n172 VDD.n171 173.148
R12 VDD.n85 VDD.n84 173.148
R13 VDD.n151 VDD.n140 144.705
R14 VDD.n66 VDD.n55 144.705
R15 VDD.n96 VDD.n94 144.705
R16 VDD.n124 VDD.t15 135.17
R17 VDD.n131 VDD.t5 135.17
R18 VDD.n33 VDD.t13 135.17
R19 VDD.n24 VDD.t7 135.17
R20 VDD.n51 VDD.n50 92.5
R21 VDD.n49 VDD.n48 92.5
R22 VDD.n47 VDD.n46 92.5
R23 VDD.n45 VDD.n44 92.5
R24 VDD.n53 VDD.n52 92.5
R25 VDD.n204 VDD.n203 92.5
R26 VDD.n202 VDD.n201 92.5
R27 VDD.n200 VDD.n199 92.5
R28 VDD.n198 VDD.n197 92.5
R29 VDD.n206 VDD.n205 92.5
R30 VDD.n161 VDD.n160 92.5
R31 VDD.n159 VDD.n158 92.5
R32 VDD.n157 VDD.n156 92.5
R33 VDD.n155 VDD.n154 92.5
R34 VDD.n163 VDD.n162 92.5
R35 VDD.n110 VDD.n109 92.5
R36 VDD.n108 VDD.n107 92.5
R37 VDD.n106 VDD.n105 92.5
R38 VDD.n104 VDD.n103 92.5
R39 VDD.n112 VDD.n111 92.5
R40 VDD.n14 VDD.n1 92.5
R41 VDD.n5 VDD.n4 92.5
R42 VDD.n7 VDD.n6 92.5
R43 VDD.n9 VDD.n8 92.5
R44 VDD.n11 VDD.n10 92.5
R45 VDD.n13 VDD.n12 92.5
R46 VDD.n21 VDD.n20 92.059
R47 VDD.n65 VDD.n64 92.059
R48 VDD.n213 VDD.n212 92.059
R49 VDD.n150 VDD.n149 92.059
R50 VDD.n118 VDD.n117 92.059
R51 VDD.n20 VDD.n16 67.194
R52 VDD.n20 VDD.n17 67.194
R53 VDD.n20 VDD.n18 67.194
R54 VDD.n20 VDD.n19 67.194
R55 VDD.n102 VDD.n101 44.141
R56 VDD.n196 VDD.n195 44.141
R57 VDD.n5 VDD.n3 44.141
R58 VDD.n195 VDD.n193 44.107
R59 VDD.n101 VDD.n99 44.107
R60 VDD.n3 VDD.n2 44.107
R61 VDD.n25  ̻Ӿ 43.472
R62 VDD.n34 ��+�
V 43.472
R63 VDD.n132  ̻Ӿ 43.472
R64 VDD.n122 @R`�
V 43.472
R65 VDD.n20 VDD.n15 41.052
R66 VDD.n59 VDD.n57 39.742
R67 VDD.n59 VDD.n58 39.742
R68 VDD.n61 VDD.n60 39.742
R69 VDD.n209 VDD.n208 39.742
R70 VDD.n114 VDD.n113 39.742
R71 VDD.n148 VDD.n145 39.742
R72 VDD.n148 VDD.n147 39.742
R73 VDD.n144 VDD.n143 39.742
R74 VDD.n195 VDD.n194 38
R75 VDD.n101 VDD.n100 38
R76 VDD.n193 VDD.n192 36.774
R77 VDD.n57 VDD.n56 36.774
R78 VDD.n147 VDD.n146 36.774
R79 VDD.n1 VDD.n0 30.923
R80 VDD.n64 VDD.n62 26.38
R81 VDD.n64 VDD.n61 26.38
R82 VDD.n64 VDD.n59 26.38
R83 VDD.n64 VDD.n63 26.38
R84 VDD.n212 VDD.n210 26.38
R85 VDD.n212 VDD.n209 26.38
R86 VDD.n212 VDD.n211 26.38
R87 VDD.n117 VDD.n115 26.38
R88 VDD.n117 VDD.n114 26.38
R89 VDD.n117 VDD.n116 26.38
R90 VDD.n149 VDD.n148 26.38
R91 VDD.n149 VDD.n144 26.38
R92 VDD.n149 VDD.n142 26.38
R93 VDD.n149 VDD.n141 26.38
R94 VDD.n120 VDD.n112 22.915
R95 VDD.n23 VDD.n14 22.915
R96 VDD.n73  ̻Ӿ 20.457
R97 VDD.n184 ��ϕ
V 20.457
R98 VDD.n86 �˻Ӿ 17.9
R99 VDD.n173 �˻Ӿ 17.9
R100 VDD.n112 VDD.n110 14.864
R101 VDD.n110 VDD.n108 14.864
R102 VDD.n108 VDD.n106 14.864
R103 VDD.n106 VDD.n104 14.864
R104 VDD.n104 VDD.n102 14.864
R105 VDD.n206 VDD.n204 14.864
R106 VDD.n204 VDD.n202 14.864
R107 VDD.n202 VDD.n200 14.864
R108 VDD.n200 VDD.n198 14.864
R109 VDD.n198 VDD.n196 14.864
R110 VDD.n53 VDD.n51 14.864
R111 VDD.n51 VDD.n49 14.864
R112 VDD.n49 VDD.n47 14.864
R113 VDD.n47 VDD.n45 14.864
R114 VDD.n45 VDD.n43 14.864
R115 VDD.n43 VDD.n42 14.864
R116 VDD.n163 VDD.n161 14.864
R117 VDD.n161 VDD.n159 14.864
R118 VDD.n159 VDD.n157 14.864
R119 VDD.n157 VDD.n155 14.864
R120 VDD.n155 VDD.n153 14.864
R121 VDD.n153 VDD.n152 14.864
R122 VDD.n14 VDD.n13 14.864
R123 VDD.n13 VDD.n11 14.864
R124 VDD.n11 VDD.n9 14.864
R125 VDD.n9 VDD.n7 14.864
R126 VDD.n7 VDD.n5 14.864
R127 VDD.n67 VDD.n54 14.864
R128 VDD.n215 VDD.n207 14.864
R129 VDD.n165 VDD.n164 14.864
R130 VDD.n171 VDD.t17 14.282
R131 VDD.n171 VDD.t19 14.282
R132 VDD.n84 VDD.t11 14.282
R133 VDD.n84 VDD.t9 14.282
R134 VDD.n23 VDD.n22 8.855
R135 VDD.n22 VDD.n21 8.855
R136 VDD.n27 VDD.n26 8.855
R137 VDD.n26 VDD.n25 8.855
R138 VDD.n31 VDD.n30 8.855
R139 VDD.n30 VDD.n29 8.855
R140 VDD.n36 VDD.n35 8.855
R141 VDD.n35 VDD.n34 8.855
R142 VDD.n40 VDD.n39 8.855
R143 VDD.n39 VDD.n38 8.855
R144 VDD.n67 VDD.n66 8.855
R145 VDD.n66 VDD.n65 8.855
R146 VDD.n71 VDD.n70 8.855
R147 VDD.n70 VDD.n69 8.855
R148 VDD.n75 VDD.n74 8.855
R149 VDD.n74 VDD.n73 8.855
R150 VDD.n78 VDD.n77 8.855
R151 VDD.n77 �˻Ӿ 8.855
R152 VDD.n82 VDD.n81 8.855
R153 VDD.n81 VDD.n80 8.855
R154 VDD.n88 VDD.n87 8.855
R155 VDD.n87 VDD.n86 8.855
R156 VDD.n92 VDD.n91 8.855
R157 VDD.n91 VDD.n90 8.855
R158 VDD.n97 VDD.n96 8.855
R159 VDD.n96 VDD.n95 8.855
R160 VDD.n215 VDD.n214 8.855
R161 VDD.n214 VDD.n213 8.855
R162 VDD.n190 VDD.n189 8.855
R163 VDD.n189 VDD.n188 8.855
R164 VDD.n186 VDD.n185 8.855
R165 VDD.n185 VDD.n184 8.855
R166 VDD.n182 VDD.n181 8.855
R167 VDD.n181 VDD.t1 8.855
R168 VDD.n179 VDD.n178 8.855
R169 VDD.n178 VDD.n177 8.855
R170 VDD.n175 VDD.n174 8.855
R171 VDD.n174 VDD.n173 8.855
R172 VDD.n169 VDD.n168 8.855
R173 VDD.n168 VDD.n167 8.855
R174 VDD.n165 VDD.n151 8.855
R175 VDD.n151 VDD.n150 8.855
R176 VDD.n138 VDD.n137 8.855
R177 VDD.n137 VDD.n136 8.855
R178 VDD.n134 VDD.n133 8.855
R179 VDD.n133 VDD.n132 8.855
R180 VDD.n129 VDD.n128 8.855
R181 VDD.n128 VDD.n127 8.855
R182 VDD.n125 VDD.n123 8.855
R183 VDD.n123 VDD.n122 8.855
R184 VDD.n120 VDD.n119 8.855
R185 VDD.n119 VDD.n118 8.855
R186 VDD.n207 VDD.n206 8.051
R187 VDD.n54 VDD.n53 8.051
R188 VDD.n164 VDD.n163 8.051
R189 VDD.n88 VDD.n85 6.193
R190 VDD.n175 VDD.n172 6.193
R191 VDD.n28 VDD.n23 4.795
R192 VDD.n28 VDD.n27 4.65
R193 VDD.n32 VDD.n31 4.65
R194 VDD.n37 VDD.n36 4.65
R195 VDD.n41 VDD.n40 4.65
R196 VDD.n68 VDD.n67 4.65
R197 VDD.n72 VDD.n71 4.65
R198 VDD.n76 VDD.n75 4.65
R199 VDD.n79 VDD.n78 4.65
R200 VDD.n83 VDD.n82 4.65
R201 VDD.n89 VDD.n88 4.65
R202 VDD.n93 VDD.n92 4.65
R203 VDD.n98 VDD.n97 4.65
R204 VDD.n216 VDD.n215 4.65
R205 VDD.n191 VDD.n190 4.65
R206 VDD.n187 VDD.n186 4.65
R207 VDD.n183 VDD.n182 4.65
R208 VDD.n180 VDD.n179 4.65
R209 VDD.n176 VDD.n175 4.65
R210 VDD.n170 VDD.n169 4.65
R211 VDD.n166 VDD.n165 4.65
R212 VDD.n139 VDD.n138 4.65
R213 VDD.n135 VDD.n134 4.65
R214 VDD.n130 VDD.n129 4.65
R215 VDD.n126 VDD.n125 4.65
R216 VDD.n121 VDD.n120 4.65
R217 VDD.n80 ��C�
V 2.557
R218 VDD.n177  ̻Ӿ 2.557
R219 VDD.n27 VDD.n24 2.064
R220 VDD.n36 VDD.n33 2.064
R221 VDD.n134 VDD.n131 2.064
R222 VDD.n125 VDD.n124 2.064
R223 VDD.n68 VDD.n41 0.29
R224 VDD.n166 VDD.n139 0.29
R225 VDD.n121 VDD 0.207
R226 VDD.n83 VDD.n79 0.181
R227 VDD.n183 VDD.n180 0.181
R228 VDD.n32 VDD.n28 0.157
R229 VDD.n37 VDD.n32 0.157
R230 VDD.n135 VDD.n130 0.157
R231 VDD.n130 VDD.n126 0.157
R232 VDD.n41 VDD.n37 0.145
R233 VDD.n72 VDD.n68 0.145
R234 VDD.n76 VDD.n72 0.145
R235 VDD.n79 VDD.n76 0.145
R236 VDD.n89 VDD.n83 0.145
R237 VDD.n93 VDD.n89 0.145
R238 VDD.n98 VDD.n93 0.145
R239 VDD VDD.n98 0.145
R240 VDD VDD.n216 0.145
R241 VDD.n216 VDD.n191 0.145
R242 VDD.n191 VDD.n187 0.145
R243 VDD.n187 VDD.n183 0.145
R244 VDD.n180 VDD.n176 0.145
R245 VDD.n176 VDD.n170 0.145
R246 VDD.n170 VDD.n166 0.145
R247 VDD.n139 VDD.n135 0.145
R248 VDD.n126 VDD.n121 0.145
R249 a_807_990.n0 a_807_990.t4 477.179
R250 a_807_990.n0 a_807_990.t3 406.485
R251 a_807_990.n5 a_807_990.t5 312.917
R252 a_807_990.n5 a_807_990.n4 244.592
R253 a_807_990.n7 a_807_990.n6 215.563
R254 a_807_990.n6 a_807_990.n0 156.869
R255 a_807_990.n6 a_807_990.n5 83.576
R256 a_807_990.n4 a_807_990.n3 30
R257 a_807_990.n2 a_807_990.n1 24.383
R258 a_807_990.n4 a_807_990.n2 23.684
R259 a_807_990.n7 a_807_990.t1 14.282
R260 a_807_990.t2 a_807_990.n7 14.282
R261 A.n2 A.t4 512.525
R262 A.n0 A.t5 480.392
R263 A.n1 A.t1 412.921
R264 A.n0 A.t3 403.272
R265 A.n2 A.t0 371.139
R266 A.n3 A.t2 366.428
R267 A.n3 A.n2 163.771
R268 A.n1 A.n0 115.947
R269 A.n4 A.n1 6.509
R270 A.n4 A.n3 4.65
R271 A.n4 A 0.046
R272 a_185_209.n0 a_185_209.t5 477.179
R273 a_185_209.n0 a_185_209.t4 406.485
R274 a_185_209.n1 a_185_209.t3 341.566
R275 a_185_209.n6 a_185_209.n5 272.451
R276 a_185_209.n7 a_185_209.n6 271.281
R277 a_185_209.n1 a_185_209.n0 199.524
R278 a_185_209.n5 a_185_209.n4 30
R279 a_185_209.n3 a_185_209.n2 24.383
R280 a_185_209.n5 a_185_209.n3 23.684
R281 a_185_209.n7 a_185_209.t1 14.282
R282 a_185_209.t2 a_185_209.n7 14.282
R283 a_185_209.n6 a_185_209.n1 13.879
R284 a_556_101.t0 a_556_101.n6 93.333
R285 a_556_101.n5 a_556_101.n4 51.907
R286 a_556_101.n5 a_556_101.n3 51.594
R287 a_556_101.n2 a_556_101.n0 41.528
R288 a_556_101.t0 a_556_101.n5 38.864
R289 a_556_101.t0 a_556_101.n7 8.137
R290 a_556_101.n2 a_556_101.n1 3.644
R291 a_556_101.t0 a_556_101.n2 1.093
R292 GND.n118 GND.n117 237.558
R293 GND.n88 GND.n87 237.558
R294 GND.n29 GND.n28 237.558
R295 GND.n26 GND.n25 210.82
R296 GND.n90 GND.n89 210.82
R297 GND.n115 GND.n114 210.82
R298 GND.n98 GND.n97 172.612
R299 GND.n48 GND.n47 151.605
R300 GND.n18 GND.n17 38.384
R301 GND.n68 GND.n67 37.582
R302 GND.n4 GND.n3 34.159
R303 GND.t0 GND.n65 32.601
R304 GND.n47 GND.n46 28.421
R305 GND.n47 GND.n45 25.263
R306 GND.n45 GND.n44 24.383
R307 GND.n65 GND.n64 21.734
R308 GND.n5 GND.n4 20.705
R309 GND.n12 GND.n11 20.705
R310 GND.n19 GND.n18 20.705
R311 GND.n80 GND.n79 20.705
R312 GND.n74 GND.n73 20.705
R313 GND.n69 GND.n68 20.705
R314 GND.n79 GND.n78 19.952
R315 GND.n3 GND.n2 19.926
R316 GND.n27 GND.n26 18.953
R317 GND.n91 GND.n90 18.953
R318 GND.n116 GND.n115 18.953
R319 GND.n17 GND.t5 15.889
R320 GND.n67 GND.t0 15.644
R321 GND.n30 GND.n27 14.864
R322 GND.n119 GND.n116 14.864
R323 GND.n92 GND.n91 14.864
R324 GND.n17 GND.n16 13.624
R325 GND.n67 GND.n66 13.541
R326 GND.n70 GND.n61 9.154
R327 GND.n76 GND.n75 9.154
R328 GND.n82 GND.n81 9.154
R329 GND.n85 GND.n84 9.154
R330 GND.n92 GND.n88 9.154
R331 GND.n95 GND.n94 9.154
R332 GND.n100 GND.n99 9.154
R333 GND.n103 GND.n102 9.154
R334 GND.n106 GND.n105 9.154
R335 GND.n109 GND.n108 9.154
R336 GND.n112 GND.n111 9.154
R337 GND.n119 GND.n118 9.154
R338 GND.n56 GND.n55 9.154
R339 GND.n53 GND.n52 9.154
R340 GND.n50 GND.n49 9.154
R341 GND.n42 GND.n41 9.154
R342 GND.n39 GND.n38 9.154
R343 GND.n36 GND.n35 9.154
R344 GND.n33 GND.n32 9.154
R345 GND.n30 GND.n29 9.154
R346 GND.n23 GND.n22 9.154
R347 GND.n20 GND.n15 9.154
R348 GND.n13 GND.n9 9.154
R349 GND.n7 GND.n6 9.154
R350 GND.n8 GND.n1 4.795
R351 GND.n60 GND.n59 4.65
R352 GND.n8 GND.n7 4.65
R353 GND.n14 GND.n13 4.65
R354 GND.n21 GND.n20 4.65
R355 GND.n24 GND.n23 4.65
R356 GND.n31 GND.n30 4.65
R357 GND.n34 GND.n33 4.65
R358 GND.n37 GND.n36 4.65
R359 GND.n40 GND.n39 4.65
R360 GND.n43 GND.n42 4.65
R361 GND.n51 GND.n50 4.65
R362 GND.n54 GND.n53 4.65
R363 GND.n57 GND.n56 4.65
R364 GND.n120 GND.n119 4.65
R365 GND.n113 GND.n112 4.65
R366 GND.n110 GND.n109 4.65
R367 GND.n107 GND.n106 4.65
R368 GND.n104 GND.n103 4.65
R369 GND.n101 GND.n100 4.65
R370 GND.n96 GND.n95 4.65
R371 GND.n93 GND.n92 4.65
R372 GND.n86 GND.n85 4.65
R373 GND.n83 GND.n82 4.65
R374 GND.n77 GND.n76 4.65
R375 GND.n71 GND.n70 4.65
R376 GND.n63 GND.n62 4.504
R377 GND.n20 GND.n19 4.129
R378 GND.n50 GND.n48 4.129
R379 GND.n100 GND.n98 4.129
R380 GND.n82 GND.n80 4.129
R381 GND.n7 GND.n5 3.716
R382 GND.n70 GND.n69 3.716
R383 GND.t0 GND.n63 2.452
R384 GND.n1 GND.n0 0.474
R385 GND.n59 GND.n58 0.474
R386 GND.n11 GND.n10 0.376
R387 GND.n73 GND.n72 0.376
R388 GND.n31 GND.n24 0.29
R389 GND.n93 GND.n86 0.29
R390 GND.n60 GND 0.207
R391 GND.n13 GND.n12 0.206
R392 GND.n76 GND.n74 0.206
R393 GND.n43 GND.n40 0.181
R394 GND.n107 GND.n104 0.181
R395 GND.n14 GND.n8 0.157
R396 GND.n21 GND.n14 0.157
R397 GND.n83 GND.n77 0.157
R398 GND.n77 GND.n71 0.157
R399 GND.n24 GND.n21 0.145
R400 GND.n34 GND.n31 0.145
R401 GND.n37 GND.n34 0.145
R402 GND.n40 GND.n37 0.145
R403 GND.n51 GND.n43 0.145
R404 GND.n54 GND.n51 0.145
R405 GND.n57 GND.n54 0.145
R406 GND GND.n57 0.145
R407 GND GND.n120 0.145
R408 GND.n120 GND.n113 0.145
R409 GND.n113 GND.n110 0.145
R410 GND.n110 GND.n107 0.145
R411 GND.n104 GND.n101 0.145
R412 GND.n101 GND.n96 0.145
R413 GND.n96 GND.n93 0.145
R414 GND.n86 GND.n83 0.145
R415 GND.n71 GND.n60 0.145
R416 Y.n8 Y.n7 327.32
R417 Y.n5 Y.n4 305.581
R418 Y.n5 Y.n0 260.107
R419 Y.n8 Y.n6 260.107
R420 Y.n4 Y.n3 30
R421 Y.n2 Y.n1 24.383
R422 Y.n4 Y.n2 23.684
R423 Y.n0 Y.t0 14.282
R424 Y.n0 Y.t2 14.282
R425 Y.n6 Y.t4 14.282
R426 Y.n6 Y.t3 14.282
R427 Y Y.n8 7.007
R428 Y.n9 Y.n5 4.65
R429 Y.n9 Y 0.046
R430 a_575_1051.n1 a_575_1051.t3 228.368
R431 a_575_1051.t1 a_575_1051.n1 219.777
R432 a_575_1051.n1 a_575_1051.n0 42.29
R433 a_575_1051.n0 a_575_1051.t2 14.282
R434 a_575_1051.n0 a_575_1051.t0 14.282
R435 a_1222_101.n3 a_1222_101.n1 42.788
R436 a_1222_101.t0 a_1222_101.n0 8.137
R437 a_1222_101.n3 a_1222_101.n2 4.665
R438 a_1222_101.t0 a_1222_101.n3 0.06
R439 a_1241_1051.t1 a_1241_1051.n1 228.371
R440 a_1241_1051.n1 a_1241_1051.t2 219.777
R441 a_1241_1051.n1 a_1241_1051.n0 42.29
R442 a_1241_1051.n0 a_1241_1051.t0 14.282
R443 a_1241_1051.n0 a_1241_1051.t3 14.282
C6 VDD GND 4.24fF
C7 a_1241_1051.n0 GND 0.22fF
C8 a_1241_1051.n1 GND 0.50fF
C9 a_1222_101.n0 GND 0.05fF
C10 a_1222_101.n1 GND 0.12fF
C11 a_1222_101.n2 GND 0.04fF
C12 a_1222_101.n3 GND 0.17fF
C13 a_575_1051.n0 GND 0.22fF
C14 a_575_1051.n1 GND 0.50fF
C15 Y.n0 GND 0.88fF
C16 Y.n1 GND 0.06fF
C17 Y.n2 GND 0.09fF
C18 Y.n3 GND 0.05fF
C19 Y.n4 GND 0.36fF
C20 Y.n5 GND 1.01fF
C21 Y.n6 GND 0.88fF
C22 Y.n7 GND 0.54fF
C23 Y.n8 GND 1.19fF
C24 Y.n9 GND 0.05fF
C25 a_556_101.n0 GND 0.08fF
C26 a_556_101.n1 GND 0.02fF
C27 a_556_101.n2 GND 0.02fF
C28 a_556_101.n3 GND 0.09fF
C29 a_556_101.n4 GND 0.07fF
C30 a_556_101.n5 GND 0.04fF
C31 a_556_101.n6 GND 0.02fF
C32 a_556_101.n7 GND 0.05fF
C33 a_185_209.n0 GND 0.45fF
C34 a_185_209.n1 GND 1.24fF
C35 a_185_209.n2 GND 0.05fF
C36 a_185_209.n3 GND 0.07fF
C37 a_185_209.n4 GND 0.04fF
C38 a_185_209.n5 GND 0.24fF
C39 a_185_209.n6 GND 1.48fF
C40 a_185_209.n7 GND 0.82fF
C41 a_807_990.n0 GND 0.54fF
C42 a_807_990.n1 GND 0.06fF
C43 a_807_990.n2 GND 0.08fF
C44 a_807_990.n3 GND 0.05fF
C45 a_807_990.n4 GND 0.24fF
C46 a_807_990.n5 GND 1.64fF
C47 a_807_990.n6 GND 2.07fF
C48 a_807_990.n7 GND 0.86fF
C49 VDD.n1 GND 0.03fF
C50 VDD.n2 GND 0.09fF
C51 VDD.n3 GND 0.03fF
C52 VDD.n4 GND 0.02fF
C53 VDD.n5 GND 0.06fF
C54 VDD.n6 GND 0.02fF
C55 VDD.n7 GND 0.02fF
C56 VDD.n8 GND 0.02fF
C57 VDD.n9 GND 0.02fF
C58 VDD.n10 GND 0.02fF
C59 VDD.n11 GND 0.02fF
C60 VDD.n12 GND 0.02fF
C61 VDD.n13 GND 0.02fF
C62 VDD.n14 GND 0.03fF
C63 VDD.n15 GND 0.01fF
C64 VDD.n20 GND 0.43fF
C65 VDD.n21 GND 0.26fF
C66 VDD.n22 GND 0.02fF
C67 VDD.n23 GND 0.03fF
C68 VDD.n24 GND 0.06fF
C69 VDD.n25 GND 0.19fF
C70 VDD.n26 GND 0.01fF
C71 VDD.n27 GND 0.01fF
C72 VDD.n28 GND 0.06fF
C73 VDD.n29 GND 0.16fF
C74 VDD.n30 GND 0.01fF
C75 VDD.n31 GND 0.02fF
C76 VDD.n32 GND 0.02fF
C77 VDD.n33 GND 0.06fF
C78 VDD.n34 GND 0.19fF
C79 VDD.n35 GND 0.01fF
C80 VDD.n36 GND 0.01fF
C81 VDD.n37 GND 0.02fF
C82 VDD.n38 GND 0.26fF
C83 VDD.n39 GND 0.01fF
C84 VDD.n40 GND 0.02fF
C85 VDD.n41 GND 0.03fF
C86 VDD.n42 GND 0.05fF
C87 VDD.n43 GND 0.02fF
C88 VDD.n44 GND 0.02fF
C89 VDD.n45 GND 0.02fF
C90 VDD.n46 GN