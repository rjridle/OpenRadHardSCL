magic
tech sky130A
magscale 1 2
timestamp 1643045510
<< error_p >>
rect 85 318 86 319
rect 86 317 87 318
rect 101 287 102 288
rect 136 287 137 288
rect 101 184 102 185
rect 136 184 137 185
<< nwell >>
rect -159 612 399 1353
<< nmos >>
rect 56 318 86 368
rect 56 288 152 318
tri 152 288 182 318 sw
rect 56 184 86 288
tri 86 272 102 288 nw
tri 136 272 152 288 ne
tri 86 184 102 200 sw
tri 136 184 152 200 se
rect 152 184 182 288
tri 56 154 86 184 ne
rect 86 154 152 184
tri 152 154 182 184 nw
<< pmos >>
rect 56 829 86 1229
rect 144 829 174 1229
<< ndiff >>
rect -7 307 56 368
rect 86 318 245 368
rect -7 273 10 307
rect 44 273 56 307
tri 152 288 182 318 ne
rect 182 307 245 318
rect -7 211 56 273
rect -7 177 10 211
rect 44 177 56 211
tri 86 272 102 288 se
rect 102 272 136 288
tri 136 272 152 288 sw
rect 86 240 152 272
rect 86 206 98 240
rect 132 206 152 240
rect 86 200 152 206
tri 86 184 102 200 ne
rect 102 184 136 200
tri 136 184 152 200 nw
rect 182 273 194 307
rect 228 273 245 307
rect 182 211 245 273
rect -7 154 56 177
tri 56 154 86 184 sw
tri 152 154 182 184 se
rect 182 177 194 211
rect 228 177 245 211
rect 182 154 245 177
rect -7 143 245 154
rect -7 109 10 143
rect 44 109 98 143
rect 132 109 194 143
rect 228 109 245 143
rect -7 101 245 109
<< pdiff >>
rect 0 1213 56 1229
rect 0 1179 10 1213
rect 44 1179 56 1213
rect 0 1145 56 1179
rect 0 1111 10 1145
rect 44 1111 56 1145
rect 0 1077 56 1111
rect 0 1043 10 1077
rect 44 1043 56 1077
rect 0 1009 56 1043
rect 0 975 10 1009
rect 44 975 56 1009
rect 0 941 56 975
rect 0 907 10 941
rect 44 907 56 941
rect 0 829 56 907
rect 86 1213 144 1229
rect 86 1179 98 1213
rect 132 1179 144 1213
rect 86 1145 144 1179
rect 86 1111 98 1145
rect 132 1111 144 1145
rect 86 1077 144 1111
rect 86 1043 98 1077
rect 132 1043 144 1077
rect 86 1009 144 1043
rect 86 975 98 1009
rect 132 975 144 1009
rect 86 941 144 975
rect 86 907 98 941
rect 132 907 144 941
rect 86 829 144 907
rect 174 1213 228 1229
rect 174 1179 186 1213
rect 220 1179 228 1213
rect 174 1145 228 1179
rect 174 1111 186 1145
rect 220 1111 228 1145
rect 174 1077 228 1111
rect 174 1043 186 1077
rect 220 1043 228 1077
rect 174 1009 228 1043
rect 174 975 186 1009
rect 220 975 228 1009
rect 174 941 228 975
rect 174 907 186 941
rect 220 907 228 941
rect 174 829 228 907
<< ndiffc >>
rect 10 273 44 307
rect 10 177 44 211
rect 98 206 132 240
rect 194 273 228 307
rect 194 177 228 211
rect 10 109 44 143
rect 98 109 132 143
rect 194 109 228 143
<< pdiffc >>
rect 10 1179 44 1213
rect 10 1111 44 1145
rect 10 1043 44 1077
rect 10 975 44 1009
rect 10 907 44 941
rect 98 1179 132 1213
rect 98 1111 132 1145
rect 98 1043 132 1077
rect 98 975 132 1009
rect 98 907 132 941
rect 186 1179 220 1213
rect 186 1111 220 1145
rect 186 1043 220 1077
rect 186 975 220 1009
rect 186 907 220 941
<< psubdiff >>
rect -123 487 361 549
rect -123 455 -61 487
rect -123 421 -108 455
rect -74 421 -61 455
rect -123 387 -61 421
rect -123 353 -108 387
rect -74 353 -61 387
rect 299 455 361 487
rect 299 421 313 455
rect 347 421 361 455
rect 299 387 361 421
rect -123 319 -61 353
rect -123 285 -108 319
rect -74 285 -61 319
rect -123 251 -61 285
rect -123 217 -108 251
rect -74 217 -61 251
rect -123 183 -61 217
rect -123 149 -108 183
rect -74 149 -61 183
rect -123 115 -61 149
rect -123 81 -109 115
rect -75 81 -61 115
rect 299 353 313 387
rect 347 353 361 387
rect 299 319 361 353
rect 299 285 313 319
rect 347 285 361 319
rect 299 251 361 285
rect 299 217 313 251
rect 347 217 361 251
rect 299 183 361 217
rect 299 149 313 183
rect 347 149 361 183
rect 299 115 361 149
rect -123 47 -61 81
rect 299 81 313 115
rect 347 81 361 115
rect 299 47 361 81
rect -123 13 -44 47
rect -10 13 24 47
rect 58 13 93 47
rect 127 13 167 47
rect 201 13 235 47
rect 269 13 361 47
rect -123 0 361 13
<< nsubdiff >>
rect -123 1283 -44 1317
rect -10 1283 24 1317
rect 58 1283 92 1317
rect 126 1283 160 1317
rect 195 1283 229 1317
rect 264 1283 363 1317
rect -123 1249 -61 1283
rect -123 1215 -109 1249
rect -74 1215 -61 1249
rect 301 1249 363 1283
rect -123 1181 -61 1215
rect -123 1147 -109 1181
rect -74 1147 -61 1181
rect -123 1113 -61 1147
rect -123 1079 -109 1113
rect -74 1079 -61 1113
rect -123 1045 -61 1079
rect -123 1011 -109 1045
rect -74 1011 -61 1045
rect -123 977 -61 1011
rect -123 943 -109 977
rect -74 943 -61 977
rect -123 909 -61 943
rect -123 875 -109 909
rect -74 875 -61 909
rect -123 841 -61 875
rect -123 807 -109 841
rect -74 807 -61 841
rect 301 1215 314 1249
rect 349 1215 363 1249
rect 301 1181 363 1215
rect 301 1147 314 1181
rect 349 1147 363 1181
rect 301 1113 363 1147
rect 301 1079 314 1113
rect 349 1079 363 1113
rect 301 1045 363 1079
rect 301 1011 314 1045
rect 349 1011 363 1045
rect 301 977 363 1011
rect 301 943 314 977
rect 349 943 363 977
rect 301 909 363 943
rect 301 875 314 909
rect 349 875 363 909
rect 301 841 363 875
rect -123 773 -61 807
rect -123 739 -109 773
rect -74 739 -61 773
rect -123 710 -61 739
rect 301 807 314 841
rect 349 807 363 841
rect 301 773 363 807
rect 301 739 314 773
rect 349 739 363 773
rect 301 710 363 739
rect -123 648 363 710
<< psubdiffcont >>
rect -108 421 -74 455
rect -108 353 -74 387
rect 313 421 347 455
rect -108 285 -74 319
rect -108 217 -74 251
rect -108 149 -74 183
rect -109 81 -75 115
rect 313 353 347 387
rect 313 285 347 319
rect 313 217 347 251
rect 313 149 347 183
rect 313 81 347 115
rect -44 13 -10 47
rect 24 13 58 47
rect 93 13 127 47
rect 167 13 201 47
rect 235 13 269 47
<< nsubdiffcont >>
rect -44 1283 -10 1317
rect 24 1283 58 1317
rect 92 1283 126 1317
rect 160 1283 195 1317
rect 229 1283 264 1317
rect -109 1215 -74 1249
rect -109 1147 -74 1181
rect -109 1079 -74 1113
rect -109 1011 -74 1045
rect -109 943 -74 977
rect -109 875 -74 909
rect -109 807 -74 841
rect 314 1215 349 1249
rect 314 1147 349 1181
rect 314 1079 349 1113
rect 314 1011 349 1045
rect 314 943 349 977
rect 314 875 349 909
rect -109 739 -74 773
rect 314 807 349 841
rect 314 739 349 773
<< poly >>
rect 56 1229 86 1255
rect 144 1229 174 1255
rect 56 802 86 829
rect 144 802 174 829
rect 56 801 174 802
rect -2 782 174 801
rect -2 748 14 782
rect 48 772 174 782
rect 48 748 64 772
rect -2 738 64 748
rect 4 449 86 465
rect 4 415 14 449
rect 48 415 86 449
rect 4 399 86 415
rect 56 368 86 399
<< polycont >>
rect 14 748 48 782
rect 14 415 48 449
<< locali >>
rect -123 1317 363 1332
rect -123 1283 -44 1317
rect -10 1283 24 1317
rect 58 1283 92 1317
rect 126 1283 160 1317
rect 195 1283 229 1317
rect 264 1283 363 1317
rect -123 1270 363 1283
rect -123 1249 -61 1270
rect -123 1215 -109 1249
rect -74 1215 -61 1249
rect -123 1181 -61 1215
rect -123 1147 -109 1181
rect -74 1147 -61 1181
rect -123 1113 -61 1147
rect -123 1079 -109 1113
rect -74 1079 -61 1113
rect -123 1045 -61 1079
rect -123 1011 -109 1045
rect -74 1011 -61 1045
rect -123 977 -61 1011
rect -123 943 -109 977
rect -74 943 -61 977
rect -123 909 -61 943
rect -123 875 -109 909
rect -74 875 -61 909
rect -123 841 -61 875
rect 10 1213 44 1270
rect 10 1145 44 1179
rect 10 1077 44 1111
rect 10 1009 44 1043
rect 10 941 44 975
rect 10 847 44 907
rect 98 1213 132 1229
rect 98 1145 132 1179
rect 98 1077 132 1111
rect 98 1009 132 1043
rect 98 941 132 975
rect 98 884 132 907
rect 186 1213 220 1270
rect 186 1145 220 1179
rect 186 1077 220 1111
rect 186 1009 220 1043
rect 186 941 220 975
rect 186 854 220 907
rect 301 1249 363 1270
rect 301 1215 314 1249
rect 349 1215 363 1249
rect 301 1181 363 1215
rect 301 1147 314 1181
rect 349 1147 363 1181
rect 301 1113 363 1147
rect 301 1079 314 1113
rect 349 1079 363 1113
rect 301 1045 363 1079
rect 301 1011 314 1045
rect 349 1011 363 1045
rect 301 977 363 1011
rect 301 943 314 977
rect 349 943 363 977
rect 301 909 363 943
rect 301 875 314 909
rect 349 875 363 909
rect -123 807 -109 841
rect -74 807 -61 841
rect -123 773 -61 807
rect -123 739 -109 773
rect -74 739 -61 773
rect -2 748 14 782
rect 48 748 64 782
rect -123 648 -61 739
rect -123 455 -61 549
rect -123 421 -108 455
rect -74 421 -61 455
rect -123 387 -61 421
rect 14 449 48 465
rect 14 399 48 415
rect -123 353 -108 387
rect -74 353 -61 387
rect -123 319 -61 353
rect -123 285 -108 319
rect -74 285 -61 319
rect -123 251 -61 285
rect -123 217 -108 251
rect -74 217 -61 251
rect -123 183 -61 217
rect -123 149 -108 183
rect -74 149 -61 183
rect -123 115 -61 149
rect 10 307 44 365
rect 10 211 44 273
rect 98 240 132 850
rect 301 841 363 875
rect 301 807 314 841
rect 349 807 363 841
rect 301 773 363 807
rect 301 739 314 773
rect 349 739 363 773
rect 301 648 363 739
rect 299 455 361 549
rect 299 421 313 455
rect 347 421 361 455
rect 299 387 361 421
rect 98 190 132 206
rect 194 307 228 358
rect 194 211 228 273
rect 10 143 44 177
rect 194 143 228 177
rect 299 353 313 387
rect 347 353 361 387
rect 299 319 361 353
rect 299 285 313 319
rect 347 285 361 319
rect 299 251 361 285
rect 299 217 313 251
rect 347 217 361 251
rect 299 183 361 217
rect 299 149 313 183
rect 347 149 361 183
rect -123 81 -109 115
rect -75 81 -61 115
rect -7 109 10 143
rect 44 109 98 143
rect 132 109 194 143
rect 228 109 245 143
rect 299 115 361 149
rect -123 62 -61 81
rect 10 62 44 109
rect 194 62 228 109
rect 299 81 313 115
rect 347 81 361 115
rect 299 62 361 81
rect -123 47 361 62
rect -123 13 -44 47
rect -10 13 24 47
rect 58 13 93 47
rect 127 13 167 47
rect 201 13 235 47
rect 269 13 361 47
rect -123 0 361 13
<< viali >>
rect -44 1283 -10 1317
rect 24 1283 58 1317
rect 92 1283 126 1317
rect 160 1283 195 1317
rect 229 1283 264 1317
rect -109 1215 -74 1249
rect -109 1147 -74 1181
rect -109 1079 -74 1113
rect -109 1011 -74 1045
rect -109 943 -74 977
rect -109 875 -74 909
rect 98 850 132 884
rect 314 1215 349 1249
rect 314 1147 349 1181
rect 314 1079 349 1113
rect 314 1011 349 1045
rect 314 943 349 977
rect 314 875 349 909
rect -109 807 -74 841
rect -109 739 -74 773
rect 14 748 48 782
rect -108 421 -74 455
rect 14 415 48 449
rect -108 353 -74 387
rect -108 285 -74 319
rect -108 217 -74 251
rect -108 149 -74 183
rect 314 807 349 841
rect 314 739 349 773
rect 313 421 347 455
rect 313 353 347 387
rect 313 285 347 319
rect 313 217 347 251
rect 313 149 347 183
rect -109 81 -75 115
rect 313 81 347 115
rect -44 13 -10 47
rect 24 13 58 47
rect 93 13 127 47
rect 167 13 201 47
rect 235 13 269 47
<< metal1 >>
rect -123 1317 363 1332
rect -123 1283 -44 1317
rect -10 1283 24 1317
rect 58 1283 92 1317
rect 126 1283 160 1317
rect 195 1283 229 1317
rect 264 1283 363 1317
rect -123 1270 363 1283
rect -123 1249 -61 1270
rect -123 1215 -109 1249
rect -74 1215 -61 1249
rect -123 1181 -61 1215
rect -123 1147 -109 1181
rect -74 1147 -61 1181
rect -123 1113 -61 1147
rect -123 1079 -109 1113
rect -74 1079 -61 1113
rect -123 1045 -61 1079
rect -123 1011 -109 1045
rect -74 1011 -61 1045
rect -123 977 -61 1011
rect -123 943 -109 977
rect -74 943 -61 977
rect -123 909 -61 943
rect -123 875 -109 909
rect -74 875 -61 909
rect 301 1249 363 1270
rect 301 1215 314 1249
rect 349 1215 363 1249
rect 301 1181 363 1215
rect 301 1147 314 1181
rect 349 1147 363 1181
rect 301 1113 363 1147
rect 301 1079 314 1113
rect 349 1079 363 1113
rect 301 1045 363 1079
rect 301 1011 314 1045
rect 349 1011 363 1045
rect 301 977 363 1011
rect 301 943 314 977
rect 349 943 363 977
rect 301 909 363 943
rect 98 890 132 896
rect -123 841 -61 875
rect 92 884 138 890
rect 92 850 98 884
rect 132 850 138 884
rect 92 844 138 850
rect 301 875 314 909
rect 349 875 363 909
rect -123 807 -109 841
rect -74 807 -61 841
rect -123 773 -61 807
rect 14 788 48 794
rect -123 739 -109 773
rect -74 739 -61 773
rect 8 782 54 788
rect 8 748 14 782
rect 48 748 54 782
rect 98 770 132 844
rect 301 841 363 875
rect 301 807 314 841
rect 349 807 363 841
rect 301 773 363 807
rect 8 742 54 748
rect -123 648 -61 739
rect -123 455 -61 549
rect 14 456 48 742
rect 301 739 314 773
rect 349 739 363 773
rect 301 648 363 739
rect -123 421 -108 455
rect -74 421 -61 455
rect -123 387 -61 421
rect 8 449 54 456
rect 8 415 14 449
rect 48 415 54 449
rect 8 408 54 415
rect 299 455 361 549
rect 299 421 313 455
rect 347 421 361 455
rect 14 392 48 408
rect -123 353 -108 387
rect -74 353 -61 387
rect -123 319 -61 353
rect -123 285 -108 319
rect -74 285 -61 319
rect -123 251 -61 285
rect -123 217 -108 251
rect -74 217 -61 251
rect -123 183 -61 217
rect -123 149 -108 183
rect -74 149 -61 183
rect -123 115 -61 149
rect -123 81 -109 115
rect -75 81 -61 115
rect -123 62 -61 81
rect 299 387 361 421
rect 299 353 313 387
rect 347 353 361 387
rect 299 319 361 353
rect 299 285 313 319
rect 347 285 361 319
rect 299 251 361 285
rect 299 217 313 251
rect 347 217 361 251
rect 299 183 361 217
rect 299 149 313 183
rect 347 149 361 183
rect 299 115 361 149
rect 299 81 313 115
rect 347 81 361 115
rect 299 62 361 81
rect -123 47 361 62
rect -123 13 -44 47
rect -10 13 24 47
rect 58 13 93 47
rect 127 13 167 47
rect 201 13 235 47
rect 269 13 361 47
rect -123 0 361 13
<< labels >>
rlabel metal1 161 1325 161 1325 1 VDD
port 1 n
rlabel metal1 98 850 132 884 1 Y
port 2 n
rlabel metal1 14 748 48 782 1 A
port 3 n
rlabel metal1 146 31 146 31 1 VSS
port 4 n
<< end >>
