magic
tech sky130A
magscale 1 2
timestamp 1643180485
<< poly >>
rect 70 449 124 465
rect 70 415 80 449
rect 114 415 124 449
rect 70 399 124 415
<< polycont >>
rect 80 415 114 449
<< locali >>
rect 80 449 114 465
rect 80 399 114 415
<< viali >>
rect 80 415 114 449
<< metal1 >>
rect 80 455 114 473
rect 74 449 120 455
rect 74 415 80 449
rect 114 415 120 449
rect 74 409 120 415
rect 80 391 114 409
<< end >>
