magic
tech sky130A
magscale 1 2
timestamp 1648505949
<< nwell >>
rect 55 1505 89 1539
<< psubdiffcont >>
rect 55 13 89 47
<< nsubdiffcont >>
rect 55 1505 89 1539
<< viali >>
rect 55 1505 89 1539
rect 55 13 89 47
<< metal1 >>
rect 1093 945 1127 979
rect 205 797 239 831
rect 4089 797 4554 831
rect 3497 723 4707 757
rect 4719 723 4753 757
rect 2055 427 2089 461
use li1_M1_contact  li1_M1_contact_2 pcells
timestamp 1648061256
transform 1 0 4736 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform -1 0 3478 0 -1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_11
timestamp 1648061256
transform -1 0 4070 0 -1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_19
timestamp 1648061256
transform 1 0 4588 0 1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform 1 0 222 0 1 814
box -53 -33 29 33
use dffsnqx1  dffsnqx1_0 pcells
timestamp 1648501217
transform 1 0 0 0 1 0
box -84 0 4968 1575
<< labels >>
rlabel metal1 4719 723 4753 757 1 Q
port 1 n
rlabel metal1 205 797 239 831 1 D
port 2 n
rlabel metal1 1093 945 1127 979 1 CLK
port 3 n
rlabel metal1 2055 427 2089 461 1 SN
port 4 n
rlabel metal1 55 1505 89 1539 1 VDD
port 6 n
rlabel metal1 55 13 89 47 1 VSS
port 7 n
<< end >>
