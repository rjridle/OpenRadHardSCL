** sch_path: /home/rjridle/OpenRadHardSCL/lib/xschem/schematics/INVX2.sch
**.subckt INVX2 A Y
*.ipin A
*.opin Y
M3 Y A VDD VDD pmos w=2u l=0.150u m=1
M2 Y A VDD VDD pmos w=2u l=0.150u m=1
M1 Y A GND GND nmos w=3u l=0.150u m=1
M4 Y A VDD VDD pmos w=2u l=0.150u m=1
M5 Y A VDD VDD pmos w=2u l=0.150u m=1
M6 Y A GND GND nmos w=3u l=0.150u m=1
**.ends
.GLOBAL GND
.GLOBAL VDD
.end
