magic
tech sky130A
magscale 1 2
timestamp 1642407040
<< error_p >>
rect 127 318 128 319
rect 311 318 312 319
rect 612 318 613 319
rect 128 317 129 318
rect 312 317 313 318
rect 613 317 614 318
rect 143 287 144 288
rect 178 287 179 288
rect 327 287 328 288
rect 362 287 363 288
rect 628 287 629 288
rect 663 287 664 288
rect 143 184 144 185
rect 178 184 179 185
rect 327 184 328 185
rect 362 184 363 185
rect 628 184 629 185
rect 663 184 664 185
<< nwell >>
rect 0 591 799 1353
<< nmos >>
rect 98 318 128 368
rect 98 288 194 318
tri 194 288 224 318 sw
rect 282 318 312 368
rect 98 184 128 288
tri 128 272 144 288 nw
tri 178 272 194 288 ne
tri 128 184 144 200 sw
tri 178 184 194 200 se
rect 194 184 224 288
rect 282 288 378 318
tri 378 288 408 318 sw
tri 98 154 128 184 ne
rect 128 154 194 184
tri 194 154 224 184 nw
rect 282 184 312 288
tri 312 272 328 288 nw
tri 362 272 378 288 ne
tri 312 184 328 200 sw
tri 362 184 378 200 se
rect 378 184 408 288
tri 282 154 312 184 ne
rect 312 154 378 184
tri 378 154 408 184 nw
rect 583 318 613 368
rect 583 288 679 318
tri 679 288 709 318 sw
rect 583 184 613 288
tri 613 272 629 288 nw
tri 663 272 679 288 ne
tri 613 184 629 200 sw
tri 663 184 679 200 se
rect 679 184 709 288
tri 583 154 613 184 ne
rect 613 154 679 184
tri 679 154 709 184 nw
<< pmos >>
rect 98 629 128 1229
rect 186 629 216 1229
rect 282 629 312 1229
rect 370 629 400 1229
rect 583 629 613 1229
rect 671 629 701 1229
<< ndiff >>
rect 36 347 98 368
rect 36 313 52 347
rect 86 313 98 347
rect 128 347 282 368
rect 128 318 236 347
rect 36 279 98 313
tri 194 288 224 318 ne
rect 224 313 236 318
rect 270 313 282 347
rect 312 347 466 368
rect 312 318 420 347
rect 36 245 52 279
rect 86 245 98 279
rect 36 211 98 245
rect 36 177 52 211
rect 86 177 98 211
tri 128 272 144 288 se
rect 144 272 178 288
tri 178 272 194 288 sw
rect 128 240 194 272
rect 128 206 140 240
rect 174 206 194 240
rect 128 200 194 206
tri 128 184 144 200 ne
rect 144 184 178 200
tri 178 184 194 200 nw
rect 224 279 282 313
tri 378 288 408 318 ne
rect 408 313 420 318
rect 454 313 466 347
rect 224 245 236 279
rect 270 245 282 279
rect 224 211 282 245
rect 36 154 98 177
tri 98 154 128 184 sw
tri 194 154 224 184 se
rect 224 177 236 211
rect 270 177 282 211
tri 312 272 328 288 se
rect 328 272 362 288
tri 362 272 378 288 sw
rect 312 240 378 272
rect 312 206 324 240
rect 358 206 378 240
rect 312 200 378 206
tri 312 184 328 200 ne
rect 328 184 362 200
tri 362 184 378 200 nw
rect 408 279 466 313
rect 408 245 420 279
rect 454 245 466 279
rect 408 211 466 245
rect 224 154 282 177
tri 282 154 312 184 sw
tri 378 154 408 184 se
rect 408 177 420 211
rect 454 177 466 211
rect 408 154 466 177
rect 36 143 466 154
rect 36 109 52 143
rect 86 109 144 143
rect 178 109 236 143
rect 270 109 328 143
rect 362 109 420 143
rect 454 109 466 143
rect 36 101 466 109
rect 520 347 583 368
rect 520 313 537 347
rect 571 313 583 347
rect 613 347 772 368
rect 613 318 721 347
rect 520 279 583 313
tri 679 288 709 318 ne
rect 709 313 721 318
rect 755 313 772 347
rect 520 245 537 279
rect 571 245 583 279
rect 520 211 583 245
rect 520 177 537 211
rect 571 177 583 211
tri 613 272 629 288 se
rect 629 272 663 288
tri 663 272 679 288 sw
rect 613 240 679 272
rect 613 206 625 240
rect 659 206 679 240
rect 613 200 679 206
tri 613 184 629 200 ne
rect 629 184 663 200
tri 663 184 679 200 nw
rect 709 279 772 313
rect 709 245 721 279
rect 755 245 772 279
rect 709 211 772 245
rect 520 154 583 177
tri 583 154 613 184 sw
tri 679 154 709 184 se
rect 709 177 721 211
rect 755 177 772 211
rect 709 154 772 177
rect 520 143 772 154
rect 520 109 537 143
rect 571 109 625 143
rect 659 109 721 143
rect 755 109 772 143
rect 520 101 772 109
<< pdiff >>
rect 40 1213 98 1229
rect 40 1179 52 1213
rect 86 1179 98 1213
rect 40 1145 98 1179
rect 40 1111 52 1145
rect 86 1111 98 1145
rect 40 1077 98 1111
rect 40 1043 52 1077
rect 86 1043 98 1077
rect 40 1009 98 1043
rect 40 975 52 1009
rect 86 975 98 1009
rect 40 941 98 975
rect 40 907 52 941
rect 86 907 98 941
rect 40 873 98 907
rect 40 839 52 873
rect 86 839 98 873
rect 40 805 98 839
rect 40 771 52 805
rect 86 771 98 805
rect 40 737 98 771
rect 40 703 52 737
rect 86 703 98 737
rect 40 629 98 703
rect 128 629 186 1229
rect 216 1213 282 1229
rect 216 1179 230 1213
rect 264 1179 282 1213
rect 216 1145 282 1179
rect 216 1111 230 1145
rect 264 1111 282 1145
rect 216 1077 282 1111
rect 216 1043 230 1077
rect 264 1043 282 1077
rect 216 1009 282 1043
rect 216 975 230 1009
rect 264 975 282 1009
rect 216 941 282 975
rect 216 907 230 941
rect 264 907 282 941
rect 216 873 282 907
rect 216 839 230 873
rect 264 839 282 873
rect 216 805 282 839
rect 216 771 230 805
rect 264 771 282 805
rect 216 737 282 771
rect 216 703 230 737
rect 264 703 282 737
rect 216 629 282 703
rect 312 629 370 1229
rect 400 1213 454 1229
rect 400 1179 412 1213
rect 446 1179 454 1213
rect 400 1145 454 1179
rect 400 1111 412 1145
rect 446 1111 454 1145
rect 400 1077 454 1111
rect 400 1043 412 1077
rect 446 1043 454 1077
rect 400 1009 454 1043
rect 400 975 412 1009
rect 446 975 454 1009
rect 400 941 454 975
rect 400 907 412 941
rect 446 907 454 941
rect 400 873 454 907
rect 400 839 412 873
rect 446 839 454 873
rect 400 805 454 839
rect 400 771 412 805
rect 446 771 454 805
rect 400 737 454 771
rect 400 703 412 737
rect 446 703 454 737
rect 400 629 454 703
rect 527 1213 583 1229
rect 527 1179 537 1213
rect 571 1179 583 1213
rect 527 1145 583 1179
rect 527 1111 537 1145
rect 571 1111 583 1145
rect 527 1077 583 1111
rect 527 1043 537 1077
rect 571 1043 583 1077
rect 527 1009 583 1043
rect 527 975 537 1009
rect 571 975 583 1009
rect 527 941 583 975
rect 527 907 537 941
rect 571 907 583 941
rect 527 873 583 907
rect 527 839 537 873
rect 571 839 583 873
rect 527 805 583 839
rect 527 771 537 805
rect 571 771 583 805
rect 527 737 583 771
rect 527 703 537 737
rect 571 703 583 737
rect 527 629 583 703
rect 613 1213 671 1229
rect 613 1179 625 1213
rect 659 1179 671 1213
rect 613 1145 671 1179
rect 613 1111 625 1145
rect 659 1111 671 1145
rect 613 1077 671 1111
rect 613 1043 625 1077
rect 659 1043 671 1077
rect 613 1009 671 1043
rect 613 975 625 1009
rect 659 975 671 1009
rect 613 941 671 975
rect 613 907 625 941
rect 659 907 671 941
rect 613 873 671 907
rect 613 839 625 873
rect 659 839 671 873
rect 613 805 671 839
rect 613 771 625 805
rect 659 771 671 805
rect 613 737 671 771
rect 613 703 625 737
rect 659 703 671 737
rect 613 629 671 703
rect 701 1213 755 1229
rect 701 1179 713 1213
rect 747 1179 755 1213
rect 701 1145 755 1179
rect 701 1111 713 1145
rect 747 1111 755 1145
rect 701 1077 755 1111
rect 701 1043 713 1077
rect 747 1043 755 1077
rect 701 1009 755 1043
rect 701 975 713 1009
rect 747 975 755 1009
rect 701 941 755 975
rect 701 907 713 941
rect 747 907 755 941
rect 701 873 755 907
rect 701 839 713 873
rect 747 839 755 873
rect 701 805 755 839
rect 701 771 713 805
rect 747 771 755 805
rect 701 737 755 771
rect 701 703 713 737
rect 747 703 755 737
rect 701 629 755 703
<< ndiffc >>
rect 52 313 86 347
rect 236 313 270 347
rect 52 245 86 279
rect 52 177 86 211
rect 140 206 174 240
rect 420 313 454 347
rect 236 245 270 279
rect 236 177 270 211
rect 324 206 358 240
rect 420 245 454 279
rect 420 177 454 211
rect 52 109 86 143
rect 144 109 178 143
rect 236 109 270 143
rect 328 109 362 143
rect 420 109 454 143
rect 537 313 571 347
rect 721 313 755 347
rect 537 245 571 279
rect 537 177 571 211
rect 625 206 659 240
rect 721 245 755 279
rect 721 177 755 211
rect 537 109 571 143
rect 625 109 659 143
rect 721 109 755 143
<< pdiffc >>
rect 52 1179 86 1213
rect 52 1111 86 1145
rect 52 1043 86 1077
rect 52 975 86 1009
rect 52 907 86 941
rect 52 839 86 873
rect 52 771 86 805
rect 52 703 86 737
rect 230 1179 264 1213
rect 230 1111 264 1145
rect 230 1043 264 1077
rect 230 975 264 1009
rect 230 907 264 941
rect 230 839 264 873
rect 230 771 264 805
rect 230 703 264 737
rect 412 1179 446 1213
rect 412 1111 446 1145
rect 412 1043 446 1077
rect 412 975 446 1009
rect 412 907 446 941
rect 412 839 446 873
rect 412 771 446 805
rect 412 703 446 737
rect 537 1179 571 1213
rect 537 1111 571 1145
rect 537 1043 571 1077
rect 537 975 571 1009
rect 537 907 571 941
rect 537 839 571 873
rect 537 771 571 805
rect 537 703 571 737
rect 625 1179 659 1213
rect 625 1111 659 1145
rect 625 1043 659 1077
rect 625 975 659 1009
rect 625 907 659 941
rect 625 839 659 873
rect 625 771 659 805
rect 625 703 659 737
rect 713 1179 747 1213
rect 713 1111 747 1145
rect 713 1043 747 1077
rect 713 975 747 1009
rect 713 907 747 941
rect 713 839 747 873
rect 713 771 747 805
rect 713 703 747 737
<< psubdiff >>
rect 36 13 60 47
rect 94 13 129 47
rect 163 13 205 47
rect 239 13 273 47
rect 307 13 342 47
rect 376 13 410 47
rect 444 13 478 47
rect 512 13 546 47
rect 580 13 614 47
rect 648 13 682 47
rect 716 13 763 47
<< nsubdiff >>
rect 36 1283 60 1317
rect 94 1283 128 1317
rect 162 1283 196 1317
rect 231 1283 265 1317
rect 299 1283 333 1317
rect 367 1283 401 1317
rect 435 1283 469 1317
rect 503 1283 537 1317
rect 571 1283 605 1317
rect 640 1283 674 1317
rect 709 1283 763 1317
<< psubdiffcont >>
rect 60 13 94 47
rect 129 13 163 47
rect 205 13 239 47
rect 273 13 307 47
rect 342 13 376 47
rect 410 13 444 47
rect 478 13 512 47
rect 546 13 580 47
rect 614 13 648 47
rect 682 13 716 47
<< nsubdiffcont >>
rect 60 1283 94 1317
rect 128 1283 162 1317
rect 196 1283 231 1317
rect 265 1283 299 1317
rect 333 1283 367 1317
rect 401 1283 435 1317
rect 469 1283 503 1317
rect 537 1283 571 1317
rect 605 1283 640 1317
rect 674 1283 709 1317
<< poly >>
rect 98 1229 128 1255
rect 186 1229 216 1255
rect 282 1229 312 1255
rect 370 1229 400 1255
rect 583 1229 613 1255
rect 671 1229 701 1255
rect 98 612 128 629
rect 186 612 216 629
rect 98 582 216 612
rect 282 612 312 629
rect 370 612 400 629
rect 282 582 400 612
rect 583 612 613 629
rect 671 612 701 629
rect 583 582 701 612
rect 98 568 128 582
rect 62 552 128 568
rect 62 518 72 552
rect 106 518 128 552
rect 62 502 128 518
rect 98 368 128 502
rect 282 494 312 582
rect 583 494 613 582
rect 249 478 312 494
rect 249 444 259 478
rect 293 444 312 478
rect 249 428 312 444
rect 547 478 613 494
rect 547 444 557 478
rect 591 444 613 478
rect 547 428 613 444
rect 282 368 312 428
rect 583 368 613 428
<< polycont >>
rect 72 518 106 552
rect 259 444 293 478
rect 557 444 591 478
<< locali >>
rect 36 1317 763 1332
rect 36 1283 60 1317
rect 94 1283 128 1317
rect 162 1283 196 1317
rect 231 1283 265 1317
rect 299 1283 333 1317
rect 367 1283 401 1317
rect 435 1283 469 1317
rect 503 1283 537 1317
rect 571 1283 605 1317
rect 640 1283 674 1317
rect 709 1283 763 1317
rect 36 1270 763 1283
rect 52 1213 86 1229
rect 52 1145 86 1179
rect 52 1077 86 1111
rect 52 1009 86 1043
rect 52 941 86 975
rect 52 873 86 907
rect 52 805 86 839
rect 52 737 86 771
rect 52 684 86 703
rect 52 629 86 650
rect 230 1213 264 1270
rect 230 1145 264 1179
rect 230 1077 264 1111
rect 230 1009 264 1043
rect 230 941 264 975
rect 230 873 264 907
rect 230 805 264 839
rect 230 737 264 771
rect 230 629 264 703
rect 412 1213 446 1229
rect 412 1145 446 1179
rect 412 1077 446 1111
rect 412 1009 446 1043
rect 412 941 446 975
rect 412 873 446 907
rect 412 805 446 839
rect 412 737 446 771
rect 412 684 446 703
rect 537 1213 571 1270
rect 537 1145 571 1179
rect 537 1077 571 1111
rect 537 1009 571 1043
rect 537 941 571 975
rect 537 873 571 907
rect 537 805 571 839
rect 537 737 571 771
rect 537 627 571 703
rect 625 1213 659 1229
rect 625 1145 659 1179
rect 625 1077 659 1111
rect 625 1009 659 1043
rect 625 941 659 975
rect 625 873 659 907
rect 625 805 659 839
rect 625 737 659 771
rect 625 684 659 703
rect 72 552 106 568
rect 72 502 106 518
rect 259 478 293 494
rect 259 428 293 444
rect 557 478 591 494
rect 557 428 591 444
rect 52 347 86 363
rect 52 279 86 313
rect 236 347 270 363
rect 52 211 86 245
rect 140 240 174 246
rect 140 190 174 206
rect 236 279 270 313
rect 420 347 454 363
rect 236 211 270 245
rect 52 143 86 177
rect 324 280 358 286
rect 324 240 358 246
rect 324 188 358 206
rect 420 279 454 313
rect 420 211 454 245
rect 236 143 270 177
rect 420 143 454 177
rect 537 347 571 363
rect 537 279 571 313
rect 537 211 571 245
rect 625 240 659 650
rect 713 1213 747 1270
rect 713 1145 747 1179
rect 713 1077 747 1111
rect 713 1009 747 1043
rect 713 941 747 975
rect 713 873 747 907
rect 713 805 747 839
rect 713 737 747 771
rect 713 627 747 703
rect 625 190 659 206
rect 721 347 755 363
rect 721 279 755 313
rect 721 211 755 245
rect 537 143 571 177
rect 721 143 755 177
rect 36 109 52 143
rect 86 109 144 143
rect 178 109 236 143
rect 270 109 328 143
rect 362 109 420 143
rect 454 109 466 143
rect 520 109 537 143
rect 571 109 625 143
rect 659 109 721 143
rect 755 109 772 143
rect 52 62 86 109
rect 144 62 178 109
rect 236 62 270 109
rect 328 62 362 109
rect 420 62 454 109
rect 537 62 571 109
rect 625 62 659 109
rect 721 62 755 109
rect 36 47 763 62
rect 36 13 60 47
rect 94 13 129 47
rect 163 13 205 47
rect 239 13 273 47
rect 307 13 342 47
rect 376 13 410 47
rect 444 13 478 47
rect 512 13 546 47
rect 580 13 614 47
rect 648 13 682 47
rect 716 13 763 47
rect 36 0 763 13
<< viali >>
rect 60 1283 94 1317
rect 128 1283 162 1317
rect 196 1283 231 1317
rect 265 1283 299 1317
rect 333 1283 367 1317
rect 401 1283 435 1317
rect 469 1283 503 1317
rect 537 1283 571 1317
rect 605 1283 640 1317
rect 674 1283 709 1317
rect 52 650 86 684
rect 412 650 446 684
rect 625 650 659 684
rect 72 518 106 552
rect 259 444 293 478
rect 557 444 591 478
rect 140 246 174 280
rect 324 246 358 280
rect 60 13 94 47
rect 129 13 163 47
rect 205 13 239 47
rect 273 13 307 47
rect 342 13 376 47
rect 410 13 444 47
rect 478 13 512 47
rect 546 13 580 47
rect 614 13 648 47
rect 682 13 716 47
<< metal1 >>
rect 36 1317 763 1332
rect 36 1283 60 1317
rect 94 1283 128 1317
rect 162 1283 196 1317
rect 231 1283 265 1317
rect 299 1283 333 1317
rect 367 1283 401 1317
rect 435 1283 469 1317
rect 503 1283 537 1317
rect 571 1283 605 1317
rect 640 1283 674 1317
rect 709 1283 763 1317
rect 36 1270 763 1283
rect 625 690 659 696
rect 46 684 92 690
rect 406 684 452 690
rect 619 684 665 690
rect 40 650 52 684
rect 86 650 412 684
rect 446 650 591 684
rect 46 644 92 650
rect 72 559 106 573
rect 62 552 112 559
rect 62 518 72 552
rect 106 518 112 552
rect 62 511 112 518
rect 72 497 106 511
rect 140 286 174 650
rect 406 644 452 650
rect 259 485 293 499
rect 557 485 591 650
rect 619 650 625 684
rect 659 650 665 684
rect 619 644 665 650
rect 625 614 659 644
rect 249 478 299 485
rect 249 444 259 478
rect 293 444 299 478
rect 249 437 299 444
rect 551 478 597 485
rect 551 444 557 478
rect 591 444 597 478
rect 551 437 597 444
rect 259 423 293 437
rect 557 421 591 437
rect 134 280 180 286
rect 318 280 364 286
rect 128 246 140 280
rect 174 246 324 280
rect 358 246 370 280
rect 134 245 364 246
rect 134 240 180 245
rect 318 240 364 245
rect 36 47 763 62
rect 36 13 60 47
rect 94 13 129 47
rect 163 13 205 47
rect 239 13 273 47
rect 307 13 342 47
rect 376 13 410 47
rect 444 13 478 47
rect 512 13 546 47
rect 580 13 614 47
rect 648 13 682 47
rect 716 13 763 47
rect 36 0 763 13
<< labels >>
rlabel metal1 197 1325 197 1325 1 VDD
rlabel metal1 184 31 184 31 1 VSS
rlabel metal1 72 518 106 552 1 A
rlabel metal1 259 444 293 478 1 B
rlabel metal1 625 650 659 684 1 Y
<< end >>
