* SPICE3 file created from INVX2.ext - technology: sky130A

.subckt INVX2 A Y VDD VSS
M1000 Y A VDD VDD pshort w=3u l=0.15u
+  ad=1.74p pd=13.16u as=2.49p ps=19.66u
M1001 Y A VSS VSS nshort w=3u l=0.15u
+  ad=0.3176p pd=3u as=1.8318p ps=12.66u
M1002 VDD A Y VDD pshort w=3u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 VDD A Y VDD pshort w=3u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A VDD VDD pshort w=3u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y A VSS VSS nshort w=3u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
.ends
