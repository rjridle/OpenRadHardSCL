magic
tech sky130A
magscale 1 2
timestamp 1649530825
<< nwell >>
rect -84 832 14958 1575
<< nmos >>
rect 147 318 177 379
tri 177 318 193 334 sw
rect 447 318 477 379
rect 147 288 253 318
tri 253 288 283 318 sw
rect 147 187 177 288
tri 177 272 193 288 nw
tri 237 272 253 288 ne
tri 177 187 193 203 sw
tri 237 187 253 203 se
rect 253 187 283 288
tri 342 288 372 318 se
rect 372 288 477 318
rect 342 194 372 288
tri 372 272 388 288 nw
tri 431 272 447 288 ne
tri 372 194 388 210 sw
tri 431 194 447 210 se
rect 447 194 477 288
tri 147 157 177 187 ne
rect 177 157 253 187
tri 253 157 283 187 nw
tri 342 164 372 194 ne
rect 372 164 447 194
tri 447 164 477 194 nw
rect 649 326 679 379
tri 679 326 695 342 sw
rect 649 296 755 326
tri 755 296 785 326 sw
rect 649 195 679 296
tri 679 280 695 296 nw
tri 739 280 755 296 ne
tri 679 195 695 211 sw
tri 739 195 755 211 se
rect 755 195 785 296
tri 649 165 679 195 ne
rect 679 165 755 195
tri 755 165 785 195 nw
rect 1130 316 1160 377
tri 1160 316 1176 332 sw
rect 1324 324 1354 377
tri 1354 324 1370 340 sw
rect 1130 286 1236 316
tri 1236 286 1266 316 sw
rect 1324 294 1430 324
tri 1430 294 1460 324 sw
rect 1130 185 1160 286
tri 1160 270 1176 286 nw
tri 1220 270 1236 286 ne
tri 1160 185 1176 201 sw
tri 1220 185 1236 201 se
rect 1236 185 1266 286
rect 1324 193 1354 294
tri 1354 278 1370 294 nw
tri 1414 278 1430 294 ne
tri 1354 193 1370 209 sw
tri 1414 193 1430 209 se
rect 1430 193 1460 294
tri 1130 155 1160 185 ne
rect 1160 155 1236 185
tri 1236 155 1266 185 nw
tri 1324 163 1354 193 ne
rect 1354 163 1430 193
tri 1430 163 1460 193 nw
rect 1796 316 1826 377
tri 1826 316 1842 332 sw
rect 1990 324 2020 377
tri 2020 324 2036 340 sw
rect 1796 286 1902 316
tri 1902 286 1932 316 sw
rect 1990 294 2096 324
tri 2096 294 2126 324 sw
rect 1796 185 1826 286
tri 1826 270 1842 286 nw
tri 1886 270 1902 286 ne
tri 1826 185 1842 201 sw
tri 1886 185 1902 201 se
rect 1902 185 1932 286
rect 1990 193 2020 294
tri 2020 278 2036 294 nw
tri 2080 278 2096 294 ne
tri 2020 193 2036 209 sw
tri 2080 193 2096 209 se
rect 2096 193 2126 294
tri 1796 155 1826 185 ne
rect 1826 155 1902 185
tri 1902 155 1932 185 nw
tri 1990 163 2020 193 ne
rect 2020 163 2096 193
tri 2096 163 2126 193 nw
rect 2462 316 2492 377
tri 2492 316 2508 332 sw
rect 2656 324 2686 377
tri 2686 324 2702 340 sw
rect 2462 286 2568 316
tri 2568 286 2598 316 sw
rect 2656 294 2762 324
tri 2762 294 2792 324 sw
rect 2462 185 2492 286
tri 2492 270 2508 286 nw
tri 2552 270 2568 286 ne
tri 2492 185 2508 201 sw
tri 2552 185 2568 201 se
rect 2568 185 2598 286
rect 2656 193 2686 294
tri 2686 278 2702 294 nw
tri 2746 278 2762 294 ne
tri 2686 193 2702 209 sw
tri 2746 193 2762 209 se
rect 2762 193 2792 294
tri 2462 155 2492 185 ne
rect 2492 155 2568 185
tri 2568 155 2598 185 nw
tri 2656 163 2686 193 ne
rect 2686 163 2762 193
tri 2762 163 2792 193 nw
rect 3128 316 3158 377
tri 3158 316 3174 332 sw
rect 3322 324 3352 377
tri 3352 324 3368 340 sw
rect 3128 286 3234 316
tri 3234 286 3264 316 sw
rect 3322 294 3428 324
tri 3428 294 3458 324 sw
rect 3128 185 3158 286
tri 3158 270 3174 286 nw
tri 3218 270 3234 286 ne
tri 3158 185 3174 201 sw
tri 3218 185 3234 201 se
rect 3234 185 3264 286
rect 3322 193 3352 294
tri 3352 278 3368 294 nw
tri 3412 278 3428 294 ne
tri 3352 193 3368 209 sw
tri 3412 193 3428 209 se
rect 3428 193 3458 294
tri 3128 155 3158 185 ne
rect 3158 155 3234 185
tri 3234 155 3264 185 nw
tri 3322 163 3352 193 ne
rect 3352 163 3428 193
tri 3428 163 3458 193 nw
rect 3794 316 3824 377
tri 3824 316 3840 332 sw
rect 3988 324 4018 377
tri 4018 324 4034 340 sw
rect 3794 286 3900 316
tri 3900 286 3930 316 sw
rect 3988 294 4094 324
tri 4094 294 4124 324 sw
rect 3794 185 3824 286
tri 3824 270 3840 286 nw
tri 3884 270 3900 286 ne
tri 3824 185 3840 201 sw
tri 3884 185 3900 201 se
rect 3900 185 3930 286
rect 3988 193 4018 294
tri 4018 278 4034 294 nw
tri 4078 278 4094 294 ne
tri 4018 193 4034 209 sw
tri 4078 193 4094 209 se
rect 4094 193 4124 294
tri 3794 155 3824 185 ne
rect 3824 155 3900 185
tri 3900 155 3930 185 nw
tri 3988 163 4018 193 ne
rect 4018 163 4094 193
tri 4094 163 4124 193 nw
rect 4439 318 4469 379
tri 4469 318 4485 334 sw
rect 4739 318 4769 379
rect 4439 288 4545 318
tri 4545 288 4575 318 sw
rect 4439 187 4469 288
tri 4469 272 4485 288 nw
tri 4529 272 4545 288 ne
tri 4469 187 4485 203 sw
tri 4529 187 4545 203 se
rect 4545 187 4575 288
tri 4634 288 4664 318 se
rect 4664 288 4769 318
rect 4634 194 4664 288
tri 4664 272 4680 288 nw
tri 4723 272 4739 288 ne
tri 4664 194 4680 210 sw
tri 4723 194 4739 210 se
rect 4739 194 4769 288
tri 4439 157 4469 187 ne
rect 4469 157 4545 187
tri 4545 157 4575 187 nw
tri 4634 164 4664 194 ne
rect 4664 164 4739 194
tri 4739 164 4769 194 nw
rect 4941 326 4971 379
tri 4971 326 4987 342 sw
rect 4941 296 5047 326
tri 5047 296 5077 326 sw
rect 4941 195 4971 296
tri 4971 280 4987 296 nw
tri 5031 280 5047 296 ne
tri 4971 195 4987 211 sw
tri 5031 195 5047 211 se
rect 5047 195 5077 296
tri 4941 165 4971 195 ne
rect 4971 165 5047 195
tri 5047 165 5077 195 nw
rect 5422 316 5452 377
tri 5452 316 5468 332 sw
rect 5616 324 5646 377
tri 5646 324 5662 340 sw
rect 5422 286 5528 316
tri 5528 286 5558 316 sw
rect 5616 294 5722 324
tri 5722 294 5752 324 sw
rect 5422 185 5452 286
tri 5452 270 5468 286 nw
tri 5512 270 5528 286 ne
tri 5452 185 5468 201 sw
tri 5512 185 5528 201 se
rect 5528 185 5558 286
rect 5616 193 5646 294
tri 5646 278 5662 294 nw
tri 5706 278 5722 294 ne
tri 5646 193 5662 209 sw
tri 5706 193 5722 209 se
rect 5722 193 5752 294
tri 5422 155 5452 185 ne
rect 5452 155 5528 185
tri 5528 155 5558 185 nw
tri 5616 163 5646 193 ne
rect 5646 163 5722 193
tri 5722 163 5752 193 nw
rect 6088 316 6118 377
tri 6118 316 6134 332 sw
rect 6282 324 6312 377
tri 6312 324 6328 340 sw
rect 6088 286 6194 316
tri 6194 286 6224 316 sw
rect 6282 294 6388 324
tri 6388 294 6418 324 sw
rect 6088 185 6118 286
tri 6118 270 6134 286 nw
tri 6178 270 6194 286 ne
tri 6118 185 6134 201 sw
tri 6178 185 6194 201 se
rect 6194 185 6224 286
rect 6282 193 6312 294
tri 6312 278 6328 294 nw
tri 6372 278 6388 294 ne
tri 6312 193 6328 209 sw
tri 6372 193 6388 209 se
rect 6388 193 6418 294
tri 6088 155 6118 185 ne
rect 6118 155 6194 185
tri 6194 155 6224 185 nw
tri 6282 163 6312 193 ne
rect 6312 163 6388 193
tri 6388 163 6418 193 nw
rect 6754 316 6784 377
tri 6784 316 6800 332 sw
rect 6948 324 6978 377
tri 6978 324 6994 340 sw
rect 6754 286 6860 316
tri 6860 286 6890 316 sw
rect 6948 294 7054 324
tri 7054 294 7084 324 sw
rect 6754 185 6784 286
tri 6784 270 6800 286 nw
tri 6844 270 6860 286 ne
tri 6784 185 6800 201 sw
tri 6844 185 6860 201 se
rect 6860 185 6890 286
rect 6948 193 6978 294
tri 6978 278 6994 294 nw
tri 7038 278 7054 294 ne
tri 6978 193 6994 209 sw
tri 7038 193 7054 209 se
rect 7054 193 7084 294
tri 6754 155 6784 185 ne
rect 6784 155 6860 185
tri 6860 155 6890 185 nw
tri 6948 163 6978 193 ne
rect 6978 163 7054 193
tri 7054 163 7084 193 nw
rect 7420 316 7450 377
tri 7450 316 7466 332 sw
rect 7614 324 7644 377
tri 7644 324 7660 340 sw
rect 7420 286 7526 316
tri 7526 286 7556 316 sw
rect 7614 294 7720 324
tri 7720 294 7750 324 sw
rect 7420 185 7450 286
tri 7450 270 7466 286 nw
tri 7510 270 7526 286 ne
tri 7450 185 7466 201 sw
tri 7510 185 7526 201 se
rect 7526 185 7556 286
rect 7614 193 7644 294
tri 7644 278 7660 294 nw
tri 7704 278 7720 294 ne
tri 7644 193 7660 209 sw
tri 7704 193 7720 209 se
rect 7720 193 7750 294
tri 7420 155 7450 185 ne
rect 7450 155 7526 185
tri 7526 155 7556 185 nw
tri 7614 163 7644 193 ne
rect 7644 163 7720 193
tri 7720 163 7750 193 nw
rect 8086 316 8116 377
tri 8116 316 8132 332 sw
rect 8280 324 8310 377
tri 8310 324 8326 340 sw
rect 8086 286 8192 316
tri 8192 286 8222 316 sw
rect 8280 294 8386 324
tri 8386 294 8416 324 sw
rect 8086 185 8116 286
tri 8116 270 8132 286 nw
tri 8176 270 8192 286 ne
tri 8116 185 8132 201 sw
tri 8176 185 8192 201 se
rect 8192 185 8222 286
rect 8280 193 8310 294
tri 8310 278 8326 294 nw
tri 8370 278 8386 294 ne
tri 8310 193 8326 209 sw
tri 8370 193 8386 209 se
rect 8386 193 8416 294
tri 8086 155 8116 185 ne
rect 8116 155 8192 185
tri 8192 155 8222 185 nw
tri 8280 163 8310 193 ne
rect 8310 163 8386 193
tri 8386 163 8416 193 nw
rect 8731 318 8761 379
tri 8761 318 8777 334 sw
rect 9031 318 9061 379
rect 8731 288 8837 318
tri 8837 288 8867 318 sw
rect 8731 187 8761 288
tri 8761 272 8777 288 nw
tri 8821 272 8837 288 ne
tri 8761 187 8777 203 sw
tri 8821 187 8837 203 se
rect 8837 187 8867 288
tri 8926 288 8956 318 se
rect 8956 288 9061 318
rect 8926 194 8956 288
tri 8956 272 8972 288 nw
tri 9015 272 9031 288 ne
tri 8956 194 8972 210 sw
tri 9015 194 9031 210 se
rect 9031 194 9061 288
tri 8731 157 8761 187 ne
rect 8761 157 8837 187
tri 8837 157 8867 187 nw
tri 8926 164 8956 194 ne
rect 8956 164 9031 194
tri 9031 164 9061 194 nw
rect 9233 326 9263 379
tri 9263 326 9279 342 sw
rect 9233 296 9339 326
tri 9339 296 9369 326 sw
rect 9233 195 9263 296
tri 9263 280 9279 296 nw
tri 9323 280 9339 296 ne
tri 9263 195 9279 211 sw
tri 9323 195 9339 211 se
rect 9339 195 9369 296
tri 9233 165 9263 195 ne
rect 9263 165 9339 195
tri 9339 165 9369 195 nw
rect 9714 316 9744 377
tri 9744 316 9760 332 sw
rect 9908 324 9938 377
tri 9938 324 9954 340 sw
rect 9714 286 9820 316
tri 9820 286 9850 316 sw
rect 9908 294 10014 324
tri 10014 294 10044 324 sw
rect 9714 185 9744 286
tri 9744 270 9760 286 nw
tri 9804 270 9820 286 ne
tri 9744 185 9760 201 sw
tri 9804 185 9820 201 se
rect 9820 185 9850 286
rect 9908 193 9938 294
tri 9938 278 9954 294 nw
tri 9998 278 10014 294 ne
tri 9938 193 9954 209 sw
tri 9998 193 10014 209 se
rect 10014 193 10044 294
tri 9714 155 9744 185 ne
rect 9744 155 9820 185
tri 9820 155 9850 185 nw
tri 9908 163 9938 193 ne
rect 9938 163 10014 193
tri 10014 163 10044 193 nw
rect 10380 316 10410 377
tri 10410 316 10426 332 sw
rect 10574 324 10604 377
tri 10604 324 10620 340 sw
rect 10380 286 10486 316
tri 10486 286 10516 316 sw
rect 10574 294 10680 324
tri 10680 294 10710 324 sw
rect 10380 185 10410 286
tri 10410 270 10426 286 nw
tri 10470 270 10486 286 ne
tri 10410 185 10426 201 sw
tri 10470 185 10486 201 se
rect 10486 185 10516 286
rect 10574 193 10604 294
tri 10604 278 10620 294 nw
tri 10664 278 10680 294 ne
tri 10604 193 10620 209 sw
tri 10664 193 10680 209 se
rect 10680 193 10710 294
tri 10380 155 10410 185 ne
rect 10410 155 10486 185
tri 10486 155 10516 185 nw
tri 10574 163 10604 193 ne
rect 10604 163 10680 193
tri 10680 163 10710 193 nw
rect 11046 316 11076 377
tri 11076 316 11092 332 sw
rect 11240 324 11270 377
tri 11270 324 11286 340 sw
rect 11046 286 11152 316
tri 11152 286 11182 316 sw
rect 11240 294 11346 324
tri 11346 294 11376 324 sw
rect 11046 185 11076 286
tri 11076 270 11092 286 nw
tri 11136 270 11152 286 ne
tri 11076 185 11092 201 sw
tri 11136 185 11152 201 se
rect 11152 185 11182 286
rect 11240 193 11270 294
tri 11270 278 11286 294 nw
tri 11330 278 11346 294 ne
tri 11270 193 11286 209 sw
tri 11330 193 11346 209 se
rect 11346 193 11376 294
tri 11046 155 11076 185 ne
rect 11076 155 11152 185
tri 11152 155 11182 185 nw
tri 11240 163 11270 193 ne
rect 11270 163 11346 193
tri 11346 163 11376 193 nw
rect 11712 316 11742 377
tri 11742 316 11758 332 sw
rect 11906 324 11936 377
tri 11936 324 11952 340 sw
rect 11712 286 11818 316
tri 11818 286 11848 316 sw
rect 11906 294 12012 324
tri 12012 294 12042 324 sw
rect 11712 185 11742 286
tri 11742 270 11758 286 nw
tri 11802 270 11818 286 ne
tri 11742 185 11758 201 sw
tri 11802 185 11818 201 se
rect 11818 185 11848 286
rect 11906 193 11936 294
tri 11936 278 11952 294 nw
tri 11996 278 12012 294 ne
tri 11936 193 11952 209 sw
tri 11996 193 12012 209 se
rect 12012 193 12042 294
tri 11712 155 11742 185 ne
rect 11742 155 11818 185
tri 11818 155 11848 185 nw
tri 11906 163 11936 193 ne
rect 11936 163 12012 193
tri 12012 163 12042 193 nw
rect 12378 316 12408 377
tri 12408 316 12424 332 sw
rect 12572 324 12602 377
tri 12602 324 12618 340 sw
rect 12378 286 12484 316
tri 12484 286 12514 316 sw
rect 12572 294 12678 324
tri 12678 294 12708 324 sw
rect 12378 185 12408 286
tri 12408 270 12424 286 nw
tri 12468 270 12484 286 ne
tri 12408 185 12424 201 sw
tri 12468 185 12484 201 se
rect 12484 185 12514 286
rect 12572 193 12602 294
tri 12602 278 12618 294 nw
tri 12662 278 12678 294 ne
tri 12602 193 12618 209 sw
tri 12662 193 12678 209 se
rect 12678 193 12708 294
tri 12378 155 12408 185 ne
rect 12408 155 12484 185
tri 12484 155 12514 185 nw
tri 12572 163 12602 193 ne
rect 12602 163 12678 193
tri 12678 163 12708 193 nw
rect 13044 316 13074 377
tri 13074 316 13090 332 sw
rect 13238 324 13268 377
tri 13268 324 13284 340 sw
rect 13044 286 13150 316
tri 13150 286 13180 316 sw
rect 13238 294 13344 324
tri 13344 294 13374 324 sw
rect 13044 185 13074 286
tri 13074 270 13090 286 nw
tri 13134 270 13150 286 ne
tri 13074 185 13090 201 sw
tri 13134 185 13150 201 se
rect 13150 185 13180 286
rect 13238 193 13268 294
tri 13268 278 13284 294 nw
tri 13328 278 13344 294 ne
tri 13268 193 13284 209 sw
tri 13328 193 13344 209 se
rect 13344 193 13374 294
tri 13044 155 13074 185 ne
rect 13074 155 13150 185
tri 13150 155 13180 185 nw
tri 13238 163 13268 193 ne
rect 13268 163 13344 193
tri 13344 163 13374 193 nw
rect 13710 316 13740 377
tri 13740 316 13756 332 sw
tri 13994 324 14010 340 se
rect 14010 324 14040 377
rect 13710 286 13816 316
tri 13816 286 13846 316 sw
tri 13904 294 13934 324 se
rect 13934 294 14040 324
rect 13710 185 13740 286
tri 13740 270 13756 286 nw
tri 13800 270 13816 286 ne
tri 13740 185 13756 201 sw
tri 13800 185 13816 201 se
rect 13816 185 13846 286
rect 13904 193 13934 294
tri 13934 278 13950 294 nw
tri 13994 278 14010 294 ne
tri 13934 193 13950 209 sw
tri 13994 193 14010 209 se
rect 14010 193 14040 294
tri 13710 155 13740 185 ne
rect 13740 155 13816 185
tri 13816 155 13846 185 nw
tri 13904 163 13934 193 ne
rect 13934 163 14010 193
tri 14010 163 14040 193 nw
rect 14376 316 14406 377
tri 14406 316 14422 332 sw
rect 14570 324 14600 377
tri 14600 324 14616 340 sw
rect 14376 286 14482 316
tri 14482 286 14512 316 sw
rect 14570 294 14676 324
tri 14676 294 14706 324 sw
rect 14376 185 14406 286
tri 14406 270 14422 286 nw
tri 14466 270 14482 286 ne
tri 14406 185 14422 201 sw
tri 14466 185 14482 201 se
rect 14482 185 14512 286
rect 14570 279 14601 294
tri 14601 279 14616 294 nw
tri 14660 279 14675 294 ne
rect 14675 279 14706 294
rect 14570 193 14600 279
tri 14600 193 14616 209 sw
tri 14660 193 14676 209 se
rect 14676 193 14706 279
tri 14376 155 14406 185 ne
rect 14406 155 14482 185
tri 14482 155 14512 185 nw
tri 14570 163 14600 193 ne
rect 14600 163 14676 193
tri 14676 163 14706 193 nw
<< pmos >>
rect 247 1050 277 1450
rect 335 1050 365 1450
rect 423 1050 453 1450
rect 511 1050 541 1450
rect 599 1050 629 1450
rect 687 1050 717 1450
rect 1149 1050 1179 1450
rect 1237 1050 1267 1450
rect 1325 1050 1355 1450
rect 1413 1050 1443 1450
rect 1815 1050 1845 1450
rect 1903 1050 1933 1450
rect 1991 1050 2021 1450
rect 2079 1050 2109 1450
rect 2481 1050 2511 1450
rect 2569 1050 2599 1450
rect 2657 1050 2687 1450
rect 2745 1050 2775 1450
rect 3147 1050 3177 1450
rect 3235 1050 3265 1450
rect 3323 1050 3353 1450
rect 3411 1050 3441 1450
rect 3813 1050 3843 1450
rect 3901 1050 3931 1450
rect 3989 1050 4019 1450
rect 4077 1050 4107 1450
rect 4539 1050 4569 1450
rect 4627 1050 4657 1450
rect 4715 1050 4745 1450
rect 4803 1050 4833 1450
rect 4891 1050 4921 1450
rect 4979 1050 5009 1450
rect 5441 1050 5471 1450
rect 5529 1050 5559 1450
rect 5617 1050 5647 1450
rect 5705 1050 5735 1450
rect 6107 1050 6137 1450
rect 6195 1050 6225 1450
rect 6283 1050 6313 1450
rect 6371 1050 6401 1450
rect 6773 1050 6803 1450
rect 6861 1050 6891 1450
rect 6949 1050 6979 1450
rect 7037 1050 7067 1450
rect 7439 1050 7469 1450
rect 7527 1050 7557 1450
rect 7615 1050 7645 1450
rect 7703 1050 7733 1450
rect 8105 1050 8135 1450
rect 8193 1050 8223 1450
rect 8281 1050 8311 1450
rect 8369 1050 8399 1450
rect 8831 1050 8861 1450
rect 8919 1050 8949 1450
rect 9007 1050 9037 1450
rect 9095 1050 9125 1450
rect 9183 1050 9213 1450
rect 9271 1050 9301 1450
rect 9733 1050 9763 1450
rect 9821 1050 9851 1450
rect 9909 1050 9939 1450
rect 9997 1050 10027 1450
rect 10399 1050 10429 1450
rect 10487 1050 10517 1450
rect 10575 1050 10605 1450
rect 10663 1050 10693 1450
rect 11065 1050 11095 1450
rect 11153 1050 11183 1450
rect 11241 1050 11271 1450
rect 11329 1050 11359 1450
rect 11731 1050 11761 1450
rect 11819 1050 11849 1450
rect 11907 1050 11937 1450
rect 11995 1050 12025 1450
rect 12397 1050 12427 1450
rect 12485 1050 12515 1450
rect 12573 1050 12603 1450
rect 12661 1050 12691 1450
rect 13063 1051 13093 1451
rect 13151 1051 13181 1451
rect 13239 1051 13269 1451
rect 13327 1051 13357 1451
rect 13727 1051 13757 1451
rect 13815 1051 13845 1451
rect 13903 1051 13933 1451
rect 13991 1051 14021 1451
rect 14395 1051 14425 1451
rect 14483 1051 14513 1451
rect 14571 1051 14601 1451
rect 14659 1051 14689 1451
<< ndiff >>
rect 91 363 147 379
rect 91 329 101 363
rect 135 329 147 363
rect 91 291 147 329
rect 177 363 447 379
rect 177 334 198 363
tri 177 318 193 334 ne
rect 193 329 198 334
rect 232 329 295 363
rect 329 329 392 363
rect 426 329 447 363
rect 193 318 447 329
rect 477 363 533 379
rect 477 329 489 363
rect 523 329 533 363
rect 91 257 101 291
rect 135 257 147 291
tri 253 288 283 318 ne
rect 283 291 342 318
rect 91 223 147 257
rect 91 189 101 223
rect 135 189 147 223
rect 91 157 147 189
tri 177 272 193 288 se
rect 193 272 237 288
tri 237 272 253 288 sw
rect 177 238 253 272
rect 177 204 198 238
rect 232 204 253 238
rect 177 203 253 204
tri 177 187 193 203 ne
rect 193 187 237 203
tri 237 187 253 203 nw
rect 283 257 295 291
rect 329 257 342 291
tri 342 288 372 318 nw
rect 283 223 342 257
rect 283 189 295 223
rect 329 189 342 223
tri 372 272 388 288 se
rect 388 272 431 288
tri 431 272 447 288 sw
rect 372 244 447 272
rect 372 210 393 244
rect 427 210 447 244
tri 372 194 388 210 ne
rect 388 194 431 210
tri 431 194 447 210 nw
tri 147 157 177 187 sw
tri 253 157 283 187 se
rect 283 164 342 189
tri 342 164 372 194 sw
tri 447 164 477 194 se
rect 477 164 533 329
rect 283 157 533 164
rect 91 153 533 157
rect 91 119 101 153
rect 135 119 295 153
rect 329 119 392 153
rect 426 119 489 153
rect 523 119 533 153
rect 91 103 533 119
rect 593 363 649 379
rect 593 329 603 363
rect 637 329 649 363
rect 593 291 649 329
rect 679 342 841 379
tri 679 326 695 342 ne
rect 695 326 841 342
tri 755 296 785 326 ne
rect 593 257 603 291
rect 637 257 649 291
rect 593 223 649 257
rect 593 189 603 223
rect 637 189 649 223
tri 679 280 695 296 se
rect 695 280 739 296
tri 739 280 755 296 sw
rect 679 247 755 280
rect 679 213 700 247
rect 734 213 755 247
rect 679 211 755 213
tri 679 195 695 211 ne
rect 695 195 739 211
tri 739 195 755 211 nw
rect 785 291 841 326
rect 785 257 797 291
rect 831 257 841 291
rect 785 223 841 257
rect 593 165 649 189
tri 649 165 679 195 sw
tri 755 165 785 195 se
rect 785 189 797 223
rect 831 189 841 223
rect 785 165 841 189
rect 593 153 841 165
rect 593 119 603 153
rect 637 119 700 153
rect 734 119 797 153
rect 831 119 841 153
rect 593 103 841 119
rect 1074 361 1130 377
rect 1074 327 1084 361
rect 1118 327 1130 361
rect 1074 289 1130 327
rect 1160 361 1324 377
rect 1160 332 1181 361
tri 1160 316 1176 332 ne
rect 1176 327 1181 332
rect 1215 327 1278 361
rect 1312 327 1324 361
rect 1176 316 1324 327
rect 1354 340 1516 377
tri 1354 324 1370 340 ne
rect 1370 324 1516 340
rect 1074 255 1084 289
rect 1118 255 1130 289
tri 1236 286 1266 316 ne
rect 1266 289 1324 316
tri 1430 294 1460 324 ne
rect 1074 221 1130 255
rect 1074 187 1084 221
rect 1118 187 1130 221
rect 1074 155 1130 187
tri 1160 270 1176 286 se
rect 1176 270 1220 286
tri 1220 270 1236 286 sw
rect 1160 236 1236 270
rect 1160 202 1181 236
rect 1215 202 1236 236
rect 1160 201 1236 202
tri 1160 185 1176 201 ne
rect 1176 185 1220 201
tri 1220 185 1236 201 nw
rect 1266 255 1278 289
rect 1312 255 1324 289
rect 1266 221 1324 255
rect 1266 187 1278 221
rect 1312 187 1324 221
tri 1354 278 1370 294 se
rect 1370 278 1414 294
tri 1414 278 1430 294 sw
rect 1354 245 1430 278
rect 1354 211 1375 245
rect 1409 211 1430 245
rect 1354 209 1430 211
tri 1354 193 1370 209 ne
rect 1370 193 1414 209
tri 1414 193 1430 209 nw
rect 1460 289 1516 324
rect 1460 255 1472 289
rect 1506 255 1516 289
rect 1460 221 1516 255
tri 1130 155 1160 185 sw
tri 1236 155 1266 185 se
rect 1266 163 1324 187
tri 1324 163 1354 193 sw
tri 1430 163 1460 193 se
rect 1460 187 1472 221
rect 1506 187 1516 221
rect 1460 163 1516 187
rect 1266 155 1516 163
rect 1074 151 1516 155
rect 1074 117 1084 151
rect 1118 117 1278 151
rect 1312 117 1375 151
rect 1409 117 1472 151
rect 1506 117 1516 151
rect 1074 101 1516 117
rect 1740 361 1796 377
rect 1740 327 1750 361
rect 1784 327 1796 361
rect 1740 289 1796 327
rect 1826 361 1990 377
rect 1826 332 1847 361
tri 1826 316 1842 332 ne
rect 1842 327 1847 332
rect 1881 327 1944 361
rect 1978 327 1990 361
rect 1842 316 1990 327
rect 2020 340 2182 377
tri 2020 324 2036 340 ne
rect 2036 324 2182 340
rect 1740 255 1750 289
rect 1784 255 1796 289
tri 1902 286 1932 316 ne
rect 1932 289 1990 316
tri 2096 294 2126 324 ne
rect 1740 221 1796 255
rect 1740 187 1750 221
rect 1784 187 1796 221
rect 1740 155 1796 187
tri 1826 270 1842 286 se
rect 1842 270 1886 286
tri 1886 270 1902 286 sw
rect 1826 236 1902 270
rect 1826 202 1847 236
rect 1881 202 1902 236
rect 1826 201 1902 202
tri 1826 185 1842 201 ne
rect 1842 185 1886 201
tri 1886 185 1902 201 nw
rect 1932 255 1944 289
rect 1978 255 1990 289
rect 1932 221 1990 255
rect 1932 187 1944 221
rect 1978 187 1990 221
tri 2020 278 2036 294 se
rect 2036 278 2080 294
tri 2080 278 2096 294 sw
rect 2020 245 2096 278
rect 2020 211 2041 245
rect 2075 211 2096 245
rect 2020 209 2096 211
tri 2020 193 2036 209 ne
rect 2036 193 2080 209
tri 2080 193 2096 209 nw
rect 2126 289 2182 324
rect 2126 255 2138 289
rect 2172 255 2182 289
rect 2126 221 2182 255
tri 1796 155 1826 185 sw
tri 1902 155 1932 185 se
rect 1932 163 1990 187
tri 1990 163 2020 193 sw
tri 2096 163 2126 193 se
rect 2126 187 2138 221
rect 2172 187 2182 221
rect 2126 163 2182 187
rect 1932 155 2182 163
rect 1740 151 2182 155
rect 1740 117 1750 151
rect 1784 117 1944 151
rect 1978 117 2041 151
rect 2075 117 2138 151
rect 2172 117 2182 151
rect 1740 101 2182 117
rect 2406 361 2462 377
rect 2406 327 2416 361
rect 2450 327 2462 361
rect 2406 289 2462 327
rect 2492 361 2656 377
rect 2492 332 2513 361
tri 2492 316 2508 332 ne
rect 2508 327 2513 332
rect 2547 327 2610 361
rect 2644 327 2656 361
rect 2508 316 2656 327
rect 2686 340 2848 377
tri 2686 324 2702 340 ne
rect 2702 324 2848 340
rect 2406 255 2416 289
rect 2450 255 2462 289
tri 2568 286 2598 316 ne
rect 2598 289 2656 316
tri 2762 294 2792 324 ne
rect 2406 221 2462 255
rect 2406 187 2416 221
rect 2450 187 2462 221
rect 2406 155 2462 187
tri 2492 270 2508 286 se
rect 2508 270 2552 286
tri 2552 270 2568 286 sw
rect 2492 236 2568 270
rect 2492 202 2513 236
rect 2547 202 2568 236
rect 2492 201 2568 202
tri 2492 185 2508 201 ne
rect 2508 185 2552 201
tri 2552 185 2568 201 nw
rect 2598 255 2610 289
rect 2644 255 2656 289
rect 2598 221 2656 255
rect 2598 187 2610 221
rect 2644 187 2656 221
tri 2686 278 2702 294 se
rect 2702 278 2746 294
tri 2746 278 2762 294 sw
rect 2686 245 2762 278
rect 2686 211 2707 245
rect 2741 211 2762 245
rect 2686 209 2762 211
tri 2686 193 2702 209 ne
rect 2702 193 2746 209
tri 2746 193 2762 209 nw
rect 2792 289 2848 324
rect 2792 255 2804 289
rect 2838 255 2848 289
rect 2792 221 2848 255
tri 2462 155 2492 185 sw
tri 2568 155 2598 185 se
rect 2598 163 2656 187
tri 2656 163 2686 193 sw
tri 2762 163 2792 193 se
rect 2792 187 2804 221
rect 2838 187 2848 221
rect 2792 163 2848 187
rect 2598 155 2848 163
rect 2406 151 2848 155
rect 2406 117 2416 151
rect 2450 117 2610 151
rect 2644 117 2707 151
rect 2741 117 2804 151
rect 2838 117 2848 151
rect 2406 101 2848 117
rect 3072 361 3128 377
rect 3072 327 3082 361
rect 3116 327 3128 361
rect 3072 289 3128 327
rect 3158 361 3322 377
rect 3158 332 3179 361
tri 3158 316 3174 332 ne
rect 3174 327 3179 332
rect 3213 327 3276 361
rect 3310 327 3322 361
rect 3174 316 3322 327
rect 3352 340 3514 377
tri 3352 324 3368 340 ne
rect 3368 324 3514 340
rect 3072 255 3082 289
rect 3116 255 3128 289
tri 3234 286 3264 316 ne
rect 3264 289 3322 316
tri 3428 294 3458 324 ne
rect 3072 221 3128 255
rect 3072 187 3082 221
rect 3116 187 3128 221
rect 3072 155 3128 187
tri 3158 270 3174 286 se
rect 3174 270 3218 286
tri 3218 270 3234 286 sw
rect 3158 236 3234 270
rect 3158 202 3179 236
rect 3213 202 3234 236
rect 3158 201 3234 202
tri 3158 185 3174 201 ne
rect 3174 185 3218 201
tri 3218 185 3234 201 nw
rect 3264 255 3276 289
rect 3310 255 3322 289
rect 3264 221 3322 255
rect 3264 187 3276 221
rect 3310 187 3322 221
tri 3352 278 3368 294 se
rect 3368 278 3412 294
tri 3412 278 3428 294 sw
rect 3352 245 3428 278
rect 3352 211 3373 245
rect 3407 211 3428 245
rect 3352 209 3428 211
tri 3352 193 3368 209 ne
rect 3368 193 3412 209
tri 3412 193 3428 209 nw
rect 3458 289 3514 324
rect 3458 255 3470 289
rect 3504 255 3514 289
rect 3458 221 3514 255
tri 3128 155 3158 185 sw
tri 3234 155 3264 185 se
rect 3264 163 3322 187
tri 3322 163 3352 193 sw
tri 3428 163 3458 193 se
rect 3458 187 3470 221
rect 3504 187 3514 221
rect 3458 163 3514 187
rect 3264 155 3514 163
rect 3072 151 3514 155
rect 3072 117 3082 151
rect 3116 117 3276 151
rect 3310 117 3373 151
rect 3407 117 3470 151
rect 3504 117 3514 151
rect 3072 101 3514 117
rect 3738 361 3794 377
rect 3738 327 3748 361
rect 3782 327 3794 361
rect 3738 289 3794 327
rect 3824 361 3988 377
rect 3824 332 3845 361
tri 3824 316 3840 332 ne
rect 3840 327 3845 332
rect 3879 327 3942 361
rect 3976 327 3988 361
rect 3840 316 3988 327
rect 4018 340 4180 377
tri 4018 324 4034 340 ne
rect 4034 324 4180 340
rect 3738 255 3748 289
rect 3782 255 3794 289
tri 3900 286 3930 316 ne
rect 3930 289 3988 316
tri 4094 294 4124 324 ne
rect 3738 221 3794 255
rect 3738 187 3748 221
rect 3782 187 3794 221
rect 3738 155 3794 187
tri 3824 270 3840 286 se
rect 3840 270 3884 286
tri 3884 270 3900 286 sw
rect 3824 236 3900 270
rect 3824 202 3845 236
rect 3879 202 3900 236
rect 3824 201 3900 202
tri 3824 185 3840 201 ne
rect 3840 185 3884 201
tri 3884 185 3900 201 nw
rect 3930 255 3942 289
rect 3976 255 3988 289
rect 3930 221 3988 255
rect 3930 187 3942 221
rect 3976 187 3988 221
tri 4018 278 4034 294 se
rect 4034 278 4078 294
tri 4078 278 4094 294 sw
rect 4018 245 4094 278
rect 4018 211 4039 245
rect 4073 211 4094 245
rect 4018 209 4094 211
tri 4018 193 4034 209 ne
rect 4034 193 4078 209
tri 4078 193 4094 209 nw
rect 4124 289 4180 324
rect 4124 255 4136 289
rect 4170 255 4180 289
rect 4124 221 4180 255
tri 3794 155 3824 185 sw
tri 3900 155 3930 185 se
rect 3930 163 3988 187
tri 3988 163 4018 193 sw
tri 4094 163 4124 193 se
rect 4124 187 4136 221
rect 4170 187 4180 221
rect 4124 163 4180 187
rect 3930 155 4180 163
rect 3738 151 4180 155
rect 3738 117 3748 151
rect 3782 117 3942 151
rect 3976 117 4039 151
rect 4073 117 4136 151
rect 4170 117 4180 151
rect 3738 101 4180 117
rect 4383 363 4439 379
rect 4383 329 4393 363
rect 4427 329 4439 363
rect 4383 291 4439 329
rect 4469 363 4739 379
rect 4469 334 4490 363
tri 4469 318 4485 334 ne
rect 4485 329 4490 334
rect 4524 329 4587 363
rect 4621 329 4684 363
rect 4718 329 4739 363
rect 4485 318 4739 329
rect 4769 363 4825 379
rect 4769 329 4781 363
rect 4815 329 4825 363
rect 4383 257 4393 291
rect 4427 257 4439 291
tri 4545 288 4575 318 ne
rect 4575 291 4634 318
rect 4383 223 4439 257
rect 4383 189 4393 223
rect 4427 189 4439 223
rect 4383 157 4439 189
tri 4469 272 4485 288 se
rect 4485 272 4529 288
tri 4529 272 4545 288 sw
rect 4469 238 4545 272
rect 4469 204 4490 238
rect 4524 204 4545 238
rect 4469 203 4545 204
tri 4469 187 4485 203 ne
rect 4485 187 4529 203
tri 4529 187 4545 203 nw
rect 4575 257 4587 291
rect 4621 257 4634 291
tri 4634 288 4664 318 nw
rect 4575 223 4634 257
rect 4575 189 4587 223
rect 4621 189 4634 223
tri 4664 272 4680 288 se
rect 4680 272 4723 288
tri 4723 272 4739 288 sw
rect 4664 244 4739 272
rect 4664 210 4685 244
rect 4719 210 4739 244
tri 4664 194 4680 210 ne
rect 4680 194 4723 210
tri 4723 194 4739 210 nw
tri 4439 157 4469 187 sw
tri 4545 157 4575 187 se
rect 4575 164 4634 189
tri 4634 164 4664 194 sw
tri 4739 164 4769 194 se
rect 4769 164 4825 329
rect 4575 157 4825 164
rect 4383 153 4825 157
rect 4383 119 4393 153
rect 4427 119 4587 153
rect 4621 119 4684 153
rect 4718 119 4781 153
rect 4815 119 4825 153
rect 4383 103 4825 119
rect 4885 363 4941 379
rect 4885 329 4895 363
rect 4929 329 4941 363
rect 4885 291 4941 329
rect 4971 342 5133 379
tri 4971 326 4987 342 ne
rect 4987 326 5133 342
tri 5047 296 5077 326 ne
rect 4885 257 4895 291
rect 4929 257 4941 291
rect 4885 223 4941 257
rect 4885 189 4895 223
rect 4929 189 4941 223
tri 4971 280 4987 296 se
rect 4987 280 5031 296
tri 5031 280 5047 296 sw
rect 4971 247 5047 280
rect 4971 213 4992 247
rect 5026 213 5047 247
rect 4971 211 5047 213
tri 4971 195 4987 211 ne
rect 4987 195 5031 211
tri 5031 195 5047 211 nw
rect 5077 291 5133 326
rect 5077 257 5089 291
rect 5123 257 5133 291
rect 5077 223 5133 257
rect 4885 165 4941 189
tri 4941 165 4971 195 sw
tri 5047 165 5077 195 se
rect 5077 189 5089 223
rect 5123 189 5133 223
rect 5077 165 5133 189
rect 4885 153 5133 165
rect 4885 119 4895 153
rect 4929 119 4992 153
rect 5026 119 5089 153
rect 5123 119 5133 153
rect 4885 103 5133 119
rect 5366 361 5422 377
rect 5366 327 5376 361
rect 5410 327 5422 361
rect 5366 289 5422 327
rect 5452 361 5616 377
rect 5452 332 5473 361
tri 5452 316 5468 332 ne
rect 5468 327 5473 332
rect 5507 327 5570 361
rect 5604 327 5616 361
rect 5468 316 5616 327
rect 5646 340 5808 377
tri 5646 324 5662 340 ne
rect 5662 324 5808 340
rect 5366 255 5376 289
rect 5410 255 5422 289
tri 5528 286 5558 316 ne
rect 5558 289 5616 316
tri 5722 294 5752 324 ne
rect 5366 221 5422 255
rect 5366 187 5376 221
rect 5410 187 5422 221
rect 5366 155 5422 187
tri 5452 270 5468 286 se
rect 5468 270 5512 286
tri 5512 270 5528 286 sw
rect 5452 236 5528 270
rect 5452 202 5473 236
rect 5507 202 5528 236
rect 5452 201 5528 202
tri 5452 185 5468 201 ne
rect 5468 185 5512 201
tri 5512 185 5528 201 nw
rect 5558 255 5570 289
rect 5604 255 5616 289
rect 5558 221 5616 255
rect 5558 187 5570 221
rect 5604 187 5616 221
tri 5646 278 5662 294 se
rect 5662 278 5706 294
tri 5706 278 5722 294 sw
rect 5646 245 5722 278
rect 5646 211 5667 245
rect 5701 211 5722 245
rect 5646 209 5722 211
tri 5646 193 5662 209 ne
rect 5662 193 5706 209
tri 5706 193 5722 209 nw
rect 5752 289 5808 324
rect 5752 255 5764 289
rect 5798 255 5808 289
rect 5752 221 5808 255
tri 5422 155 5452 185 sw
tri 5528 155 5558 185 se
rect 5558 163 5616 187
tri 5616 163 5646 193 sw
tri 5722 163 5752 193 se
rect 5752 187 5764 221
rect 5798 187 5808 221
rect 5752 163 5808 187
rect 5558 155 5808 163
rect 5366 151 5808 155
rect 5366 117 5376 151
rect 5410 117 5570 151
rect 5604 117 5667 151
rect 5701 117 5764 151
rect 5798 117 5808 151
rect 5366 101 5808 117
rect 6032 361 6088 377
rect 6032 327 6042 361
rect 6076 327 6088 361
rect 6032 289 6088 327
rect 6118 361 6282 377
rect 6118 332 6139 361
tri 6118 316 6134 332 ne
rect 6134 327 6139 332
rect 6173 327 6236 361
rect 6270 327 6282 361
rect 6134 316 6282 327
rect 6312 340 6474 377
tri 6312 324 6328 340 ne
rect 6328 324 6474 340
rect 6032 255 6042 289
rect 6076 255 6088 289
tri 6194 286 6224 316 ne
rect 6224 289 6282 316
tri 6388 294 6418 324 ne
rect 6032 221 6088 255
rect 6032 187 6042 221
rect 6076 187 6088 221
rect 6032 155 6088 187
tri 6118 270 6134 286 se
rect 6134 270 6178 286
tri 6178 270 6194 286 sw
rect 6118 236 6194 270
rect 6118 202 6139 236
rect 6173 202 6194 236
rect 6118 201 6194 202
tri 6118 185 6134 201 ne
rect 6134 185 6178 201
tri 6178 185 6194 201 nw
rect 6224 255 6236 289
rect 6270 255 6282 289
rect 6224 221 6282 255
rect 6224 187 6236 221
rect 6270 187 6282 221
tri 6312 278 6328 294 se
rect 6328 278 6372 294
tri 6372 278 6388 294 sw
rect 6312 245 6388 278
rect 6312 211 6333 245
rect 6367 211 6388 245
rect 6312 209 6388 211
tri 6312 193 6328 209 ne
rect 6328 193 6372 209
tri 6372 193 6388 209 nw
rect 6418 289 6474 324
rect 6418 255 6430 289
rect 6464 255 6474 289
rect 6418 221 6474 255
tri 6088 155 6118 185 sw
tri 6194 155 6224 185 se
rect 6224 163 6282 187
tri 6282 163 6312 193 sw
tri 6388 163 6418 193 se
rect 6418 187 6430 221
rect 6464 187 6474 221
rect 6418 163 6474 187
rect 6224 155 6474 163
rect 6032 151 6474 155
rect 6032 117 6042 151
rect 6076 117 6236 151
rect 6270 117 6333 151
rect 6367 117 6430 151
rect 6464 117 6474 151
rect 6032 101 6474 117
rect 6698 361 6754 377
rect 6698 327 6708 361
rect 6742 327 6754 361
rect 6698 289 6754 327
rect 6784 361 6948 377
rect 6784 332 6805 361
tri 6784 316 6800 332 ne
rect 6800 327 6805 332
rect 6839 327 6902 361
rect 6936 327 6948 361
rect 6800 316 6948 327
rect 6978 340 7140 377
tri 6978 324 6994 340 ne
rect 6994 324 7140 340
rect 6698 255 6708 289
rect 6742 255 6754 289
tri 6860 286 6890 316 ne
rect 6890 289 6948 316
tri 7054 294 7084 324 ne
rect 6698 221 6754 255
rect 6698 187 6708 221
rect 6742 187 6754 221
rect 6698 155 6754 187
tri 6784 270 6800 286 se
rect 6800 270 6844 286
tri 6844 270 6860 286 sw
rect 6784 236 6860 270
rect 6784 202 6805 236
rect 6839 202 6860 236
rect 6784 201 6860 202
tri 6784 185 6800 201 ne
rect 6800 185 6844 201
tri 6844 185 6860 201 nw
rect 6890 255 6902 289
rect 6936 255 6948 289
rect 6890 221 6948 255
rect 6890 187 6902 221
rect 6936 187 6948 221
tri 6978 278 6994 294 se
rect 6994 278 7038 294
tri 7038 278 7054 294 sw
rect 6978 245 7054 278
rect 6978 211 6999 245
rect 7033 211 7054 245
rect 6978 209 7054 211
tri 6978 193 6994 209 ne
rect 6994 193 7038 209
tri 7038 193 7054 209 nw
rect 7084 289 7140 324
rect 7084 255 7096 289
rect 7130 255 7140 289
rect 7084 221 7140 255
tri 6754 155 6784 185 sw
tri 6860 155 6890 185 se
rect 6890 163 6948 187
tri 6948 163 6978 193 sw
tri 7054 163 7084 193 se
rect 7084 187 7096 221
rect 7130 187 7140 221
rect 7084 163 7140 187
rect 6890 155 7140 163
rect 6698 151 7140 155
rect 6698 117 6708 151
rect 6742 117 6902 151
rect 6936 117 6999 151
rect 7033 117 7096 151
rect 7130 117 7140 151
rect 6698 101 7140 117
rect 7364 361 7420 377
rect 7364 327 7374 361
rect 7408 327 7420 361
rect 7364 289 7420 327
rect 7450 361 7614 377
rect 7450 332 7471 361
tri 7450 316 7466 332 ne
rect 7466 327 7471 332
rect 7505 327 7568 361
rect 7602 327 7614 361
rect 7466 316 7614 327
rect 7644 340 7806 377
tri 7644 324 7660 340 ne
rect 7660 324 7806 340
rect 7364 255 7374 289
rect 7408 255 7420 289
tri 7526 286 7556 316 ne
rect 7556 289 7614 316
tri 7720 294 7750 324 ne
rect 7364 221 7420 255
rect 7364 187 7374 221
rect 7408 187 7420 221
rect 7364 155 7420 187
tri 7450 270 7466 286 se
rect 7466 270 7510 286
tri 7510 270 7526 286 sw
rect 7450 236 7526 270
rect 7450 202 7471 236
rect 7505 202 7526 236
rect 7450 201 7526 202
tri 7450 185 7466 201 ne
rect 7466 185 7510 201
tri 7510 185 7526 201 nw
rect 7556 255 7568 289
rect 7602 255 7614 289
rect 7556 221 7614 255
rect 7556 187 7568 221
rect 7602 187 7614 221
tri 7644 278 7660 294 se
rect 7660 278 7704 294
tri 7704 278 7720 294 sw
rect 7644 245 7720 278
rect 7644 211 7665 245
rect 7699 211 7720 245
rect 7644 209 7720 211
tri 7644 193 7660 209 ne
rect 7660 193 7704 209
tri 7704 193 7720 209 nw
rect 7750 289 7806 324
rect 7750 255 7762 289
rect 7796 255 7806 289
rect 7750 221 7806 255
tri 7420 155 7450 185 sw
tri 7526 155 7556 185 se
rect 7556 163 7614 187
tri 7614 163 7644 193 sw
tri 7720 163 7750 193 se
rect 7750 187 7762 221
rect 7796 187 7806 221
rect 7750 163 7806 187
rect 7556 155 7806 163
rect 7364 151 7806 155
rect 7364 117 7374 151
rect 7408 117 7568 151
rect 7602 117 7665 151
rect 7699 117 7762 151
rect 7796 117 7806 151
rect 7364 101 7806 117
rect 8030 361 8086 377
rect 8030 327 8040 361
rect 8074 327 8086 361
rect 8030 289 8086 327
rect 8116 361 8280 377
rect 8116 332 8137 361
tri 8116 316 8132 332 ne
rect 8132 327 8137 332
rect 8171 327 8234 361
rect 8268 327 8280 361
rect 8132 316 8280 327
rect 8310 340 8472 377
tri 8310 324 8326 340 ne
rect 8326 324 8472 340
rect 8030 255 8040 289
rect 8074 255 8086 289
tri 8192 286 8222 316 ne
rect 8222 289 8280 316
tri 8386 294 8416 324 ne
rect 8030 221 8086 255
rect 8030 187 8040 221
rect 8074 187 8086 221
rect 8030 155 8086 187
tri 8116 270 8132 286 se
rect 8132 270 8176 286
tri 8176 270 8192 286 sw
rect 8116 236 8192 270
rect 8116 202 8137 236
rect 8171 202 8192 236
rect 8116 201 8192 202
tri 8116 185 8132 201 ne
rect 8132 185 8176 201
tri 8176 185 8192 201 nw
rect 8222 255 8234 289
rect 8268 255 8280 289
rect 8222 221 8280 255
rect 8222 187 8234 221
rect 8268 187 8280 221
tri 8310 278 8326 294 se
rect 8326 278 8370 294
tri 8370 278 8386 294 sw
rect 8310 245 8386 278
rect 8310 211 8331 245
rect 8365 211 8386 245
rect 8310 209 8386 211
tri 8310 193 8326 209 ne
rect 8326 193 8370 209
tri 8370 193 8386 209 nw
rect 8416 289 8472 324
rect 8416 255 8428 289
rect 8462 255 8472 289
rect 8416 221 8472 255
tri 8086 155 8116 185 sw
tri 8192 155 8222 185 se
rect 8222 163 8280 187
tri 8280 163 8310 193 sw
tri 8386 163 8416 193 se
rect 8416 187 8428 221
rect 8462 187 8472 221
rect 8416 163 8472 187
rect 8222 155 8472 163
rect 8030 151 8472 155
rect 8030 117 8040 151
rect 8074 117 8234 151
rect 8268 117 8331 151
rect 8365 117 8428 151
rect 8462 117 8472 151
rect 8030 101 8472 117
rect 8675 363 8731 379
rect 8675 329 8685 363
rect 8719 329 8731 363
rect 8675 291 8731 329
rect 8761 363 9031 379
rect 8761 334 8782 363
tri 8761 318 8777 334 ne
rect 8777 329 8782 334
rect 8816 329 8879 363
rect 8913 329 8976 363
rect 9010 329 9031 363
rect 8777 318 9031 329
rect 9061 363 9117 379
rect 9061 329 9073 363
rect 9107 329 9117 363
rect 8675 257 8685 291
rect 8719 257 8731 291
tri 8837 288 8867 318 ne
rect 8867 291 8926 318
rect 8675 223 8731 257
rect 8675 189 8685 223
rect 8719 189 8731 223
rect 8675 157 8731 189
tri 8761 272 8777 288 se
rect 8777 272 8821 288
tri 8821 272 8837 288 sw
rect 8761 238 8837 272
rect 8761 204 8782 238
rect 8816 204 8837 238
rect 8761 203 8837 204
tri 8761 187 8777 203 ne
rect 8777 187 8821 203
tri 8821 187 8837 203 nw
rect 8867 257 8879 291
rect 8913 257 8926 291
tri 8926 288 8956 318 nw
rect 8867 223 8926 257
rect 8867 189 8879 223
rect 8913 189 8926 223
tri 8956 272 8972 288 se
rect 8972 272 9015 288
tri 9015 272 9031 288 sw
rect 8956 244 9031 272
rect 8956 210 8977 244
rect 9011 210 9031 244
tri 8956 194 8972 210 ne
rect 8972 194 9015 210
tri 9015 194 9031 210 nw
tri 8731 157 8761 187 sw
tri 8837 157 8867 187 se
rect 8867 164 8926 189
tri 8926 164 8956 194 sw
tri 9031 164 9061 194 se
rect 9061 164 9117 329
rect 8867 157 9117 164
rect 8675 153 9117 157
rect 8675 119 8685 153
rect 8719 119 8879 153
rect 8913 119 8976 153
rect 9010 119 9073 153
rect 9107 119 9117 153
rect 8675 103 9117 119
rect 9177 363 9233 379
rect 9177 329 9187 363
rect 9221 329 9233 363
rect 9177 291 9233 329
rect 9263 342 9425 379
tri 9263 326 9279 342 ne
rect 9279 326 9425 342
tri 9339 296 9369 326 ne
rect 9177 257 9187 291
rect 9221 257 9233 291
rect 9177 223 9233 257
rect 9177 189 9187 223
rect 9221 189 9233 223
tri 9263 280 9279 296 se
rect 9279 280 9323 296
tri 9323 280 9339 296 sw
rect 9263 247 9339 280
rect 9263 213 9284 247
rect 9318 213 9339 247
rect 9263 211 9339 213
tri 9263 195 9279 211 ne
rect 9279 195 9323 211
tri 9323 195 9339 211 nw
rect 9369 291 9425 326
rect 9369 257 9381 291
rect 9415 257 9425 291
rect 9369 223 9425 257
rect 9177 165 9233 189
tri 9233 165 9263 195 sw
tri 9339 165 9369 195 se
rect 9369 189 9381 223
rect 9415 189 9425 223
rect 9369 165 9425 189
rect 9177 153 9425 165
rect 9177 119 9187 153
rect 9221 119 9284 153
rect 9318 119 9381 153
rect 9415 119 9425 153
rect 9177 103 9425 119
rect 9658 361 9714 377
rect 9658 327 9668 361
rect 9702 327 9714 361
rect 9658 289 9714 327
rect 9744 361 9908 377
rect 9744 332 9765 361
tri 9744 316 9760 332 ne
rect 9760 327 9765 332
rect 9799 327 9862 361
rect 9896 327 9908 361
rect 9760 316 9908 327
rect 9938 340 10100 377
tri 9938 324 9954 340 ne
rect 9954 324 10100 340
rect 9658 255 9668 289
rect 9702 255 9714 289
tri 9820 286 9850 316 ne
rect 9850 289 9908 316
tri 10014 294 10044 324 ne
rect 9658 221 9714 255
rect 9658 187 9668 221
rect 9702 187 9714 221
rect 9658 155 9714 187
tri 9744 270 9760 286 se
rect 9760 270 9804 286
tri 9804 270 9820 286 sw
rect 9744 236 9820 270
rect 9744 202 9765 236
rect 9799 202 9820 236
rect 9744 201 9820 202
tri 9744 185 9760 201 ne
rect 9760 185 9804 201
tri 9804 185 9820 201 nw
rect 9850 255 9862 289
rect 9896 255 9908 289
rect 9850 221 9908 255
rect 9850 187 9862 221
rect 9896 187 9908 221
tri 9938 278 9954 294 se
rect 9954 278 9998 294
tri 9998 278 10014 294 sw
rect 9938 245 10014 278
rect 9938 211 9959 245
rect 9993 211 10014 245
rect 9938 209 10014 211
tri 9938 193 9954 209 ne
rect 9954 193 9998 209
tri 9998 193 10014 209 nw
rect 10044 289 10100 324
rect 10044 255 10056 289
rect 10090 255 10100 289
rect 10044 221 10100 255
tri 9714 155 9744 185 sw
tri 9820 155 9850 185 se
rect 9850 163 9908 187
tri 9908 163 9938 193 sw
tri 10014 163 10044 193 se
rect 10044 187 10056 221
rect 10090 187 10100 221
rect 10044 163 10100 187
rect 9850 155 10100 163
rect 9658 151 10100 155
rect 9658 117 9668 151
rect 9702 117 9862 151
rect 9896 117 9959 151
rect 9993 117 10056 151
rect 10090 117 10100 151
rect 9658 101 10100 117
rect 10324 361 10380 377
rect 10324 327 10334 361
rect 10368 327 10380 361
rect 10324 289 10380 327
rect 10410 361 10574 377
rect 10410 332 10431 361
tri 10410 316 10426 332 ne
rect 10426 327 10431 332
rect 10465 327 10528 361
rect 10562 327 10574 361
rect 10426 316 10574 327
rect 10604 340 10766 377
tri 10604 324 10620 340 ne
rect 10620 324 10766 340
rect 10324 255 10334 289
rect 10368 255 10380 289
tri 10486 286 10516 316 ne
rect 10516 289 10574 316
tri 10680 294 10710 324 ne
rect 10324 221 10380 255
rect 10324 187 10334 221
rect 10368 187 10380 221
rect 10324 155 10380 187
tri 10410 270 10426 286 se
rect 10426 270 10470 286
tri 10470 270 10486 286 sw
rect 10410 236 10486 270
rect 10410 202 10431 236
rect 10465 202 10486 236
rect 10410 201 10486 202
tri 10410 185 10426 201 ne
rect 10426 185 10470 201
tri 10470 185 10486 201 nw
rect 10516 255 10528 289
rect 10562 255 10574 289
rect 10516 221 10574 255
rect 10516 187 10528 221
rect 10562 187 10574 221
tri 10604 278 10620 294 se
rect 10620 278 10664 294
tri 10664 278 10680 294 sw
rect 10604 245 10680 278
rect 10604 211 10625 245
rect 10659 211 10680 245
rect 10604 209 10680 211
tri 10604 193 10620 209 ne
rect 10620 193 10664 209
tri 10664 193 10680 209 nw
rect 10710 289 10766 324
rect 10710 255 10722 289
rect 10756 255 10766 289
rect 10710 221 10766 255
tri 10380 155 10410 185 sw
tri 10486 155 10516 185 se
rect 10516 163 10574 187
tri 10574 163 10604 193 sw
tri 10680 163 10710 193 se
rect 10710 187 10722 221
rect 10756 187 10766 221
rect 10710 163 10766 187
rect 10516 155 10766 163
rect 10324 151 10766 155
rect 10324 117 10334 151
rect 10368 117 10528 151
rect 10562 117 10625 151
rect 10659 117 10722 151
rect 10756 117 10766 151
rect 10324 101 10766 117
rect 10990 361 11046 377
rect 10990 327 11000 361
rect 11034 327 11046 361
rect 10990 289 11046 327
rect 11076 361 11240 377
rect 11076 332 11097 361
tri 11076 316 11092 332 ne
rect 11092 327 11097 332
rect 11131 327 11194 361
rect 11228 327 11240 361
rect 11092 316 11240 327
rect 11270 340 11432 377
tri 11270 324 11286 340 ne
rect 11286 324 11432 340
rect 10990 255 11000 289
rect 11034 255 11046 289
tri 11152 286 11182 316 ne
rect 11182 289 11240 316
tri 11346 294 11376 324 ne
rect 10990 221 11046 255
rect 10990 187 11000 221
rect 11034 187 11046 221
rect 10990 155 11046 187
tri 11076 270 11092 286 se
rect 11092 270 11136 286
tri 11136 270 11152 286 sw
rect 11076 236 11152 270
rect 11076 202 11097 236
rect 11131 202 11152 236
rect 11076 201 11152 202
tri 11076 185 11092 201 ne
rect 11092 185 11136 201
tri 11136 185 11152 201 nw
rect 11182 255 11194 289
rect 11228 255 11240 289
rect 11182 221 11240 255
rect 11182 187 11194 221
rect 11228 187 11240 221
tri 11270 278 11286 294 se
rect 11286 278 11330 294
tri 11330 278 11346 294 sw
rect 11270 245 11346 278
rect 11270 211 11291 245
rect 11325 211 11346 245
rect 11270 209 11346 211
tri 11270 193 11286 209 ne
rect 11286 193 11330 209
tri 11330 193 11346 209 nw
rect 11376 289 11432 324
rect 11376 255 11388 289
rect 11422 255 11432 289
rect 11376 221 11432 255
tri 11046 155 11076 185 sw
tri 11152 155 11182 185 se
rect 11182 163 11240 187
tri 11240 163 11270 193 sw
tri 11346 163 11376 193 se
rect 11376 187 11388 221
rect 11422 187 11432 221
rect 11376 163 11432 187
rect 11182 155 11432 163
rect 10990 151 11432 155
rect 10990 117 11000 151
rect 11034 117 11194 151
rect 11228 117 11291 151
rect 11325 117 11388 151
rect 11422 117 11432 151
rect 10990 101 11432 117
rect 11656 361 11712 377
rect 11656 327 11666 361
rect 11700 327 11712 361
rect 11656 289 11712 327
rect 11742 361 11906 377
rect 11742 332 11763 361
tri 11742 316 11758 332 ne
rect 11758 327 11763 332
rect 11797 327 11860 361
rect 11894 327 11906 361
rect 11758 316 11906 327
rect 11936 340 12098 377
tri 11936 324 11952 340 ne
rect 11952 324 12098 340
rect 11656 255 11666 289
rect 11700 255 11712 289
tri 11818 286 11848 316 ne
rect 11848 289 11906 316
tri 12012 294 12042 324 ne
rect 11656 221 11712 255
rect 11656 187 11666 221
rect 11700 187 11712 221
rect 11656 155 11712 187
tri 11742 270 11758 286 se
rect 11758 270 11802 286
tri 11802 270 11818 286 sw
rect 11742 236 11818 270
rect 11742 202 11763 236
rect 11797 202 11818 236
rect 11742 201 11818 202
tri 11742 185 11758 201 ne
rect 11758 185 11802 201
tri 11802 185 11818 201 nw
rect 11848 255 11860 289
rect 11894 255 11906 289
rect 11848 221 11906 255
rect 11848 187 11860 221
rect 11894 187 11906 221
tri 11936 278 11952 294 se
rect 11952 278 11996 294
tri 11996 278 12012 294 sw
rect 11936 245 12012 278
rect 11936 211 11957 245
rect 11991 211 12012 245
rect 11936 209 12012 211
tri 11936 193 11952 209 ne
rect 11952 193 11996 209
tri 11996 193 12012 209 nw
rect 12042 289 12098 324
rect 12042 255 12054 289
rect 12088 255 12098 289
rect 12042 221 12098 255
tri 11712 155 11742 185 sw
tri 11818 155 11848 185 se
rect 11848 163 11906 187
tri 11906 163 11936 193 sw
tri 12012 163 12042 193 se
rect 12042 187 12054 221
rect 12088 187 12098 221
rect 12042 163 12098 187
rect 11848 155 12098 163
rect 11656 151 12098 155
rect 11656 117 11666 151
rect 11700 117 11860 151
rect 11894 117 11957 151
rect 11991 117 12054 151
rect 12088 117 12098 151
rect 11656 101 12098 117
rect 12322 361 12378 377
rect 12322 327 12332 361
rect 12366 327 12378 361
rect 12322 289 12378 327
rect 12408 361 12572 377
rect 12408 332 12429 361
tri 12408 316 12424 332 ne
rect 12424 327 12429 332
rect 12463 327 12526 361
rect 12560 327 12572 361
rect 12424 316 12572 327
rect 12602 340 12764 377
tri 12602 324 12618 340 ne
rect 12618 324 12764 340
rect 12322 255 12332 289
rect 12366 255 12378 289
tri 12484 286 12514 316 ne
rect 12514 289 12572 316
tri 12678 294 12708 324 ne
rect 12322 221 12378 255
rect 12322 187 12332 221
rect 12366 187 12378 221
rect 12322 155 12378 187
tri 12408 270 12424 286 se
rect 12424 270 12468 286
tri 12468 270 12484 286 sw
rect 12408 236 12484 270
rect 12408 202 12429 236
rect 12463 202 12484 236
rect 12408 201 12484 202
tri 12408 185 12424 201 ne
rect 12424 185 12468 201
tri 12468 185 12484 201 nw
rect 12514 255 12526 289
rect 12560 255 12572 289
rect 12514 221 12572 255
rect 12514 187 12526 221
rect 12560 187 12572 221
tri 12602 278 12618 294 se
rect 12618 278 12662 294
tri 12662 278 12678 294 sw
rect 12602 245 12678 278
rect 12602 211 12623 245
rect 12657 211 12678 245
rect 12602 209 12678 211
tri 12602 193 12618 209 ne
rect 12618 193 12662 209
tri 12662 193 12678 209 nw
rect 12708 289 12764 324
rect 12708 255 12720 289
rect 12754 255 12764 289
rect 12708 221 12764 255
tri 12378 155 12408 185 sw
tri 12484 155 12514 185 se
rect 12514 163 12572 187
tri 12572 163 12602 193 sw
tri 12678 163 12708 193 se
rect 12708 187 12720 221
rect 12754 187 12764 221
rect 12708 163 12764 187
rect 12514 155 12764 163
rect 12322 151 12764 155
rect 12322 117 12332 151
rect 12366 117 12526 151
rect 12560 117 12623 151
rect 12657 117 12720 151
rect 12754 117 12764 151
rect 12322 101 12764 117
rect 12988 361 13044 377
rect 12988 327 12998 361
rect 13032 327 13044 361
rect 12988 289 13044 327
rect 13074 361 13238 377
rect 13074 332 13095 361
tri 13074 316 13090 332 ne
rect 13090 327 13095 332
rect 13129 327 13192 361
rect 13226 327 13238 361
rect 13090 316 13238 327
rect 13268 361 13428 377
rect 13268 340 13386 361
tri 13268 324 13284 340 ne
rect 13284 327 13386 340
rect 13420 327 13428 361
rect 13284 324 13428 327
rect 12988 255 12998 289
rect 13032 255 13044 289
tri 13150 286 13180 316 ne
rect 13180 289 13238 316
tri 13344 294 13374 324 ne
rect 12988 221 13044 255
rect 12988 187 12998 221
rect 13032 187 13044 221
rect 12988 155 13044 187
tri 13074 270 13090 286 se
rect 13090 270 13134 286
tri 13134 270 13150 286 sw
rect 13074 236 13150 270
rect 13074 202 13095 236
rect 13129 202 13150 236
rect 13074 201 13150 202
tri 13074 185 13090 201 ne
rect 13090 185 13134 201
tri 13134 185 13150 201 nw
rect 13180 255 13192 289
rect 13226 255 13238 289
rect 13180 221 13238 255
rect 13180 187 13192 221
rect 13226 187 13238 221
tri 13268 278 13284 294 se
rect 13284 278 13328 294
tri 13328 278 13344 294 sw
rect 13268 245 13344 278
rect 13268 211 13288 245
rect 13322 211 13344 245
rect 13268 209 13344 211
tri 13268 193 13284 209 ne
rect 13284 193 13328 209
tri 13328 193 13344 209 nw
rect 13374 289 13428 324
rect 13374 255 13386 289
rect 13420 255 13428 289
rect 13374 221 13428 255
tri 13044 155 13074 185 sw
tri 13150 155 13180 185 se
rect 13180 163 13238 187
tri 13238 163 13268 193 sw
tri 13344 163 13374 193 se
rect 13374 187 13386 221
rect 13420 187 13428 221
rect 13374 163 13428 187
rect 13180 155 13428 163
rect 12988 151 13428 155
rect 12988 117 12998 151
rect 13032 117 13192 151
rect 13226 117 13288 151
rect 13322 117 13386 151
rect 13420 117 13428 151
rect 12988 101 13428 117
rect 13654 361 13710 377
rect 13654 327 13664 361
rect 13698 327 13710 361
rect 13654 289 13710 327
rect 13740 361 14010 377
rect 13740 332 13761 361
tri 13740 316 13756 332 ne
rect 13756 327 13761 332
rect 13795 327 13858 361
rect 13892 340 14010 361
rect 13892 327 13994 340
rect 13756 324 13994 327
tri 13994 324 14010 340 nw
rect 14040 361 14096 377
rect 14040 327 14052 361
rect 14086 327 14096 361
rect 13756 316 13904 324
rect 13654 255 13664 289
rect 13698 255 13710 289
tri 13816 286 13846 316 ne
rect 13846 289 13904 316
tri 13904 294 13934 324 nw
rect 13654 221 13710 255
rect 13654 187 13664 221
rect 13698 187 13710 221
rect 13654 155 13710 187
tri 13740 270 13756 286 se
rect 13756 270 13800 286
tri 13800 270 13816 286 sw
rect 13740 236 13816 270
rect 13740 202 13761 236
rect 13795 202 13816 236
rect 13740 201 13816 202
tri 13740 185 13756 201 ne
rect 13756 185 13800 201
tri 13800 185 13816 201 nw
rect 13846 255 13858 289
rect 13892 255 13904 289
rect 13846 221 13904 255
rect 13846 187 13858 221
rect 13892 187 13904 221
tri 13934 278 13950 294 se
rect 13950 278 13994 294
tri 13994 278 14010 294 sw
rect 13934 245 14010 278
rect 13934 211 13955 245
rect 13989 211 14010 245
rect 13934 209 14010 211
tri 13934 193 13950 209 ne
rect 13950 193 13994 209
tri 13994 193 14010 209 nw
rect 14040 289 14096 327
rect 14040 255 14052 289
rect 14086 255 14096 289
rect 14040 221 14096 255
tri 13710 155 13740 185 sw
tri 13816 155 13846 185 se
rect 13846 163 13904 187
tri 13904 163 13934 193 sw
tri 14010 163 14040 193 se
rect 14040 187 14052 221
rect 14086 187 14096 221
rect 14040 163 14096 187
rect 13846 155 14096 163
rect 13654 151 14096 155
rect 13654 117 13664 151
rect 13698 117 13858 151
rect 13892 117 13955 151
rect 13989 117 14052 151
rect 14086 117 14096 151
rect 13654 101 14096 117
rect 14320 361 14376 377
rect 14320 327 14330 361
rect 14364 327 14376 361
rect 14320 289 14376 327
rect 14406 361 14570 377
rect 14406 332 14427 361
tri 14406 316 14422 332 ne
rect 14422 327 14427 332
rect 14461 327 14524 361
rect 14558 327 14570 361
rect 14422 316 14570 327
rect 14600 340 14762 377
tri 14600 324 14616 340 ne
rect 14616 324 14762 340
rect 14320 255 14330 289
rect 14364 255 14376 289
tri 14482 286 14512 316 ne
rect 14512 289 14570 316
tri 14676 294 14706 324 ne
rect 14320 221 14376 255
rect 14320 187 14330 221
rect 14364 187 14376 221
rect 14320 155 14376 187
tri 14406 270 14422 286 se
rect 14422 270 14466 286
tri 14466 270 14482 286 sw
rect 14406 236 14482 270
rect 14406 202 14427 236
rect 14461 202 14482 236
rect 14406 201 14482 202
tri 14406 185 14422 201 ne
rect 14422 185 14466 201
tri 14466 185 14482 201 nw
rect 14512 255 14524 289
rect 14558 255 14570 289
tri 14601 279 14616 294 se
rect 14616 279 14660 294
tri 14660 279 14675 294 sw
rect 14706 289 14762 324
rect 14512 221 14570 255
rect 14512 187 14524 221
rect 14558 187 14570 221
rect 14600 245 14676 279
rect 14600 211 14621 245
rect 14655 211 14676 245
rect 14600 209 14676 211
tri 14600 193 14616 209 ne
rect 14616 193 14660 209
tri 14660 193 14676 209 nw
rect 14706 255 14718 289
rect 14752 255 14762 289
rect 14706 221 14762 255
tri 14376 155 14406 185 sw
tri 14482 155 14512 185 se
rect 14512 163 14570 187
tri 14570 163 14600 193 sw
tri 14676 163 14706 193 se
rect 14706 187 14718 221
rect 14752 187 14762 221
rect 14706 163 14762 187
rect 14512 155 14762 163
rect 14320 151 14762 155
rect 14320 117 14330 151
rect 14364 117 14524 151
rect 14558 117 14621 151
rect 14655 117 14718 151
rect 14752 117 14762 151
rect 14320 101 14762 117
<< pdiff >>
rect 191 1412 247 1450
rect 191 1378 201 1412
rect 235 1378 247 1412
rect 191 1344 247 1378
rect 191 1310 201 1344
rect 235 1310 247 1344
rect 191 1276 247 1310
rect 191 1242 201 1276
rect 235 1242 247 1276
rect 191 1208 247 1242
rect 191 1174 201 1208
rect 235 1174 247 1208
rect 191 1139 247 1174
rect 191 1105 201 1139
rect 235 1105 247 1139
rect 191 1050 247 1105
rect 277 1412 335 1450
rect 277 1378 289 1412
rect 323 1378 335 1412
rect 277 1344 335 1378
rect 277 1310 289 1344
rect 323 1310 335 1344
rect 277 1276 335 1310
rect 277 1242 289 1276
rect 323 1242 335 1276
rect 277 1208 335 1242
rect 277 1174 289 1208
rect 323 1174 335 1208
rect 277 1139 335 1174
rect 277 1105 289 1139
rect 323 1105 335 1139
rect 277 1050 335 1105
rect 365 1412 423 1450
rect 365 1378 377 1412
rect 411 1378 423 1412
rect 365 1344 423 1378
rect 365 1310 377 1344
rect 411 1310 423 1344
rect 365 1276 423 1310
rect 365 1242 377 1276
rect 411 1242 423 1276
rect 365 1208 423 1242
rect 365 1174 377 1208
rect 411 1174 423 1208
rect 365 1050 423 1174
rect 453 1412 511 1450
rect 453 1378 465 1412
rect 499 1378 511 1412
rect 453 1344 511 1378
rect 453 1310 465 1344
rect 499 1310 511 1344
rect 453 1276 511 1310
rect 453 1242 465 1276
rect 499 1242 511 1276
rect 453 1208 511 1242
rect 453 1174 465 1208
rect 499 1174 511 1208
rect 453 1139 511 1174
rect 453 1105 465 1139
rect 499 1105 511 1139
rect 453 1050 511 1105
rect 541 1412 599 1450
rect 541 1378 553 1412
rect 587 1378 599 1412
rect 541 1344 599 1378
rect 541 1310 553 1344
rect 587 1310 599 1344
rect 541 1276 599 1310
rect 541 1242 553 1276
rect 587 1242 599 1276
rect 541 1208 599 1242
rect 541 1174 553 1208
rect 587 1174 599 1208
rect 541 1050 599 1174
rect 629 1412 687 1450
rect 629 1378 641 1412
rect 675 1378 687 1412
rect 629 1344 687 1378
rect 629 1310 641 1344
rect 675 1310 687 1344
rect 629 1276 687 1310
rect 629 1242 641 1276
rect 675 1242 687 1276
rect 629 1208 687 1242
rect 629 1174 641 1208
rect 675 1174 687 1208
rect 629 1139 687 1174
rect 629 1105 641 1139
rect 675 1105 687 1139
rect 629 1050 687 1105
rect 717 1412 771 1450
rect 717 1378 729 1412
rect 763 1378 771 1412
rect 717 1344 771 1378
rect 717 1310 729 1344
rect 763 1310 771 1344
rect 717 1276 771 1310
rect 717 1242 729 1276
rect 763 1242 771 1276
rect 717 1208 771 1242
rect 717 1174 729 1208
rect 763 1174 771 1208
rect 717 1050 771 1174
rect 1093 1412 1149 1450
rect 1093 1378 1103 1412
rect 1137 1378 1149 1412
rect 1093 1344 1149 1378
rect 1093 1310 1103 1344
rect 1137 1310 1149 1344
rect 1093 1276 1149 1310
rect 1093 1242 1103 1276
rect 1137 1242 1149 1276
rect 1093 1208 1149 1242
rect 1093 1174 1103 1208
rect 1137 1174 1149 1208
rect 1093 1139 1149 1174
rect 1093 1105 1103 1139
rect 1137 1105 1149 1139
rect 1093 1050 1149 1105
rect 1179 1412 1237 1450
rect 1179 1378 1191 1412
rect 1225 1378 1237 1412
rect 1179 1344 1237 1378
rect 1179 1310 1191 1344
rect 1225 1310 1237 1344
rect 1179 1276 1237 1310
rect 1179 1242 1191 1276
rect 1225 1242 1237 1276
rect 1179 1208 1237 1242
rect 1179 1174 1191 1208
rect 1225 1174 1237 1208
rect 1179 1139 1237 1174
rect 1179 1105 1191 1139
rect 1225 1105 1237 1139
rect 1179 1050 1237 1105
rect 1267 1412 1325 1450
rect 1267 1378 1279 1412
rect 1313 1378 1325 1412
rect 1267 1344 1325 1378
rect 1267 1310 1279 1344
rect 1313 1310 1325 1344
rect 1267 1276 1325 1310
rect 1267 1242 1279 1276
rect 1313 1242 1325 1276
rect 1267 1208 1325 1242
rect 1267 1174 1279 1208
rect 1313 1174 1325 1208
rect 1267 1050 1325 1174
rect 1355 1412 1413 1450
rect 1355 1378 1367 1412
rect 1401 1378 1413 1412
rect 1355 1344 1413 1378
rect 1355 1310 1367 1344
rect 1401 1310 1413 1344
rect 1355 1276 1413 1310
rect 1355 1242 1367 1276
rect 1401 1242 1413 1276
rect 1355 1208 1413 1242
rect 1355 1174 1367 1208
rect 1401 1174 1413 1208
rect 1355 1139 1413 1174
rect 1355 1105 1367 1139
rect 1401 1105 1413 1139
rect 1355 1050 1413 1105
rect 1443 1412 1497 1450
rect 1443 1378 1455 1412
rect 1489 1378 1497 1412
rect 1443 1344 1497 1378
rect 1443 1310 1455 1344
rect 1489 1310 1497 1344
rect 1443 1276 1497 1310
rect 1443 1242 1455 1276
rect 1489 1242 1497 1276
rect 1443 1208 1497 1242
rect 1443 1174 1455 1208
rect 1489 1174 1497 1208
rect 1443 1050 1497 1174
rect 1759 1412 1815 1450
rect 1759 1378 1769 1412
rect 1803 1378 1815 1412
rect 1759 1344 1815 1378
rect 1759 1310 1769 1344
rect 1803 1310 1815 1344
rect 1759 1276 1815 1310
rect 1759 1242 1769 1276
rect 1803 1242 1815 1276
rect 1759 1208 1815 1242
rect 1759 1174 1769 1208
rect 1803 1174 1815 1208
rect 1759 1139 1815 1174
rect 1759 1105 1769 1139
rect 1803 1105 1815 1139
rect 1759 1050 1815 1105
rect 1845 1412 1903 1450
rect 1845 1378 1857 1412
rect 1891 1378 1903 1412
rect 1845 1344 1903 1378
rect 1845 1310 1857 1344
rect 1891 1310 1903 1344
rect 1845 1276 1903 1310
rect 1845 1242 1857 1276
rect 1891 1242 1903 1276
rect 1845 1208 1903 1242
rect 1845 1174 1857 1208
rect 1891 1174 1903 1208
rect 1845 1139 1903 1174
rect 1845 1105 1857 1139
rect 1891 1105 1903 1139
rect 1845 1050 1903 1105
rect 1933 1412 1991 1450
rect 1933 1378 1945 1412
rect 1979 1378 1991 1412
rect 1933 1344 1991 1378
rect 1933 1310 1945 1344
rect 1979 1310 1991 1344
rect 1933 1276 1991 1310
rect 1933 1242 1945 1276
rect 1979 1242 1991 1276
rect 1933 1208 1991 1242
rect 1933 1174 1945 1208
rect 1979 1174 1991 1208
rect 1933 1050 1991 1174
rect 2021 1412 2079 1450
rect 2021 1378 2033 1412
rect 2067 1378 2079 1412
rect 2021 1344 2079 1378
rect 2021 1310 2033 1344
rect 2067 1310 2079 1344
rect 2021 1276 2079 1310
rect 2021 1242 2033 1276
rect 2067 1242 2079 1276
rect 2021 1208 2079 1242
rect 2021 1174 2033 1208
rect 2067 1174 2079 1208
rect 2021 1139 2079 1174
rect 2021 1105 2033 1139
rect 2067 1105 2079 1139
rect 2021 1050 2079 1105
rect 2109 1412 2163 1450
rect 2109 1378 2121 1412
rect 2155 1378 2163 1412
rect 2109 1344 2163 1378
rect 2109 1310 2121 1344
rect 2155 1310 2163 1344
rect 2109 1276 2163 1310
rect 2109 1242 2121 1276
rect 2155 1242 2163 1276
rect 2109 1208 2163 1242
rect 2109 1174 2121 1208
rect 2155 1174 2163 1208
rect 2109 1050 2163 1174
rect 2425 1412 2481 1450
rect 2425 1378 2435 1412
rect 2469 1378 2481 1412
rect 2425 1344 2481 1378
rect 2425 1310 2435 1344
rect 2469 1310 2481 1344
rect 2425 1276 2481 1310
rect 2425 1242 2435 1276
rect 2469 1242 2481 1276
rect 2425 1208 2481 1242
rect 2425 1174 2435 1208
rect 2469 1174 2481 1208
rect 2425 1139 2481 1174
rect 2425 1105 2435 1139
rect 2469 1105 2481 1139
rect 2425 1050 2481 1105
rect 2511 1412 2569 1450
rect 2511 1378 2523 1412
rect 2557 1378 2569 1412
rect 2511 1344 2569 1378
rect 2511 1310 2523 1344
rect 2557 1310 2569 1344
rect 2511 1276 2569 1310
rect 2511 1242 2523 1276
rect 2557 1242 2569 1276
rect 2511 1208 2569 1242
rect 2511 1174 2523 1208
rect 2557 1174 2569 1208
rect 2511 1139 2569 1174
rect 2511 1105 2523 1139
rect 2557 1105 2569 1139
rect 2511 1050 2569 1105
rect 2599 1412 2657 1450
rect 2599 1378 2611 1412
rect 2645 1378 2657 1412
rect 2599 1344 2657 1378
rect 2599 1310 2611 1344
rect 2645 1310 2657 1344
rect 2599 1276 2657 1310
rect 2599 1242 2611 1276
rect 2645 1242 2657 1276
rect 2599 1208 2657 1242
rect 2599 1174 2611 1208
rect 2645 1174 2657 1208
rect 2599 1050 2657 1174
rect 2687 1412 2745 1450
rect 2687 1378 2699 1412
rect 2733 1378 2745 1412
rect 2687 1344 2745 1378
rect 2687 1310 2699 1344
rect 2733 1310 2745 1344
rect 2687 1276 2745 1310
rect 2687 1242 2699 1276
rect 2733 1242 2745 1276
rect 2687 1208 2745 1242
rect 2687 1174 2699 1208
rect 2733 1174 2745 1208
rect 2687 1139 2745 1174
rect 2687 1105 2699 1139
rect 2733 1105 2745 1139
rect 2687 1050 2745 1105
rect 2775 1412 2829 1450
rect 2775 1378 2787 1412
rect 2821 1378 2829 1412
rect 2775 1344 2829 1378
rect 2775 1310 2787 1344
rect 2821 1310 2829 1344
rect 2775 1276 2829 1310
rect 2775 1242 2787 1276
rect 2821 1242 2829 1276
rect 2775 1208 2829 1242
rect 2775 1174 2787 1208
rect 2821 1174 2829 1208
rect 2775 1050 2829 1174
rect 3091 1412 3147 1450
rect 3091 1378 3101 1412
rect 3135 1378 3147 1412
rect 3091 1344 3147 1378
rect 3091 1310 3101 1344
rect 3135 1310 3147 1344
rect 3091 1276 3147 1310
rect 3091 1242 3101 1276
rect 3135 1242 3147 1276
rect 3091 1208 3147 1242
rect 3091 1174 3101 1208
rect 3135 1174 3147 1208
rect 3091 1139 3147 1174
rect 3091 1105 3101 1139
rect 3135 1105 3147 1139
rect 3091 1050 3147 1105
rect 3177 1412 3235 1450
rect 3177 1378 3189 1412
rect 3223 1378 3235 1412
rect 3177 1344 3235 1378
rect 3177 1310 3189 1344
rect 3223 1310 3235 1344
rect 3177 1276 3235 1310
rect 3177 1242 3189 1276
rect 3223 1242 3235 1276
rect 3177 1208 3235 1242
rect 3177 1174 3189 1208
rect 3223 1174 3235 1208
rect 3177 1139 3235 1174
rect 3177 1105 3189 1139
rect 3223 1105 3235 1139
rect 3177 1050 3235 1105
rect 3265 1412 3323 1450
rect 3265 1378 3277 1412
rect 3311 1378 3323 1412
rect 3265 1344 3323 1378
rect 3265 1310 3277 1344
rect 3311 1310 3323 1344
rect 3265 1276 3323 1310
rect 3265 1242 3277 1276
rect 3311 1242 3323 1276
rect 3265 1208 3323 1242
rect 3265 1174 3277 1208
rect 3311 1174 3323 1208
rect 3265 1050 3323 1174
rect 3353 1412 3411 1450
rect 3353 1378 3365 1412
rect 3399 1378 3411 1412
rect 3353 1344 3411 1378
rect 3353 1310 3365 1344
rect 3399 1310 3411 1344
rect 3353 1276 3411 1310
rect 3353 1242 3365 1276
rect 3399 1242 3411 1276
rect 3353 1208 3411 1242
rect 3353 1174 3365 1208
rect 3399 1174 3411 1208
rect 3353 1139 3411 1174
rect 3353 1105 3365 1139
rect 3399 1105 3411 1139
rect 3353 1050 3411 1105
rect 3441 1412 3495 1450
rect 3441 1378 3453 1412
rect 3487 1378 3495 1412
rect 3441 1344 3495 1378
rect 3441 1310 3453 1344
rect 3487 1310 3495 1344
rect 3441 1276 3495 1310
rect 3441 1242 3453 1276
rect 3487 1242 3495 1276
rect 3441 1208 3495 1242
rect 3441 1174 3453 1208
rect 3487 1174 3495 1208
rect 3441 1050 3495 1174
rect 3757 1412 3813 1450
rect 3757 1378 3767 1412
rect 3801 1378 3813 1412
rect 3757 1344 3813 1378
rect 3757 1310 3767 1344
rect 3801 1310 3813 1344
rect 3757 1276 3813 1310
rect 3757 1242 3767 1276
rect 3801 1242 3813 1276
rect 3757 1208 3813 1242
rect 3757 1174 3767 1208
rect 3801 1174 3813 1208
rect 3757 1139 3813 1174
rect 3757 1105 3767 1139
rect 3801 1105 3813 1139
rect 3757 1050 3813 1105
rect 3843 1412 3901 1450
rect 3843 1378 3855 1412
rect 3889 1378 3901 1412
rect 3843 1344 3901 1378
rect 3843 1310 3855 1344
rect 3889 1310 3901 1344
rect 3843 1276 3901 1310
rect 3843 1242 3855 1276
rect 3889 1242 3901 1276
rect 3843 1208 3901 1242
rect 3843 1174 3855 1208
rect 3889 1174 3901 1208
rect 3843 1139 3901 1174
rect 3843 1105 3855 1139
rect 3889 1105 3901 1139
rect 3843 1050 3901 1105
rect 3931 1412 3989 1450
rect 3931 1378 3943 1412
rect 3977 1378 3989 1412
rect 3931 1344 3989 1378
rect 3931 1310 3943 1344
rect 3977 1310 3989 1344
rect 3931 1276 3989 1310
rect 3931 1242 3943 1276
rect 3977 1242 3989 1276
rect 3931 1208 3989 1242
rect 3931 1174 3943 1208
rect 3977 1174 3989 1208
rect 3931 1050 3989 1174
rect 4019 1412 4077 1450
rect 4019 1378 4031 1412
rect 4065 1378 4077 1412
rect 4019 1344 4077 1378
rect 4019 1310 4031 1344
rect 4065 1310 4077 1344
rect 4019 1276 4077 1310
rect 4019 1242 4031 1276
rect 4065 1242 4077 1276
rect 4019 1208 4077 1242
rect 4019 1174 4031 1208
rect 4065 1174 4077 1208
rect 4019 1139 4077 1174
rect 4019 1105 4031 1139
rect 4065 1105 4077 1139
rect 4019 1050 4077 1105
rect 4107 1412 4161 1450
rect 4107 1378 4119 1412
rect 4153 1378 4161 1412
rect 4107 1344 4161 1378
rect 4107 1310 4119 1344
rect 4153 1310 4161 1344
rect 4107 1276 4161 1310
rect 4107 1242 4119 1276
rect 4153 1242 4161 1276
rect 4107 1208 4161 1242
rect 4107 1174 4119 1208
rect 4153 1174 4161 1208
rect 4107 1050 4161 1174
rect 4483 1412 4539 1450
rect 4483 1378 4493 1412
rect 4527 1378 4539 1412
rect 4483 1344 4539 1378
rect 4483 1310 4493 1344
rect 4527 1310 4539 1344
rect 4483 1276 4539 1310
rect 4483 1242 4493 1276
rect 4527 1242 4539 1276
rect 4483 1208 4539 1242
rect 4483 1174 4493 1208
rect 4527 1174 4539 1208
rect 4483 1139 4539 1174
rect 4483 1105 4493 1139
rect 4527 1105 4539 1139
rect 4483 1050 4539 1105
rect 4569 1412 4627 1450
rect 4569 1378 4581 1412
rect 4615 1378 4627 1412
rect 4569 1344 4627 1378
rect 4569 1310 4581 1344
rect 4615 1310 4627 1344
rect 4569 1276 4627 1310
rect 4569 1242 4581 1276
rect 4615 1242 4627 1276
rect 4569 1208 4627 1242
rect 4569 1174 4581 1208
rect 4615 1174 4627 1208
rect 4569 1139 4627 1174
rect 4569 1105 4581 1139
rect 4615 1105 4627 1139
rect 4569 1050 4627 1105
rect 4657 1412 4715 1450
rect 4657 1378 4669 1412
rect 4703 1378 4715 1412
rect 4657 1344 4715 1378
rect 4657 1310 4669 1344
rect 4703 1310 4715 1344
rect 4657 1276 4715 1310
rect 4657 1242 4669 1276
rect 4703 1242 4715 1276
rect 4657 1208 4715 1242
rect 4657 1174 4669 1208
rect 4703 1174 4715 1208
rect 4657 1050 4715 1174
rect 4745 1412 4803 1450
rect 4745 1378 4757 1412
rect 4791 1378 4803 1412
rect 4745 1344 4803 1378
rect 4745 1310 4757 1344
rect 4791 1310 4803 1344
rect 4745 1276 4803 1310
rect 4745 1242 4757 1276
rect 4791 1242 4803 1276
rect 4745 1208 4803 1242
rect 4745 1174 4757 1208
rect 4791 1174 4803 1208
rect 4745 1139 4803 1174
rect 4745 1105 4757 1139
rect 4791 1105 4803 1139
rect 4745 1050 4803 1105
rect 4833 1412 4891 1450
rect 4833 1378 4845 1412
rect 4879 1378 4891 1412
rect 4833 1344 4891 1378
rect 4833 1310 4845 1344
rect 4879 1310 4891 1344
rect 4833 1276 4891 1310
rect 4833 1242 4845 1276
rect 4879 1242 4891 1276
rect 4833 1208 4891 1242
rect 4833 1174 4845 1208
rect 4879 1174 4891 1208
rect 4833 1050 4891 1174
rect 4921 1412 4979 1450
rect 4921 1378 4933 1412
rect 4967 1378 4979 1412
rect 4921 1344 4979 1378
rect 4921 1310 4933 1344
rect 4967 1310 4979 1344
rect 4921 1276 4979 1310
rect 4921 1242 4933 1276
rect 4967 1242 4979 1276
rect 4921 1208 4979 1242
rect 4921 1174 4933 1208
rect 4967 1174 4979 1208
rect 4921 1139 4979 1174
rect 4921 1105 4933 1139
rect 4967 1105 4979 1139
rect 4921 1050 4979 1105
rect 5009 1412 5063 1450
rect 5009 1378 5021 1412
rect 5055 1378 5063 1412
rect 5009 1344 5063 1378
rect 5009 1310 5021 1344
rect 5055 1310 5063 1344
rect 5009 1276 5063 1310
rect 5009 1242 5021 1276
rect 5055 1242 5063 1276
rect 5009 1208 5063 1242
rect 5009 1174 5021 1208
rect 5055 1174 5063 1208
rect 5009 1050 5063 1174
rect 5385 1412 5441 1450
rect 5385 1378 5395 1412
rect 5429 1378 5441 1412
rect 5385 1344 5441 1378
rect 5385 1310 5395 1344
rect 5429 1310 5441 1344
rect 5385 1276 5441 1310
rect 5385 1242 5395 1276
rect 5429 1242 5441 1276
rect 5385 1208 5441 1242
rect 5385 1174 5395 1208
rect 5429 1174 5441 1208
rect 5385 1139 5441 1174
rect 5385 1105 5395 1139
rect 5429 1105 5441 1139
rect 5385 1050 5441 1105
rect 5471 1412 5529 1450
rect 5471 1378 5483 1412
rect 5517 1378 5529 1412
rect 5471 1344 5529 1378
rect 5471 1310 5483 1344
rect 5517 1310 5529 1344
rect 5471 1276 5529 1310
rect 5471 1242 5483 1276
rect 5517 1242 5529 1276
rect 5471 1208 5529 1242
rect 5471 1174 5483 1208
rect 5517 1174 5529 1208
rect 5471 1139 5529 1174
rect 5471 1105 5483 1139
rect 5517 1105 5529 1139
rect 5471 1050 5529 1105
rect 5559 1412 5617 1450
rect 5559 1378 5571 1412
rect 5605 1378 5617 1412
rect 5559 1344 5617 1378
rect 5559 1310 5571 1344
rect 5605 1310 5617 1344
rect 5559 1276 5617 1310
rect 5559 1242 5571 1276
rect 5605 1242 5617 1276
rect 5559 1208 5617 1242
rect 5559 1174 5571 1208
rect 5605 1174 5617 1208
rect 5559 1050 5617 1174
rect 5647 1412 5705 1450
rect 5647 1378 5659 1412
rect 5693 1378 5705 1412
rect 5647 1344 5705 1378
rect 5647 1310 5659 1344
rect 5693 1310 5705 1344
rect 5647 1276 5705 1310
rect 5647 1242 5659 1276
rect 5693 1242 5705 1276
rect 5647 1208 5705 1242
rect 5647 1174 5659 1208
rect 5693 1174 5705 1208
rect 5647 1139 5705 1174
rect 5647 1105 5659 1139
rect 5693 1105 5705 1139
rect 5647 1050 5705 1105
rect 5735 1412 5789 1450
rect 5735 1378 5747 1412
rect 5781 1378 5789 1412
rect 5735 1344 5789 1378
rect 5735 1310 5747 1344
rect 5781 1310 5789 1344
rect 5735 1276 5789 1310
rect 5735 1242 5747 1276
rect 5781 1242 5789 1276
rect 5735 1208 5789 1242
rect 5735 1174 5747 1208
rect 5781 1174 5789 1208
rect 5735 1050 5789 1174
rect 6051 1412 6107 1450
rect 6051 1378 6061 1412
rect 6095 1378 6107 1412
rect 6051 1344 6107 1378
rect 6051 1310 6061 1344
rect 6095 1310 6107 1344
rect 6051 1276 6107 1310
rect 6051 1242 6061 1276
rect 6095 1242 6107 1276
rect 6051 1208 6107 1242
rect 6051 1174 6061 1208
rect 6095 1174 6107 1208
rect 6051 1139 6107 1174
rect 6051 1105 6061 1139
rect 6095 1105 6107 1139
rect 6051 1050 6107 1105
rect 6137 1412 6195 1450
rect 6137 1378 6149 1412
rect 6183 1378 6195 1412
rect 6137 1344 6195 1378
rect 6137 1310 6149 1344
rect 6183 1310 6195 1344
rect 6137 1276 6195 1310
rect 6137 1242 6149 1276
rect 6183 1242 6195 1276
rect 6137 1208 6195 1242
rect 6137 1174 6149 1208
rect 6183 1174 6195 1208
rect 6137 1139 6195 1174
rect 6137 1105 6149 1139
rect 6183 1105 6195 1139
rect 6137 1050 6195 1105
rect 6225 1412 6283 1450
rect 6225 1378 6237 1412
rect 6271 1378 6283 1412
rect 6225 1344 6283 1378
rect 6225 1310 6237 1344
rect 6271 1310 6283 1344
rect 6225 1276 6283 1310
rect 6225 1242 6237 1276
rect 6271 1242 6283 1276
rect 6225 1208 6283 1242
rect 6225 1174 6237 1208
rect 6271 1174 6283 1208
rect 6225 1050 6283 1174
rect 6313 1412 6371 1450
rect 6313 1378 6325 1412
rect 6359 1378 6371 1412
rect 6313 1344 6371 1378
rect 6313 1310 6325 1344
rect 6359 1310 6371 1344
rect 6313 1276 6371 1310
rect 6313 1242 6325 1276
rect 6359 1242 6371 1276
rect 6313 1208 6371 1242
rect 6313 1174 6325 1208
rect 6359 1174 6371 1208
rect 6313 1139 6371 1174
rect 6313 1105 6325 1139
rect 6359 1105 6371 1139
rect 6313 1050 6371 1105
rect 6401 1412 6455 1450
rect 6401 1378 6413 1412
rect 6447 1378 6455 1412
rect 6401 1344 6455 1378
rect 6401 1310 6413 1344
rect 6447 1310 6455 1344
rect 6401 1276 6455 1310
rect 6401 1242 6413 1276
rect 6447 1242 6455 1276
rect 6401 1208 6455 1242
rect 6401 1174 6413 1208
rect 6447 1174 6455 1208
rect 6401 1050 6455 1174
rect 6717 1412 6773 1450
rect 6717 1378 6727 1412
rect 6761 1378 6773 1412
rect 6717 1344 6773 1378
rect 6717 1310 6727 1344
rect 6761 1310 6773 1344
rect 6717 1276 6773 1310
rect 6717 1242 6727 1276
rect 6761 1242 6773 1276
rect 6717 1208 6773 1242
rect 6717 1174 6727 1208
rect 6761 1174 6773 1208
rect 6717 1139 6773 1174
rect 6717 1105 6727 1139
rect 6761 1105 6773 1139
rect 6717 1050 6773 1105
rect 6803 1412 6861 1450
rect 6803 1378 6815 1412
rect 6849 1378 6861 1412
rect 6803 1344 6861 1378
rect 6803 1310 6815 1344
rect 6849 1310 6861 1344
rect 6803 1276 6861 1310
rect 6803 1242 6815 1276
rect 6849 1242 6861 1276
rect 6803 1208 6861 1242
rect 6803 1174 6815 1208
rect 6849 1174 6861 1208
rect 6803 1139 6861 1174
rect 6803 1105 6815 1139
rect 6849 1105 6861 1139
rect 6803 1050 6861 1105
rect 6891 1412 6949 1450
rect 6891 1378 6903 1412
rect 6937 1378 6949 1412
rect 6891 1344 6949 1378
rect 6891 1310 6903 1344
rect 6937 1310 6949 1344
rect 6891 1276 6949 1310
rect 6891 1242 6903 1276
rect 6937 1242 6949 1276
rect 6891 1208 6949 1242
rect 6891 1174 6903 1208
rect 6937 1174 6949 1208
rect 6891 1050 6949 1174
rect 6979 1412 7037 1450
rect 6979 1378 6991 1412
rect 7025 1378 7037 1412
rect 6979 1344 7037 1378
rect 6979 1310 6991 1344
rect 7025 1310 7037 1344
rect 6979 1276 7037 1310
rect 6979 1242 6991 1276
rect 7025 1242 7037 1276
rect 6979 1208 7037 1242
rect 6979 1174 6991 1208
rect 7025 1174 7037 1208
rect 6979 1139 7037 1174
rect 6979 1105 6991 1139
rect 7025 1105 7037 1139
rect 6979 1050 7037 1105
rect 7067 1412 7121 1450
rect 7067 1378 7079 1412
rect 7113 1378 7121 1412
rect 7067 1344 7121 1378
rect 7067 1310 7079 1344
rect 7113 1310 7121 1344
rect 7067 1276 7121 1310
rect 7067 1242 7079 1276
rect 7113 1242 7121 1276
rect 7067 1208 7121 1242
rect 7067 1174 7079 1208
rect 7113 1174 7121 1208
rect 7067 1050 7121 1174
rect 7383 1412 7439 1450
rect 7383 1378 7393 1412
rect 7427 1378 7439 1412
rect 7383 1344 7439 1378
rect 7383 1310 7393 1344
rect 7427 1310 7439 1344
rect 7383 1276 7439 1310
rect 7383 1242 7393 1276
rect 7427 1242 7439 1276
rect 7383 1208 7439 1242
rect 7383 1174 7393 1208
rect 7427 1174 7439 1208
rect 7383 1139 7439 1174
rect 7383 1105 7393 1139
rect 7427 1105 7439 1139
rect 7383 1050 7439 1105
rect 7469 1412 7527 1450
rect 7469 1378 7481 1412
rect 7515 1378 7527 1412
rect 7469 1344 7527 1378
rect 7469 1310 7481 1344
rect 7515 1310 7527 1344
rect 7469 1276 7527 1310
rect 7469 1242 7481 1276
rect 7515 1242 7527 1276
rect 7469 1208 7527 1242
rect 7469 1174 7481 1208
rect 7515 1174 7527 1208
rect 7469 1139 7527 1174
rect 7469 1105 7481 1139
rect 7515 1105 7527 1139
rect 7469 1050 7527 1105
rect 7557 1412 7615 1450
rect 7557 1378 7569 1412
rect 7603 1378 7615 1412
rect 7557 1344 7615 1378
rect 7557 1310 7569 1344
rect 7603 1310 7615 1344
rect 7557 1276 7615 1310
rect 7557 1242 7569 1276
rect 7603 1242 7615 1276
rect 7557 1208 7615 1242
rect 7557 1174 7569 1208
rect 7603 1174 7615 1208
rect 7557 1050 7615 1174
rect 7645 1412 7703 1450
rect 7645 1378 7657 1412
rect 7691 1378 7703 1412
rect 7645 1344 7703 1378
rect 7645 1310 7657 1344
rect 7691 1310 7703 1344
rect 7645 1276 7703 1310
rect 7645 1242 7657 1276
rect 7691 1242 7703 1276
rect 7645 1208 7703 1242
rect 7645 1174 7657 1208
rect 7691 1174 7703 1208
rect 7645 1139 7703 1174
rect 7645 1105 7657 1139
rect 7691 1105 7703 1139
rect 7645 1050 7703 1105
rect 7733 1412 7787 1450
rect 7733 1378 7745 1412
rect 7779 1378 7787 1412
rect 7733 1344 7787 1378
rect 7733 1310 7745 1344
rect 7779 1310 7787 1344
rect 7733 1276 7787 1310
rect 7733 1242 7745 1276
rect 7779 1242 7787 1276
rect 7733 1208 7787 1242
rect 7733 1174 7745 1208
rect 7779 1174 7787 1208
rect 7733 1050 7787 1174
rect 8049 1412 8105 1450
rect 8049 1378 8059 1412
rect 8093 1378 8105 1412
rect 8049 1344 8105 1378
rect 8049 1310 8059 1344
rect 8093 1310 8105 1344
rect 8049 1276 8105 1310
rect 8049 1242 8059 1276
rect 8093 1242 8105 1276
rect 8049 1208 8105 1242
rect 8049 1174 8059 1208
rect 8093 1174 8105 1208
rect 8049 1139 8105 1174
rect 8049 1105 8059 1139
rect 8093 1105 8105 1139
rect 8049 1050 8105 1105
rect 8135 1412 8193 1450
rect 8135 1378 8147 1412
rect 8181 1378 8193 1412
rect 8135 1344 8193 1378
rect 8135 1310 8147 1344
rect 8181 1310 8193 1344
rect 8135 1276 8193 1310
rect 8135 1242 8147 1276
rect 8181 1242 8193 1276
rect 8135 1208 8193 1242
rect 8135 1174 8147 1208
rect 8181 1174 8193 1208
rect 8135 1139 8193 1174
rect 8135 1105 8147 1139
rect 8181 1105 8193 1139
rect 8135 1050 8193 1105
rect 8223 1412 8281 1450
rect 8223 1378 8235 1412
rect 8269 1378 8281 1412
rect 8223 1344 8281 1378
rect 8223 1310 8235 1344
rect 8269 1310 8281 1344
rect 8223 1276 8281 1310
rect 8223 1242 8235 1276
rect 8269 1242 8281 1276
rect 8223 1208 8281 1242
rect 8223 1174 8235 1208
rect 8269 1174 8281 1208
rect 8223 1050 8281 1174
rect 8311 1412 8369 1450
rect 8311 1378 8323 1412
rect 8357 1378 8369 1412
rect 8311 1344 8369 1378
rect 8311 1310 8323 1344
rect 8357 1310 8369 1344
rect 8311 1276 8369 1310
rect 8311 1242 8323 1276
rect 8357 1242 8369 1276
rect 8311 1208 8369 1242
rect 8311 1174 8323 1208
rect 8357 1174 8369 1208
rect 8311 1139 8369 1174
rect 8311 1105 8323 1139
rect 8357 1105 8369 1139
rect 8311 1050 8369 1105
rect 8399 1412 8453 1450
rect 8399 1378 8411 1412
rect 8445 1378 8453 1412
rect 8399 1344 8453 1378
rect 8399 1310 8411 1344
rect 8445 1310 8453 1344
rect 8399 1276 8453 1310
rect 8399 1242 8411 1276
rect 8445 1242 8453 1276
rect 8399 1208 8453 1242
rect 8399 1174 8411 1208
rect 8445 1174 8453 1208
rect 8399 1050 8453 1174
rect 8775 1412 8831 1450
rect 8775 1378 8785 1412
rect 8819 1378 8831 1412
rect 8775 1344 8831 1378
rect 8775 1310 8785 1344
rect 8819 1310 8831 1344
rect 8775 1276 8831 1310
rect 8775 1242 8785 1276
rect 8819 1242 8831 1276
rect 8775 1208 8831 1242
rect 8775 1174 8785 1208
rect 8819 1174 8831 1208
rect 8775 1139 8831 1174
rect 8775 1105 8785 1139
rect 8819 1105 8831 1139
rect 8775 1050 8831 1105
rect 8861 1412 8919 1450
rect 8861 1378 8873 1412
rect 8907 1378 8919 1412
rect 8861 1344 8919 1378
rect 8861 1310 8873 1344
rect 8907 1310 8919 1344
rect 8861 1276 8919 1310
rect 8861 1242 8873 1276
rect 8907 1242 8919 1276
rect 8861 1208 8919 1242
rect 8861 1174 8873 1208
rect 8907 1174 8919 1208
rect 8861 1139 8919 1174
rect 8861 1105 8873 1139
rect 8907 1105 8919 1139
rect 8861 1050 8919 1105
rect 8949 1412 9007 1450
rect 8949 1378 8961 1412
rect 8995 1378 9007 1412
rect 8949 1344 9007 1378
rect 8949 1310 8961 1344
rect 8995 1310 9007 1344
rect 8949 1276 9007 1310
rect 8949 1242 8961 1276
rect 8995 1242 9007 1276
rect 8949 1208 9007 1242
rect 8949 1174 8961 1208
rect 8995 1174 9007 1208
rect 8949 1050 9007 1174
rect 9037 1412 9095 1450
rect 9037 1378 9049 1412
rect 9083 1378 9095 1412
rect 9037 1344 9095 1378
rect 9037 1310 9049 1344
rect 9083 1310 9095 1344
rect 9037 1276 9095 1310
rect 9037 1242 9049 1276
rect 9083 1242 9095 1276
rect 9037 1208 9095 1242
rect 9037 1174 9049 1208
rect 9083 1174 9095 1208
rect 9037 1139 9095 1174
rect 9037 1105 9049 1139
rect 9083 1105 9095 1139
rect 9037 1050 9095 1105
rect 9125 1412 9183 1450
rect 9125 1378 9137 1412
rect 9171 1378 9183 1412
rect 9125 1344 9183 1378
rect 9125 1310 9137 1344
rect 9171 1310 9183 1344
rect 9125 1276 9183 1310
rect 9125 1242 9137 1276
rect 9171 1242 9183 1276
rect 9125 1208 9183 1242
rect 9125 1174 9137 1208
rect 9171 1174 9183 1208
rect 9125 1050 9183 1174
rect 9213 1412 9271 1450
rect 9213 1378 9225 1412
rect 9259 1378 9271 1412
rect 9213 1344 9271 1378
rect 9213 1310 9225 1344
rect 9259 1310 9271 1344
rect 9213 1276 9271 1310
rect 9213 1242 9225 1276
rect 9259 1242 9271 1276
rect 9213 1208 9271 1242
rect 9213 1174 9225 1208
rect 9259 1174 9271 1208
rect 9213 1139 9271 1174
rect 9213 1105 9225 1139
rect 9259 1105 9271 1139
rect 9213 1050 9271 1105
rect 9301 1412 9355 1450
rect 9301 1378 9313 1412
rect 9347 1378 9355 1412
rect 9301 1344 9355 1378
rect 9301 1310 9313 1344
rect 9347 1310 9355 1344
rect 9301 1276 9355 1310
rect 9301 1242 9313 1276
rect 9347 1242 9355 1276
rect 9301 1208 9355 1242
rect 9301 1174 9313 1208
rect 9347 1174 9355 1208
rect 9301 1050 9355 1174
rect 9677 1412 9733 1450
rect 9677 1378 9687 1412
rect 9721 1378 9733 1412
rect 9677 1344 9733 1378
rect 9677 1310 9687 1344
rect 9721 1310 9733 1344
rect 9677 1276 9733 1310
rect 9677 1242 9687 1276
rect 9721 1242 9733 1276
rect 9677 1208 9733 1242
rect 9677 1174 9687 1208
rect 9721 1174 9733 1208
rect 9677 1139 9733 1174
rect 9677 1105 9687 1139
rect 9721 1105 9733 1139
rect 9677 1050 9733 1105
rect 9763 1412 9821 1450
rect 9763 1378 9775 1412
rect 9809 1378 9821 1412
rect 9763 1344 9821 1378
rect 9763 1310 9775 1344
rect 9809 1310 9821 1344
rect 9763 1276 9821 1310
rect 9763 1242 9775 1276
rect 9809 1242 9821 1276
rect 9763 1208 9821 1242
rect 9763 1174 9775 1208
rect 9809 1174 9821 1208
rect 9763 1139 9821 1174
rect 9763 1105 9775 1139
rect 9809 1105 9821 1139
rect 9763 1050 9821 1105
rect 9851 1412 9909 1450
rect 9851 1378 9863 1412
rect 9897 1378 9909 1412
rect 9851 1344 9909 1378
rect 9851 1310 9863 1344
rect 9897 1310 9909 1344
rect 9851 1276 9909 1310
rect 9851 1242 9863 1276
rect 9897 1242 9909 1276
rect 9851 1208 9909 1242
rect 9851 1174 9863 1208
rect 9897 1174 9909 1208
rect 9851 1050 9909 1174
rect 9939 1412 9997 1450
rect 9939 1378 9951 1412
rect 9985 1378 9997 1412
rect 9939 1344 9997 1378
rect 9939 1310 9951 1344
rect 9985 1310 9997 1344
rect 9939 1276 9997 1310
rect 9939 1242 9951 1276
rect 9985 1242 9997 1276
rect 9939 1208 9997 1242
rect 9939 1174 9951 1208
rect 9985 1174 9997 1208
rect 9939 1139 9997 1174
rect 9939 1105 9951 1139
rect 9985 1105 9997 1139
rect 9939 1050 9997 1105
rect 10027 1412 10081 1450
rect 10027 1378 10039 1412
rect 10073 1378 10081 1412
rect 10027 1344 10081 1378
rect 10027 1310 10039 1344
rect 10073 1310 10081 1344
rect 10027 1276 10081 1310
rect 10027 1242 10039 1276
rect 10073 1242 10081 1276
rect 10027 1208 10081 1242
rect 10027 1174 10039 1208
rect 10073 1174 10081 1208
rect 10027 1050 10081 1174
rect 10343 1412 10399 1450
rect 10343 1378 10353 1412
rect 10387 1378 10399 1412
rect 10343 1344 10399 1378
rect 10343 1310 10353 1344
rect 10387 1310 10399 1344
rect 10343 1276 10399 1310
rect 10343 1242 10353 1276
rect 10387 1242 10399 1276
rect 10343 1208 10399 1242
rect 10343 1174 10353 1208
rect 10387 1174 10399 1208
rect 10343 1139 10399 1174
rect 10343 1105 10353 1139
rect 10387 1105 10399 1139
rect 10343 1050 10399 1105
rect 10429 1412 10487 1450
rect 10429 1378 10441 1412
rect 10475 1378 10487 1412
rect 10429 1344 10487 1378
rect 10429 1310 10441 1344
rect 10475 1310 10487 1344
rect 10429 1276 10487 1310
rect 10429 1242 10441 1276
rect 10475 1242 10487 1276
rect 10429 1208 10487 1242
rect 10429 1174 10441 1208
rect 10475 1174 10487 1208
rect 10429 1139 10487 1174
rect 10429 1105 10441 1139
rect 10475 1105 10487 1139
rect 10429 1050 10487 1105
rect 10517 1412 10575 1450
rect 10517 1378 10529 1412
rect 10563 1378 10575 1412
rect 10517 1344 10575 1378
rect 10517 1310 10529 1344
rect 10563 1310 10575 1344
rect 10517 1276 10575 1310
rect 10517 1242 10529 1276
rect 10563 1242 10575 1276
rect 10517 1208 10575 1242
rect 10517 1174 10529 1208
rect 10563 1174 10575 1208
rect 10517 1050 10575 1174
rect 10605 1412 10663 1450
rect 10605 1378 10617 1412
rect 10651 1378 10663 1412
rect 10605 1344 10663 1378
rect 10605 1310 10617 1344
rect 10651 1310 10663 1344
rect 10605 1276 10663 1310
rect 10605 1242 10617 1276
rect 10651 1242 10663 1276
rect 10605 1208 10663 1242
rect 10605 1174 10617 1208
rect 10651 1174 10663 1208
rect 10605 1139 10663 1174
rect 10605 1105 10617 1139
rect 10651 1105 10663 1139
rect 10605 1050 10663 1105
rect 10693 1412 10747 1450
rect 10693 1378 10705 1412
rect 10739 1378 10747 1412
rect 10693 1344 10747 1378
rect 10693 1310 10705 1344
rect 10739 1310 10747 1344
rect 10693 1276 10747 1310
rect 10693 1242 10705 1276
rect 10739 1242 10747 1276
rect 10693 1208 10747 1242
rect 10693 1174 10705 1208
rect 10739 1174 10747 1208
rect 10693 1050 10747 1174
rect 11009 1412 11065 1450
rect 11009 1378 11019 1412
rect 11053 1378 11065 1412
rect 11009 1344 11065 1378
rect 11009 1310 11019 1344
rect 11053 1310 11065 1344
rect 11009 1276 11065 1310
rect 11009 1242 11019 1276
rect 11053 1242 11065 1276
rect 11009 1208 11065 1242
rect 11009 1174 11019 1208
rect 11053 1174 11065 1208
rect 11009 1139 11065 1174
rect 11009 1105 11019 1139
rect 11053 1105 11065 1139
rect 11009 1050 11065 1105
rect 11095 1412 11153 1450
rect 11095 1378 11107 1412
rect 11141 1378 11153 1412
rect 11095 1344 11153 1378
rect 11095 1310 11107 1344
rect 11141 1310 11153 1344
rect 11095 1276 11153 1310
rect 11095 1242 11107 1276
rect 11141 1242 11153 1276
rect 11095 1208 11153 1242
rect 11095 1174 11107 1208
rect 11141 1174 11153 1208
rect 11095 1139 11153 1174
rect 11095 1105 11107 1139
rect 11141 1105 11153 1139
rect 11095 1050 11153 1105
rect 11183 1412 11241 1450
rect 11183 1378 11195 1412
rect 11229 1378 11241 1412
rect 11183 1344 11241 1378
rect 11183 1310 11195 1344
rect 11229 1310 11241 1344
rect 11183 1276 11241 1310
rect 11183 1242 11195 1276
rect 11229 1242 11241 1276
rect 11183 1208 11241 1242
rect 11183 1174 11195 1208
rect 11229 1174 11241 1208
rect 11183 1050 11241 1174
rect 11271 1412 11329 1450
rect 11271 1378 11283 1412
rect 11317 1378 11329 1412
rect 11271 1344 11329 1378
rect 11271 1310 11283 1344
rect 11317 1310 11329 1344
rect 11271 1276 11329 1310
rect 11271 1242 11283 1276
rect 11317 1242 11329 1276
rect 11271 1208 11329 1242
rect 11271 1174 11283 1208
rect 11317 1174 11329 1208
rect 11271 1139 11329 1174
rect 11271 1105 11283 1139
rect 11317 1105 11329 1139
rect 11271 1050 11329 1105
rect 11359 1412 11413 1450
rect 11359 1378 11371 1412
rect 11405 1378 11413 1412
rect 11359 1344 11413 1378
rect 11359 1310 11371 1344
rect 11405 1310 11413 1344
rect 11359 1276 11413 1310
rect 11359 1242 11371 1276
rect 11405 1242 11413 1276
rect 11359 1208 11413 1242
rect 11359 1174 11371 1208
rect 11405 1174 11413 1208
rect 11359 1050 11413 1174
rect 11675 1412 11731 1450
rect 11675 1378 11685 1412
rect 11719 1378 11731 1412
rect 11675 1344 11731 1378
rect 11675 1310 11685 1344
rect 11719 1310 11731 1344
rect 11675 1276 11731 1310
rect 11675 1242 11685 1276
rect 11719 1242 11731 1276
rect 11675 1208 11731 1242
rect 11675 1174 11685 1208
rect 11719 1174 11731 1208
rect 11675 1139 11731 1174
rect 11675 1105 11685 1139
rect 11719 1105 11731 1139
rect 11675 1050 11731 1105
rect 11761 1412 11819 1450
rect 11761 1378 11773 1412
rect 11807 1378 11819 1412
rect 11761 1344 11819 1378
rect 11761 1310 11773 1344
rect 11807 1310 11819 1344
rect 11761 1276 11819 1310
rect 11761 1242 11773 1276
rect 11807 1242 11819 1276
rect 11761 1208 11819 1242
rect 11761 1174 11773 1208
rect 11807 1174 11819 1208
rect 11761 1139 11819 1174
rect 11761 1105 11773 1139
rect 11807 1105 11819 1139
rect 11761 1050 11819 1105
rect 11849 1412 11907 1450
rect 11849 1378 11861 1412
rect 11895 1378 11907 1412
rect 11849 1344 11907 1378
rect 11849 1310 11861 1344
rect 11895 1310 11907 1344
rect 11849 1276 11907 1310
rect 11849 1242 11861 1276
rect 11895 1242 11907 1276
rect 11849 1208 11907 1242
rect 11849 1174 11861 1208
rect 11895 1174 11907 1208
rect 11849 1050 11907 1174
rect 11937 1412 11995 1450
rect 11937 1378 11949 1412
rect 11983 1378 11995 1412
rect 11937 1344 11995 1378
rect 11937 1310 11949 1344
rect 11983 1310 11995 1344
rect 11937 1276 11995 1310
rect 11937 1242 11949 1276
rect 11983 1242 11995 1276
rect 11937 1208 11995 1242
rect 11937 1174 11949 1208
rect 11983 1174 11995 1208
rect 11937 1139 11995 1174
rect 11937 1105 11949 1139
rect 11983 1105 11995 1139
rect 11937 1050 11995 1105
rect 12025 1412 12079 1450
rect 12025 1378 12037 1412
rect 12071 1378 12079 1412
rect 12025 1344 12079 1378
rect 12025 1310 12037 1344
rect 12071 1310 12079 1344
rect 12025 1276 12079 1310
rect 12025 1242 12037 1276
rect 12071 1242 12079 1276
rect 12025 1208 12079 1242
rect 12025 1174 12037 1208
rect 12071 1174 12079 1208
rect 12025 1050 12079 1174
rect 12341 1412 12397 1450
rect 12341 1378 12351 1412
rect 12385 1378 12397 1412
rect 12341 1344 12397 1378
rect 12341 1310 12351 1344
rect 12385 1310 12397 1344
rect 12341 1276 12397 1310
rect 12341 1242 12351 1276
rect 12385 1242 12397 1276
rect 12341 1208 12397 1242
rect 12341 1174 12351 1208
rect 12385 1174 12397 1208
rect 12341 1139 12397 1174
rect 12341 1105 12351 1139
rect 12385 1105 12397 1139
rect 12341 1050 12397 1105
rect 12427 1412 12485 1450
rect 12427 1378 12439 1412
rect 12473 1378 12485 1412
rect 12427 1344 12485 1378
rect 12427 1310 12439 1344
rect 12473 1310 12485 1344
rect 12427 1276 12485 1310
rect 12427 1242 12439 1276
rect 12473 1242 12485 1276
rect 12427 1208 12485 1242
rect 12427 1174 12439 1208
rect 12473 1174 12485 1208
rect 12427 1139 12485 1174
rect 12427 1105 12439 1139
rect 12473 1105 12485 1139
rect 12427 1050 12485 1105
rect 12515 1412 12573 1450
rect 12515 1378 12527 1412
rect 12561 1378 12573 1412
rect 12515 1344 12573 1378
rect 12515 1310 12527 1344
rect 12561 1310 12573 1344
rect 12515 1276 12573 1310
rect 12515 1242 12527 1276
rect 12561 1242 12573 1276
rect 12515 1208 12573 1242
rect 12515 1174 12527 1208
rect 12561 1174 12573 1208
rect 12515 1050 12573 1174
rect 12603 1412 12661 1450
rect 12603 1378 12615 1412
rect 12649 1378 12661 1412
rect 12603 1344 12661 1378
rect 12603 1310 12615 1344
rect 12649 1310 12661 1344
rect 12603 1276 12661 1310
rect 12603 1242 12615 1276
rect 12649 1242 12661 1276
rect 12603 1208 12661 1242
rect 12603 1174 12615 1208
rect 12649 1174 12661 1208
rect 12603 1139 12661 1174
rect 12603 1105 12615 1139
rect 12649 1105 12661 1139
rect 12603 1050 12661 1105
rect 12691 1412 12745 1450
rect 12691 1378 12703 1412
rect 12737 1378 12745 1412
rect 12691 1344 12745 1378
rect 12691 1310 12703 1344
rect 12737 1310 12745 1344
rect 12691 1276 12745 1310
rect 12691 1242 12703 1276
rect 12737 1242 12745 1276
rect 12691 1208 12745 1242
rect 12691 1174 12703 1208
rect 12737 1174 12745 1208
rect 12691 1050 12745 1174
rect 13007 1411 13063 1451
rect 13007 1377 13017 1411
rect 13051 1377 13063 1411
rect 13007 1343 13063 1377
rect 13007 1309 13017 1343
rect 13051 1309 13063 1343
rect 13007 1275 13063 1309
rect 13007 1241 13017 1275
rect 13051 1241 13063 1275
rect 13007 1207 13063 1241
rect 13007 1173 13017 1207
rect 13051 1173 13063 1207
rect 13007 1139 13063 1173
rect 13007 1105 13017 1139
rect 13051 1105 13063 1139
rect 13007 1051 13063 1105
rect 13093 1411 13151 1451
rect 13093 1377 13105 1411
rect 13139 1377 13151 1411
rect 13093 1343 13151 1377
rect 13093 1309 13105 1343
rect 13139 1309 13151 1343
rect 13093 1275 13151 1309
rect 13093 1241 13105 1275
rect 13139 1241 13151 1275
rect 13093 1207 13151 1241
rect 13093 1173 13105 1207
rect 13139 1173 13151 1207
rect 13093 1139 13151 1173
rect 13093 1105 13105 1139
rect 13139 1105 13151 1139
rect 13093 1051 13151 1105
rect 13181 1411 13239 1451
rect 13181 1377 13193 1411
rect 13227 1377 13239 1411
rect 13181 1343 13239 1377
rect 13181 1309 13193 1343
rect 13227 1309 13239 1343
rect 13181 1275 13239 1309
rect 13181 1241 13193 1275
rect 13227 1241 13239 1275
rect 13181 1207 13239 1241
rect 13181 1173 13193 1207
rect 13227 1173 13239 1207
rect 13181 1051 13239 1173
rect 13269 1411 13327 1451
rect 13269 1377 13281 1411
rect 13315 1377 13327 1411
rect 13269 1343 13327 1377
rect 13269 1309 13281 1343
rect 13315 1309 13327 1343
rect 13269 1275 13327 1309
rect 13269 1241 13281 1275
rect 13315 1241 13327 1275
rect 13269 1207 13327 1241
rect 13269 1173 13281 1207
rect 13315 1173 13327 1207
rect 13269 1051 13327 1173
rect 13357 1411 13411 1451
rect 13357 1377 13369 1411
rect 13403 1377 13411 1411
rect 13357 1343 13411 1377
rect 13357 1309 13369 1343
rect 13403 1309 13411 1343
rect 13357 1275 13411 1309
rect 13357 1241 13369 1275
rect 13403 1241 13411 1275
rect 13357 1207 13411 1241
rect 13357 1173 13369 1207
rect 13403 1173 13411 1207
rect 13357 1139 13411 1173
rect 13357 1105 13369 1139
rect 13403 1105 13411 1139
rect 13357 1051 13411 1105
rect 13673 1411 13727 1451
rect 13673 1377 13681 1411
rect 13715 1377 13727 1411
rect 13673 1343 13727 1377
rect 13673 1309 13681 1343
rect 13715 1309 13727 1343
rect 13673 1275 13727 1309
rect 13673 1241 13681 1275
rect 13715 1241 13727 1275
rect 13673 1207 13727 1241
rect 13673 1173 13681 1207
rect 13715 1173 13727 1207
rect 13673 1051 13727 1173
rect 13757 1343 13815 1451
rect 13757 1309 13769 1343
rect 13803 1309 13815 1343
rect 13757 1275 13815 1309
rect 13757 1241 13769 1275
rect 13803 1241 13815 1275
rect 13757 1207 13815 1241
rect 13757 1173 13769 1207
rect 13803 1173 13815 1207
rect 13757 1139 13815 1173
rect 13757 1105 13769 1139
rect 13803 1105 13815 1139
rect 13757 1051 13815 1105
rect 13845 1411 13903 1451
rect 13845 1377 13857 1411
rect 13891 1377 13903 1411
rect 13845 1343 13903 1377
rect 13845 1309 13857 1343
rect 13891 1309 13903 1343
rect 13845 1275 13903 1309
rect 13845 1241 13857 1275
rect 13891 1241 13903 1275
rect 13845 1207 13903 1241
rect 13845 1173 13857 1207
rect 13891 1173 13903 1207
rect 13845 1051 13903 1173
rect 13933 1343 13991 1451
rect 13933 1309 13945 1343
rect 13979 1309 13991 1343
rect 13933 1275 13991 1309
rect 13933 1241 13945 1275
rect 13979 1241 13991 1275
rect 13933 1207 13991 1241
rect 13933 1173 13945 1207
rect 13979 1173 13991 1207
rect 13933 1051 13991 1173
rect 14021 1411 14077 1451
rect 14021 1377 14033 1411
rect 14067 1377 14077 1411
rect 14021 1343 14077 1377
rect 14021 1309 14033 1343
rect 14067 1309 14077 1343
rect 14021 1275 14077 1309
rect 14021 1241 14033 1275
rect 14067 1241 14077 1275
rect 14021 1207 14077 1241
rect 14021 1173 14033 1207
rect 14067 1173 14077 1207
rect 14021 1051 14077 1173
rect 14339 1411 14395 1451
rect 14339 1377 14349 1411
rect 14383 1377 14395 1411
rect 14339 1343 14395 1377
rect 14339 1309 14349 1343
rect 14383 1309 14395 1343
rect 14339 1275 14395 1309
rect 14339 1241 14349 1275
rect 14383 1241 14395 1275
rect 14339 1207 14395 1241
rect 14339 1173 14349 1207
rect 14383 1173 14395 1207
rect 14339 1051 14395 1173
rect 14425 1343 14483 1451
rect 14425 1309 14437 1343
rect 14471 1309 14483 1343
rect 14425 1275 14483 1309
rect 14425 1241 14437 1275
rect 14471 1241 14483 1275
rect 14425 1207 14483 1241
rect 14425 1173 14437 1207
rect 14471 1173 14483 1207
rect 14425 1139 14483 1173
rect 14425 1105 14437 1139
rect 14471 1105 14483 1139
rect 14425 1051 14483 1105
rect 14513 1411 14571 1451
rect 14513 1377 14525 1411
rect 14559 1377 14571 1411
rect 14513 1343 14571 1377
rect 14513 1309 14525 1343
rect 14559 1309 14571 1343
rect 14513 1275 14571 1309
rect 14513 1241 14525 1275
rect 14559 1241 14571 1275
rect 14513 1207 14571 1241
rect 14513 1173 14525 1207
rect 14559 1173 14571 1207
rect 14513 1051 14571 1173
rect 14601 1343 14659 1451
rect 14601 1309 14613 1343
rect 14647 1309 14659 1343
rect 14601 1275 14659 1309
rect 14601 1241 14613 1275
rect 14647 1241 14659 1275
rect 14601 1207 14659 1241
rect 14601 1173 14613 1207
rect 14647 1173 14659 1207
rect 14601 1139 14659 1173
rect 14601 1105 14613 1139
rect 14647 1105 14659 1139
rect 14601 1051 14659 1105
rect 14689 1411 14743 1451
rect 14689 1377 14701 1411
rect 14735 1377 14743 1411
rect 14689 1343 14743 1377
rect 14689 1309 14701 1343
rect 14735 1309 14743 1343
rect 14689 1275 14743 1309
rect 14689 1241 14701 1275
rect 14735 1241 14743 1275
rect 14689 1207 14743 1241
rect 14689 1173 14701 1207
rect 14735 1173 14743 1207
rect 14689 1051 14743 1173
<< ndiffc >>
rect 101 329 135 363
rect 198 329 232 363
rect 295 329 329 363
rect 392 329 426 363
rect 489 329 523 363
rect 101 257 135 291
rect 101 189 135 223
rect 198 204 232 238
rect 295 257 329 291
rect 295 189 329 223
rect 393 210 427 244
rect 101 119 135 153
rect 295 119 329 153
rect 392 119 426 153
rect 489 119 523 153
rect 603 329 637 363
rect 603 257 637 291
rect 603 189 637 223
rect 700 213 734 247
rect 797 257 831 291
rect 797 189 831 223
rect 603 119 637 153
rect 700 119 734 153
rect 797 119 831 153
rect 1084 327 1118 361
rect 1181 327 1215 361
rect 1278 327 1312 361
rect 1084 255 1118 289
rect 1084 187 1118 221
rect 1181 202 1215 236
rect 1278 255 1312 289
rect 1278 187 1312 221
rect 1375 211 1409 245
rect 1472 255 1506 289
rect 1472 187 1506 221
rect 1084 117 1118 151
rect 1278 117 1312 151
rect 1375 117 1409 151
rect 1472 117 1506 151
rect 1750 327 1784 361
rect 1847 327 1881 361
rect 1944 327 1978 361
rect 1750 255 1784 289
rect 1750 187 1784 221
rect 1847 202 1881 236
rect 1944 255 1978 289
rect 1944 187 1978 221
rect 2041 211 2075 245
rect 2138 255 2172 289
rect 2138 187 2172 221
rect 1750 117 1784 151
rect 1944 117 1978 151
rect 2041 117 2075 151
rect 2138 117 2172 151
rect 2416 327 2450 361
rect 2513 327 2547 361
rect 2610 327 2644 361
rect 2416 255 2450 289
rect 2416 187 2450 221
rect 2513 202 2547 236
rect 2610 255 2644 289
rect 2610 187 2644 221
rect 2707 211 2741 245
rect 2804 255 2838 289
rect 2804 187 2838 221
rect 2416 117 2450 151
rect 2610 117 2644 151
rect 2707 117 2741 151
rect 2804 117 2838 151
rect 3082 327 3116 361
rect 3179 327 3213 361
rect 3276 327 3310 361
rect 3082 255 3116 289
rect 3082 187 3116 221
rect 3179 202 3213 236
rect 3276 255 3310 289
rect 3276 187 3310 221
rect 3373 211 3407 245
rect 3470 255 3504 289
rect 3470 187 3504 221
rect 3082 117 3116 151
rect 3276 117 3310 151
rect 3373 117 3407 151
rect 3470 117 3504 151
rect 3748 327 3782 361
rect 3845 327 3879 361
rect 3942 327 3976 361
rect 3748 255 3782 289
rect 3748 187 3782 221
rect 3845 202 3879 236
rect 3942 255 3976 289
rect 3942 187 3976 221
rect 4039 211 4073 245
rect 4136 255 4170 289
rect 4136 187 4170 221
rect 3748 117 3782 151
rect 3942 117 3976 151
rect 4039 117 4073 151
rect 4136 117 4170 151
rect 4393 329 4427 363
rect 4490 329 4524 363
rect 4587 329 4621 363
rect 4684 329 4718 363
rect 4781 329 4815 363
rect 4393 257 4427 291
rect 4393 189 4427 223
rect 4490 204 4524 238
rect 4587 257 4621 291
rect 4587 189 4621 223
rect 4685 210 4719 244
rect 4393 119 4427 153
rect 4587 119 4621 153
rect 4684 119 4718 153
rect 4781 119 4815 153
rect 4895 329 4929 363
rect 4895 257 4929 291
rect 4895 189 4929 223
rect 4992 213 5026 247
rect 5089 257 5123 291
rect 5089 189 5123 223
rect 4895 119 4929 153
rect 4992 119 5026 153
rect 5089 119 5123 153
rect 5376 327 5410 361
rect 5473 327 5507 361
rect 5570 327 5604 361
rect 5376 255 5410 289
rect 5376 187 5410 221
rect 5473 202 5507 236
rect 5570 255 5604 289
rect 5570 187 5604 221
rect 5667 211 5701 245
rect 5764 255 5798 289
rect 5764 187 5798 221
rect 5376 117 5410 151
rect 5570 117 5604 151
rect 5667 117 5701 151
rect 5764 117 5798 151
rect 6042 327 6076 361
rect 6139 327 6173 361
rect 6236 327 6270 361
rect 6042 255 6076 289
rect 6042 187 6076 221
rect 6139 202 6173 236
rect 6236 255 6270 289
rect 6236 187 6270 221
rect 6333 211 6367 245
rect 6430 255 6464 289
rect 6430 187 6464 221
rect 6042 117 6076 151
rect 6236 117 6270 151
rect 6333 117 6367 151
rect 6430 117 6464 151
rect 6708 327 6742 361
rect 6805 327 6839 361
rect 6902 327 6936 361
rect 6708 255 6742 289
rect 6708 187 6742 221
rect 6805 202 6839 236
rect 6902 255 6936 289
rect 6902 187 6936 221
rect 6999 211 7033 245
rect 7096 255 7130 289
rect 7096 187 7130 221
rect 6708 117 6742 151
rect 6902 117 6936 151
rect 6999 117 7033 151
rect 7096 117 7130 151
rect 7374 327 7408 361
rect 7471 327 7505 361
rect 7568 327 7602 361
rect 7374 255 7408 289
rect 7374 187 7408 221
rect 7471 202 7505 236
rect 7568 255 7602 289
rect 7568 187 7602 221
rect 7665 211 7699 245
rect 7762 255 7796 289
rect 7762 187 7796 221
rect 7374 117 7408 151
rect 7568 117 7602 151
rect 7665 117 7699 151
rect 7762 117 7796 151
rect 8040 327 8074 361
rect 8137 327 8171 361
rect 8234 327 8268 361
rect 8040 255 8074 289
rect 8040 187 8074 221
rect 8137 202 8171 236
rect 8234 255 8268 289
rect 8234 187 8268 221
rect 8331 211 8365 245
rect 8428 255 8462 289
rect 8428 187 8462 221
rect 8040 117 8074 151
rect 8234 117 8268 151
rect 8331 117 8365 151
rect 8428 117 8462 151
rect 8685 329 8719 363
rect 8782 329 8816 363
rect 8879 329 8913 363
rect 8976 329 9010 363
rect 9073 329 9107 363
rect 8685 257 8719 291
rect 8685 189 8719 223
rect 8782 204 8816 238
rect 8879 257 8913 291
rect 8879 189 8913 223
rect 8977 210 9011 244
rect 8685 119 8719 153
rect 8879 119 8913 153
rect 8976 119 9010 153
rect 9073 119 9107 153
rect 9187 329 9221 363
rect 9187 257 9221 291
rect 9187 189 9221 223
rect 9284 213 9318 247
rect 9381 257 9415 291
rect 9381 189 9415 223
rect 9187 119 9221 153
rect 9284 119 9318 153
rect 9381 119 9415 153
rect 9668 327 9702 361
rect 9765 327 9799 361
rect 9862 327 9896 361
rect 9668 255 9702 289
rect 9668 187 9702 221
rect 9765 202 9799 236
rect 9862 255 9896 289
rect 9862 187 9896 221
rect 9959 211 9993 245
rect 10056 255 10090 289
rect 10056 187 10090 221
rect 9668 117 9702 151
rect 9862 117 9896 151
rect 9959 117 9993 151
rect 10056 117 10090 151
rect 10334 327 10368 361
rect 10431 327 10465 361
rect 10528 327 10562 361
rect 10334 255 10368 289
rect 10334 187 10368 221
rect 10431 202 10465 236
rect 10528 255 10562 289
rect 10528 187 10562 221
rect 10625 211 10659 245
rect 10722 255 10756 289
rect 10722 187 10756 221
rect 10334 117 10368 151
rect 10528 117 10562 151
rect 10625 117 10659 151
rect 10722 117 10756 151
rect 11000 327 11034 361
rect 11097 327 11131 361
rect 11194 327 11228 361
rect 11000 255 11034 289
rect 11000 187 11034 221
rect 11097 202 11131 236
rect 11194 255 11228 289
rect 11194 187 11228 221
rect 11291 211 11325 245
rect 11388 255 11422 289
rect 11388 187 11422 221
rect 11000 117 11034 151
rect 11194 117 11228 151
rect 11291 117 11325 151
rect 11388 117 11422 151
rect 11666 327 11700 361
rect 11763 327 11797 361
rect 11860 327 11894 361
rect 11666 255 11700 289
rect 11666 187 11700 221
rect 11763 202 11797 236
rect 11860 255 11894 289
rect 11860 187 11894 221
rect 11957 211 11991 245
rect 12054 255 12088 289
rect 12054 187 12088 221
rect 11666 117 11700 151
rect 11860 117 11894 151
rect 11957 117 11991 151
rect 12054 117 12088 151
rect 12332 327 12366 361
rect 12429 327 12463 361
rect 12526 327 12560 361
rect 12332 255 12366 289
rect 12332 187 12366 221
rect 12429 202 12463 236
rect 12526 255 12560 289
rect 12526 187 12560 221
rect 12623 211 12657 245
rect 12720 255 12754 289
rect 12720 187 12754 221
rect 12332 117 12366 151
rect 12526 117 12560 151
rect 12623 117 12657 151
rect 12720 117 12754 151
rect 12998 327 13032 361
rect 13095 327 13129 361
rect 13192 327 13226 361
rect 13386 327 13420 361
rect 12998 255 13032 289
rect 12998 187 13032 221
rect 13095 202 13129 236
rect 13192 255 13226 289
rect 13192 187 13226 221
rect 13288 211 13322 245
rect 13386 255 13420 289
rect 13386 187 13420 221
rect 12998 117 13032 151
rect 13192 117 13226 151
rect 13288 117 13322 151
rect 13386 117 13420 151
rect 13664 327 13698 361
rect 13761 327 13795 361
rect 13858 327 13892 361
rect 14052 327 14086 361
rect 13664 255 13698 289
rect 13664 187 13698 221
rect 13761 202 13795 236
rect 13858 255 13892 289
rect 13858 187 13892 221
rect 13955 211 13989 245
rect 14052 255 14086 289
rect 14052 187 14086 221
rect 13664 117 13698 151
rect 13858 117 13892 151
rect 13955 117 13989 151
rect 14052 117 14086 151
rect 14330 327 14364 361
rect 14427 327 14461 361
rect 14524 327 14558 361
rect 14330 255 14364 289
rect 14330 187 14364 221
rect 14427 202 14461 236
rect 14524 255 14558 289
rect 14524 187 14558 221
rect 14621 211 14655 245
rect 14718 255 14752 289
rect 14718 187 14752 221
rect 14330 117 14364 151
rect 14524 117 14558 151
rect 14621 117 14655 151
rect 14718 117 14752 151
<< pdiffc >>
rect 201 1378 235 1412
rect 201 1310 235 1344
rect 201 1242 235 1276
rect 201 1174 235 1208
rect 201 1105 235 1139
rect 289 1378 323 1412
rect 289 1310 323 1344
rect 289 1242 323 1276
rect 289 1174 323 1208
rect 289 1105 323 1139
rect 377 1378 411 1412
rect 377 1310 411 1344
rect 377 1242 411 1276
rect 377 1174 411 1208
rect 465 1378 499 1412
rect 465 1310 499 1344
rect 465 1242 499 1276
rect 465 1174 499 1208
rect 465 1105 499 1139
rect 553 1378 587 1412
rect 553 1310 587 1344
rect 553 1242 587 1276
rect 553 1174 587 1208
rect 641 1378 675 1412
rect 641 1310 675 1344
rect 641 1242 675 1276
rect 641 1174 675 1208
rect 641 1105 675 1139
rect 729 1378 763 1412
rect 729 1310 763 1344
rect 729 1242 763 1276
rect 729 1174 763 1208
rect 1103 1378 1137 1412
rect 1103 1310 1137 1344
rect 1103 1242 1137 1276
rect 1103 1174 1137 1208
rect 1103 1105 1137 1139
rect 1191 1378 1225 1412
rect 1191 1310 1225 1344
rect 1191 1242 1225 1276
rect 1191 1174 1225 1208
rect 1191 1105 1225 1139
rect 1279 1378 1313 1412
rect 1279 1310 1313 1344
rect 1279 1242 1313 1276
rect 1279 1174 1313 1208
rect 1367 1378 1401 1412
rect 1367 1310 1401 1344
rect 1367 1242 1401 1276
rect 1367 1174 1401 1208
rect 1367 1105 1401 1139
rect 1455 1378 1489 1412
rect 1455 1310 1489 1344
rect 1455 1242 1489 1276
rect 1455 1174 1489 1208
rect 1769 1378 1803 1412
rect 1769 1310 1803 1344
rect 1769 1242 1803 1276
rect 1769 1174 1803 1208
rect 1769 1105 1803 1139
rect 1857 1378 1891 1412
rect 1857 1310 1891 1344
rect 1857 1242 1891 1276
rect 1857 1174 1891 1208
rect 1857 1105 1891 1139
rect 1945 1378 1979 1412
rect 1945 1310 1979 1344
rect 1945 1242 1979 1276
rect 1945 1174 1979 1208
rect 2033 1378 2067 1412
rect 2033 1310 2067 1344
rect 2033 1242 2067 1276
rect 2033 1174 2067 1208
rect 2033 1105 2067 1139
rect 2121 1378 2155 1412
rect 2121 1310 2155 1344
rect 2121 1242 2155 1276
rect 2121 1174 2155 1208
rect 2435 1378 2469 1412
rect 2435 1310 2469 1344
rect 2435 1242 2469 1276
rect 2435 1174 2469 1208
rect 2435 1105 2469 1139
rect 2523 1378 2557 1412
rect 2523 1310 2557 1344
rect 2523 1242 2557 1276
rect 2523 1174 2557 1208
rect 2523 1105 2557 1139
rect 2611 1378 2645 1412
rect 2611 1310 2645 1344
rect 2611 1242 2645 1276
rect 2611 1174 2645 1208
rect 2699 1378 2733 1412
rect 2699 1310 2733 1344
rect 2699 1242 2733 1276
rect 2699 1174 2733 1208
rect 2699 1105 2733 1139
rect 2787 1378 2821 1412
rect 2787 1310 2821 1344
rect 2787 1242 2821 1276
rect 2787 1174 2821 1208
rect 3101 1378 3135 1412
rect 3101 1310 3135 1344
rect 3101 1242 3135 1276
rect 3101 1174 3135 1208
rect 3101 1105 3135 1139
rect 3189 1378 3223 1412
rect 3189 1310 3223 1344
rect 3189 1242 3223 1276
rect 3189 1174 3223 1208
rect 3189 1105 3223 1139
rect 3277 1378 3311 1412
rect 3277 1310 3311 1344
rect 3277 1242 3311 1276
rect 3277 1174 3311 1208
rect 3365 1378 3399 1412
rect 3365 1310 3399 1344
rect 3365 1242 3399 1276
rect 3365 1174 3399 1208
rect 3365 1105 3399 1139
rect 3453 1378 3487 1412
rect 3453 1310 3487 1344
rect 3453 1242 3487 1276
rect 3453 1174 3487 1208
rect 3767 1378 3801 1412
rect 3767 1310 3801 1344
rect 3767 1242 3801 1276
rect 3767 1174 3801 1208
rect 3767 1105 3801 1139
rect 3855 1378 3889 1412
rect 3855 1310 3889 1344
rect 3855 1242 3889 1276
rect 3855 1174 3889 1208
rect 3855 1105 3889 1139
rect 3943 1378 3977 1412
rect 3943 1310 3977 1344
rect 3943 1242 3977 1276
rect 3943 1174 3977 1208
rect 4031 1378 4065 1412
rect 4031 1310 4065 1344
rect 4031 1242 4065 1276
rect 4031 1174 4065 1208
rect 4031 1105 4065 1139
rect 4119 1378 4153 1412
rect 4119 1310 4153 1344
rect 4119 1242 4153 1276
rect 4119 1174 4153 1208
rect 4493 1378 4527 1412
rect 4493 1310 4527 1344
rect 4493 1242 4527 1276
rect 4493 1174 4527 1208
rect 4493 1105 4527 1139
rect 4581 1378 4615 1412
rect 4581 1310 4615 1344
rect 4581 1242 4615 1276
rect 4581 1174 4615 1208
rect 4581 1105 4615 1139
rect 4669 1378 4703 1412
rect 4669 1310 4703 1344
rect 4669 1242 4703 1276
rect 4669 1174 4703 1208
rect 4757 1378 4791 1412
rect 4757 1310 4791 1344
rect 4757 1242 4791 1276
rect 4757 1174 4791 1208
rect 4757 1105 4791 1139
rect 4845 1378 4879 1412
rect 4845 1310 4879 1344
rect 4845 1242 4879 1276
rect 4845 1174 4879 1208
rect 4933 1378 4967 1412
rect 4933 1310 4967 1344
rect 4933 1242 4967 1276
rect 4933 1174 4967 1208
rect 4933 1105 4967 1139
rect 5021 1378 5055 1412
rect 5021 1310 5055 1344
rect 5021 1242 5055 1276
rect 5021 1174 5055 1208
rect 5395 1378 5429 1412
rect 5395 1310 5429 1344
rect 5395 1242 5429 1276
rect 5395 1174 5429 1208
rect 5395 1105 5429 1139
rect 5483 1378 5517 1412
rect 5483 1310 5517 1344
rect 5483 1242 5517 1276
rect 5483 1174 5517 1208
rect 5483 1105 5517 1139
rect 5571 1378 5605 1412
rect 5571 1310 5605 1344
rect 5571 1242 5605 1276
rect 5571 1174 5605 1208
rect 5659 1378 5693 1412
rect 5659 1310 5693 1344
rect 5659 1242 5693 1276
rect 5659 1174 5693 1208
rect 5659 1105 5693 1139
rect 5747 1378 5781 1412
rect 5747 1310 5781 1344
rect 5747 1242 5781 1276
rect 5747 1174 5781 1208
rect 6061 1378 6095 1412
rect 6061 1310 6095 1344
rect 6061 1242 6095 1276
rect 6061 1174 6095 1208
rect 6061 1105 6095 1139
rect 6149 1378 6183 1412
rect 6149 1310 6183 1344
rect 6149 1242 6183 1276
rect 6149 1174 6183 1208
rect 6149 1105 6183 1139
rect 6237 1378 6271 1412
rect 6237 1310 6271 1344
rect 6237 1242 6271 1276
rect 6237 1174 6271 1208
rect 6325 1378 6359 1412
rect 6325 1310 6359 1344
rect 6325 1242 6359 1276
rect 6325 1174 6359 1208
rect 6325 1105 6359 1139
rect 6413 1378 6447 1412
rect 6413 1310 6447 1344
rect 6413 1242 6447 1276
rect 6413 1174 6447 1208
rect 6727 1378 6761 1412
rect 6727 1310 6761 1344
rect 6727 1242 6761 1276
rect 6727 1174 6761 1208
rect 6727 1105 6761 1139
rect 6815 1378 6849 1412
rect 6815 1310 6849 1344
rect 6815 1242 6849 1276
rect 6815 1174 6849 1208
rect 6815 1105 6849 1139
rect 6903 1378 6937 1412
rect 6903 1310 6937 1344
rect 6903 1242 6937 1276
rect 6903 1174 6937 1208
rect 6991 1378 7025 1412
rect 6991 1310 7025 1344
rect 6991 1242 7025 1276
rect 6991 1174 7025 1208
rect 6991 1105 7025 1139
rect 7079 1378 7113 1412
rect 7079 1310 7113 1344
rect 7079 1242 7113 1276
rect 7079 1174 7113 1208
rect 7393 1378 7427 1412
rect 7393 1310 7427 1344
rect 7393 1242 7427 1276
rect 7393 1174 7427 1208
rect 7393 1105 7427 1139
rect 7481 1378 7515 1412
rect 7481 1310 7515 1344
rect 7481 1242 7515 1276
rect 7481 1174 7515 1208
rect 7481 1105 7515 1139
rect 7569 1378 7603 1412
rect 7569 1310 7603 1344
rect 7569 1242 7603 1276
rect 7569 1174 7603 1208
rect 7657 1378 7691 1412
rect 7657 1310 7691 1344
rect 7657 1242 7691 1276
rect 7657 1174 7691 1208
rect 7657 1105 7691 1139
rect 7745 1378 7779 1412
rect 7745 1310 7779 1344
rect 7745 1242 7779 1276
rect 7745 1174 7779 1208
rect 8059 1378 8093 1412
rect 8059 1310 8093 1344
rect 8059 1242 8093 1276
rect 8059 1174 8093 1208
rect 8059 1105 8093 1139
rect 8147 1378 8181 1412
rect 8147 1310 8181 1344
rect 8147 1242 8181 1276
rect 8147 1174 8181 1208
rect 8147 1105 8181 1139
rect 8235 1378 8269 1412
rect 8235 1310 8269 1344
rect 8235 1242 8269 1276
rect 8235 1174 8269 1208
rect 8323 1378 8357 1412
rect 8323 1310 8357 1344
rect 8323 1242 8357 1276
rect 8323 1174 8357 1208
rect 8323 1105 8357 1139
rect 8411 1378 8445 1412
rect 8411 1310 8445 1344
rect 8411 1242 8445 1276
rect 8411 1174 8445 1208
rect 8785 1378 8819 1412
rect 8785 1310 8819 1344
rect 8785 1242 8819 1276
rect 8785 1174 8819 1208
rect 8785 1105 8819 1139
rect 8873 1378 8907 1412
rect 8873 1310 8907 1344
rect 8873 1242 8907 1276
rect 8873 1174 8907 1208
rect 8873 1105 8907 1139
rect 8961 1378 8995 1412
rect 8961 1310 8995 1344
rect 8961 1242 8995 1276
rect 8961 1174 8995 1208
rect 9049 1378 9083 1412
rect 9049 1310 9083 1344
rect 9049 1242 9083 1276
rect 9049 1174 9083 1208
rect 9049 1105 9083 1139
rect 9137 1378 9171 1412
rect 9137 1310 9171 1344
rect 9137 1242 9171 1276
rect 9137 1174 9171 1208
rect 9225 1378 9259 1412
rect 9225 1310 9259 1344
rect 9225 1242 9259 1276
rect 9225 1174 9259 1208
rect 9225 1105 9259 1139
rect 9313 1378 9347 1412
rect 9313 1310 9347 1344
rect 9313 1242 9347 1276
rect 9313 1174 9347 1208
rect 9687 1378 9721 1412
rect 9687 1310 9721 1344
rect 9687 1242 9721 1276
rect 9687 1174 9721 1208
rect 9687 1105 9721 1139
rect 9775 1378 9809 1412
rect 9775 1310 9809 1344
rect 9775 1242 9809 1276
rect 9775 1174 9809 1208
rect 9775 1105 9809 1139
rect 9863 1378 9897 1412
rect 9863 1310 9897 1344
rect 9863 1242 9897 1276
rect 9863 1174 9897 1208
rect 9951 1378 9985 1412
rect 9951 1310 9985 1344
rect 9951 1242 9985 1276
rect 9951 1174 9985 1208
rect 9951 1105 9985 1139
rect 10039 1378 10073 1412
rect 10039 1310 10073 1344
rect 10039 1242 10073 1276
rect 10039 1174 10073 1208
rect 10353 1378 10387 1412
rect 10353 1310 10387 1344
rect 10353 1242 10387 1276
rect 10353 1174 10387 1208
rect 10353 1105 10387 1139
rect 10441 1378 10475 1412
rect 10441 1310 10475 1344
rect 10441 1242 10475 1276
rect 10441 1174 10475 1208
rect 10441 1105 10475 1139
rect 10529 1378 10563 1412
rect 10529 1310 10563 1344
rect 10529 1242 10563 1276
rect 10529 1174 10563 1208
rect 10617 1378 10651 1412
rect 10617 1310 10651 1344
rect 10617 1242 10651 1276
rect 10617 1174 10651 1208
rect 10617 1105 10651 1139
rect 10705 1378 10739 1412
rect 10705 1310 10739 1344
rect 10705 1242 10739 1276
rect 10705 1174 10739 1208
rect 11019 1378 11053 1412
rect 11019 1310 11053 1344
rect 11019 1242 11053 1276
rect 11019 1174 11053 1208
rect 11019 1105 11053 1139
rect 11107 1378 11141 1412
rect 11107 1310 11141 1344
rect 11107 1242 11141 1276
rect 11107 1174 11141 1208
rect 11107 1105 11141 1139
rect 11195 1378 11229 1412
rect 11195 1310 11229 1344
rect 11195 1242 11229 1276
rect 11195 1174 11229 1208
rect 11283 1378 11317 1412
rect 11283 1310 11317 1344
rect 11283 1242 11317 1276
rect 11283 1174 11317 1208
rect 11283 1105 11317 1139
rect 11371 1378 11405 1412
rect 11371 1310 11405 1344
rect 11371 1242 11405 1276
rect 11371 1174 11405 1208
rect 11685 1378 11719 1412
rect 11685 1310 11719 1344
rect 11685 1242 11719 1276
rect 11685 1174 11719 1208
rect 11685 1105 11719 1139
rect 11773 1378 11807 1412
rect 11773 1310 11807 1344
rect 11773 1242 11807 1276
rect 11773 1174 11807 1208
rect 11773 1105 11807 1139
rect 11861 1378 11895 1412
rect 11861 1310 11895 1344
rect 11861 1242 11895 1276
rect 11861 1174 11895 1208
rect 11949 1378 11983 1412
rect 11949 1310 11983 1344
rect 11949 1242 11983 1276
rect 11949 1174 11983 1208
rect 11949 1105 11983 1139
rect 12037 1378 12071 1412
rect 12037 1310 12071 1344
rect 12037 1242 12071 1276
rect 12037 1174 12071 1208
rect 12351 1378 12385 1412
rect 12351 1310 12385 1344
rect 12351 1242 12385 1276
rect 12351 1174 12385 1208
rect 12351 1105 12385 1139
rect 12439 1378 12473 1412
rect 12439 1310 12473 1344
rect 12439 1242 12473 1276
rect 12439 1174 12473 1208
rect 12439 1105 12473 1139
rect 12527 1378 12561 1412
rect 12527 1310 12561 1344
rect 12527 1242 12561 1276
rect 12527 1174 12561 1208
rect 12615 1378 12649 1412
rect 12615 1310 12649 1344
rect 12615 1242 12649 1276
rect 12615 1174 12649 1208
rect 12615 1105 12649 1139
rect 12703 1378 12737 1412
rect 12703 1310 12737 1344
rect 12703 1242 12737 1276
rect 12703 1174 12737 1208
rect 13017 1377 13051 1411
rect 13017 1309 13051 1343
rect 13017 1241 13051 1275
rect 13017 1173 13051 1207
rect 13017 1105 13051 1139
rect 13105 1377 13139 1411
rect 13105 1309 13139 1343
rect 13105 1241 13139 1275
rect 13105 1173 13139 1207
rect 13105 1105 13139 1139
rect 13193 1377 13227 1411
rect 13193 1309 13227 1343
rect 13193 1241 13227 1275
rect 13193 1173 13227 1207
rect 13281 1377 13315 1411
rect 13281 1309 13315 1343
rect 13281 1241 13315 1275
rect 13281 1173 13315 1207
rect 13369 1377 13403 1411
rect 13369 1309 13403 1343
rect 13369 1241 13403 1275
rect 13369 1173 13403 1207
rect 13369 1105 13403 1139
rect 13681 1377 13715 1411
rect 13681 1309 13715 1343
rect 13681 1241 13715 1275
rect 13681 1173 13715 1207
rect 13769 1309 13803 1343
rect 13769 1241 13803 1275
rect 13769 1173 13803 1207
rect 13769 1105 13803 1139
rect 13857 1377 13891 1411
rect 13857 1309 13891 1343
rect 13857 1241 13891 1275
rect 13857 1173 13891 1207
rect 13945 1309 13979 1343
rect 13945 1241 13979 1275
rect 13945 1173 13979 1207
rect 14033 1377 14067 1411
rect 14033 1309 14067 1343
rect 14033 1241 14067 1275
rect 14033 1173 14067 1207
rect 14349 1377 14383 1411
rect 14349 1309 14383 1343
rect 14349 1241 14383 1275
rect 14349 1173 14383 1207
rect 14437 1309 14471 1343
rect 14437 1241 14471 1275
rect 14437 1173 14471 1207
rect 14437 1105 14471 1139
rect 14525 1377 14559 1411
rect 14525 1309 14559 1343
rect 14525 1241 14559 1275
rect 14525 1173 14559 1207
rect 14613 1309 14647 1343
rect 14613 1241 14647 1275
rect 14613 1173 14647 1207
rect 14613 1105 14647 1139
rect 14701 1377 14735 1411
rect 14701 1309 14735 1343
rect 14701 1241 14735 1275
rect 14701 1173 14735 1207
<< psubdiff >>
rect -31 546 14905 572
rect -31 512 -17 546
rect 17 512 945 546
rect 979 512 1611 546
rect 1645 512 2277 546
rect 2311 512 2943 546
rect 2977 512 3609 546
rect 3643 512 4275 546
rect 4309 512 5237 546
rect 5271 512 5903 546
rect 5937 512 6569 546
rect 6603 512 7235 546
rect 7269 512 7901 546
rect 7935 512 8567 546
rect 8601 512 9529 546
rect 9563 512 10195 546
rect 10229 512 10861 546
rect 10895 512 11527 546
rect 11561 512 12193 546
rect 12227 512 12859 546
rect 12893 512 13525 546
rect 13559 512 14191 546
rect 14225 512 14857 546
rect 14891 512 14905 546
rect -31 510 14905 512
rect -31 474 31 510
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect -31 368 -17 402
rect 17 368 31 402
rect 931 474 993 510
rect 931 440 945 474
rect 979 440 993 474
rect 931 402 993 440
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect 931 368 945 402
rect 979 368 993 402
rect 1597 474 1659 510
rect 1597 440 1611 474
rect 1645 440 1659 474
rect 1597 402 1659 440
rect 931 330 993 368
rect 931 296 945 330
rect 979 296 993 330
rect 931 258 993 296
rect 931 224 945 258
rect 979 224 993 258
rect 931 186 993 224
rect 931 152 945 186
rect 979 152 993 186
rect 931 114 993 152
rect -31 47 31 80
rect 931 80 945 114
rect 979 80 993 114
rect 1597 368 1611 402
rect 1645 368 1659 402
rect 2263 474 2325 510
rect 2263 440 2277 474
rect 2311 440 2325 474
rect 2263 402 2325 440
rect 1597 330 1659 368
rect 1597 296 1611 330
rect 1645 296 1659 330
rect 1597 258 1659 296
rect 1597 224 1611 258
rect 1645 224 1659 258
rect 1597 186 1659 224
rect 1597 152 1611 186
rect 1645 152 1659 186
rect 1597 114 1659 152
rect 931 47 993 80
rect 1597 80 1611 114
rect 1645 80 1659 114
rect 2263 368 2277 402
rect 2311 368 2325 402
rect 2929 474 2991 510
rect 2929 440 2943 474
rect 2977 440 2991 474
rect 2929 402 2991 440
rect 2263 330 2325 368
rect 2263 296 2277 330
rect 2311 296 2325 330
rect 2263 258 2325 296
rect 2263 224 2277 258
rect 2311 224 2325 258
rect 2263 186 2325 224
rect 2263 152 2277 186
rect 2311 152 2325 186
rect 2263 114 2325 152
rect 1597 47 1659 80
rect 2263 80 2277 114
rect 2311 80 2325 114
rect 2929 368 2943 402
rect 2977 368 2991 402
rect 3595 474 3657 510
rect 3595 440 3609 474
rect 3643 440 3657 474
rect 3595 402 3657 440
rect 2929 330 2991 368
rect 2929 296 2943 330
rect 2977 296 2991 330
rect 2929 258 2991 296
rect 2929 224 2943 258
rect 2977 224 2991 258
rect 2929 186 2991 224
rect 2929 152 2943 186
rect 2977 152 2991 186
rect 2929 114 2991 152
rect 2263 47 2325 80
rect 2929 80 2943 114
rect 2977 80 2991 114
rect 3595 368 3609 402
rect 3643 368 3657 402
rect 4261 474 4323 510
rect 4261 440 4275 474
rect 4309 440 4323 474
rect 4261 402 4323 440
rect 3595 330 3657 368
rect 3595 296 3609 330
rect 3643 296 3657 330
rect 3595 258 3657 296
rect 3595 224 3609 258
rect 3643 224 3657 258
rect 3595 186 3657 224
rect 3595 152 3609 186
rect 3643 152 3657 186
rect 3595 114 3657 152
rect 2929 47 2991 80
rect 3595 80 3609 114
rect 3643 80 3657 114
rect 4261 368 4275 402
rect 4309 368 4323 402
rect 5223 474 5285 510
rect 5223 440 5237 474
rect 5271 440 5285 474
rect 5223 402 5285 440
rect 4261 330 4323 368
rect 4261 296 4275 330
rect 4309 296 4323 330
rect 4261 258 4323 296
rect 4261 224 4275 258
rect 4309 224 4323 258
rect 4261 186 4323 224
rect 4261 152 4275 186
rect 4309 152 4323 186
rect 4261 114 4323 152
rect 3595 47 3657 80
rect 4261 80 4275 114
rect 4309 80 4323 114
rect 5223 368 5237 402
rect 5271 368 5285 402
rect 5889 474 5951 510
rect 5889 440 5903 474
rect 5937 440 5951 474
rect 5889 402 5951 440
rect 5223 330 5285 368
rect 5223 296 5237 330
rect 5271 296 5285 330
rect 5223 258 5285 296
rect 5223 224 5237 258
rect 5271 224 5285 258
rect 5223 186 5285 224
rect 5223 152 5237 186
rect 5271 152 5285 186
rect 5223 114 5285 152
rect 4261 47 4323 80
rect 5223 80 5237 114
rect 5271 80 5285 114
rect 5889 368 5903 402
rect 5937 368 5951 402
rect 6555 474 6617 510
rect 6555 440 6569 474
rect 6603 440 6617 474
rect 6555 402 6617 440
rect 5889 330 5951 368
rect 5889 296 5903 330
rect 5937 296 5951 330
rect 5889 258 5951 296
rect 5889 224 5903 258
rect 5937 224 5951 258
rect 5889 186 5951 224
rect 5889 152 5903 186
rect 5937 152 5951 186
rect 5889 114 5951 152
rect 5223 47 5285 80
rect 5889 80 5903 114
rect 5937 80 5951 114
rect 6555 368 6569 402
rect 6603 368 6617 402
rect 7221 474 7283 510
rect 7221 440 7235 474
rect 7269 440 7283 474
rect 7221 402 7283 440
rect 6555 330 6617 368
rect 6555 296 6569 330
rect 6603 296 6617 330
rect 6555 258 6617 296
rect 6555 224 6569 258
rect 6603 224 6617 258
rect 6555 186 6617 224
rect 6555 152 6569 186
rect 6603 152 6617 186
rect 6555 114 6617 152
rect 5889 47 5951 80
rect 6555 80 6569 114
rect 6603 80 6617 114
rect 7221 368 7235 402
rect 7269 368 7283 402
rect 7887 474 7949 510
rect 7887 440 7901 474
rect 7935 440 7949 474
rect 7887 402 7949 440
rect 7221 330 7283 368
rect 7221 296 7235 330
rect 7269 296 7283 330
rect 7221 258 7283 296
rect 7221 224 7235 258
rect 7269 224 7283 258
rect 7221 186 7283 224
rect 7221 152 7235 186
rect 7269 152 7283 186
rect 7221 114 7283 152
rect 6555 47 6617 80
rect 7221 80 7235 114
rect 7269 80 7283 114
rect 7887 368 7901 402
rect 7935 368 7949 402
rect 8553 474 8615 510
rect 8553 440 8567 474
rect 8601 440 8615 474
rect 8553 402 8615 440
rect 7887 330 7949 368
rect 7887 296 7901 330
rect 7935 296 7949 330
rect 7887 258 7949 296
rect 7887 224 7901 258
rect 7935 224 7949 258
rect 7887 186 7949 224
rect 7887 152 7901 186
rect 7935 152 7949 186
rect 7887 114 7949 152
rect 7221 47 7283 80
rect 7887 80 7901 114
rect 7935 80 7949 114
rect 8553 368 8567 402
rect 8601 368 8615 402
rect 9515 474 9577 510
rect 9515 440 9529 474
rect 9563 440 9577 474
rect 9515 402 9577 440
rect 8553 330 8615 368
rect 8553 296 8567 330
rect 8601 296 8615 330
rect 8553 258 8615 296
rect 8553 224 8567 258
rect 8601 224 8615 258
rect 8553 186 8615 224
rect 8553 152 8567 186
rect 8601 152 8615 186
rect 8553 114 8615 152
rect 7887 47 7949 80
rect 8553 80 8567 114
rect 8601 80 8615 114
rect 9515 368 9529 402
rect 9563 368 9577 402
rect 10181 474 10243 510
rect 10181 440 10195 474
rect 10229 440 10243 474
rect 10181 402 10243 440
rect 9515 330 9577 368
rect 9515 296 9529 330
rect 9563 296 9577 330
rect 9515 258 9577 296
rect 9515 224 9529 258
rect 9563 224 9577 258
rect 9515 186 9577 224
rect 9515 152 9529 186
rect 9563 152 9577 186
rect 9515 114 9577 152
rect 8553 47 8615 80
rect 9515 80 9529 114
rect 9563 80 9577 114
rect 10181 368 10195 402
rect 10229 368 10243 402
rect 10847 474 10909 510
rect 10847 440 10861 474
rect 10895 440 10909 474
rect 10847 402 10909 440
rect 10181 330 10243 368
rect 10181 296 10195 330
rect 10229 296 10243 330
rect 10181 258 10243 296
rect 10181 224 10195 258
rect 10229 224 10243 258
rect 10181 186 10243 224
rect 10181 152 10195 186
rect 10229 152 10243 186
rect 10181 114 10243 152
rect 9515 47 9577 80
rect 10181 80 10195 114
rect 10229 80 10243 114
rect 10847 368 10861 402
rect 10895 368 10909 402
rect 11513 474 11575 510
rect 11513 440 11527 474
rect 11561 440 11575 474
rect 11513 402 11575 440
rect 10847 330 10909 368
rect 10847 296 10861 330
rect 10895 296 10909 330
rect 10847 258 10909 296
rect 10847 224 10861 258
rect 10895 224 10909 258
rect 10847 186 10909 224
rect 10847 152 10861 186
rect 10895 152 10909 186
rect 10847 114 10909 152
rect 10181 47 10243 80
rect 10847 80 10861 114
rect 10895 80 10909 114
rect 11513 368 11527 402
rect 11561 368 11575 402
rect 12179 474 12241 510
rect 12179 440 12193 474
rect 12227 440 12241 474
rect 12179 402 12241 440
rect 11513 330 11575 368
rect 11513 296 11527 330
rect 11561 296 11575 330
rect 11513 258 11575 296
rect 11513 224 11527 258
rect 11561 224 11575 258
rect 11513 186 11575 224
rect 11513 152 11527 186
rect 11561 152 11575 186
rect 11513 114 11575 152
rect 10847 47 10909 80
rect 11513 80 11527 114
rect 11561 80 11575 114
rect 12179 368 12193 402
rect 12227 368 12241 402
rect 12845 474 12907 510
rect 12845 440 12859 474
rect 12893 440 12907 474
rect 12845 402 12907 440
rect 13511 474 13573 510
rect 13511 440 13525 474
rect 13559 440 13573 474
rect 12179 330 12241 368
rect 12179 296 12193 330
rect 12227 296 12241 330
rect 12179 258 12241 296
rect 12179 224 12193 258
rect 12227 224 12241 258
rect 12179 186 12241 224
rect 12179 152 12193 186
rect 12227 152 12241 186
rect 12179 114 12241 152
rect 11513 47 11575 80
rect 12179 80 12193 114
rect 12227 80 12241 114
rect 12845 368 12859 402
rect 12893 368 12907 402
rect 13511 402 13573 440
rect 12845 330 12907 368
rect 12845 296 12859 330
rect 12893 296 12907 330
rect 12845 258 12907 296
rect 12845 224 12859 258
rect 12893 224 12907 258
rect 12845 186 12907 224
rect 12845 152 12859 186
rect 12893 152 12907 186
rect 12845 114 12907 152
rect 12179 47 12241 80
rect 12845 80 12859 114
rect 12893 80 12907 114
rect 13511 368 13525 402
rect 13559 368 13573 402
rect 14177 474 14239 510
rect 14177 440 14191 474
rect 14225 440 14239 474
rect 14177 402 14239 440
rect 14843 474 14905 510
rect 14843 440 14857 474
rect 14891 440 14905 474
rect 13511 330 13573 368
rect 13511 296 13525 330
rect 13559 296 13573 330
rect 13511 258 13573 296
rect 13511 224 13525 258
rect 13559 224 13573 258
rect 13511 186 13573 224
rect 13511 152 13525 186
rect 13559 152 13573 186
rect 13511 114 13573 152
rect 12845 47 12907 80
rect 13511 80 13525 114
rect 13559 80 13573 114
rect 14177 368 14191 402
rect 14225 368 14239 402
rect 14843 402 14905 440
rect 14177 330 14239 368
rect 14177 296 14191 330
rect 14225 296 14239 330
rect 14177 258 14239 296
rect 14177 224 14191 258
rect 14225 224 14239 258
rect 14177 186 14239 224
rect 14177 152 14191 186
rect 14225 152 14239 186
rect 14177 114 14239 152
rect 13511 47 13573 80
rect 14177 80 14191 114
rect 14225 80 14239 114
rect 14843 368 14857 402
rect 14891 368 14905 402
rect 14843 330 14905 368
rect 14843 296 14857 330
rect 14891 296 14905 330
rect 14843 258 14905 296
rect 14843 224 14857 258
rect 14891 224 14905 258
rect 14843 186 14905 224
rect 14843 152 14857 186
rect 14891 152 14905 186
rect 14843 114 14905 152
rect 14177 47 14239 80
rect 14843 80 14857 114
rect 14891 80 14905 114
rect 14843 47 14905 80
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 343 47
rect 377 13 415 47
rect 449 13 513 47
rect 547 13 585 47
rect 619 13 657 47
rect 691 13 729 47
rect 763 13 801 47
rect 835 13 873 47
rect 907 13 1017 47
rect 1051 13 1089 47
rect 1123 13 1161 47
rect 1195 13 1233 47
rect 1267 13 1323 47
rect 1357 13 1395 47
rect 1429 13 1467 47
rect 1501 13 1539 47
rect 1573 13 1683 47
rect 1717 13 1755 47
rect 1789 13 1827 47
rect 1861 13 1899 47
rect 1933 13 1989 47
rect 2023 13 2061 47
rect 2095 13 2133 47
rect 2167 13 2205 47
rect 2239 13 2349 47
rect 2383 13 2421 47
rect 2455 13 2493 47
rect 2527 13 2565 47
rect 2599 13 2655 47
rect 2689 13 2727 47
rect 2761 13 2799 47
rect 2833 13 2871 47
rect 2905 13 3015 47
rect 3049 13 3087 47
rect 3121 13 3159 47
rect 3193 13 3231 47
rect 3265 13 3321 47
rect 3355 13 3393 47
rect 3427 13 3465 47
rect 3499 13 3537 47
rect 3571 13 3681 47
rect 3715 13 3753 47
rect 3787 13 3825 47
rect 3859 13 3897 47
rect 3931 13 3987 47
rect 4021 13 4059 47
rect 4093 13 4131 47
rect 4165 13 4203 47
rect 4237 13 4347 47
rect 4381 13 4419 47
rect 4453 13 4491 47
rect 4525 13 4563 47
rect 4597 13 4635 47
rect 4669 13 4707 47
rect 4741 13 4805 47
rect 4839 13 4877 47
rect 4911 13 4949 47
rect 4983 13 5021 47
rect 5055 13 5093 47
rect 5127 13 5165 47
rect 5199 13 5309 47
rect 5343 13 5381 47
rect 5415 13 5453 47
rect 5487 13 5525 47
rect 5559 13 5615 47
rect 5649 13 5687 47
rect 5721 13 5759 47
rect 5793 13 5831 47
rect 5865 13 5975 47
rect 6009 13 6047 47
rect 6081 13 6119 47
rect 6153 13 6191 47
rect 6225 13 6281 47
rect 6315 13 6353 47
rect 6387 13 6425 47
rect 6459 13 6497 47
rect 6531 13 6641 47
rect 6675 13 6713 47
rect 6747 13 6785 47
rect 6819 13 6857 47
rect 6891 13 6947 47
rect 6981 13 7019 47
rect 7053 13 7091 47
rect 7125 13 7163 47
rect 7197 13 7307 47
rect 7341 13 7379 47
rect 7413 13 7451 47
rect 7485 13 7523 47
rect 7557 13 7613 47
rect 7647 13 7685 47
rect 7719 13 7757 47
rect 7791 13 7829 47
rect 7863 13 7973 47
rect 8007 13 8045 47
rect 8079 13 8117 47
rect 8151 13 8189 47
rect 8223 13 8279 47
rect 8313 13 8351 47
rect 8385 13 8423 47
rect 8457 13 8495 47
rect 8529 13 8639 47
rect 8673 13 8711 47
rect 8745 13 8783 47
rect 8817 13 8855 47
rect 8889 13 8927 47
rect 8961 13 8999 47
rect 9033 13 9097 47
rect 9131 13 9169 47
rect 9203 13 9241 47
rect 9275 13 9313 47
rect 9347 13 9385 47
rect 9419 13 9457 47
rect 9491 13 9601 47
rect 9635 13 9673 47
rect 9707 13 9745 47
rect 9779 13 9817 47
rect 9851 13 9907 47
rect 9941 13 9979 47
rect 10013 13 10051 47
rect 10085 13 10123 47
rect 10157 13 10267 47
rect 10301 13 10339 47
rect 10373 13 10411 47
rect 10445 13 10483 47
rect 10517 13 10573 47
rect 10607 13 10645 47
rect 10679 13 10717 47
rect 10751 13 10789 47
rect 10823 13 10933 47
rect 10967 13 11005 47
rect 11039 13 11077 47
rect 11111 13 11149 47
rect 11183 13 11239 47
rect 11273 13 11311 47
rect 11345 13 11383 47
rect 11417 13 11455 47
rect 11489 13 11599 47
rect 11633 13 11671 47
rect 11705 13 11743 47
rect 11777 13 11815 47
rect 11849 13 11905 47
rect 11939 13 11977 47
rect 12011 13 12049 47
rect 12083 13 12121 47
rect 12155 13 12265 47
rect 12299 13 12337 47
rect 12371 13 12409 47
rect 12443 13 12481 47
rect 12515 13 12571 47
rect 12605 13 12643 47
rect 12677 13 12715 47
rect 12749 13 12787 47
rect 12821 13 12931 47
rect 12965 13 13003 47
rect 13037 13 13075 47
rect 13109 13 13147 47
rect 13181 13 13237 47
rect 13271 13 13309 47
rect 13343 13 13381 47
rect 13415 13 13453 47
rect 13487 13 13597 47
rect 13631 13 13669 47
rect 13703 13 13741 47
rect 13775 13 13813 47
rect 13847 13 13903 47
rect 13937 13 13975 47
rect 14009 13 14047 47
rect 14081 13 14119 47
rect 14153 13 14263 47
rect 14297 13 14335 47
rect 14369 13 14407 47
rect 14441 13 14479 47
rect 14513 13 14569 47
rect 14603 13 14641 47
rect 14675 13 14713 47
rect 14747 13 14785 47
rect 14819 13 14905 47
rect -31 11 31 13
rect 931 11 993 13
rect 1597 11 1659 13
rect 2263 11 2325 13
rect 2929 11 2991 13
rect 3595 11 3657 13
rect 4261 11 4323 13
rect 5223 11 5285 13
rect 5889 11 5951 13
rect 6555 11 6617 13
rect 7221 11 7283 13
rect 7887 11 7949 13
rect 8553 11 8615 13
rect 9515 11 9577 13
rect 10181 11 10243 13
rect 10847 11 10909 13
rect 11513 11 11575 13
rect 12179 11 12241 13
rect 12845 11 12907 13
rect 13511 11 13573 13
rect 14177 11 14239 13
rect 14843 11 14905 13
<< nsubdiff >>
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 343 1539
rect 377 1505 415 1539
rect 449 1505 513 1539
rect 547 1505 585 1539
rect 619 1505 657 1539
rect 691 1505 729 1539
rect 763 1505 801 1539
rect 835 1505 873 1539
rect 907 1505 1017 1539
rect 1051 1505 1089 1539
rect 1123 1505 1161 1539
rect 1195 1505 1233 1539
rect 1267 1505 1323 1539
rect 1357 1505 1395 1539
rect 1429 1505 1467 1539
rect 1501 1505 1539 1539
rect 1573 1505 1683 1539
rect 1717 1505 1755 1539
rect 1789 1505 1827 1539
rect 1861 1505 1899 1539
rect 1933 1505 1989 1539
rect 2023 1505 2061 1539
rect 2095 1505 2133 1539
rect 2167 1505 2205 1539
rect 2239 1505 2349 1539
rect 2383 1505 2421 1539
rect 2455 1505 2493 1539
rect 2527 1505 2565 1539
rect 2599 1505 2655 1539
rect 2689 1505 2727 1539
rect 2761 1505 2799 1539
rect 2833 1505 2871 1539
rect 2905 1505 3015 1539
rect 3049 1505 3087 1539
rect 3121 1505 3159 1539
rect 3193 1505 3231 1539
rect 3265 1505 3321 1539
rect 3355 1505 3393 1539
rect 3427 1505 3465 1539
rect 3499 1505 3537 1539
rect 3571 1505 3681 1539
rect 3715 1505 3753 1539
rect 3787 1505 3825 1539
rect 3859 1505 3897 1539
rect 3931 1505 3987 1539
rect 4021 1505 4059 1539
rect 4093 1505 4131 1539
rect 4165 1505 4203 1539
rect 4237 1505 4347 1539
rect 4381 1505 4419 1539
rect 4453 1505 4491 1539
rect 4525 1505 4563 1539
rect 4597 1505 4635 1539
rect 4669 1505 4707 1539
rect 4741 1505 4805 1539
rect 4839 1505 4877 1539
rect 4911 1505 4949 1539
rect 4983 1505 5021 1539
rect 5055 1505 5093 1539
rect 5127 1505 5165 1539
rect 5199 1505 5309 1539
rect 5343 1505 5381 1539
rect 5415 1505 5453 1539
rect 5487 1505 5525 1539
rect 5559 1505 5615 1539
rect 5649 1505 5687 1539
rect 5721 1505 5759 1539
rect 5793 1505 5831 1539
rect 5865 1505 5975 1539
rect 6009 1505 6047 1539
rect 6081 1505 6119 1539
rect 6153 1505 6191 1539
rect 6225 1505 6281 1539
rect 6315 1505 6353 1539
rect 6387 1505 6425 1539
rect 6459 1505 6497 1539
rect 6531 1505 6641 1539
rect 6675 1505 6713 1539
rect 6747 1505 6785 1539
rect 6819 1505 6857 1539
rect 6891 1505 6947 1539
rect 6981 1505 7019 1539
rect 7053 1505 7091 1539
rect 7125 1505 7163 1539
rect 7197 1505 7307 1539
rect 7341 1505 7379 1539
rect 7413 1505 7451 1539
rect 7485 1505 7523 1539
rect 7557 1505 7613 1539
rect 7647 1505 7685 1539
rect 7719 1505 7757 1539
rect 7791 1505 7829 1539
rect 7863 1505 7973 1539
rect 8007 1505 8045 1539
rect 8079 1505 8117 1539
rect 8151 1505 8189 1539
rect 8223 1505 8279 1539
rect 8313 1505 8351 1539
rect 8385 1505 8423 1539
rect 8457 1505 8495 1539
rect 8529 1505 8639 1539
rect 8673 1505 8711 1539
rect 8745 1505 8783 1539
rect 8817 1505 8855 1539
rect 8889 1505 8927 1539
rect 8961 1505 8999 1539
rect 9033 1505 9097 1539
rect 9131 1505 9169 1539
rect 9203 1505 9241 1539
rect 9275 1505 9313 1539
rect 9347 1505 9385 1539
rect 9419 1505 9457 1539
rect 9491 1505 9601 1539
rect 9635 1505 9673 1539
rect 9707 1505 9745 1539
rect 9779 1505 9817 1539
rect 9851 1505 9907 1539
rect 9941 1505 9979 1539
rect 10013 1505 10051 1539
rect 10085 1505 10123 1539
rect 10157 1505 10267 1539
rect 10301 1505 10339 1539
rect 10373 1505 10411 1539
rect 10445 1505 10483 1539
rect 10517 1505 10573 1539
rect 10607 1505 10645 1539
rect 10679 1505 10717 1539
rect 10751 1505 10789 1539
rect 10823 1505 10933 1539
rect 10967 1505 11005 1539
rect 11039 1505 11077 1539
rect 11111 1505 11149 1539
rect 11183 1505 11239 1539
rect 11273 1505 11311 1539
rect 11345 1505 11383 1539
rect 11417 1505 11455 1539
rect 11489 1505 11599 1539
rect 11633 1505 11671 1539
rect 11705 1505 11743 1539
rect 11777 1505 11815 1539
rect 11849 1505 11905 1539
rect 11939 1505 11977 1539
rect 12011 1505 12049 1539
rect 12083 1505 12121 1539
rect 12155 1505 12265 1539
rect 12299 1505 12337 1539
rect 12371 1505 12409 1539
rect 12443 1505 12481 1539
rect 12515 1505 12571 1539
rect 12605 1505 12643 1539
rect 12677 1505 12715 1539
rect 12749 1505 12787 1539
rect 12821 1505 12931 1539
rect 12965 1505 13003 1539
rect 13037 1505 13075 1539
rect 13109 1505 13147 1539
rect 13181 1505 13237 1539
rect 13271 1505 13309 1539
rect 13343 1505 13381 1539
rect 13415 1505 13453 1539
rect 13487 1505 13597 1539
rect 13631 1505 13669 1539
rect 13703 1505 13741 1539
rect 13775 1505 13813 1539
rect 13847 1505 13903 1539
rect 13937 1505 13975 1539
rect 14009 1505 14047 1539
rect 14081 1505 14119 1539
rect 14153 1505 14263 1539
rect 14297 1505 14335 1539
rect 14369 1505 14407 1539
rect 14441 1505 14479 1539
rect 14513 1505 14569 1539
rect 14603 1505 14641 1539
rect 14675 1505 14713 1539
rect 14747 1505 14785 1539
rect 14819 1505 14905 1539
rect -31 1470 31 1505
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect 931 1470 993 1505
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect -31 1038 31 1076
rect 931 1436 945 1470
rect 979 1436 993 1470
rect 1597 1470 1659 1505
rect 931 1398 993 1436
rect 931 1364 945 1398
rect 979 1364 993 1398
rect 931 1326 993 1364
rect 931 1292 945 1326
rect 979 1292 993 1326
rect 931 1254 993 1292
rect 931 1220 945 1254
rect 979 1220 993 1254
rect 931 1182 993 1220
rect 931 1148 945 1182
rect 979 1148 993 1182
rect 931 1110 993 1148
rect 931 1076 945 1110
rect 979 1076 993 1110
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect 931 1038 993 1076
rect 1597 1436 1611 1470
rect 1645 1436 1659 1470
rect 2263 1470 2325 1505
rect 1597 1398 1659 1436
rect 1597 1364 1611 1398
rect 1645 1364 1659 1398
rect 1597 1326 1659 1364
rect 1597 1292 1611 1326
rect 1645 1292 1659 1326
rect 1597 1254 1659 1292
rect 1597 1220 1611 1254
rect 1645 1220 1659 1254
rect 1597 1182 1659 1220
rect 1597 1148 1611 1182
rect 1645 1148 1659 1182
rect 1597 1110 1659 1148
rect 1597 1076 1611 1110
rect 1645 1076 1659 1110
rect 931 1004 945 1038
rect 979 1004 993 1038
rect 931 966 993 1004
rect -31 930 31 932
rect 931 932 945 966
rect 979 932 993 966
rect 1597 1038 1659 1076
rect 2263 1436 2277 1470
rect 2311 1436 2325 1470
rect 2929 1470 2991 1505
rect 2263 1398 2325 1436
rect 2263 1364 2277 1398
rect 2311 1364 2325 1398
rect 2263 1326 2325 1364
rect 2263 1292 2277 1326
rect 2311 1292 2325 1326
rect 2263 1254 2325 1292
rect 2263 1220 2277 1254
rect 2311 1220 2325 1254
rect 2263 1182 2325 1220
rect 2263 1148 2277 1182
rect 2311 1148 2325 1182
rect 2263 1110 2325 1148
rect 2263 1076 2277 1110
rect 2311 1076 2325 1110
rect 1597 1004 1611 1038
rect 1645 1004 1659 1038
rect 1597 966 1659 1004
rect 931 930 993 932
rect 1597 932 1611 966
rect 1645 932 1659 966
rect 2263 1038 2325 1076
rect 2929 1436 2943 1470
rect 2977 1436 2991 1470
rect 3595 1470 3657 1505
rect 2929 1398 2991 1436
rect 2929 1364 2943 1398
rect 2977 1364 2991 1398
rect 2929 1326 2991 1364
rect 2929 1292 2943 1326
rect 2977 1292 2991 1326
rect 2929 1254 2991 1292
rect 2929 1220 2943 1254
rect 2977 1220 2991 1254
rect 2929 1182 2991 1220
rect 2929 1148 2943 1182
rect 2977 1148 2991 1182
rect 2929 1110 2991 1148
rect 2929 1076 2943 1110
rect 2977 1076 2991 1110
rect 2263 1004 2277 1038
rect 2311 1004 2325 1038
rect 2263 966 2325 1004
rect 1597 930 1659 932
rect 2263 932 2277 966
rect 2311 932 2325 966
rect 2929 1038 2991 1076
rect 3595 1436 3609 1470
rect 3643 1436 3657 1470
rect 4261 1470 4323 1505
rect 3595 1398 3657 1436
rect 3595 1364 3609 1398
rect 3643 1364 3657 1398
rect 3595 1326 3657 1364
rect 3595 1292 3609 1326
rect 3643 1292 3657 1326
rect 3595 1254 3657 1292
rect 3595 1220 3609 1254
rect 3643 1220 3657 1254
rect 3595 1182 3657 1220
rect 3595 1148 3609 1182
rect 3643 1148 3657 1182
rect 3595 1110 3657 1148
rect 3595 1076 3609 1110
rect 3643 1076 3657 1110
rect 2929 1004 2943 1038
rect 2977 1004 2991 1038
rect 2929 966 2991 1004
rect 2263 930 2325 932
rect 2929 932 2943 966
rect 2977 932 2991 966
rect 3595 1038 3657 1076
rect 4261 1436 4275 1470
rect 4309 1436 4323 1470
rect 5223 1470 5285 1505
rect 4261 1398 4323 1436
rect 4261 1364 4275 1398
rect 4309 1364 4323 1398
rect 4261 1326 4323 1364
rect 4261 1292 4275 1326
rect 4309 1292 4323 1326
rect 4261 1254 4323 1292
rect 4261 1220 4275 1254
rect 4309 1220 4323 1254
rect 4261 1182 4323 1220
rect 4261 1148 4275 1182
rect 4309 1148 4323 1182
rect 4261 1110 4323 1148
rect 4261 1076 4275 1110
rect 4309 1076 4323 1110
rect 3595 1004 3609 1038
rect 3643 1004 3657 1038
rect 3595 966 3657 1004
rect 2929 930 2991 932
rect 3595 932 3609 966
rect 3643 932 3657 966
rect 4261 1038 4323 1076
rect 5223 1436 5237 1470
rect 5271 1436 5285 1470
rect 5889 1470 5951 1505
rect 5223 1398 5285 1436
rect 5223 1364 5237 1398
rect 5271 1364 5285 1398
rect 5223 1326 5285 1364
rect 5223 1292 5237 1326
rect 5271 1292 5285 1326
rect 5223 1254 5285 1292
rect 5223 1220 5237 1254
rect 5271 1220 5285 1254
rect 5223 1182 5285 1220
rect 5223 1148 5237 1182
rect 5271 1148 5285 1182
rect 5223 1110 5285 1148
rect 5223 1076 5237 1110
rect 5271 1076 5285 1110
rect 4261 1004 4275 1038
rect 4309 1004 4323 1038
rect 4261 966 4323 1004
rect 3595 930 3657 932
rect 4261 932 4275 966
rect 4309 932 4323 966
rect 5223 1038 5285 1076
rect 5889 1436 5903 1470
rect 5937 1436 5951 1470
rect 6555 1470 6617 1505
rect 5889 1398 5951 1436
rect 5889 1364 5903 1398
rect 5937 1364 5951 1398
rect 5889 1326 5951 1364
rect 5889 1292 5903 1326
rect 5937 1292 5951 1326
rect 5889 1254 5951 1292
rect 5889 1220 5903 1254
rect 5937 1220 5951 1254
rect 5889 1182 5951 1220
rect 5889 1148 5903 1182
rect 5937 1148 5951 1182
rect 5889 1110 5951 1148
rect 5889 1076 5903 1110
rect 5937 1076 5951 1110
rect 5223 1004 5237 1038
rect 5271 1004 5285 1038
rect 5223 966 5285 1004
rect 4261 930 4323 932
rect 5223 932 5237 966
rect 5271 932 5285 966
rect 5889 1038 5951 1076
rect 6555 1436 6569 1470
rect 6603 1436 6617 1470
rect 7221 1470 7283 1505
rect 6555 1398 6617 1436
rect 6555 1364 6569 1398
rect 6603 1364 6617 1398
rect 6555 1326 6617 1364
rect 6555 1292 6569 1326
rect 6603 1292 6617 1326
rect 6555 1254 6617 1292
rect 6555 1220 6569 1254
rect 6603 1220 6617 1254
rect 6555 1182 6617 1220
rect 6555 1148 6569 1182
rect 6603 1148 6617 1182
rect 6555 1110 6617 1148
rect 6555 1076 6569 1110
rect 6603 1076 6617 1110
rect 5889 1004 5903 1038
rect 5937 1004 5951 1038
rect 5889 966 5951 1004
rect 5223 930 5285 932
rect 5889 932 5903 966
rect 5937 932 5951 966
rect 6555 1038 6617 1076
rect 7221 1436 7235 1470
rect 7269 1436 7283 1470
rect 7887 1470 7949 1505
rect 7221 1398 7283 1436
rect 7221 1364 7235 1398
rect 7269 1364 7283 1398
rect 7221 1326 7283 1364
rect 7221 1292 7235 1326
rect 7269 1292 7283 1326
rect 7221 1254 7283 1292
rect 7221 1220 7235 1254
rect 7269 1220 7283 1254
rect 7221 1182 7283 1220
rect 7221 1148 7235 1182
rect 7269 1148 7283 1182
rect 7221 1110 7283 1148
rect 7221 1076 7235 1110
rect 7269 1076 7283 1110
rect 6555 1004 6569 1038
rect 6603 1004 6617 1038
rect 6555 966 6617 1004
rect 5889 930 5951 932
rect 6555 932 6569 966
rect 6603 932 6617 966
rect 7221 1038 7283 1076
rect 7887 1436 7901 1470
rect 7935 1436 7949 1470
rect 8553 1470 8615 1505
rect 7887 1398 7949 1436
rect 7887 1364 7901 1398
rect 7935 1364 7949 1398
rect 7887 1326 7949 1364
rect 7887 1292 7901 1326
rect 7935 1292 7949 1326
rect 7887 1254 7949 1292
rect 7887 1220 7901 1254
rect 7935 1220 7949 1254
rect 7887 1182 7949 1220
rect 7887 1148 7901 1182
rect 7935 1148 7949 1182
rect 7887 1110 7949 1148
rect 7887 1076 7901 1110
rect 7935 1076 7949 1110
rect 7221 1004 7235 1038
rect 7269 1004 7283 1038
rect 7221 966 7283 1004
rect 6555 930 6617 932
rect 7221 932 7235 966
rect 7269 932 7283 966
rect 7887 1038 7949 1076
rect 8553 1436 8567 1470
rect 8601 1436 8615 1470
rect 9515 1470 9577 1505
rect 8553 1398 8615 1436
rect 8553 1364 8567 1398
rect 8601 1364 8615 1398
rect 8553 1326 8615 1364
rect 8553 1292 8567 1326
rect 8601 1292 8615 1326
rect 8553 1254 8615 1292
rect 8553 1220 8567 1254
rect 8601 1220 8615 1254
rect 8553 1182 8615 1220
rect 8553 1148 8567 1182
rect 8601 1148 8615 1182
rect 8553 1110 8615 1148
rect 8553 1076 8567 1110
rect 8601 1076 8615 1110
rect 7887 1004 7901 1038
rect 7935 1004 7949 1038
rect 7887 966 7949 1004
rect 7221 930 7283 932
rect 7887 932 7901 966
rect 7935 932 7949 966
rect 8553 1038 8615 1076
rect 9515 1436 9529 1470
rect 9563 1436 9577 1470
rect 10181 1470 10243 1505
rect 9515 1398 9577 1436
rect 9515 1364 9529 1398
rect 9563 1364 9577 1398
rect 9515 1326 9577 1364
rect 9515 1292 9529 1326
rect 9563 1292 9577 1326
rect 9515 1254 9577 1292
rect 9515 1220 9529 1254
rect 9563 1220 9577 1254
rect 9515 1182 9577 1220
rect 9515 1148 9529 1182
rect 9563 1148 9577 1182
rect 9515 1110 9577 1148
rect 9515 1076 9529 1110
rect 9563 1076 9577 1110
rect 8553 1004 8567 1038
rect 8601 1004 8615 1038
rect 8553 966 8615 1004
rect 7887 930 7949 932
rect 8553 932 8567 966
rect 8601 932 8615 966
rect 9515 1038 9577 1076
rect 10181 1436 10195 1470
rect 10229 1436 10243 1470
rect 10847 1470 10909 1505
rect 10181 1398 10243 1436
rect 10181 1364 10195 1398
rect 10229 1364 10243 1398
rect 10181 1326 10243 1364
rect 10181 1292 10195 1326
rect 10229 1292 10243 1326
rect 10181 1254 10243 1292
rect 10181 1220 10195 1254
rect 10229 1220 10243 1254
rect 10181 1182 10243 1220
rect 10181 1148 10195 1182
rect 10229 1148 10243 1182
rect 10181 1110 10243 1148
rect 10181 1076 10195 1110
rect 10229 1076 10243 1110
rect 9515 1004 9529 1038
rect 9563 1004 9577 1038
rect 9515 966 9577 1004
rect 8553 930 8615 932
rect 9515 932 9529 966
rect 9563 932 9577 966
rect 10181 1038 10243 1076
rect 10847 1436 10861 1470
rect 10895 1436 10909 1470
rect 11513 1470 11575 1505
rect 10847 1398 10909 1436
rect 10847 1364 10861 1398
rect 10895 1364 10909 1398
rect 10847 1326 10909 1364
rect 10847 1292 10861 1326
rect 10895 1292 10909 1326
rect 10847 1254 10909 1292
rect 10847 1220 10861 1254
rect 10895 1220 10909 1254
rect 10847 1182 10909 1220
rect 10847 1148 10861 1182
rect 10895 1148 10909 1182
rect 10847 1110 10909 1148
rect 10847 1076 10861 1110
rect 10895 1076 10909 1110
rect 10181 1004 10195 1038
rect 10229 1004 10243 1038
rect 10181 966 10243 1004
rect 9515 930 9577 932
rect 10181 932 10195 966
rect 10229 932 10243 966
rect 10847 1038 10909 1076
rect 11513 1436 11527 1470
rect 11561 1436 11575 1470
rect 12179 1470 12241 1505
rect 11513 1398 11575 1436
rect 11513 1364 11527 1398
rect 11561 1364 11575 1398
rect 11513 1326 11575 1364
rect 11513 1292 11527 1326
rect 11561 1292 11575 1326
rect 11513 1254 11575 1292
rect 11513 1220 11527 1254
rect 11561 1220 11575 1254
rect 11513 1182 11575 1220
rect 11513 1148 11527 1182
rect 11561 1148 11575 1182
rect 11513 1110 11575 1148
rect 11513 1076 11527 1110
rect 11561 1076 11575 1110
rect 10847 1004 10861 1038
rect 10895 1004 10909 1038
rect 10847 966 10909 1004
rect 10181 930 10243 932
rect 10847 932 10861 966
rect 10895 932 10909 966
rect 11513 1038 11575 1076
rect 12179 1436 12193 1470
rect 12227 1436 12241 1470
rect 12845 1470 12907 1505
rect 12179 1398 12241 1436
rect 12179 1364 12193 1398
rect 12227 1364 12241 1398
rect 12179 1326 12241 1364
rect 12179 1292 12193 1326
rect 12227 1292 12241 1326
rect 12179 1254 12241 1292
rect 12179 1220 12193 1254
rect 12227 1220 12241 1254
rect 12179 1182 12241 1220
rect 12179 1148 12193 1182
rect 12227 1148 12241 1182
rect 12179 1110 12241 1148
rect 12179 1076 12193 1110
rect 12227 1076 12241 1110
rect 11513 1004 11527 1038
rect 11561 1004 11575 1038
rect 11513 966 11575 1004
rect 10847 930 10909 932
rect 11513 932 11527 966
rect 11561 932 11575 966
rect 12179 1038 12241 1076
rect 12845 1436 12859 1470
rect 12893 1436 12907 1470
rect 13511 1470 13573 1505
rect 12845 1398 12907 1436
rect 12845 1364 12859 1398
rect 12893 1364 12907 1398
rect 12845 1326 12907 1364
rect 12845 1292 12859 1326
rect 12893 1292 12907 1326
rect 12845 1254 12907 1292
rect 12845 1220 12859 1254
rect 12893 1220 12907 1254
rect 12845 1182 12907 1220
rect 12845 1148 12859 1182
rect 12893 1148 12907 1182
rect 12845 1110 12907 1148
rect 12845 1076 12859 1110
rect 12893 1076 12907 1110
rect 12179 1004 12193 1038
rect 12227 1004 12241 1038
rect 12179 966 12241 1004
rect 11513 930 11575 932
rect 12179 932 12193 966
rect 12227 932 12241 966
rect 12845 1038 12907 1076
rect 13511 1436 13525 1470
rect 13559 1436 13573 1470
rect 14177 1470 14239 1505
rect 13511 1398 13573 1436
rect 13511 1364 13525 1398
rect 13559 1364 13573 1398
rect 13511 1326 13573 1364
rect 13511 1292 13525 1326
rect 13559 1292 13573 1326
rect 13511 1254 13573 1292
rect 13511 1220 13525 1254
rect 13559 1220 13573 1254
rect 13511 1182 13573 1220
rect 13511 1148 13525 1182
rect 13559 1148 13573 1182
rect 13511 1110 13573 1148
rect 13511 1076 13525 1110
rect 13559 1076 13573 1110
rect 12845 1004 12859 1038
rect 12893 1004 12907 1038
rect 12845 966 12907 1004
rect 12179 930 12241 932
rect 12845 932 12859 966
rect 12893 932 12907 966
rect 13511 1038 13573 1076
rect 14177 1436 14191 1470
rect 14225 1436 14239 1470
rect 14843 1470 14905 1505
rect 14177 1398 14239 1436
rect 14177 1364 14191 1398
rect 14225 1364 14239 1398
rect 14177 1326 14239 1364
rect 14177 1292 14191 1326
rect 14225 1292 14239 1326
rect 14177 1254 14239 1292
rect 14177 1220 14191 1254
rect 14225 1220 14239 1254
rect 14177 1182 14239 1220
rect 14177 1148 14191 1182
rect 14225 1148 14239 1182
rect 14177 1110 14239 1148
rect 14177 1076 14191 1110
rect 14225 1076 14239 1110
rect 13511 1004 13525 1038
rect 13559 1004 13573 1038
rect 13511 966 13573 1004
rect 12845 930 12907 932
rect 13511 932 13525 966
rect 13559 932 13573 966
rect 14177 1038 14239 1076
rect 14843 1436 14857 1470
rect 14891 1436 14905 1470
rect 14843 1398 14905 1436
rect 14843 1364 14857 1398
rect 14891 1364 14905 1398
rect 14843 1326 14905 1364
rect 14843 1292 14857 1326
rect 14891 1292 14905 1326
rect 14843 1254 14905 1292
rect 14843 1220 14857 1254
rect 14891 1220 14905 1254
rect 14843 1182 14905 1220
rect 14843 1148 14857 1182
rect 14891 1148 14905 1182
rect 14843 1110 14905 1148
rect 14843 1076 14857 1110
rect 14891 1076 14905 1110
rect 14177 1004 14191 1038
rect 14225 1004 14239 1038
rect 14177 966 14239 1004
rect 13511 930 13573 932
rect 14177 932 14191 966
rect 14225 932 14239 966
rect 14843 1038 14905 1076
rect 14843 1004 14857 1038
rect 14891 1004 14905 1038
rect 14843 966 14905 1004
rect 14177 930 14239 932
rect 14843 932 14857 966
rect 14891 932 14905 966
rect 14843 930 14905 932
rect -31 868 14905 930
<< psubdiffcont >>
rect -17 512 17 546
rect 945 512 979 546
rect 1611 512 1645 546
rect 2277 512 2311 546
rect 2943 512 2977 546
rect 3609 512 3643 546
rect 4275 512 4309 546
rect 5237 512 5271 546
rect 5903 512 5937 546
rect 6569 512 6603 546
rect 7235 512 7269 546
rect 7901 512 7935 546
rect 8567 512 8601 546
rect 9529 512 9563 546
rect 10195 512 10229 546
rect 10861 512 10895 546
rect 11527 512 11561 546
rect 12193 512 12227 546
rect 12859 512 12893 546
rect 13525 512 13559 546
rect 14191 512 14225 546
rect 14857 512 14891 546
rect -17 440 17 474
rect -17 368 17 402
rect 945 440 979 474
rect -17 296 17 330
rect -17 224 17 258
rect -17 152 17 186
rect -17 80 17 114
rect 945 368 979 402
rect 1611 440 1645 474
rect 945 296 979 330
rect 945 224 979 258
rect 945 152 979 186
rect 945 80 979 114
rect 1611 368 1645 402
rect 2277 440 2311 474
rect 1611 296 1645 330
rect 1611 224 1645 258
rect 1611 152 1645 186
rect 1611 80 1645 114
rect 2277 368 2311 402
rect 2943 440 2977 474
rect 2277 296 2311 330
rect 2277 224 2311 258
rect 2277 152 2311 186
rect 2277 80 2311 114
rect 2943 368 2977 402
rect 3609 440 3643 474
rect 2943 296 2977 330
rect 2943 224 2977 258
rect 2943 152 2977 186
rect 2943 80 2977 114
rect 3609 368 3643 402
rect 4275 440 4309 474
rect 3609 296 3643 330
rect 3609 224 3643 258
rect 3609 152 3643 186
rect 3609 80 3643 114
rect 4275 368 4309 402
rect 5237 440 5271 474
rect 4275 296 4309 330
rect 4275 224 4309 258
rect 4275 152 4309 186
rect 4275 80 4309 114
rect 5237 368 5271 402
rect 5903 440 5937 474
rect 5237 296 5271 330
rect 5237 224 5271 258
rect 5237 152 5271 186
rect 5237 80 5271 114
rect 5903 368 5937 402
rect 6569 440 6603 474
rect 5903 296 5937 330
rect 5903 224 5937 258
rect 5903 152 5937 186
rect 5903 80 5937 114
rect 6569 368 6603 402
rect 7235 440 7269 474
rect 6569 296 6603 330
rect 6569 224 6603 258
rect 6569 152 6603 186
rect 6569 80 6603 114
rect 7235 368 7269 402
rect 7901 440 7935 474
rect 7235 296 7269 330
rect 7235 224 7269 258
rect 7235 152 7269 186
rect 7235 80 7269 114
rect 7901 368 7935 402
rect 8567 440 8601 474
rect 7901 296 7935 330
rect 7901 224 7935 258
rect 7901 152 7935 186
rect 7901 80 7935 114
rect 8567 368 8601 402
rect 9529 440 9563 474
rect 8567 296 8601 330
rect 8567 224 8601 258
rect 8567 152 8601 186
rect 8567 80 8601 114
rect 9529 368 9563 402
rect 10195 440 10229 474
rect 9529 296 9563 330
rect 9529 224 9563 258
rect 9529 152 9563 186
rect 9529 80 9563 114
rect 10195 368 10229 402
rect 10861 440 10895 474
rect 10195 296 10229 330
rect 10195 224 10229 258
rect 10195 152 10229 186
rect 10195 80 10229 114
rect 10861 368 10895 402
rect 11527 440 11561 474
rect 10861 296 10895 330
rect 10861 224 10895 258
rect 10861 152 10895 186
rect 10861 80 10895 114
rect 11527 368 11561 402
rect 12193 440 12227 474
rect 11527 296 11561 330
rect 11527 224 11561 258
rect 11527 152 11561 186
rect 11527 80 11561 114
rect 12193 368 12227 402
rect 12859 440 12893 474
rect 13525 440 13559 474
rect 12193 296 12227 330
rect 12193 224 12227 258
rect 12193 152 12227 186
rect 12193 80 12227 114
rect 12859 368 12893 402
rect 12859 296 12893 330
rect 12859 224 12893 258
rect 12859 152 12893 186
rect 12859 80 12893 114
rect 13525 368 13559 402
rect 14191 440 14225 474
rect 14857 440 14891 474
rect 13525 296 13559 330
rect 13525 224 13559 258
rect 13525 152 13559 186
rect 13525 80 13559 114
rect 14191 368 14225 402
rect 14191 296 14225 330
rect 14191 224 14225 258
rect 14191 152 14225 186
rect 14191 80 14225 114
rect 14857 368 14891 402
rect 14857 296 14891 330
rect 14857 224 14891 258
rect 14857 152 14891 186
rect 14857 80 14891 114
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 343 13 377 47
rect 415 13 449 47
rect 513 13 547 47
rect 585 13 619 47
rect 657 13 691 47
rect 729 13 763 47
rect 801 13 835 47
rect 873 13 907 47
rect 1017 13 1051 47
rect 1089 13 1123 47
rect 1161 13 1195 47
rect 1233 13 1267 47
rect 1323 13 1357 47
rect 1395 13 1429 47
rect 1467 13 1501 47
rect 1539 13 1573 47
rect 1683 13 1717 47
rect 1755 13 1789 47
rect 1827 13 1861 47
rect 1899 13 1933 47
rect 1989 13 2023 47
rect 2061 13 2095 47
rect 2133 13 2167 47
rect 2205 13 2239 47
rect 2349 13 2383 47
rect 2421 13 2455 47
rect 2493 13 2527 47
rect 2565 13 2599 47
rect 2655 13 2689 47
rect 2727 13 2761 47
rect 2799 13 2833 47
rect 2871 13 2905 47
rect 3015 13 3049 47
rect 3087 13 3121 47
rect 3159 13 3193 47
rect 3231 13 3265 47
rect 3321 13 3355 47
rect 3393 13 3427 47
rect 3465 13 3499 47
rect 3537 13 3571 47
rect 3681 13 3715 47
rect 3753 13 3787 47
rect 3825 13 3859 47
rect 3897 13 3931 47
rect 3987 13 4021 47
rect 4059 13 4093 47
rect 4131 13 4165 47
rect 4203 13 4237 47
rect 4347 13 4381 47
rect 4419 13 4453 47
rect 4491 13 4525 47
rect 4563 13 4597 47
rect 4635 13 4669 47
rect 4707 13 4741 47
rect 4805 13 4839 47
rect 4877 13 4911 47
rect 4949 13 4983 47
rect 5021 13 5055 47
rect 5093 13 5127 47
rect 5165 13 5199 47
rect 5309 13 5343 47
rect 5381 13 5415 47
rect 5453 13 5487 47
rect 5525 13 5559 47
rect 5615 13 5649 47
rect 5687 13 5721 47
rect 5759 13 5793 47
rect 5831 13 5865 47
rect 5975 13 6009 47
rect 6047 13 6081 47
rect 6119 13 6153 47
rect 6191 13 6225 47
rect 6281 13 6315 47
rect 6353 13 6387 47
rect 6425 13 6459 47
rect 6497 13 6531 47
rect 6641 13 6675 47
rect 6713 13 6747 47
rect 6785 13 6819 47
rect 6857 13 6891 47
rect 6947 13 6981 47
rect 7019 13 7053 47
rect 7091 13 7125 47
rect 7163 13 7197 47
rect 7307 13 7341 47
rect 7379 13 7413 47
rect 7451 13 7485 47
rect 7523 13 7557 47
rect 7613 13 7647 47
rect 7685 13 7719 47
rect 7757 13 7791 47
rect 7829 13 7863 47
rect 7973 13 8007 47
rect 8045 13 8079 47
rect 8117 13 8151 47
rect 8189 13 8223 47
rect 8279 13 8313 47
rect 8351 13 8385 47
rect 8423 13 8457 47
rect 8495 13 8529 47
rect 8639 13 8673 47
rect 8711 13 8745 47
rect 8783 13 8817 47
rect 8855 13 8889 47
rect 8927 13 8961 47
rect 8999 13 9033 47
rect 9097 13 9131 47
rect 9169 13 9203 47
rect 9241 13 9275 47
rect 9313 13 9347 47
rect 9385 13 9419 47
rect 9457 13 9491 47
rect 9601 13 9635 47
rect 9673 13 9707 47
rect 9745 13 9779 47
rect 9817 13 9851 47
rect 9907 13 9941 47
rect 9979 13 10013 47
rect 10051 13 10085 47
rect 10123 13 10157 47
rect 10267 13 10301 47
rect 10339 13 10373 47
rect 10411 13 10445 47
rect 10483 13 10517 47
rect 10573 13 10607 47
rect 10645 13 10679 47
rect 10717 13 10751 47
rect 10789 13 10823 47
rect 10933 13 10967 47
rect 11005 13 11039 47
rect 11077 13 11111 47
rect 11149 13 11183 47
rect 11239 13 11273 47
rect 11311 13 11345 47
rect 11383 13 11417 47
rect 11455 13 11489 47
rect 11599 13 11633 47
rect 11671 13 11705 47
rect 11743 13 11777 47
rect 11815 13 11849 47
rect 11905 13 11939 47
rect 11977 13 12011 47
rect 12049 13 12083 47
rect 12121 13 12155 47
rect 12265 13 12299 47
rect 12337 13 12371 47
rect 12409 13 12443 47
rect 12481 13 12515 47
rect 12571 13 12605 47
rect 12643 13 12677 47
rect 12715 13 12749 47
rect 12787 13 12821 47
rect 12931 13 12965 47
rect 13003 13 13037 47
rect 13075 13 13109 47
rect 13147 13 13181 47
rect 13237 13 13271 47
rect 13309 13 13343 47
rect 13381 13 13415 47
rect 13453 13 13487 47
rect 13597 13 13631 47
rect 13669 13 13703 47
rect 13741 13 13775 47
rect 13813 13 13847 47
rect 13903 13 13937 47
rect 13975 13 14009 47
rect 14047 13 14081 47
rect 14119 13 14153 47
rect 14263 13 14297 47
rect 14335 13 14369 47
rect 14407 13 14441 47
rect 14479 13 14513 47
rect 14569 13 14603 47
rect 14641 13 14675 47
rect 14713 13 14747 47
rect 14785 13 14819 47
<< nsubdiffcont >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 343 1505 377 1539
rect 415 1505 449 1539
rect 513 1505 547 1539
rect 585 1505 619 1539
rect 657 1505 691 1539
rect 729 1505 763 1539
rect 801 1505 835 1539
rect 873 1505 907 1539
rect 1017 1505 1051 1539
rect 1089 1505 1123 1539
rect 1161 1505 1195 1539
rect 1233 1505 1267 1539
rect 1323 1505 1357 1539
rect 1395 1505 1429 1539
rect 1467 1505 1501 1539
rect 1539 1505 1573 1539
rect 1683 1505 1717 1539
rect 1755 1505 1789 1539
rect 1827 1505 1861 1539
rect 1899 1505 1933 1539
rect 1989 1505 2023 1539
rect 2061 1505 2095 1539
rect 2133 1505 2167 1539
rect 2205 1505 2239 1539
rect 2349 1505 2383 1539
rect 2421 1505 2455 1539
rect 2493 1505 2527 1539
rect 2565 1505 2599 1539
rect 2655 1505 2689 1539
rect 2727 1505 2761 1539
rect 2799 1505 2833 1539
rect 2871 1505 2905 1539
rect 3015 1505 3049 1539
rect 3087 1505 3121 1539
rect 3159 1505 3193 1539
rect 3231 1505 3265 1539
rect 3321 1505 3355 1539
rect 3393 1505 3427 1539
rect 3465 1505 3499 1539
rect 3537 1505 3571 1539
rect 3681 1505 3715 1539
rect 3753 1505 3787 1539
rect 3825 1505 3859 1539
rect 3897 1505 3931 1539
rect 3987 1505 4021 1539
rect 4059 1505 4093 1539
rect 4131 1505 4165 1539
rect 4203 1505 4237 1539
rect 4347 1505 4381 1539
rect 4419 1505 4453 1539
rect 4491 1505 4525 1539
rect 4563 1505 4597 1539
rect 4635 1505 4669 1539
rect 4707 1505 4741 1539
rect 4805 1505 4839 1539
rect 4877 1505 4911 1539
rect 4949 1505 4983 1539
rect 5021 1505 5055 1539
rect 5093 1505 5127 1539
rect 5165 1505 5199 1539
rect 5309 1505 5343 1539
rect 5381 1505 5415 1539
rect 5453 1505 5487 1539
rect 5525 1505 5559 1539
rect 5615 1505 5649 1539
rect 5687 1505 5721 1539
rect 5759 1505 5793 1539
rect 5831 1505 5865 1539
rect 5975 1505 6009 1539
rect 6047 1505 6081 1539
rect 6119 1505 6153 1539
rect 6191 1505 6225 1539
rect 6281 1505 6315 1539
rect 6353 1505 6387 1539
rect 6425 1505 6459 1539
rect 6497 1505 6531 1539
rect 6641 1505 6675 1539
rect 6713 1505 6747 1539
rect 6785 1505 6819 1539
rect 6857 1505 6891 1539
rect 6947 1505 6981 1539
rect 7019 1505 7053 1539
rect 7091 1505 7125 1539
rect 7163 1505 7197 1539
rect 7307 1505 7341 1539
rect 7379 1505 7413 1539
rect 7451 1505 7485 1539
rect 7523 1505 7557 1539
rect 7613 1505 7647 1539
rect 7685 1505 7719 1539
rect 7757 1505 7791 1539
rect 7829 1505 7863 1539
rect 7973 1505 8007 1539
rect 8045 1505 8079 1539
rect 8117 1505 8151 1539
rect 8189 1505 8223 1539
rect 8279 1505 8313 1539
rect 8351 1505 8385 1539
rect 8423 1505 8457 1539
rect 8495 1505 8529 1539
rect 8639 1505 8673 1539
rect 8711 1505 8745 1539
rect 8783 1505 8817 1539
rect 8855 1505 8889 1539
rect 8927 1505 8961 1539
rect 8999 1505 9033 1539
rect 9097 1505 9131 1539
rect 9169 1505 9203 1539
rect 9241 1505 9275 1539
rect 9313 1505 9347 1539
rect 9385 1505 9419 1539
rect 9457 1505 9491 1539
rect 9601 1505 9635 1539
rect 9673 1505 9707 1539
rect 9745 1505 9779 1539
rect 9817 1505 9851 1539
rect 9907 1505 9941 1539
rect 9979 1505 10013 1539
rect 10051 1505 10085 1539
rect 10123 1505 10157 1539
rect 10267 1505 10301 1539
rect 10339 1505 10373 1539
rect 10411 1505 10445 1539
rect 10483 1505 10517 1539
rect 10573 1505 10607 1539
rect 10645 1505 10679 1539
rect 10717 1505 10751 1539
rect 10789 1505 10823 1539
rect 10933 1505 10967 1539
rect 11005 1505 11039 1539
rect 11077 1505 11111 1539
rect 11149 1505 11183 1539
rect 11239 1505 11273 1539
rect 11311 1505 11345 1539
rect 11383 1505 11417 1539
rect 11455 1505 11489 1539
rect 11599 1505 11633 1539
rect 11671 1505 11705 1539
rect 11743 1505 11777 1539
rect 11815 1505 11849 1539
rect 11905 1505 11939 1539
rect 11977 1505 12011 1539
rect 12049 1505 12083 1539
rect 12121 1505 12155 1539
rect 12265 1505 12299 1539
rect 12337 1505 12371 1539
rect 12409 1505 12443 1539
rect 12481 1505 12515 1539
rect 12571 1505 12605 1539
rect 12643 1505 12677 1539
rect 12715 1505 12749 1539
rect 12787 1505 12821 1539
rect 12931 1505 12965 1539
rect 13003 1505 13037 1539
rect 13075 1505 13109 1539
rect 13147 1505 13181 1539
rect 13237 1505 13271 1539
rect 13309 1505 13343 1539
rect 13381 1505 13415 1539
rect 13453 1505 13487 1539
rect 13597 1505 13631 1539
rect 13669 1505 13703 1539
rect 13741 1505 13775 1539
rect 13813 1505 13847 1539
rect 13903 1505 13937 1539
rect 13975 1505 14009 1539
rect 14047 1505 14081 1539
rect 14119 1505 14153 1539
rect 14263 1505 14297 1539
rect 14335 1505 14369 1539
rect 14407 1505 14441 1539
rect 14479 1505 14513 1539
rect 14569 1505 14603 1539
rect 14641 1505 14675 1539
rect 14713 1505 14747 1539
rect 14785 1505 14819 1539
rect -17 1436 17 1470
rect -17 1364 17 1398
rect -17 1292 17 1326
rect -17 1220 17 1254
rect -17 1148 17 1182
rect -17 1076 17 1110
rect 945 1436 979 1470
rect 945 1364 979 1398
rect 945 1292 979 1326
rect 945 1220 979 1254
rect 945 1148 979 1182
rect 945 1076 979 1110
rect -17 1004 17 1038
rect -17 932 17 966
rect 1611 1436 1645 1470
rect 1611 1364 1645 1398
rect 1611 1292 1645 1326
rect 1611 1220 1645 1254
rect 1611 1148 1645 1182
rect 1611 1076 1645 1110
rect 945 1004 979 1038
rect 945 932 979 966
rect 2277 1436 2311 1470
rect 2277 1364 2311 1398
rect 2277 1292 2311 1326
rect 2277 1220 2311 1254
rect 2277 1148 2311 1182
rect 2277 1076 2311 1110
rect 1611 1004 1645 1038
rect 1611 932 1645 966
rect 2943 1436 2977 1470
rect 2943 1364 2977 1398
rect 2943 1292 2977 1326
rect 2943 1220 2977 1254
rect 2943 1148 2977 1182
rect 2943 1076 2977 1110
rect 2277 1004 2311 1038
rect 2277 932 2311 966
rect 3609 1436 3643 1470
rect 3609 1364 3643 1398
rect 3609 1292 3643 1326
rect 3609 1220 3643 1254
rect 3609 1148 3643 1182
rect 3609 1076 3643 1110
rect 2943 1004 2977 1038
rect 2943 932 2977 966
rect 4275 1436 4309 1470
rect 4275 1364 4309 1398
rect 4275 1292 4309 1326
rect 4275 1220 4309 1254
rect 4275 1148 4309 1182
rect 4275 1076 4309 1110
rect 3609 1004 3643 1038
rect 3609 932 3643 966
rect 5237 1436 5271 1470
rect 5237 1364 5271 1398
rect 5237 1292 5271 1326
rect 5237 1220 5271 1254
rect 5237 1148 5271 1182
rect 5237 1076 5271 1110
rect 4275 1004 4309 1038
rect 4275 932 4309 966
rect 5903 1436 5937 1470
rect 5903 1364 5937 1398
rect 5903 1292 5937 1326
rect 5903 1220 5937 1254
rect 5903 1148 5937 1182
rect 5903 1076 5937 1110
rect 5237 1004 5271 1038
rect 5237 932 5271 966
rect 6569 1436 6603 1470
rect 6569 1364 6603 1398
rect 6569 1292 6603 1326
rect 6569 1220 6603 1254
rect 6569 1148 6603 1182
rect 6569 1076 6603 1110
rect 5903 1004 5937 1038
rect 5903 932 5937 966
rect 7235 1436 7269 1470
rect 7235 1364 7269 1398
rect 7235 1292 7269 1326
rect 7235 1220 7269 1254
rect 7235 1148 7269 1182
rect 7235 1076 7269 1110
rect 6569 1004 6603 1038
rect 6569 932 6603 966
rect 7901 1436 7935 1470
rect 7901 1364 7935 1398
rect 7901 1292 7935 1326
rect 7901 1220 7935 1254
rect 7901 1148 7935 1182
rect 7901 1076 7935 1110
rect 7235 1004 7269 1038
rect 7235 932 7269 966
rect 8567 1436 8601 1470
rect 8567 1364 8601 1398
rect 8567 1292 8601 1326
rect 8567 1220 8601 1254
rect 8567 1148 8601 1182
rect 8567 1076 8601 1110
rect 7901 1004 7935 1038
rect 7901 932 7935 966
rect 9529 1436 9563 1470
rect 9529 1364 9563 1398
rect 9529 1292 9563 1326
rect 9529 1220 9563 1254
rect 9529 1148 9563 1182
rect 9529 1076 9563 1110
rect 8567 1004 8601 1038
rect 8567 932 8601 966
rect 10195 1436 10229 1470
rect 10195 1364 10229 1398
rect 10195 1292 10229 1326
rect 10195 1220 10229 1254
rect 10195 1148 10229 1182
rect 10195 1076 10229 1110
rect 9529 1004 9563 1038
rect 9529 932 9563 966
rect 10861 1436 10895 1470
rect 10861 1364 10895 1398
rect 10861 1292 10895 1326
rect 10861 1220 10895 1254
rect 10861 1148 10895 1182
rect 10861 1076 10895 1110
rect 10195 1004 10229 1038
rect 10195 932 10229 966
rect 11527 1436 11561 1470
rect 11527 1364 11561 1398
rect 11527 1292 11561 1326
rect 11527 1220 11561 1254
rect 11527 1148 11561 1182
rect 11527 1076 11561 1110
rect 10861 1004 10895 1038
rect 10861 932 10895 966
rect 12193 1436 12227 1470
rect 12193 1364 12227 1398
rect 12193 1292 12227 1326
rect 12193 1220 12227 1254
rect 12193 1148 12227 1182
rect 12193 1076 12227 1110
rect 11527 1004 11561 1038
rect 11527 932 11561 966
rect 12859 1436 12893 1470
rect 12859 1364 12893 1398
rect 12859 1292 12893 1326
rect 12859 1220 12893 1254
rect 12859 1148 12893 1182
rect 12859 1076 12893 1110
rect 12193 1004 12227 1038
rect 12193 932 12227 966
rect 13525 1436 13559 1470
rect 13525 1364 13559 1398
rect 13525 1292 13559 1326
rect 13525 1220 13559 1254
rect 13525 1148 13559 1182
rect 13525 1076 13559 1110
rect 12859 1004 12893 1038
rect 12859 932 12893 966
rect 14191 1436 14225 1470
rect 14191 1364 14225 1398
rect 14191 1292 14225 1326
rect 14191 1220 14225 1254
rect 14191 1148 14225 1182
rect 14191 1076 14225 1110
rect 13525 1004 13559 1038
rect 13525 932 13559 966
rect 14857 1436 14891 1470
rect 14857 1364 14891 1398
rect 14857 1292 14891 1326
rect 14857 1220 14891 1254
rect 14857 1148 14891 1182
rect 14857 1076 14891 1110
rect 14191 1004 14225 1038
rect 14191 932 14225 966
rect 14857 1004 14891 1038
rect 14857 932 14891 966
<< poly >>
rect 247 1450 277 1476
rect 335 1450 365 1476
rect 423 1450 453 1476
rect 511 1450 541 1476
rect 599 1450 629 1476
rect 687 1450 717 1476
rect 1149 1450 1179 1476
rect 1237 1450 1267 1476
rect 1325 1450 1355 1476
rect 1413 1450 1443 1476
rect 247 1019 277 1050
rect 335 1019 365 1050
rect 423 1019 453 1050
rect 511 1019 541 1050
rect 195 1003 365 1019
rect 195 969 205 1003
rect 239 989 365 1003
rect 417 1003 541 1019
rect 239 969 249 989
rect 195 953 249 969
rect 417 969 427 1003
rect 461 989 541 1003
rect 599 1019 629 1050
rect 687 1019 717 1050
rect 599 1003 717 1019
rect 599 989 649 1003
rect 461 969 471 989
rect 417 953 471 969
rect 639 969 649 989
rect 683 989 717 1003
rect 1815 1450 1845 1476
rect 1903 1450 1933 1476
rect 1991 1450 2021 1476
rect 2079 1450 2109 1476
rect 683 969 693 989
rect 639 953 693 969
rect 1149 1019 1179 1050
rect 1237 1019 1267 1050
rect 1325 1019 1355 1050
rect 1413 1019 1443 1050
rect 1149 1003 1267 1019
rect 1149 989 1167 1003
rect 1157 969 1167 989
rect 1201 989 1267 1003
rect 1311 1003 1443 1019
rect 1201 969 1211 989
rect 1157 953 1211 969
rect 1311 969 1321 1003
rect 1355 989 1443 1003
rect 2481 1450 2511 1476
rect 2569 1450 2599 1476
rect 2657 1450 2687 1476
rect 2745 1450 2775 1476
rect 1355 969 1365 989
rect 1311 953 1365 969
rect 1815 1019 1845 1050
rect 1903 1019 1933 1050
rect 1991 1019 2021 1050
rect 2079 1019 2109 1050
rect 1815 1003 1933 1019
rect 1815 989 1833 1003
rect 1823 969 1833 989
rect 1867 989 1933 1003
rect 1977 1003 2109 1019
rect 1867 969 1877 989
rect 1823 953 1877 969
rect 1977 969 1987 1003
rect 2021 989 2109 1003
rect 3147 1450 3177 1476
rect 3235 1450 3265 1476
rect 3323 1450 3353 1476
rect 3411 1450 3441 1476
rect 2021 969 2031 989
rect 1977 953 2031 969
rect 2481 1019 2511 1050
rect 2569 1019 2599 1050
rect 2657 1019 2687 1050
rect 2745 1019 2775 1050
rect 2481 1003 2599 1019
rect 2481 989 2499 1003
rect 2489 969 2499 989
rect 2533 989 2599 1003
rect 2643 1003 2775 1019
rect 2533 969 2543 989
rect 2489 953 2543 969
rect 2643 969 2653 1003
rect 2687 989 2775 1003
rect 3813 1450 3843 1476
rect 3901 1450 3931 1476
rect 3989 1450 4019 1476
rect 4077 1450 4107 1476
rect 2687 969 2697 989
rect 2643 953 2697 969
rect 3147 1019 3177 1050
rect 3235 1019 3265 1050
rect 3323 1019 3353 1050
rect 3411 1019 3441 1050
rect 3147 1003 3265 1019
rect 3147 989 3165 1003
rect 3155 969 3165 989
rect 3199 989 3265 1003
rect 3309 1003 3441 1019
rect 3199 969 3209 989
rect 3155 953 3209 969
rect 3309 969 3319 1003
rect 3353 989 3441 1003
rect 4539 1450 4569 1476
rect 4627 1450 4657 1476
rect 4715 1450 4745 1476
rect 4803 1450 4833 1476
rect 4891 1450 4921 1476
rect 4979 1450 5009 1476
rect 3353 969 3363 989
rect 3309 953 3363 969
rect 3813 1019 3843 1050
rect 3901 1019 3931 1050
rect 3989 1019 4019 1050
rect 4077 1019 4107 1050
rect 3813 1003 3931 1019
rect 3813 989 3831 1003
rect 3821 969 3831 989
rect 3865 989 3931 1003
rect 3975 1003 4107 1019
rect 3865 969 3875 989
rect 3821 953 3875 969
rect 3975 969 3985 1003
rect 4019 989 4107 1003
rect 5441 1450 5471 1476
rect 5529 1450 5559 1476
rect 5617 1450 5647 1476
rect 5705 1450 5735 1476
rect 4539 1019 4569 1050
rect 4627 1019 4657 1050
rect 4715 1019 4745 1050
rect 4803 1019 4833 1050
rect 4019 969 4029 989
rect 3975 953 4029 969
rect 4487 1003 4657 1019
rect 4487 969 4497 1003
rect 4531 989 4657 1003
rect 4709 1003 4833 1019
rect 4531 969 4541 989
rect 4487 953 4541 969
rect 4709 969 4719 1003
rect 4753 989 4833 1003
rect 4891 1019 4921 1050
rect 4979 1019 5009 1050
rect 4891 1003 5009 1019
rect 4891 989 4941 1003
rect 4753 969 4763 989
rect 4709 953 4763 969
rect 4931 969 4941 989
rect 4975 989 5009 1003
rect 6107 1450 6137 1476
rect 6195 1450 6225 1476
rect 6283 1450 6313 1476
rect 6371 1450 6401 1476
rect 4975 969 4985 989
rect 4931 953 4985 969
rect 5441 1019 5471 1050
rect 5529 1019 5559 1050
rect 5617 1019 5647 1050
rect 5705 1019 5735 1050
rect 5441 1003 5559 1019
rect 5441 989 5459 1003
rect 5449 969 5459 989
rect 5493 989 5559 1003
rect 5603 1003 5735 1019
rect 5493 969 5503 989
rect 5449 953 5503 969
rect 5603 969 5613 1003
rect 5647 989 5735 1003
rect 6773 1450 6803 1476
rect 6861 1450 6891 1476
rect 6949 1450 6979 1476
rect 7037 1450 7067 1476
rect 5647 969 5657 989
rect 5603 953 5657 969
rect 6107 1019 6137 1050
rect 6195 1019 6225 1050
rect 6283 1019 6313 1050
rect 6371 1019 6401 1050
rect 6107 1003 6225 1019
rect 6107 989 6125 1003
rect 6115 969 6125 989
rect 6159 989 6225 1003
rect 6269 1003 6401 1019
rect 6159 969 6169 989
rect 6115 953 6169 969
rect 6269 969 6279 1003
rect 6313 989 6401 1003
rect 7439 1450 7469 1476
rect 7527 1450 7557 1476
rect 7615 1450 7645 1476
rect 7703 1450 7733 1476
rect 6313 969 6323 989
rect 6269 953 6323 969
rect 6773 1019 6803 1050
rect 6861 1019 6891 1050
rect 6949 1019 6979 1050
rect 7037 1019 7067 1050
rect 6773 1003 6891 1019
rect 6773 989 6791 1003
rect 6781 969 6791 989
rect 6825 989 6891 1003
rect 6935 1003 7067 1019
rect 6825 969 6835 989
rect 6781 953 6835 969
rect 6935 969 6945 1003
rect 6979 989 7067 1003
rect 8105 1450 8135 1476
rect 8193 1450 8223 1476
rect 8281 1450 8311 1476
rect 8369 1450 8399 1476
rect 6979 969 6989 989
rect 6935 953 6989 969
rect 7439 1019 7469 1050
rect 7527 1019 7557 1050
rect 7615 1019 7645 1050
rect 7703 1019 7733 1050
rect 7439 1003 7557 1019
rect 7439 989 7457 1003
rect 7447 969 7457 989
rect 7491 989 7557 1003
rect 7601 1003 7733 1019
rect 7491 969 7501 989
rect 7447 953 7501 969
rect 7601 969 7611 1003
rect 7645 989 7733 1003
rect 8831 1450 8861 1476
rect 8919 1450 8949 1476
rect 9007 1450 9037 1476
rect 9095 1450 9125 1476
rect 9183 1450 9213 1476
rect 9271 1450 9301 1476
rect 7645 969 7655 989
rect 7601 953 7655 969
rect 8105 1019 8135 1050
rect 8193 1019 8223 1050
rect 8281 1019 8311 1050
rect 8369 1019 8399 1050
rect 8105 1003 8223 1019
rect 8105 989 8123 1003
rect 8113 969 8123 989
rect 8157 989 8223 1003
rect 8267 1003 8399 1019
rect 8157 969 8167 989
rect 8113 953 8167 969
rect 8267 969 8277 1003
rect 8311 989 8399 1003
rect 9733 1450 9763 1476
rect 9821 1450 9851 1476
rect 9909 1450 9939 1476
rect 9997 1450 10027 1476
rect 8831 1019 8861 1050
rect 8919 1019 8949 1050
rect 9007 1019 9037 1050
rect 9095 1019 9125 1050
rect 8311 969 8321 989
rect 8267 953 8321 969
rect 8779 1003 8949 1019
rect 8779 969 8789 1003
rect 8823 989 8949 1003
rect 9001 1003 9125 1019
rect 8823 969 8833 989
rect 8779 953 8833 969
rect 9001 969 9011 1003
rect 9045 989 9125 1003
rect 9183 1019 9213 1050
rect 9271 1019 9301 1050
rect 9183 1003 9301 1019
rect 9183 989 9233 1003
rect 9045 969 9055 989
rect 9001 953 9055 969
rect 9223 969 9233 989
rect 9267 989 9301 1003
rect 10399 1450 10429 1476
rect 10487 1450 10517 1476
rect 10575 1450 10605 1476
rect 10663 1450 10693 1476
rect 9267 969 9277 989
rect 9223 953 9277 969
rect 9733 1019 9763 1050
rect 9821 1019 9851 1050
rect 9909 1019 9939 1050
rect 9997 1019 10027 1050
rect 9733 1003 9851 1019
rect 9733 989 9751 1003
rect 9741 969 9751 989
rect 9785 989 9851 1003
rect 9895 1003 10027 1019
rect 9785 969 9795 989
rect 9741 953 9795 969
rect 9895 969 9905 1003
rect 9939 989 10027 1003
rect 11065 1450 11095 1476
rect 11153 1450 11183 1476
rect 11241 1450 11271 1476
rect 11329 1450 11359 1476
rect 9939 969 9949 989
rect 9895 953 9949 969
rect 10399 1019 10429 1050
rect 10487 1019 10517 1050
rect 10575 1019 10605 1050
rect 10663 1019 10693 1050
rect 10399 1003 10517 1019
rect 10399 989 10417 1003
rect 10407 969 10417 989
rect 10451 989 10517 1003
rect 10561 1003 10693 1019
rect 10451 969 10461 989
rect 10407 953 10461 969
rect 10561 969 10571 1003
rect 10605 989 10693 1003
rect 11731 1450 11761 1476
rect 11819 1450 11849 1476
rect 11907 1450 11937 1476
rect 11995 1450 12025 1476
rect 10605 969 10615 989
rect 10561 953 10615 969
rect 11065 1019 11095 1050
rect 11153 1019 11183 1050
rect 11241 1019 11271 1050
rect 11329 1019 11359 1050
rect 11065 1003 11183 1019
rect 11065 989 11083 1003
rect 11073 969 11083 989
rect 11117 989 11183 1003
rect 11227 1003 11359 1019
rect 11117 969 11127 989
rect 11073 953 11127 969
rect 11227 969 11237 1003
rect 11271 989 11359 1003
rect 12397 1450 12427 1476
rect 12485 1450 12515 1476
rect 12573 1450 12603 1476
rect 12661 1450 12691 1476
rect 11271 969 11281 989
rect 11227 953 11281 969
rect 11731 1019 11761 1050
rect 11819 1019 11849 1050
rect 11907 1019 11937 1050
rect 11995 1019 12025 1050
rect 11731 1003 11849 1019
rect 11731 989 11749 1003
rect 11739 969 11749 989
rect 11783 989 11849 1003
rect 11893 1003 12025 1019
rect 11783 969 11793 989
rect 11739 953 11793 969
rect 11893 969 11903 1003
rect 11937 989 12025 1003
rect 13063 1451 13093 1477
rect 13151 1451 13181 1477
rect 13239 1451 13269 1477
rect 13327 1451 13357 1477
rect 11937 969 11947 989
rect 11893 953 11947 969
rect 12397 1019 12427 1050
rect 12485 1019 12515 1050
rect 12573 1019 12603 1050
rect 12661 1019 12691 1050
rect 12397 1003 12515 1019
rect 12397 989 12415 1003
rect 12405 969 12415 989
rect 12449 989 12515 1003
rect 12559 1003 12691 1019
rect 12449 969 12459 989
rect 12405 953 12459 969
rect 12559 969 12569 1003
rect 12603 989 12691 1003
rect 13727 1451 13757 1477
rect 13815 1451 13845 1477
rect 13903 1451 13933 1477
rect 13991 1451 14021 1477
rect 13063 1020 13093 1051
rect 13151 1020 13181 1051
rect 13239 1020 13269 1051
rect 13327 1020 13357 1051
rect 12603 969 12613 989
rect 12559 953 12613 969
rect 12997 1004 13181 1020
rect 12997 970 13007 1004
rect 13041 990 13181 1004
rect 13227 1004 13357 1020
rect 13041 970 13051 990
rect 12997 954 13051 970
rect 13227 970 13237 1004
rect 13271 990 13357 1004
rect 14395 1451 14425 1477
rect 14483 1451 14513 1477
rect 14571 1451 14601 1477
rect 14659 1451 14689 1477
rect 13271 970 13281 990
rect 13227 954 13281 970
rect 13727 1020 13757 1051
rect 13815 1020 13845 1051
rect 13727 1004 13845 1020
rect 13727 990 13747 1004
rect 13737 970 13747 990
rect 13781 990 13845 1004
rect 13903 1020 13933 1051
rect 13991 1020 14021 1051
rect 13903 1004 14087 1020
rect 13903 990 14043 1004
rect 13781 970 13791 990
rect 13737 954 13791 970
rect 14033 970 14043 990
rect 14077 970 14087 1004
rect 14033 954 14087 970
rect 14395 1020 14425 1051
rect 14483 1020 14513 1051
rect 14571 1020 14601 1051
rect 14659 1020 14689 1051
rect 14329 1004 14513 1020
rect 14329 970 14339 1004
rect 14373 990 14513 1004
rect 14555 1004 14689 1020
rect 14373 970 14383 990
rect 14329 954 14383 970
rect 14555 970 14565 1004
rect 14599 990 14689 1004
rect 14599 970 14609 990
rect 14555 954 14609 970
rect 195 461 249 477
rect 195 441 205 461
rect 147 427 205 441
rect 239 427 249 461
rect 147 411 249 427
rect 417 461 471 477
rect 417 427 427 461
rect 461 441 471 461
rect 639 461 693 477
rect 461 427 477 441
rect 417 411 477 427
rect 639 427 649 461
rect 683 427 693 461
rect 639 411 693 427
rect 1157 461 1211 477
rect 1157 441 1167 461
rect 147 379 177 411
rect 447 379 477 411
rect 649 379 679 411
rect 1130 427 1167 441
rect 1201 427 1211 461
rect 1130 411 1211 427
rect 1305 461 1359 477
rect 1305 427 1315 461
rect 1349 427 1359 461
rect 1305 411 1359 427
rect 1823 461 1877 477
rect 1823 441 1833 461
rect 1130 377 1160 411
rect 1324 377 1354 411
rect 1796 427 1833 441
rect 1867 427 1877 461
rect 1796 411 1877 427
rect 1971 461 2025 477
rect 1971 427 1981 461
rect 2015 427 2025 461
rect 1971 411 2025 427
rect 2489 461 2543 477
rect 2489 441 2499 461
rect 1796 377 1826 411
rect 1990 377 2020 411
rect 2462 427 2499 441
rect 2533 427 2543 461
rect 2462 411 2543 427
rect 2637 461 2691 477
rect 2637 427 2647 461
rect 2681 427 2691 461
rect 2637 411 2691 427
rect 3155 461 3209 477
rect 3155 441 3165 461
rect 2462 377 2492 411
rect 2656 377 2686 411
rect 3128 427 3165 441
rect 3199 427 3209 461
rect 3128 411 3209 427
rect 3303 461 3357 477
rect 3303 427 3313 461
rect 3347 427 3357 461
rect 3303 411 3357 427
rect 3821 461 3875 477
rect 3821 441 3831 461
rect 3128 377 3158 411
rect 3322 377 3352 411
rect 3794 427 3831 441
rect 3865 427 3875 461
rect 3794 411 3875 427
rect 3969 461 4023 477
rect 3969 427 3979 461
rect 4013 427 4023 461
rect 3969 411 4023 427
rect 4487 461 4541 477
rect 4487 441 4497 461
rect 3794 377 3824 411
rect 3988 377 4018 411
rect 4439 427 4497 441
rect 4531 427 4541 461
rect 4439 411 4541 427
rect 4709 461 4763 477
rect 4709 427 4719 461
rect 4753 441 4763 461
rect 4931 461 4985 477
rect 4753 427 4769 441
rect 4709 411 4769 427
rect 4931 427 4941 461
rect 4975 427 4985 461
rect 4931 411 4985 427
rect 5449 461 5503 477
rect 5449 441 5459 461
rect 4439 379 4469 411
rect 4739 379 4769 411
rect 4941 379 4971 411
rect 5422 427 5459 441
rect 5493 427 5503 461
rect 5422 411 5503 427
rect 5597 461 5651 477
rect 5597 427 5607 461
rect 5641 427 5651 461
rect 5597 411 5651 427
rect 6115 461 6169 477
rect 6115 441 6125 461
rect 5422 377 5452 411
rect 5616 377 5646 411
rect 6088 427 6125 441
rect 6159 427 6169 461
rect 6088 411 6169 427
rect 6263 461 6317 477
rect 6263 427 6273 461
rect 6307 427 6317 461
rect 6263 411 6317 427
rect 6781 461 6835 477
rect 6781 441 6791 461
rect 6088 377 6118 411
rect 6282 377 6312 411
rect 6754 427 6791 441
rect 6825 427 6835 461
rect 6754 411 6835 427
rect 6929 461 6983 477
rect 6929 427 6939 461
rect 6973 427 6983 461
rect 6929 411 6983 427
rect 7447 461 7501 477
rect 7447 441 7457 461
rect 6754 377 6784 411
rect 6948 377 6978 411
rect 7420 427 7457 441
rect 7491 427 7501 461
rect 7420 411 7501 427
rect 7595 461 7649 477
rect 7595 427 7605 461
rect 7639 427 7649 461
rect 7595 411 7649 427
rect 8113 461 8167 477
rect 8113 441 8123 461
rect 7420 377 7450 411
rect 7614 377 7644 411
rect 8086 427 8123 441
rect 8157 427 8167 461
rect 8086 411 8167 427
rect 8261 461 8315 477
rect 8261 427 8271 461
rect 8305 427 8315 461
rect 8261 411 8315 427
rect 8779 461 8833 477
rect 8779 441 8789 461
rect 8086 377 8116 411
rect 8280 377 8310 411
rect 8731 427 8789 441
rect 8823 427 8833 461
rect 8731 411 8833 427
rect 9001 461 9055 477
rect 9001 427 9011 461
rect 9045 441 9055 461
rect 9223 461 9277 477
rect 9045 427 9061 441
rect 9001 411 9061 427
rect 9223 427 9233 461
rect 9267 427 9277 461
rect 9223 411 9277 427
rect 9741 461 9795 477
rect 9741 441 9751 461
rect 8731 379 8761 411
rect 9031 379 9061 411
rect 9233 379 9263 411
rect 9714 427 9751 441
rect 9785 427 9795 461
rect 9714 411 9795 427
rect 9889 461 9943 477
rect 9889 427 9899 461
rect 9933 427 9943 461
rect 9889 411 9943 427
rect 10407 461 10461 477
rect 10407 441 10417 461
rect 9714 377 9744 411
rect 9908 377 9938 411
rect 10380 427 10417 441
rect 10451 427 10461 461
rect 10380 411 10461 427
rect 10555 461 10609 477
rect 10555 427 10565 461
rect 10599 427 10609 461
rect 10555 411 10609 427
rect 11073 461 11127 477
rect 11073 441 11083 461
rect 10380 377 10410 411
rect 10574 377 10604 411
rect 11046 427 11083 441
rect 11117 427 11127 461
rect 11046 411 11127 427
rect 11221 461 11275 477
rect 11221 427 11231 461
rect 11265 427 11275 461
rect 11221 411 11275 427
rect 11739 461 11793 477
rect 11739 441 11749 461
rect 11046 377 11076 411
rect 11240 377 11270 411
rect 11712 427 11749 441
rect 11783 427 11793 461
rect 11712 411 11793 427
rect 11887 461 11941 477
rect 11887 427 11897 461
rect 11931 427 11941 461
rect 11887 411 11941 427
rect 12405 461 12459 477
rect 12405 441 12415 461
rect 11712 377 11742 411
rect 11906 377 11936 411
rect 12378 427 12415 441
rect 12449 427 12459 461
rect 12378 411 12459 427
rect 12553 461 12607 477
rect 12553 427 12563 461
rect 12597 427 12607 461
rect 12553 411 12607 427
rect 12378 377 12408 411
rect 12572 377 12602 411
rect 12997 461 13051 477
rect 12997 427 13007 461
rect 13041 441 13051 461
rect 13219 461 13273 477
rect 13041 427 13074 441
rect 12997 411 13074 427
rect 13219 427 13229 461
rect 13263 427 13273 461
rect 13219 411 13273 427
rect 13737 461 13791 477
rect 13737 441 13747 461
rect 13044 377 13074 411
rect 13238 377 13268 411
rect 13710 427 13747 441
rect 13781 427 13791 461
rect 14033 461 14087 477
rect 14033 441 14043 461
rect 13710 411 13791 427
rect 14010 427 14043 441
rect 14077 427 14087 461
rect 14010 411 14087 427
rect 13710 377 13740 411
rect 14010 377 14040 411
rect 14329 461 14383 477
rect 14329 427 14339 461
rect 14373 441 14383 461
rect 14551 461 14605 477
rect 14373 427 14406 441
rect 14329 411 14406 427
rect 14551 427 14561 461
rect 14595 427 14605 461
rect 14551 411 14605 427
rect 14376 377 14406 411
rect 14570 377 14600 411
<< polycont >>
rect 205 969 239 1003
rect 427 969 461 1003
rect 649 969 683 1003
rect 1167 969 1201 1003
rect 1321 969 1355 1003
rect 1833 969 1867 1003
rect 1987 969 2021 1003
rect 2499 969 2533 1003
rect 2653 969 2687 1003
rect 3165 969 3199 1003
rect 3319 969 3353 1003
rect 3831 969 3865 1003
rect 3985 969 4019 1003
rect 4497 969 4531 1003
rect 4719 969 4753 1003
rect 4941 969 4975 1003
rect 5459 969 5493 1003
rect 5613 969 5647 1003
rect 6125 969 6159 1003
rect 6279 969 6313 1003
rect 6791 969 6825 1003
rect 6945 969 6979 1003
rect 7457 969 7491 1003
rect 7611 969 7645 1003
rect 8123 969 8157 1003
rect 8277 969 8311 1003
rect 8789 969 8823 1003
rect 9011 969 9045 1003
rect 9233 969 9267 1003
rect 9751 969 9785 1003
rect 9905 969 9939 1003
rect 10417 969 10451 1003
rect 10571 969 10605 1003
rect 11083 969 11117 1003
rect 11237 969 11271 1003
rect 11749 969 11783 1003
rect 11903 969 11937 1003
rect 12415 969 12449 1003
rect 12569 969 12603 1003
rect 13007 970 13041 1004
rect 13237 970 13271 1004
rect 13747 970 13781 1004
rect 14043 970 14077 1004
rect 14339 970 14373 1004
rect 14565 970 14599 1004
rect 205 427 239 461
rect 427 427 461 461
rect 649 427 683 461
rect 1167 427 1201 461
rect 1315 427 1349 461
rect 1833 427 1867 461
rect 1981 427 2015 461
rect 2499 427 2533 461
rect 2647 427 2681 461
rect 3165 427 3199 461
rect 3313 427 3347 461
rect 3831 427 3865 461
rect 3979 427 4013 461
rect 4497 427 4531 461
rect 4719 427 4753 461
rect 4941 427 4975 461
rect 5459 427 5493 461
rect 5607 427 5641 461
rect 6125 427 6159 461
rect 6273 427 6307 461
rect 6791 427 6825 461
rect 6939 427 6973 461
rect 7457 427 7491 461
rect 7605 427 7639 461
rect 8123 427 8157 461
rect 8271 427 8305 461
rect 8789 427 8823 461
rect 9011 427 9045 461
rect 9233 427 9267 461
rect 9751 427 9785 461
rect 9899 427 9933 461
rect 10417 427 10451 461
rect 10565 427 10599 461
rect 11083 427 11117 461
rect 11231 427 11265 461
rect 11749 427 11783 461
rect 11897 427 11931 461
rect 12415 427 12449 461
rect 12563 427 12597 461
rect 13007 427 13041 461
rect 13229 427 13263 461
rect 13747 427 13781 461
rect 14043 427 14077 461
rect 14339 427 14373 461
rect 14561 427 14595 461
<< locali >>
rect -31 1539 14905 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 343 1539
rect 377 1505 415 1539
rect 449 1505 513 1539
rect 547 1505 585 1539
rect 619 1505 657 1539
rect 691 1505 729 1539
rect 763 1505 801 1539
rect 835 1505 873 1539
rect 907 1505 1017 1539
rect 1051 1505 1089 1539
rect 1123 1505 1161 1539
rect 1195 1505 1233 1539
rect 1267 1505 1323 1539
rect 1357 1505 1395 1539
rect 1429 1505 1467 1539
rect 1501 1505 1539 1539
rect 1573 1505 1683 1539
rect 1717 1505 1755 1539
rect 1789 1505 1827 1539
rect 1861 1505 1899 1539
rect 1933 1505 1989 1539
rect 2023 1505 2061 1539
rect 2095 1505 2133 1539
rect 2167 1505 2205 1539
rect 2239 1505 2349 1539
rect 2383 1505 2421 1539
rect 2455 1505 2493 1539
rect 2527 1505 2565 1539
rect 2599 1505 2655 1539
rect 2689 1505 2727 1539
rect 2761 1505 2799 1539
rect 2833 1505 2871 1539
rect 2905 1505 3015 1539
rect 3049 1505 3087 1539
rect 3121 1505 3159 1539
rect 3193 1505 3231 1539
rect 3265 1505 3321 1539
rect 3355 1505 3393 1539
rect 3427 1505 3465 1539
rect 3499 1505 3537 1539
rect 3571 1505 3681 1539
rect 3715 1505 3753 1539
rect 3787 1505 3825 1539
rect 3859 1505 3897 1539
rect 3931 1505 3987 1539
rect 4021 1505 4059 1539
rect 4093 1505 4131 1539
rect 4165 1505 4203 1539
rect 4237 1505 4347 1539
rect 4381 1505 4419 1539
rect 4453 1505 4491 1539
rect 4525 1505 4563 1539
rect 4597 1505 4635 1539
rect 4669 1505 4707 1539
rect 4741 1505 4805 1539
rect 4839 1505 4877 1539
rect 4911 1505 4949 1539
rect 4983 1505 5021 1539
rect 5055 1505 5093 1539
rect 5127 1505 5165 1539
rect 5199 1505 5309 1539
rect 5343 1505 5381 1539
rect 5415 1505 5453 1539
rect 5487 1505 5525 1539
rect 5559 1505 5615 1539
rect 5649 1505 5687 1539
rect 5721 1505 5759 1539
rect 5793 1505 5831 1539
rect 5865 1505 5975 1539
rect 6009 1505 6047 1539
rect 6081 1505 6119 1539
rect 6153 1505 6191 1539
rect 6225 1505 6281 1539
rect 6315 1505 6353 1539
rect 6387 1505 6425 1539
rect 6459 1505 6497 1539
rect 6531 1505 6641 1539
rect 6675 1505 6713 1539
rect 6747 1505 6785 1539
rect 6819 1505 6857 1539
rect 6891 1505 6947 1539
rect 6981 1505 7019 1539
rect 7053 1505 7091 1539
rect 7125 1505 7163 1539
rect 7197 1505 7307 1539
rect 7341 1505 7379 1539
rect 7413 1505 7451 1539
rect 7485 1505 7523 1539
rect 7557 1505 7613 1539
rect 7647 1505 7685 1539
rect 7719 1505 7757 1539
rect 7791 1505 7829 1539
rect 7863 1505 7973 1539
rect 8007 1505 8045 1539
rect 8079 1505 8117 1539
rect 8151 1505 8189 1539
rect 8223 1505 8279 1539
rect 8313 1505 8351 1539
rect 8385 1505 8423 1539
rect 8457 1505 8495 1539
rect 8529 1505 8639 1539
rect 8673 1505 8711 1539
rect 8745 1505 8783 1539
rect 8817 1505 8855 1539
rect 8889 1505 8927 1539
rect 8961 1505 8999 1539
rect 9033 1505 9097 1539
rect 9131 1505 9169 1539
rect 9203 1505 9241 1539
rect 9275 1505 9313 1539
rect 9347 1505 9385 1539
rect 9419 1505 9457 1539
rect 9491 1505 9601 1539
rect 9635 1505 9673 1539
rect 9707 1505 9745 1539
rect 9779 1505 9817 1539
rect 9851 1505 9907 1539
rect 9941 1505 9979 1539
rect 10013 1505 10051 1539
rect 10085 1505 10123 1539
rect 10157 1505 10267 1539
rect 10301 1505 10339 1539
rect 10373 1505 10411 1539
rect 10445 1505 10483 1539
rect 10517 1505 10573 1539
rect 10607 1505 10645 1539
rect 10679 1505 10717 1539
rect 10751 1505 10789 1539
rect 10823 1505 10933 1539
rect 10967 1505 11005 1539
rect 11039 1505 11077 1539
rect 11111 1505 11149 1539
rect 11183 1505 11239 1539
rect 11273 1505 11311 1539
rect 11345 1505 11383 1539
rect 11417 1505 11455 1539
rect 11489 1505 11599 1539
rect 11633 1505 11671 1539
rect 11705 1505 11743 1539
rect 11777 1505 11815 1539
rect 11849 1505 11905 1539
rect 11939 1505 11977 1539
rect 12011 1505 12049 1539
rect 12083 1505 12121 1539
rect 12155 1505 12265 1539
rect 12299 1505 12337 1539
rect 12371 1505 12409 1539
rect 12443 1505 12481 1539
rect 12515 1505 12571 1539
rect 12605 1505 12643 1539
rect 12677 1505 12715 1539
rect 12749 1505 12787 1539
rect 12821 1505 12931 1539
rect 12965 1505 13003 1539
rect 13037 1505 13075 1539
rect 13109 1505 13147 1539
rect 13181 1505 13237 1539
rect 13271 1505 13309 1539
rect 13343 1505 13381 1539
rect 13415 1505 13453 1539
rect 13487 1505 13597 1539
rect 13631 1505 13669 1539
rect 13703 1505 13741 1539
rect 13775 1505 13813 1539
rect 13847 1505 13903 1539
rect 13937 1505 13975 1539
rect 14009 1505 14047 1539
rect 14081 1505 14119 1539
rect 14153 1505 14263 1539
rect 14297 1505 14335 1539
rect 14369 1505 14407 1539
rect 14441 1505 14479 1539
rect 14513 1505 14569 1539
rect 14603 1505 14641 1539
rect 14675 1505 14713 1539
rect 14747 1505 14785 1539
rect 14819 1505 14905 1539
rect -31 1492 14905 1505
rect -31 1470 31 1492
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect 201 1412 235 1492
rect 201 1344 235 1378
rect 201 1276 235 1310
rect 201 1208 235 1242
rect 201 1139 235 1174
rect 201 1089 235 1105
rect 289 1412 323 1450
rect 289 1344 323 1378
rect 289 1276 323 1310
rect 289 1208 323 1242
rect 289 1139 323 1174
rect 377 1412 411 1492
rect 377 1344 411 1378
rect 377 1276 411 1310
rect 377 1208 411 1242
rect 377 1157 411 1174
rect 465 1412 499 1450
rect 465 1344 499 1378
rect 465 1276 499 1310
rect 465 1208 499 1242
rect 289 1094 323 1105
rect 465 1139 499 1174
rect 553 1412 587 1492
rect 553 1344 587 1378
rect 553 1276 587 1310
rect 553 1208 587 1242
rect 553 1157 587 1174
rect 641 1412 675 1450
rect 641 1344 675 1378
rect 641 1276 675 1310
rect 641 1208 675 1242
rect 465 1094 499 1105
rect 641 1139 675 1174
rect 729 1412 763 1492
rect 729 1344 763 1378
rect 729 1276 763 1310
rect 729 1208 763 1242
rect 729 1157 763 1174
rect 931 1470 993 1492
rect 931 1436 945 1470
rect 979 1436 993 1470
rect 931 1398 993 1436
rect 931 1364 945 1398
rect 979 1364 993 1398
rect 931 1326 993 1364
rect 931 1292 945 1326
rect 979 1292 993 1326
rect 931 1254 993 1292
rect 931 1220 945 1254
rect 979 1220 993 1254
rect 931 1182 993 1220
rect 641 1094 675 1105
rect 931 1148 945 1182
rect 979 1148 993 1182
rect 931 1110 993 1148
rect -31 1038 31 1076
rect 289 1060 831 1094
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect -31 868 31 932
rect 205 1003 239 1019
rect 205 905 239 969
rect -31 546 31 572
rect -31 512 -17 546
rect 17 512 31 546
rect -31 474 31 512
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect 205 461 239 871
rect 205 411 239 427
rect 427 1003 461 1019
rect 427 461 461 945
rect 427 411 461 427
rect 649 1003 683 1019
rect 649 757 683 969
rect 649 461 683 723
rect 649 411 683 427
rect 797 831 831 1060
rect 931 1076 945 1110
rect 979 1076 993 1110
rect 931 1038 993 1076
rect 1103 1412 1137 1492
rect 1103 1344 1137 1378
rect 1103 1276 1137 1310
rect 1103 1208 1137 1242
rect 1103 1139 1137 1174
rect 1103 1073 1137 1105
rect 1191 1412 1225 1450
rect 1191 1344 1225 1378
rect 1191 1276 1225 1310
rect 1191 1208 1225 1242
rect 1191 1139 1225 1174
rect 1279 1412 1313 1492
rect 1279 1344 1313 1378
rect 1279 1276 1313 1310
rect 1279 1208 1313 1242
rect 1279 1157 1313 1174
rect 1367 1412 1401 1450
rect 1367 1344 1401 1378
rect 1367 1276 1401 1310
rect 1367 1208 1401 1242
rect 1191 1103 1225 1105
rect 1367 1139 1401 1174
rect 1455 1412 1489 1492
rect 1455 1344 1489 1378
rect 1455 1276 1489 1310
rect 1455 1208 1489 1242
rect 1455 1157 1489 1174
rect 1597 1470 1659 1492
rect 1597 1436 1611 1470
rect 1645 1436 1659 1470
rect 1597 1398 1659 1436
rect 1597 1364 1611 1398
rect 1645 1364 1659 1398
rect 1597 1326 1659 1364
rect 1597 1292 1611 1326
rect 1645 1292 1659 1326
rect 1597 1254 1659 1292
rect 1597 1220 1611 1254
rect 1645 1220 1659 1254
rect 1597 1182 1659 1220
rect 1367 1103 1401 1105
rect 1597 1148 1611 1182
rect 1645 1148 1659 1182
rect 1597 1110 1659 1148
rect 1191 1069 1497 1103
rect 931 1004 945 1038
rect 979 1004 993 1038
rect 931 966 993 1004
rect 931 932 945 966
rect 979 932 993 966
rect 931 868 993 932
rect 1167 1003 1201 1019
rect 1321 1003 1355 1019
rect -31 368 -17 402
rect 17 368 31 402
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect 101 363 135 379
rect 295 363 329 379
rect 489 363 523 379
rect 135 329 198 363
rect 232 329 295 363
rect 329 329 392 363
rect 426 329 489 363
rect 101 291 135 329
rect 101 223 135 257
rect 295 291 329 329
rect 489 313 523 329
rect 603 363 637 379
rect 797 378 831 797
rect 1167 831 1201 969
rect 603 291 637 329
rect 101 153 135 189
rect 101 103 135 119
rect 198 238 232 254
rect -31 62 31 80
rect 198 62 232 204
rect 295 223 329 257
rect 393 244 427 260
rect 603 244 637 257
rect 427 223 637 244
rect 427 210 603 223
rect 393 194 427 210
rect 295 153 329 189
rect 700 344 831 378
rect 931 546 993 572
rect 931 512 945 546
rect 979 512 993 546
rect 931 474 993 512
rect 931 440 945 474
rect 979 440 993 474
rect 931 402 993 440
rect 1167 461 1201 797
rect 1167 411 1201 427
rect 1315 969 1321 988
rect 1315 953 1355 969
rect 1315 461 1349 953
rect 1315 411 1349 427
rect 1463 757 1497 1069
rect 1597 1076 1611 1110
rect 1645 1076 1659 1110
rect 1597 1038 1659 1076
rect 1769 1412 1803 1492
rect 1769 1344 1803 1378
rect 1769 1276 1803 1310
rect 1769 1208 1803 1242
rect 1769 1139 1803 1174
rect 1769 1073 1803 1105
rect 1857 1412 1891 1450
rect 1857 1344 1891 1378
rect 1857 1276 1891 1310
rect 1857 1208 1891 1242
rect 1857 1139 1891 1174
rect 1945 1412 1979 1492
rect 1945 1344 1979 1378
rect 1945 1276 1979 1310
rect 1945 1208 1979 1242
rect 1945 1157 1979 1174
rect 2033 1412 2067 1450
rect 2033 1344 2067 1378
rect 2033 1276 2067 1310
rect 2033 1208 2067 1242
rect 1857 1103 1891 1105
rect 2033 1139 2067 1174
rect 2121 1412 2155 1492
rect 2121 1344 2155 1378
rect 2121 1276 2155 1310
rect 2121 1208 2155 1242
rect 2121 1157 2155 1174
rect 2263 1470 2325 1492
rect 2263 1436 2277 1470
rect 2311 1436 2325 1470
rect 2263 1398 2325 1436
rect 2263 1364 2277 1398
rect 2311 1364 2325 1398
rect 2263 1326 2325 1364
rect 2263 1292 2277 1326
rect 2311 1292 2325 1326
rect 2263 1254 2325 1292
rect 2263 1220 2277 1254
rect 2311 1220 2325 1254
rect 2263 1182 2325 1220
rect 2033 1103 2067 1105
rect 2263 1148 2277 1182
rect 2311 1148 2325 1182
rect 2263 1110 2325 1148
rect 1857 1069 2163 1103
rect 1597 1004 1611 1038
rect 1645 1004 1659 1038
rect 1597 966 1659 1004
rect 1597 932 1611 966
rect 1645 932 1659 966
rect 1597 868 1659 932
rect 1833 1003 1867 1019
rect 1987 1003 2021 1019
rect 931 368 945 402
rect 979 368 993 402
rect 700 247 734 344
rect 931 330 993 368
rect 700 197 734 213
rect 797 291 831 307
rect 797 223 831 257
rect 489 153 523 169
rect 329 119 392 153
rect 426 119 489 153
rect 295 103 329 119
rect 489 103 523 119
rect 603 153 637 189
rect 797 153 831 189
rect 637 119 700 153
rect 734 119 797 153
rect 603 103 637 119
rect 797 103 831 119
rect 931 296 945 330
rect 979 296 993 330
rect 931 258 993 296
rect 931 224 945 258
rect 979 224 993 258
rect 931 186 993 224
rect 931 152 945 186
rect 979 152 993 186
rect 931 114 993 152
rect 931 80 945 114
rect 979 80 993 114
rect 1084 361 1118 377
rect 1278 361 1312 377
rect 1463 376 1497 723
rect 1833 757 1867 969
rect 1118 327 1181 361
rect 1215 327 1278 361
rect 1084 289 1118 327
rect 1084 221 1118 255
rect 1278 289 1312 327
rect 1084 151 1118 187
rect 1084 101 1118 117
rect 1181 236 1215 252
rect 931 62 993 80
rect 1181 62 1215 202
rect 1278 221 1312 255
rect 1375 342 1497 376
rect 1597 546 1659 572
rect 1597 512 1611 546
rect 1645 512 1659 546
rect 1597 474 1659 512
rect 1597 440 1611 474
rect 1645 440 1659 474
rect 1597 402 1659 440
rect 1833 461 1867 723
rect 1833 411 1867 427
rect 1981 969 1987 988
rect 1981 953 2021 969
rect 1981 905 2015 953
rect 1981 461 2015 871
rect 1981 411 2015 427
rect 2129 757 2163 1069
rect 2263 1076 2277 1110
rect 2311 1076 2325 1110
rect 2263 1038 2325 1076
rect 2435 1412 2469 1492
rect 2435 1344 2469 1378
rect 2435 1276 2469 1310
rect 2435 1208 2469 1242
rect 2435 1139 2469 1174
rect 2435 1073 2469 1105
rect 2523 1412 2557 1450
rect 2523 1344 2557 1378
rect 2523 1276 2557 1310
rect 2523 1208 2557 1242
rect 2523 1139 2557 1174
rect 2611 1412 2645 1492
rect 2611 1344 2645 1378
rect 2611 1276 2645 1310
rect 2611 1208 2645 1242
rect 2611 1157 2645 1174
rect 2699 1412 2733 1450
rect 2699 1344 2733 1378
rect 2699 1276 2733 1310
rect 2699 1208 2733 1242
rect 2523 1103 2557 1105
rect 2699 1139 2733 1174
rect 2787 1412 2821 1492
rect 2787 1344 2821 1378
rect 2787 1276 2821 1310
rect 2787 1208 2821 1242
rect 2787 1157 2821 1174
rect 2929 1470 2991 1492
rect 2929 1436 2943 1470
rect 2977 1436 2991 1470
rect 2929 1398 2991 1436
rect 2929 1364 2943 1398
rect 2977 1364 2991 1398
rect 2929 1326 2991 1364
rect 2929 1292 2943 1326
rect 2977 1292 2991 1326
rect 2929 1254 2991 1292
rect 2929 1220 2943 1254
rect 2977 1220 2991 1254
rect 2929 1182 2991 1220
rect 2699 1103 2733 1105
rect 2929 1148 2943 1182
rect 2977 1148 2991 1182
rect 2929 1110 2991 1148
rect 2523 1069 2829 1103
rect 2263 1004 2277 1038
rect 2311 1004 2325 1038
rect 2263 966 2325 1004
rect 2263 932 2277 966
rect 2311 932 2325 966
rect 2263 868 2325 932
rect 2499 1003 2533 1019
rect 2653 1003 2687 1019
rect 1597 368 1611 402
rect 1645 368 1659 402
rect 1375 245 1409 342
rect 1597 330 1659 368
rect 1375 195 1409 211
rect 1472 289 1506 305
rect 1472 221 1506 255
rect 1278 151 1312 187
rect 1472 151 1506 187
rect 1312 117 1375 151
rect 1409 117 1472 151
rect 1278 101 1312 117
rect 1472 101 1506 117
rect 1597 296 1611 330
rect 1645 296 1659 330
rect 1597 258 1659 296
rect 1597 224 1611 258
rect 1645 224 1659 258
rect 1597 186 1659 224
rect 1597 152 1611 186
rect 1645 152 1659 186
rect 1597 114 1659 152
rect 1597 80 1611 114
rect 1645 80 1659 114
rect 1750 361 1784 377
rect 1944 361 1978 377
rect 2129 376 2163 723
rect 2499 757 2533 969
rect 1784 327 1847 361
rect 1881 327 1944 361
rect 1750 289 1784 327
rect 1750 221 1784 255
rect 1944 289 1978 327
rect 1750 151 1784 187
rect 1750 101 1784 117
rect 1847 236 1881 252
rect 1597 62 1659 80
rect 1847 62 1881 202
rect 1944 221 1978 255
rect 2041 342 2163 376
rect 2263 546 2325 572
rect 2263 512 2277 546
rect 2311 512 2325 546
rect 2263 474 2325 512
rect 2263 440 2277 474
rect 2311 440 2325 474
rect 2263 402 2325 440
rect 2499 461 2533 723
rect 2499 411 2533 427
rect 2647 979 2653 995
rect 2681 953 2687 969
rect 2647 461 2681 945
rect 2647 411 2681 427
rect 2795 905 2829 1069
rect 2263 368 2277 402
rect 2311 368 2325 402
rect 2041 245 2075 342
rect 2263 330 2325 368
rect 2041 195 2075 211
rect 2138 289 2172 305
rect 2138 221 2172 255
rect 1944 151 1978 187
rect 2138 151 2172 187
rect 1978 117 2041 151
rect 2075 117 2138 151
rect 1944 101 1978 117
rect 2138 101 2172 117
rect 2263 296 2277 330
rect 2311 296 2325 330
rect 2263 258 2325 296
rect 2263 224 2277 258
rect 2311 224 2325 258
rect 2263 186 2325 224
rect 2263 152 2277 186
rect 2311 152 2325 186
rect 2263 114 2325 152
rect 2263 80 2277 114
rect 2311 80 2325 114
rect 2416 361 2450 377
rect 2610 361 2644 377
rect 2795 376 2829 871
rect 2929 1076 2943 1110
rect 2977 1076 2991 1110
rect 2929 1038 2991 1076
rect 3101 1412 3135 1492
rect 3101 1344 3135 1378
rect 3101 1276 3135 1310
rect 3101 1208 3135 1242
rect 3101 1139 3135 1174
rect 3101 1073 3135 1105
rect 3189 1412 3223 1450
rect 3189 1344 3223 1378
rect 3189 1276 3223 1310
rect 3189 1208 3223 1242
rect 3189 1139 3223 1174
rect 3277 1412 3311 1492
rect 3277 1344 3311 1378
rect 3277 1276 3311 1310
rect 3277 1208 3311 1242
rect 3277 1157 3311 1174
rect 3365 1412 3399 1450
rect 3365 1344 3399 1378
rect 3365 1276 3399 1310
rect 3365 1208 3399 1242
rect 3189 1103 3223 1105
rect 3365 1139 3399 1174
rect 3453 1412 3487 1492
rect 3453 1344 3487 1378
rect 3453 1276 3487 1310
rect 3453 1208 3487 1242
rect 3453 1157 3487 1174
rect 3595 1470 3657 1492
rect 3595 1436 3609 1470
rect 3643 1436 3657 1470
rect 3595 1398 3657 1436
rect 3595 1364 3609 1398
rect 3643 1364 3657 1398
rect 3595 1326 3657 1364
rect 3595 1292 3609 1326
rect 3643 1292 3657 1326
rect 3595 1254 3657 1292
rect 3595 1220 3609 1254
rect 3643 1220 3657 1254
rect 3595 1182 3657 1220
rect 3365 1103 3399 1105
rect 3595 1148 3609 1182
rect 3643 1148 3657 1182
rect 3595 1110 3657 1148
rect 3189 1069 3495 1103
rect 2929 1004 2943 1038
rect 2977 1004 2991 1038
rect 2929 966 2991 1004
rect 2929 932 2943 966
rect 2977 932 2991 966
rect 2929 868 2991 932
rect 3165 1003 3199 1019
rect 3319 1003 3353 1019
rect 3165 831 3199 969
rect 2450 327 2513 361
rect 2547 327 2610 361
rect 2416 289 2450 327
rect 2416 221 2450 255
rect 2610 289 2644 327
rect 2416 151 2450 187
rect 2416 101 2450 117
rect 2513 236 2547 252
rect 2263 62 2325 80
rect 2513 62 2547 202
rect 2610 221 2644 255
rect 2707 342 2829 376
rect 2929 546 2991 572
rect 2929 512 2943 546
rect 2977 512 2991 546
rect 2929 474 2991 512
rect 2929 440 2943 474
rect 2977 440 2991 474
rect 2929 402 2991 440
rect 3165 461 3199 797
rect 3165 411 3199 427
rect 3313 969 3319 988
rect 3313 953 3353 969
rect 3313 683 3347 953
rect 3313 461 3347 649
rect 3313 411 3347 427
rect 3461 831 3495 1069
rect 3595 1076 3609 1110
rect 3643 1076 3657 1110
rect 3595 1038 3657 1076
rect 3767 1412 3801 1492
rect 3767 1344 3801 1378
rect 3767 1276 3801 1310
rect 3767 1208 3801 1242
rect 3767 1139 3801 1174
rect 3767 1073 3801 1105
rect 3855 1412 3889 1450
rect 3855 1344 3889 1378
rect 3855 1276 3889 1310
rect 3855 1208 3889 1242
rect 3855 1139 3889 1174
rect 3943 1412 3977 1492
rect 3943 1344 3977 1378
rect 3943 1276 3977 1310
rect 3943 1208 3977 1242
rect 3943 1157 3977 1174
rect 4031 1412 4065 1450
rect 4031 1344 4065 1378
rect 4031 1276 4065 1310
rect 4031 1208 4065 1242
rect 3855 1103 3889 1105
rect 4031 1139 4065 1174
rect 4119 1412 4153 1492
rect 4119 1344 4153 1378
rect 4119 1276 4153 1310
rect 4119 1208 4153 1242
rect 4119 1157 4153 1174
rect 4261 1470 4323 1492
rect 4261 1436 4275 1470
rect 4309 1436 4323 1470
rect 4261 1398 4323 1436
rect 4261 1364 4275 1398
rect 4309 1364 4323 1398
rect 4261 1326 4323 1364
rect 4261 1292 4275 1326
rect 4309 1292 4323 1326
rect 4261 1254 4323 1292
rect 4261 1220 4275 1254
rect 4309 1220 4323 1254
rect 4261 1182 4323 1220
rect 4031 1103 4065 1105
rect 4261 1148 4275 1182
rect 4309 1148 4323 1182
rect 4261 1110 4323 1148
rect 3855 1069 4161 1103
rect 3595 1004 3609 1038
rect 3643 1004 3657 1038
rect 3595 966 3657 1004
rect 3595 932 3609 966
rect 3643 932 3657 966
rect 3595 868 3657 932
rect 3831 1003 3865 1019
rect 3985 1003 4019 1019
rect 2929 368 2943 402
rect 2977 368 2991 402
rect 2707 245 2741 342
rect 2929 330 2991 368
rect 2707 195 2741 211
rect 2804 289 2838 305
rect 2804 221 2838 255
rect 2610 151 2644 187
rect 2804 151 2838 187
rect 2644 117 2707 151
rect 2741 117 2804 151
rect 2610 101 2644 117
rect 2804 101 2838 117
rect 2929 296 2943 330
rect 2977 296 2991 330
rect 2929 258 2991 296
rect 2929 224 2943 258
rect 2977 224 2991 258
rect 2929 186 2991 224
rect 2929 152 2943 186
rect 2977 152 2991 186
rect 2929 114 2991 152
rect 2929 80 2943 114
rect 2977 80 2991 114
rect 3082 361 3116 377
rect 3276 361 3310 377
rect 3461 376 3495 797
rect 3831 831 3865 969
rect 3116 327 3179 361
rect 3213 327 3276 361
rect 3082 289 3116 327
rect 3082 221 3116 255
rect 3276 289 3310 327
rect 3082 151 3116 187
rect 3082 101 3116 117
rect 3179 236 3213 252
rect 2929 62 2991 80
rect 3179 62 3213 202
rect 3276 221 3310 255
rect 3373 342 3495 376
rect 3595 546 3657 572
rect 3595 512 3609 546
rect 3643 512 3657 546
rect 3595 474 3657 512
rect 3595 440 3609 474
rect 3643 440 3657 474
rect 3595 402 3657 440
rect 3831 461 3865 797
rect 3831 411 3865 427
rect 3979 969 3985 988
rect 3979 953 4019 969
rect 3979 905 4013 953
rect 3979 461 4013 871
rect 3979 411 4013 427
rect 4127 683 4161 1069
rect 4261 1076 4275 1110
rect 4309 1076 4323 1110
rect 4493 1412 4527 1492
rect 4493 1344 4527 1378
rect 4493 1276 4527 1310
rect 4493 1208 4527 1242
rect 4493 1139 4527 1174
rect 4493 1089 4527 1105
rect 4581 1412 4615 1450
rect 4581 1344 4615 1378
rect 4581 1276 4615 1310
rect 4581 1208 4615 1242
rect 4581 1139 4615 1174
rect 4669 1412 4703 1492
rect 4669 1344 4703 1378
rect 4669 1276 4703 1310
rect 4669 1208 4703 1242
rect 4669 1157 4703 1174
rect 4757 1412 4791 1450
rect 4757 1344 4791 1378
rect 4757 1276 4791 1310
rect 4757 1208 4791 1242
rect 4581 1094 4615 1105
rect 4757 1139 4791 1174
rect 4845 1412 4879 1492
rect 4845 1344 4879 1378
rect 4845 1276 4879 1310
rect 4845 1208 4879 1242
rect 4845 1157 4879 1174
rect 4933 1412 4967 1450
rect 4933 1344 4967 1378
rect 4933 1276 4967 1310
rect 4933 1208 4967 1242
rect 4757 1094 4791 1105
rect 4933 1139 4967 1174
rect 5021 1412 5055 1492
rect 5021 1344 5055 1378
rect 5021 1276 5055 1310
rect 5021 1208 5055 1242
rect 5021 1157 5055 1174
rect 5223 1470 5285 1492
rect 5223 1436 5237 1470
rect 5271 1436 5285 1470
rect 5223 1398 5285 1436
rect 5223 1364 5237 1398
rect 5271 1364 5285 1398
rect 5223 1326 5285 1364
rect 5223 1292 5237 1326
rect 5271 1292 5285 1326
rect 5223 1254 5285 1292
rect 5223 1220 5237 1254
rect 5271 1220 5285 1254
rect 5223 1182 5285 1220
rect 4933 1094 4967 1105
rect 5223 1148 5237 1182
rect 5271 1148 5285 1182
rect 5223 1110 5285 1148
rect 4261 1038 4323 1076
rect 4581 1060 5123 1094
rect 4261 1004 4275 1038
rect 4309 1004 4323 1038
rect 4261 966 4323 1004
rect 4261 932 4275 966
rect 4309 932 4323 966
rect 4261 868 4323 932
rect 4497 1003 4531 1019
rect 4497 905 4531 969
rect 3595 368 3609 402
rect 3643 368 3657 402
rect 3373 245 3407 342
rect 3595 330 3657 368
rect 3373 195 3407 211
rect 3470 289 3504 305
rect 3470 221 3504 255
rect 3276 151 3310 187
rect 3470 151 3504 187
rect 3310 117 3373 151
rect 3407 117 3470 151
rect 3276 101 3310 117
rect 3470 101 3504 117
rect 3595 296 3609 330
rect 3643 296 3657 330
rect 3595 258 3657 296
rect 3595 224 3609 258
rect 3643 224 3657 258
rect 3595 186 3657 224
rect 3595 152 3609 186
rect 3643 152 3657 186
rect 3595 114 3657 152
rect 3595 80 3609 114
rect 3643 80 3657 114
rect 3748 361 3782 377
rect 3942 361 3976 377
rect 4127 376 4161 649
rect 3782 327 3845 361
rect 3879 327 3942 361
rect 3748 289 3782 327
rect 3748 221 3782 255
rect 3942 289 3976 327
rect 3748 151 3782 187
rect 3748 101 3782 117
rect 3845 236 3879 252
rect 3595 62 3657 80
rect 3845 62 3879 202
rect 3942 221 3976 255
rect 4039 342 4161 376
rect 4261 546 4323 572
rect 4261 512 4275 546
rect 4309 512 4323 546
rect 4261 474 4323 512
rect 4261 440 4275 474
rect 4309 440 4323 474
rect 4261 402 4323 440
rect 4497 461 4531 871
rect 4497 411 4531 427
rect 4719 1003 4753 1019
rect 4719 461 4753 945
rect 4719 411 4753 427
rect 4941 1003 4975 1019
rect 4941 757 4975 969
rect 4941 461 4975 723
rect 4941 411 4975 427
rect 5089 831 5123 1060
rect 5223 1076 5237 1110
rect 5271 1076 5285 1110
rect 5223 1038 5285 1076
rect 5395 1412 5429 1492
rect 5395 1344 5429 1378
rect 5395 1276 5429 1310
rect 5395 1208 5429 1242
rect 5395 1139 5429 1174
rect 5395 1073 5429 1105
rect 5483 1412 5517 1450
rect 5483 1344 5517 1378
rect 5483 1276 5517 1310
rect 5483 1208 5517 1242
rect 5483 1139 5517 1174
rect 5571 1412 5605 1492
rect 5571 1344 5605 1378
rect 5571 1276 5605 1310
rect 5571 1208 5605 1242
rect 5571 1157 5605 1174
rect 5659 1412 5693 1450
rect 5659 1344 5693 1378
rect 5659 1276 5693 1310
rect 5659 1208 5693 1242
rect 5483 1103 5517 1105
rect 5659 1139 5693 1174
rect 5747 1412 5781 1492
rect 5747 1344 5781 1378
rect 5747 1276 5781 1310
rect 5747 1208 5781 1242
rect 5747 1157 5781 1174
rect 5889 1470 5951 1492
rect 5889 1436 5903 1470
rect 5937 1436 5951 1470
rect 5889 1398 5951 1436
rect 5889 1364 5903 1398
rect 5937 1364 5951 1398
rect 5889 1326 5951 1364
rect 5889 1292 5903 1326
rect 5937 1292 5951 1326
rect 5889 1254 5951 1292
rect 5889 1220 5903 1254
rect 5937 1220 5951 1254
rect 5889 1182 5951 1220
rect 5659 1103 5693 1105
rect 5889 1148 5903 1182
rect 5937 1148 5951 1182
rect 5889 1110 5951 1148
rect 5483 1069 5789 1103
rect 5223 1004 5237 1038
rect 5271 1004 5285 1038
rect 5223 966 5285 1004
rect 5223 932 5237 966
rect 5271 932 5285 966
rect 5223 868 5285 932
rect 5459 1003 5493 1019
rect 5613 1003 5647 1019
rect 4261 368 4275 402
rect 4309 368 4323 402
rect 4039 245 4073 342
rect 4261 330 4323 368
rect 4039 195 4073 211
rect 4136 289 4170 305
rect 4136 221 4170 255
rect 3942 151 3976 187
rect 4136 151 4170 187
rect 3976 117 4039 151
rect 4073 117 4136 151
rect 3942 101 3976 117
rect 4136 101 4170 117
rect 4261 296 4275 330
rect 4309 296 4323 330
rect 4261 258 4323 296
rect 4261 224 4275 258
rect 4309 224 4323 258
rect 4261 186 4323 224
rect 4261 152 4275 186
rect 4309 152 4323 186
rect 4261 114 4323 152
rect 4261 80 4275 114
rect 4309 80 4323 114
rect 4393 363 4427 379
rect 4587 363 4621 379
rect 4781 363 4815 379
rect 4427 329 4490 363
rect 4524 329 4587 363
rect 4621 329 4684 363
rect 4718 329 4781 363
rect 4393 291 4427 329
rect 4393 223 4427 257
rect 4587 291 4621 329
rect 4781 313 4815 329
rect 4895 363 4929 379
rect 5089 378 5123 797
rect 5459 831 5493 969
rect 4895 291 4929 329
rect 4393 153 4427 189
rect 4393 103 4427 119
rect 4490 238 4524 254
rect 4261 62 4323 80
rect 4490 62 4524 204
rect 4587 223 4621 257
rect 4685 244 4719 260
rect 4895 244 4929 257
rect 4719 223 4929 244
rect 4719 210 4895 223
rect 4685 194 4719 210
rect 4587 153 4621 189
rect 4992 344 5123 378
rect 5223 546 5285 572
rect 5223 512 5237 546
rect 5271 512 5285 546
rect 5223 474 5285 512
rect 5223 440 5237 474
rect 5271 440 5285 474
rect 5223 402 5285 440
rect 5459 461 5493 797
rect 5459 411 5493 427
rect 5607 969 5613 988
rect 5607 953 5647 969
rect 5607 461 5641 953
rect 5607 411 5641 427
rect 5755 757 5789 1069
rect 5889 1076 5903 1110
rect 5937 1076 5951 1110
rect 5889 1038 5951 1076
rect 6061 1412 6095 1492
rect 6061 1344 6095 1378
rect 6061 1276 6095 1310
rect 6061 1208 6095 1242
rect 6061 1139 6095 1174
rect 6061 1073 6095 1105
rect 6149 1412 6183 1450
rect 6149 1344 6183 1378
rect 6149 1276 6183 1310
rect 6149 1208 6183 1242
rect 6149 1139 6183 1174
rect 6237 1412 6271 1492
rect 6237 1344 6271 1378
rect 6237 1276 6271 1310
rect 6237 1208 6271 1242
rect 6237 1157 6271 1174
rect 6325 1412 6359 1450
rect 6325 1344 6359 1378
rect 6325 1276 6359 1310
rect 6325 1208 6359 1242
rect 6149 1103 6183 1105
rect 6325 1139 6359 1174
rect 6413 1412 6447 1492
rect 6413 1344 6447 1378
rect 6413 1276 6447 1310
rect 6413 1208 6447 1242
rect 6413 1157 6447 1174
rect 6555 1470 6617 1492
rect 6555 1436 6569 1470
rect 6603 1436 6617 1470
rect 6555 1398 6617 1436
rect 6555 1364 6569 1398
rect 6603 1364 6617 1398
rect 6555 1326 6617 1364
rect 6555 1292 6569 1326
rect 6603 1292 6617 1326
rect 6555 1254 6617 1292
rect 6555 1220 6569 1254
rect 6603 1220 6617 1254
rect 6555 1182 6617 1220
rect 6325 1103 6359 1105
rect 6555 1148 6569 1182
rect 6603 1148 6617 1182
rect 6555 1110 6617 1148
rect 6149 1069 6455 1103
rect 5889 1004 5903 1038
rect 5937 1004 5951 1038
rect 5889 966 5951 1004
rect 5889 932 5903 966
rect 5937 932 5951 966
rect 5889 868 5951 932
rect 6125 1003 6159 1019
rect 6279 1003 6313 1019
rect 5223 368 5237 402
rect 5271 368 5285 402
rect 4992 247 5026 344
rect 5223 330 5285 368
rect 4992 197 5026 213
rect 5089 291 5123 307
rect 5089 223 5123 257
rect 4781 153 4815 169
rect 4621 119 4684 153
rect 4718 119 4781 153
rect 4587 103 4621 119
rect 4781 103 4815 119
rect 4895 153 4929 189
rect 5089 153 5123 189
rect 4929 119 4992 153
rect 5026 119 5089 153
rect 4895 103 4929 119
rect 5089 103 5123 119
rect 5223 296 5237 330
rect 5271 296 5285 330
rect 5223 258 5285 296
rect 5223 224 5237 258
rect 5271 224 5285 258
rect 5223 186 5285 224
rect 5223 152 5237 186
rect 5271 152 5285 186
rect 5223 114 5285 152
rect 5223 80 5237 114
rect 5271 80 5285 114
rect 5376 361 5410 377
rect 5570 361 5604 377
rect 5755 376 5789 723
rect 6125 757 6159 969
rect 5410 327 5473 361
rect 5507 327 5570 361
rect 5376 289 5410 327
rect 5376 221 5410 255
rect 5570 289 5604 327
rect 5376 151 5410 187
rect 5376 101 5410 117
rect 5473 236 5507 252
rect 5223 62 5285 80
rect 5473 62 5507 202
rect 5570 221 5604 255
rect 5667 342 5789 376
rect 5889 546 5951 572
rect 5889 512 5903 546
rect 5937 512 5951 546
rect 5889 474 5951 512
rect 5889 440 5903 474
rect 5937 440 5951 474
rect 5889 402 5951 440
rect 6125 461 6159 723
rect 6125 411 6159 427
rect 6273 969 6279 988
rect 6273 953 6313 969
rect 6273 905 6307 953
rect 6273 461 6307 871
rect 6273 411 6307 427
rect 6421 757 6455 1069
rect 6555 1076 6569 1110
rect 6603 1076 6617 1110
rect 6555 1038 6617 1076
rect 6727 1412 6761 1492
rect 6727 1344 6761 1378
rect 6727 1276 6761 1310
rect 6727 1208 6761 1242
rect 6727 1139 6761 1174
rect 6727 1073 6761 1105
rect 6815 1412 6849 1450
rect 6815 1344 6849 1378
rect 6815 1276 6849 1310
rect 6815 1208 6849 1242
rect 6815 1139 6849 1174
rect 6903 1412 6937 1492
rect 6903 1344 6937 1378
rect 6903 1276 6937 1310
rect 6903 1208 6937 1242
rect 6903 1157 6937 1174
rect 6991 1412 7025 1450
rect 6991 1344 7025 1378
rect 6991 1276 7025 1310
rect 6991 1208 7025 1242
rect 6815 1103 6849 1105
rect 6991 1139 7025 1174
rect 7079 1412 7113 1492
rect 7079 1344 7113 1378
rect 7079 1276 7113 1310
rect 7079 1208 7113 1242
rect 7079 1157 7113 1174
rect 7221 1470 7283 1492
rect 7221 1436 7235 1470
rect 7269 1436 7283 1470
rect 7221 1398 7283 1436
rect 7221 1364 7235 1398
rect 7269 1364 7283 1398
rect 7221 1326 7283 1364
rect 7221 1292 7235 1326
rect 7269 1292 7283 1326
rect 7221 1254 7283 1292
rect 7221 1220 7235 1254
rect 7269 1220 7283 1254
rect 7221 1182 7283 1220
rect 6991 1103 7025 1105
rect 7221 1148 7235 1182
rect 7269 1148 7283 1182
rect 7221 1110 7283 1148
rect 6815 1069 7121 1103
rect 6555 1004 6569 1038
rect 6603 1004 6617 1038
rect 6555 966 6617 1004
rect 6555 932 6569 966
rect 6603 932 6617 966
rect 6555 868 6617 932
rect 6791 1003 6825 1019
rect 6945 1003 6979 1019
rect 5889 368 5903 402
rect 5937 368 5951 402
rect 5667 245 5701 342
rect 5889 330 5951 368
rect 5667 195 5701 211
rect 5764 289 5798 305
rect 5764 221 5798 255
rect 5570 151 5604 187
rect 5764 151 5798 187
rect 5604 117 5667 151
rect 5701 117 5764 151
rect 5570 101 5604 117
rect 5764 101 5798 117
rect 5889 296 5903 330
rect 5937 296 5951 330
rect 5889 258 5951 296
rect 5889 224 5903 258
rect 5937 224 5951 258
rect 5889 186 5951 224
rect 5889 152 5903 186
rect 5937 152 5951 186
rect 5889 114 5951 152
rect 5889 80 5903 114
rect 5937 80 5951 114
rect 6042 361 6076 377
rect 6236 361 6270 377
rect 6421 376 6455 723
rect 6791 757 6825 969
rect 6076 327 6139 361
rect 6173 327 6236 361
rect 6042 289 6076 327
rect 6042 221 6076 255
rect 6236 289 6270 327
rect 6042 151 6076 187
rect 6042 101 6076 117
rect 6139 236 6173 252
rect 5889 62 5951 80
rect 6139 62 6173 202
rect 6236 221 6270 255
rect 6333 342 6455 376
rect 6555 546 6617 572
rect 6555 512 6569 546
rect 6603 512 6617 546
rect 6555 474 6617 512
rect 6555 440 6569 474
rect 6603 440 6617 474
rect 6555 402 6617 440
rect 6791 461 6825 723
rect 6791 411 6825 427
rect 6939 979 6945 995
rect 6973 953 6979 969
rect 6939 461 6973 945
rect 6939 411 6973 427
rect 7087 905 7121 1069
rect 6555 368 6569 402
rect 6603 368 6617 402
rect 6333 245 6367 342
rect 6555 330 6617 368
rect 6333 195 6367 211
rect 6430 289 6464 305
rect 6430 221 6464 255
rect 6236 151 6270 187
rect 6430 151 6464 187
rect 6270 117 6333 151
rect 6367 117 6430 151
rect 6236 101 6270 117
rect 6430 101 6464 117
rect 6555 296 6569 330
rect 6603 296 6617 330
rect 6555 258 6617 296
rect 6555 224 6569 258
rect 6603 224 6617 258
rect 6555 186 6617 224
rect 6555 152 6569 186
rect 6603 152 6617 186
rect 6555 114 6617 152
rect 6555 80 6569 114
rect 6603 80 6617 114
rect 6708 361 6742 377
rect 6902 361 6936 377
rect 7087 376 7121 871
rect 7221 1076 7235 1110
rect 7269 1076 7283 1110
rect 7221 1038 7283 1076
rect 7393 1412 7427 1492
rect 7393 1344 7427 1378
rect 7393 1276 7427 1310
rect 7393 1208 7427 1242
rect 7393 1139 7427 1174
rect 7393 1073 7427 1105
rect 7481 1412 7515 1450
rect 7481 1344 7515 1378
rect 7481 1276 7515 1310
rect 7481 1208 7515 1242
rect 7481 1139 7515 1174
rect 7569 1412 7603 1492
rect 7569 1344 7603 1378
rect 7569 1276 7603 1310
rect 7569 1208 7603 1242
rect 7569 1157 7603 1174
rect 7657 1412 7691 1450
rect 7657 1344 7691 1378
rect 7657 1276 7691 1310
rect 7657 1208 7691 1242
rect 7481 1103 7515 1105
rect 7657 1139 7691 1174
rect 7745 1412 7779 1492
rect 7745 1344 7779 1378
rect 7745 1276 7779 1310
rect 7745 1208 7779 1242
rect 7745 1157 7779 1174
rect 7887 1470 7949 1492
rect 7887 1436 7901 1470
rect 7935 1436 7949 1470
rect 7887 1398 7949 1436
rect 7887 1364 7901 1398
rect 7935 1364 7949 1398
rect 7887 1326 7949 1364
rect 7887 1292 7901 1326
rect 7935 1292 7949 1326
rect 7887 1254 7949 1292
rect 7887 1220 7901 1254
rect 7935 1220 7949 1254
rect 7887 1182 7949 1220
rect 7657 1103 7691 1105
rect 7887 1148 7901 1182
rect 7935 1148 7949 1182
rect 7887 1110 7949 1148
rect 7481 1069 7787 1103
rect 7221 1004 7235 1038
rect 7269 1004 7283 1038
rect 7221 966 7283 1004
rect 7221 932 7235 966
rect 7269 932 7283 966
rect 7221 868 7283 932
rect 7457 1003 7491 1019
rect 7611 1003 7645 1019
rect 7457 831 7491 969
rect 6742 327 6805 361
rect 6839 327 6902 361
rect 6708 289 6742 327
rect 6708 221 6742 255
rect 6902 289 6936 327
rect 6708 151 6742 187
rect 6708 101 6742 117
rect 6805 236 6839 252
rect 6555 62 6617 80
rect 6805 62 6839 202
rect 6902 221 6936 255
rect 6999 342 7121 376
rect 7221 546 7283 572
rect 7221 512 7235 546
rect 7269 512 7283 546
rect 7221 474 7283 512
rect 7221 440 7235 474
rect 7269 440 7283 474
rect 7221 402 7283 440
rect 7457 461 7491 797
rect 7457 411 7491 427
rect 7605 969 7611 988
rect 7605 953 7645 969
rect 7605 535 7639 953
rect 7605 461 7639 501
rect 7605 411 7639 427
rect 7753 831 7787 1069
rect 7887 1076 7901 1110
rect 7935 1076 7949 1110
rect 7887 1038 7949 1076
rect 8059 1412 8093 1492
rect 8059 1344 8093 1378
rect 8059 1276 8093 1310
rect 8059 1208 8093 1242
rect 8059 1139 8093 1174
rect 8059 1073 8093 1105
rect 8147 1412 8181 1450
rect 8147 1344 8181 1378
rect 8147 1276 8181 1310
rect 8147 1208 8181 1242
rect 8147 1139 8181 1174
rect 8235 1412 8269 1492
rect 8235 1344 8269 1378
rect 8235 1276 8269 1310
rect 8235 1208 8269 1242
rect 8235 1157 8269 1174
rect 8323 1412 8357 1450
rect 8323 1344 8357 1378
rect 8323 1276 8357 1310
rect 8323 1208 8357 1242
rect 8147 1103 8181 1105
rect 8323 1139 8357 1174
rect 8411 1412 8445 1492
rect 8411 1344 8445 1378
rect 8411 1276 8445 1310
rect 8411 1208 8445 1242
rect 8411 1157 8445 1174
rect 8553 1470 8615 1492
rect 8553 1436 8567 1470
rect 8601 1436 8615 1470
rect 8553 1398 8615 1436
rect 8553 1364 8567 1398
rect 8601 1364 8615 1398
rect 8553 1326 8615 1364
rect 8553 1292 8567 1326
rect 8601 1292 8615 1326
rect 8553 1254 8615 1292
rect 8553 1220 8567 1254
rect 8601 1220 8615 1254
rect 8553 1182 8615 1220
rect 8323 1103 8357 1105
rect 8553 1148 8567 1182
rect 8601 1148 8615 1182
rect 8553 1110 8615 1148
rect 8147 1069 8453 1103
rect 7887 1004 7901 1038
rect 7935 1004 7949 1038
rect 7887 966 7949 1004
rect 7887 932 7901 966
rect 7935 932 7949 966
rect 7887 868 7949 932
rect 8123 1003 8157 1019
rect 8277 1003 8311 1019
rect 7221 368 7235 402
rect 7269 368 7283 402
rect 6999 245 7033 342
rect 7221 330 7283 368
rect 6999 195 7033 211
rect 7096 289 7130 305
rect 7096 221 7130 255
rect 6902 151 6936 187
rect 7096 151 7130 187
rect 6936 117 6999 151
rect 7033 117 7096 151
rect 6902 101 6936 117
rect 7096 101 7130 117
rect 7221 296 7235 330
rect 7269 296 7283 330
rect 7221 258 7283 296
rect 7221 224 7235 258
rect 7269 224 7283 258
rect 7221 186 7283 224
rect 7221 152 7235 186
rect 7269 152 7283 186
rect 7221 114 7283 152
rect 7221 80 7235 114
rect 7269 80 7283 114
rect 7374 361 7408 377
rect 7568 361 7602 377
rect 7753 376 7787 797
rect 8123 831 8157 969
rect 7408 327 7471 361
rect 7505 327 7568 361
rect 7374 289 7408 327
rect 7374 221 7408 255
rect 7568 289 7602 327
rect 7374 151 7408 187
rect 7374 101 7408 117
rect 7471 236 7505 252
rect 7221 62 7283 80
rect 7471 62 7505 202
rect 7568 221 7602 255
rect 7665 342 7787 376
rect 7887 546 7949 572
rect 7887 512 7901 546
rect 7935 512 7949 546
rect 7887 474 7949 512
rect 7887 440 7901 474
rect 7935 440 7949 474
rect 7887 402 7949 440
rect 8123 461 8157 797
rect 8123 411 8157 427
rect 8271 969 8277 988
rect 8271 953 8311 969
rect 8271 905 8305 953
rect 8271 461 8305 871
rect 8271 411 8305 427
rect 8419 535 8453 1069
rect 8553 1076 8567 1110
rect 8601 1076 8615 1110
rect 8785 1412 8819 1492
rect 8785 1344 8819 1378
rect 8785 1276 8819 1310
rect 8785 1208 8819 1242
rect 8785 1139 8819 1174
rect 8785 1089 8819 1105
rect 8873 1412 8907 1450
rect 8873 1344 8907 1378
rect 8873 1276 8907 1310
rect 8873 1208 8907 1242
rect 8873 1139 8907 1174
rect 8961 1412 8995 1492
rect 8961 1344 8995 1378
rect 8961 1276 8995 1310
rect 8961 1208 8995 1242
rect 8961 1157 8995 1174
rect 9049 1412 9083 1450
rect 9049 1344 9083 1378
rect 9049 1276 9083 1310
rect 9049 1208 9083 1242
rect 8873 1094 8907 1105
rect 9049 1139 9083 1174
rect 9137 1412 9171 1492
rect 9137 1344 9171 1378
rect 9137 1276 9171 1310
rect 9137 1208 9171 1242
rect 9137 1157 9171 1174
rect 9225 1412 9259 1450
rect 9225 1344 9259 1378
rect 9225 1276 9259 1310
rect 9225 1208 9259 1242
rect 9049 1094 9083 1105
rect 9225 1139 9259 1174
rect 9313 1412 9347 1492
rect 9313 1344 9347 1378
rect 9313 1276 9347 1310
rect 9313 1208 9347 1242
rect 9313 1157 9347 1174
rect 9515 1470 9577 1492
rect 9515 1436 9529 1470
rect 9563 1436 9577 1470
rect 9515 1398 9577 1436
rect 9515 1364 9529 1398
rect 9563 1364 9577 1398
rect 9515 1326 9577 1364
rect 9515 1292 9529 1326
rect 9563 1292 9577 1326
rect 9515 1254 9577 1292
rect 9515 1220 9529 1254
rect 9563 1220 9577 1254
rect 9515 1182 9577 1220
rect 9225 1094 9259 1105
rect 9515 1148 9529 1182
rect 9563 1148 9577 1182
rect 9515 1110 9577 1148
rect 8553 1038 8615 1076
rect 8873 1060 9415 1094
rect 8553 1004 8567 1038
rect 8601 1004 8615 1038
rect 8553 966 8615 1004
rect 8553 932 8567 966
rect 8601 932 8615 966
rect 8553 868 8615 932
rect 8789 1003 8823 1019
rect 8789 905 8823 969
rect 7887 368 7901 402
rect 7935 368 7949 402
rect 7665 245 7699 342
rect 7887 330 7949 368
rect 7665 195 7699 211
rect 7762 289 7796 305
rect 7762 221 7796 255
rect 7568 151 7602 187
rect 7762 151 7796 187
rect 7602 117 7665 151
rect 7699 117 7762 151
rect 7568 101 7602 117
rect 7762 101 7796 117
rect 7887 296 7901 330
rect 7935 296 7949 330
rect 7887 258 7949 296
rect 7887 224 7901 258
rect 7935 224 7949 258
rect 7887 186 7949 224
rect 7887 152 7901 186
rect 7935 152 7949 186
rect 7887 114 7949 152
rect 7887 80 7901 114
rect 7935 80 7949 114
rect 8040 361 8074 377
rect 8234 361 8268 377
rect 8419 376 8453 501
rect 8074 327 8137 361
rect 8171 327 8234 361
rect 8040 289 8074 327
rect 8040 221 8074 255
rect 8234 289 8268 327
rect 8040 151 8074 187
rect 8040 101 8074 117
rect 8137 236 8171 252
rect 7887 62 7949 80
rect 8137 62 8171 202
rect 8234 221 8268 255
rect 8331 342 8453 376
rect 8553 546 8615 572
rect 8553 512 8567 546
rect 8601 512 8615 546
rect 8553 474 8615 512
rect 8553 440 8567 474
rect 8601 440 8615 474
rect 8553 402 8615 440
rect 8789 461 8823 871
rect 8789 411 8823 427
rect 9011 1003 9045 1019
rect 9011 461 9045 945
rect 9011 411 9045 427
rect 9233 1003 9267 1019
rect 9233 757 9267 969
rect 9233 461 9267 723
rect 9233 411 9267 427
rect 9381 831 9415 1060
rect 9515 1076 9529 1110
rect 9563 1076 9577 1110
rect 9515 1038 9577 1076
rect 9687 1412 9721 1492
rect 9687 1344 9721 1378
rect 9687 1276 9721 1310
rect 9687 1208 9721 1242
rect 9687 1139 9721 1174
rect 9687 1073 9721 1105
rect 9775 1412 9809 1450
rect 9775 1344 9809 1378
rect 9775 1276 9809 1310
rect 9775 1208 9809 1242
rect 9775 1139 9809 1174
rect 9863 1412 9897 1492
rect 9863 1344 9897 1378
rect 9863 1276 9897 1310
rect 9863 1208 9897 1242
rect 9863 1157 9897 1174
rect 9951 1412 9985 1450
rect 9951 1344 9985 1378
rect 9951 1276 9985 1310
rect 9951 1208 9985 1242
rect 9775 1103 9809 1105
rect 9951 1139 9985 1174
rect 10039 1412 10073 1492
rect 10039 1344 10073 1378
rect 10039 1276 10073 1310
rect 10039 1208 10073 1242
rect 10039 1157 10073 1174
rect 10181 1470 10243 1492
rect 10181 1436 10195 1470
rect 10229 1436 10243 1470
rect 10181 1398 10243 1436
rect 10181 1364 10195 1398
rect 10229 1364 10243 1398
rect 10181 1326 10243 1364
rect 10181 1292 10195 1326
rect 10229 1292 10243 1326
rect 10181 1254 10243 1292
rect 10181 1220 10195 1254
rect 10229 1220 10243 1254
rect 10181 1182 10243 1220
rect 9951 1103 9985 1105
rect 10181 1148 10195 1182
rect 10229 1148 10243 1182
rect 10181 1110 10243 1148
rect 9775 1069 10081 1103
rect 9515 1004 9529 1038
rect 9563 1004 9577 1038
rect 9515 966 9577 1004
rect 9515 932 9529 966
rect 9563 932 9577 966
rect 9515 868 9577 932
rect 9751 1003 9785 1019
rect 9905 1003 9939 1019
rect 8553 368 8567 402
rect 8601 368 8615 402
rect 8331 245 8365 342
rect 8553 330 8615 368
rect 8331 195 8365 211
rect 8428 289 8462 305
rect 8428 221 8462 255
rect 8234 151 8268 187
rect 8428 151 8462 187
rect 8268 117 8331 151
rect 8365 117 8428 151
rect 8234 101 8268 117
rect 8428 101 8462 117
rect 8553 296 8567 330
rect 8601 296 8615 330
rect 8553 258 8615 296
rect 8553 224 8567 258
rect 8601 224 8615 258
rect 8553 186 8615 224
rect 8553 152 8567 186
rect 8601 152 8615 186
rect 8553 114 8615 152
rect 8553 80 8567 114
rect 8601 80 8615 114
rect 8685 363 8719 379
rect 8879 363 8913 379
rect 9073 363 9107 379
rect 8719 329 8782 363
rect 8816 329 8879 363
rect 8913 329 8976 363
rect 9010 329 9073 363
rect 8685 291 8719 329
rect 8685 223 8719 257
rect 8879 291 8913 329
rect 9073 313 9107 329
rect 9187 363 9221 379
rect 9381 378 9415 797
rect 9751 831 9785 969
rect 9187 291 9221 329
rect 8685 153 8719 189
rect 8685 103 8719 119
rect 8782 238 8816 254
rect 8553 62 8615 80
rect 8782 62 8816 204
rect 8879 223 8913 257
rect 8977 244 9011 260
rect 9187 244 9221 257
rect 9011 223 9221 244
rect 9011 210 9187 223
rect 8977 194 9011 210
rect 8879 153 8913 189
rect 9284 344 9415 378
rect 9515 546 9577 572
rect 9515 512 9529 546
rect 9563 512 9577 546
rect 9515 474 9577 512
rect 9515 440 9529 474
rect 9563 440 9577 474
rect 9515 402 9577 440
rect 9751 461 9785 797
rect 9751 411 9785 427
rect 9899 969 9905 988
rect 9899 953 9939 969
rect 9899 461 9933 953
rect 9899 411 9933 427
rect 10047 757 10081 1069
rect 10181 1076 10195 1110
rect 10229 1076 10243 1110
rect 10181 1038 10243 1076
rect 10353 1412 10387 1492
rect 10353 1344 10387 1378
rect 10353 1276 10387 1310
rect 10353 1208 10387 1242
rect 10353 1139 10387 1174
rect 10353 1073 10387 1105
rect 10441 1412 10475 1450
rect 10441 1344 10475 1378
rect 10441 1276 10475 1310
rect 10441 1208 10475 1242
rect 10441 1139 10475 1174
rect 10529 1412 10563 1492
rect 10529 1344 10563 1378
rect 10529 1276 10563 1310
rect 10529 1208 10563 1242
rect 10529 1157 10563 1174
rect 10617 1412 10651 1450
rect 10617 1344 10651 1378
rect 10617 1276 10651 1310
rect 10617 1208 10651 1242
rect 10441 1103 10475 1105
rect 10617 1139 10651 1174
rect 10705 1412 10739 1492
rect 10705 1344 10739 1378
rect 10705 1276 10739 1310
rect 10705 1208 10739 1242
rect 10705 1157 10739 1174
rect 10847 1470 10909 1492
rect 10847 1436 10861 1470
rect 10895 1436 10909 1470
rect 10847 1398 10909 1436
rect 10847 1364 10861 1398
rect 10895 1364 10909 1398
rect 10847 1326 10909 1364
rect 10847 1292 10861 1326
rect 10895 1292 10909 1326
rect 10847 1254 10909 1292
rect 10847 1220 10861 1254
rect 10895 1220 10909 1254
rect 10847 1182 10909 1220
rect 10617 1103 10651 1105
rect 10847 1148 10861 1182
rect 10895 1148 10909 1182
rect 10847 1110 10909 1148
rect 10441 1069 10747 1103
rect 10181 1004 10195 1038
rect 10229 1004 10243 1038
rect 10181 966 10243 1004
rect 10181 932 10195 966
rect 10229 932 10243 966
rect 10181 868 10243 932
rect 10417 1003 10451 1019
rect 10571 1003 10605 1019
rect 9515 368 9529 402
rect 9563 368 9577 402
rect 9284 247 9318 344
rect 9515 330 9577 368
rect 9284 197 9318 213
rect 9381 291 9415 307
rect 9381 223 9415 257
rect 9073 153 9107 169
rect 8913 119 8976 153
rect 9010 119 9073 153
rect 8879 103 8913 119
rect 9073 103 9107 119
rect 9187 153 9221 189
rect 9381 153 9415 189
rect 9221 119 9284 153
rect 9318 119 9381 153
rect 9187 103 9221 119
rect 9381 103 9415 119
rect 9515 296 9529 330
rect 9563 296 9577 330
rect 9515 258 9577 296
rect 9515 224 9529 258
rect 9563 224 9577 258
rect 9515 186 9577 224
rect 9515 152 9529 186
rect 9563 152 9577 186
rect 9515 114 9577 152
rect 9515 80 9529 114
rect 9563 80 9577 114
rect 9668 361 9702 377
rect 9862 361 9896 377
rect 10047 376 10081 723
rect 10417 757 10451 969
rect 9702 327 9765 361
rect 9799 327 9862 361
rect 9668 289 9702 327
rect 9668 221 9702 255
rect 9862 289 9896 327
rect 9668 151 9702 187
rect 9668 101 9702 117
rect 9765 236 9799 252
rect 9515 62 9577 80
rect 9765 62 9799 202
rect 9862 221 9896 255
rect 9959 342 10081 376
rect 10181 546 10243 572
rect 10181 512 10195 546
rect 10229 512 10243 546
rect 10181 474 10243 512
rect 10181 440 10195 474
rect 10229 440 10243 474
rect 10181 402 10243 440
rect 10417 461 10451 723
rect 10417 411 10451 427
rect 10565 969 10571 988
rect 10565 953 10605 969
rect 10565 905 10599 953
rect 10565 461 10599 871
rect 10565 411 10599 427
rect 10713 757 10747 1069
rect 10847 1076 10861 1110
rect 10895 1076 10909 1110
rect 10847 1038 10909 1076
rect 11019 1412 11053 1492
rect 11019 1344 11053 1378
rect 11019 1276 11053 1310
rect 11019 1208 11053 1242
rect 11019 1139 11053 1174
rect 11019 1073 11053 1105
rect 11107 1412 11141 1450
rect 11107 1344 11141 1378
rect 11107 1276 11141 1310
rect 11107 1208 11141 1242
rect 11107 1139 11141 1174
rect 11195 1412 11229 1492
rect 11195 1344 11229 1378
rect 11195 1276 11229 1310
rect 11195 1208 11229 1242
rect 11195 1157 11229 1174
rect 11283 1412 11317 1450
rect 11283 1344 11317 1378
rect 11283 1276 11317 1310
rect 11283 1208 11317 1242
rect 11107 1103 11141 1105
rect 11283 1139 11317 1174
rect 11371 1412 11405 1492
rect 11371 1344 11405 1378
rect 11371 1276 11405 1310
rect 11371 1208 11405 1242
rect 11371 1157 11405 1174
rect 11513 1470 11575 1492
rect 11513 1436 11527 1470
rect 11561 1436 11575 1470
rect 11513 1398 11575 1436
rect 11513 1364 11527 1398
rect 11561 1364 11575 1398
rect 11513 1326 11575 1364
rect 11513 1292 11527 1326
rect 11561 1292 11575 1326
rect 11513 1254 11575 1292
rect 11513 1220 11527 1254
rect 11561 1220 11575 1254
rect 11513 1182 11575 1220
rect 11283 1103 11317 1105
rect 11513 1148 11527 1182
rect 11561 1148 11575 1182
rect 11513 1110 11575 1148
rect 11107 1069 11413 1103
rect 10847 1004 10861 1038
rect 10895 1004 10909 1038
rect 10847 966 10909 1004
rect 10847 932 10861 966
rect 10895 932 10909 966
rect 10847 868 10909 932
rect 11083 1003 11117 1019
rect 11237 1003 11271 1019
rect 10181 368 10195 402
rect 10229 368 10243 402
rect 9959 245 9993 342
rect 10181 330 10243 368
rect 9959 195 9993 211
rect 10056 289 10090 305
rect 10056 221 10090 255
rect 9862 151 9896 187
rect 10056 151 10090 187
rect 9896 117 9959 151
rect 9993 117 10056 151
rect 9862 101 9896 117
rect 10056 101 10090 117
rect 10181 296 10195 330
rect 10229 296 10243 330
rect 10181 258 10243 296
rect 10181 224 10195 258
rect 10229 224 10243 258
rect 10181 186 10243 224
rect 10181 152 10195 186
rect 10229 152 10243 186
rect 10181 114 10243 152
rect 10181 80 10195 114
rect 10229 80 10243 114
rect 10334 361 10368 377
rect 10528 361 10562 377
rect 10713 376 10747 723
rect 11083 757 11117 969
rect 10368 327 10431 361
rect 10465 327 10528 361
rect 10334 289 10368 327
rect 10334 221 10368 255
rect 10528 289 10562 327
rect 10334 151 10368 187
rect 10334 101 10368 117
rect 10431 236 10465 252
rect 10181 62 10243 80
rect 10431 62 10465 202
rect 10528 221 10562 255
rect 10625 342 10747 376
rect 10847 546 10909 572
rect 10847 512 10861 546
rect 10895 512 10909 546
rect 10847 474 10909 512
rect 10847 440 10861 474
rect 10895 440 10909 474
rect 10847 402 10909 440
rect 11083 461 11117 723
rect 11083 411 11117 427
rect 11231 979 11237 995
rect 11265 953 11271 969
rect 11231 461 11265 945
rect 11231 411 11265 427
rect 11379 905 11413 1069
rect 10847 368 10861 402
rect 10895 368 10909 402
rect 10625 245 10659 342
rect 10847 330 10909 368
rect 10625 195 10659 211
rect 10722 289 10756 305
rect 10722 221 10756 255
rect 10528 151 10562 187
rect 10722 151 10756 187
rect 10562 117 10625 151
rect 10659 117 10722 151
rect 10528 101 10562 117
rect 10722 101 10756 117
rect 10847 296 10861 330
rect 10895 296 10909 330
rect 10847 258 10909 296
rect 10847 224 10861 258
rect 10895 224 10909 258
rect 10847 186 10909 224
rect 10847 152 10861 186
rect 10895 152 10909 186
rect 10847 114 10909 152
rect 10847 80 10861 114
rect 10895 80 10909 114
rect 11000 361 11034 377
rect 11194 361 11228 377
rect 11379 376 11413 871
rect 11513 1076 11527 1110
rect 11561 1076 11575 1110
rect 11513 1038 11575 1076
rect 11685 1412 11719 1492
rect 11685 1344 11719 1378
rect 11685 1276 11719 1310
rect 11685 1208 11719 1242
rect 11685 1139 11719 1174
rect 11685 1073 11719 1105
rect 11773 1412 11807 1450
rect 11773 1344 11807 1378
rect 11773 1276 11807 1310
rect 11773 1208 11807 1242
rect 11773 1139 11807 1174
rect 11861 1412 11895 1492
rect 11861 1344 11895 1378
rect 11861 1276 11895 1310
rect 11861 1208 11895 1242
rect 11861 1157 11895 1174
rect 11949 1412 11983 1450
rect 11949 1344 11983 1378
rect 11949 1276 11983 1310
rect 11949 1208 11983 1242
rect 11773 1103 11807 1105
rect 11949 1139 11983 1174
rect 12037 1412 12071 1492
rect 12037 1344 12071 1378
rect 12037 1276 12071 1310
rect 12037 1208 12071 1242
rect 12037 1157 12071 1174
rect 12179 1470 12241 1492
rect 12179 1436 12193 1470
rect 12227 1436 12241 1470
rect 12179 1398 12241 1436
rect 12179 1364 12193 1398
rect 12227 1364 12241 1398
rect 12179 1326 12241 1364
rect 12179 1292 12193 1326
rect 12227 1292 12241 1326
rect 12179 1254 12241 1292
rect 12179 1220 12193 1254
rect 12227 1220 12241 1254
rect 12179 1182 12241 1220
rect 11949 1103 11983 1105
rect 12179 1148 12193 1182
rect 12227 1148 12241 1182
rect 12179 1110 12241 1148
rect 11773 1069 12079 1103
rect 11513 1004 11527 1038
rect 11561 1004 11575 1038
rect 11513 966 11575 1004
rect 11513 932 11527 966
rect 11561 932 11575 966
rect 11513 868 11575 932
rect 11749 1003 11783 1019
rect 11903 1003 11937 1019
rect 11749 831 11783 969
rect 11034 327 11097 361
rect 11131 327 11194 361
rect 11000 289 11034 327
rect 11000 221 11034 255
rect 11194 289 11228 327
rect 11000 151 11034 187
rect 11000 101 11034 117
rect 11097 236 11131 252
rect 10847 62 10909 80
rect 11097 62 11131 202
rect 11194 221 11228 255
rect 11291 342 11413 376
rect 11513 546 11575 572
rect 11513 512 11527 546
rect 11561 512 11575 546
rect 11513 474 11575 512
rect 11513 440 11527 474
rect 11561 440 11575 474
rect 11513 402 11575 440
rect 11749 461 11783 797
rect 11749 411 11783 427
rect 11897 969 11903 988
rect 11897 953 11937 969
rect 12045 979 12079 1069
rect 11897 831 11931 953
rect 11897 461 11931 797
rect 11897 411 11931 427
rect 11513 368 11527 402
rect 11561 368 11575 402
rect 11291 245 11325 342
rect 11513 330 11575 368
rect 11291 195 11325 211
rect 11388 289 11422 305
rect 11388 221 11422 255
rect 11194 151 11228 187
rect 11388 151 11422 187
rect 11228 117 11291 151
rect 11325 117 11388 151
rect 11194 101 11228 117
rect 11388 101 11422 117
rect 11513 296 11527 330
rect 11561 296 11575 330
rect 11513 258 11575 296
rect 11513 224 11527 258
rect 11561 224 11575 258
rect 11513 186 11575 224
rect 11513 152 11527 186
rect 11561 152 11575 186
rect 11513 114 11575 152
rect 11513 80 11527 114
rect 11561 80 11575 114
rect 11666 361 11700 377
rect 11860 361 11894 377
rect 12045 376 12079 945
rect 12179 1076 12193 1110
rect 12227 1076 12241 1110
rect 12179 1038 12241 1076
rect 12351 1412 12385 1492
rect 12351 1344 12385 1378
rect 12351 1276 12385 1310
rect 12351 1208 12385 1242
rect 12351 1139 12385 1174
rect 12351 1073 12385 1105
rect 12439 1412 12473 1450
rect 12439 1344 12473 1378
rect 12439 1276 12473 1310
rect 12439 1208 12473 1242
rect 12439 1139 12473 1174
rect 12527 1412 12561 1492
rect 12527 1344 12561 1378
rect 12527 1276 12561 1310
rect 12527 1208 12561 1242
rect 12527 1157 12561 1174
rect 12615 1412 12649 1450
rect 12615 1344 12649 1378
rect 12615 1276 12649 1310
rect 12615 1208 12649 1242
rect 12439 1103 12473 1105
rect 12615 1139 12649 1174
rect 12703 1412 12737 1492
rect 12703 1344 12737 1378
rect 12703 1276 12737 1310
rect 12703 1208 12737 1242
rect 12703 1157 12737 1174
rect 12845 1470 12907 1492
rect 12845 1436 12859 1470
rect 12893 1436 12907 1470
rect 12845 1398 12907 1436
rect 12845 1364 12859 1398
rect 12893 1364 12907 1398
rect 12845 1326 12907 1364
rect 12845 1292 12859 1326
rect 12893 1292 12907 1326
rect 12845 1254 12907 1292
rect 12845 1220 12859 1254
rect 12893 1220 12907 1254
rect 12845 1182 12907 1220
rect 12615 1103 12649 1105
rect 12845 1148 12859 1182
rect 12893 1148 12907 1182
rect 12845 1110 12907 1148
rect 12439 1069 12745 1103
rect 12179 1004 12193 1038
rect 12227 1004 12241 1038
rect 12179 966 12241 1004
rect 12179 932 12193 966
rect 12227 932 12241 966
rect 12179 868 12241 932
rect 12415 1003 12449 1019
rect 12569 1003 12603 1019
rect 11700 327 11763 361
rect 11797 327 11860 361
rect 11666 289 11700 327
rect 11666 221 11700 255
rect 11860 289 11894 327
rect 11666 151 11700 187
rect 11666 101 11700 117
rect 11763 236 11797 252
rect 11513 62 11575 80
rect 11763 62 11797 202
rect 11860 221 11894 255
rect 11957 342 12079 376
rect 12179 546 12241 572
rect 12179 512 12193 546
rect 12227 512 12241 546
rect 12179 474 12241 512
rect 12179 440 12193 474
rect 12227 440 12241 474
rect 12179 402 12241 440
rect 12415 461 12449 945
rect 12415 411 12449 427
rect 12563 969 12569 988
rect 12563 953 12603 969
rect 12563 905 12597 953
rect 12563 461 12597 871
rect 12563 411 12597 427
rect 12711 831 12745 1069
rect 12845 1076 12859 1110
rect 12893 1076 12907 1110
rect 12845 1038 12907 1076
rect 13017 1411 13051 1492
rect 13017 1343 13051 1377
rect 13017 1275 13051 1309
rect 13017 1207 13051 1241
rect 13017 1139 13051 1173
rect 13017 1071 13051 1105
rect 13105 1411 13141 1445
rect 13193 1411 13227 1492
rect 13105 1343 13139 1377
rect 13105 1275 13139 1309
rect 13105 1207 13139 1241
rect 13105 1139 13139 1173
rect 13193 1343 13227 1377
rect 13193 1275 13227 1309
rect 13193 1207 13227 1241
rect 13193 1157 13227 1173
rect 13281 1411 13315 1445
rect 13281 1343 13315 1377
rect 13281 1275 13315 1309
rect 13281 1207 13315 1241
rect 13281 1105 13315 1173
rect 13105 1071 13281 1105
rect 13369 1411 13403 1492
rect 13369 1343 13403 1377
rect 13369 1275 13403 1309
rect 13369 1207 13403 1241
rect 13369 1139 13403 1173
rect 13369 1071 13403 1105
rect 13511 1470 13573 1492
rect 13511 1436 13525 1470
rect 13559 1436 13573 1470
rect 14177 1470 14239 1492
rect 13511 1398 13573 1436
rect 13511 1364 13525 1398
rect 13559 1364 13573 1398
rect 13511 1326 13573 1364
rect 13511 1292 13525 1326
rect 13559 1292 13573 1326
rect 13511 1254 13573 1292
rect 13511 1220 13525 1254
rect 13559 1220 13573 1254
rect 13511 1182 13573 1220
rect 13511 1148 13525 1182
rect 13559 1148 13573 1182
rect 13511 1110 13573 1148
rect 13511 1076 13525 1110
rect 13559 1076 13573 1110
rect 13281 1055 13315 1071
rect 12845 1004 12859 1038
rect 12893 1004 12907 1038
rect 13511 1038 13573 1076
rect 13681 1411 14067 1445
rect 13681 1343 13715 1377
rect 13681 1275 13715 1309
rect 13681 1207 13715 1241
rect 13681 1105 13715 1173
rect 13769 1343 13803 1359
rect 13769 1275 13803 1309
rect 13769 1207 13803 1241
rect 13769 1139 13803 1173
rect 13857 1343 13891 1377
rect 13857 1275 13891 1309
rect 13857 1207 13891 1241
rect 13857 1157 13891 1173
rect 13945 1343 13979 1359
rect 13945 1275 13979 1309
rect 13945 1207 13979 1241
rect 13945 1105 13979 1173
rect 14033 1343 14067 1377
rect 14033 1275 14067 1309
rect 14033 1207 14067 1241
rect 14033 1121 14067 1173
rect 14177 1436 14191 1470
rect 14225 1436 14239 1470
rect 14843 1470 14905 1492
rect 14177 1398 14239 1436
rect 14177 1364 14191 1398
rect 14225 1364 14239 1398
rect 14177 1326 14239 1364
rect 14177 1292 14191 1326
rect 14225 1292 14239 1326
rect 14177 1254 14239 1292
rect 14177 1220 14191 1254
rect 14225 1220 14239 1254
rect 14177 1182 14239 1220
rect 14177 1148 14191 1182
rect 14225 1148 14239 1182
rect 13769 1071 13945 1105
rect 13681 1055 13715 1071
rect 13945 1055 13979 1071
rect 14177 1110 14239 1148
rect 14177 1076 14191 1110
rect 14225 1076 14239 1110
rect 12845 966 12907 1004
rect 12845 932 12859 966
rect 12893 932 12907 966
rect 12845 868 12907 932
rect 13007 1004 13041 1020
rect 13237 1004 13271 1020
rect 12179 368 12193 402
rect 12227 368 12241 402
rect 11957 245 11991 342
rect 12179 330 12241 368
rect 11957 195 11991 211
rect 12054 289 12088 305
rect 12054 221 12088 255
rect 11860 151 11894 187
rect 12054 151 12088 187
rect 11894 117 11957 151
rect 11991 117 12054 151
rect 11860 101 11894 117
rect 12054 101 12088 117
rect 12179 296 12193 330
rect 12227 296 12241 330
rect 12179 258 12241 296
rect 12179 224 12193 258
rect 12227 224 12241 258
rect 12179 186 12241 224
rect 12179 152 12193 186
rect 12227 152 12241 186
rect 12179 114 12241 152
rect 12179 80 12193 114
rect 12227 80 12241 114
rect 12332 361 12366 377
rect 12526 361 12560 377
rect 12711 376 12745 797
rect 13007 831 13041 945
rect 12366 327 12429 361
rect 12463 327 12526 361
rect 12332 289 12366 327
rect 12332 221 12366 255
rect 12526 289 12560 327
rect 12332 151 12366 187
rect 12332 101 12366 117
rect 12429 236 12463 252
rect 12179 62 12241 80
rect 12429 62 12463 202
rect 12526 221 12560 255
rect 12623 342 12745 376
rect 12845 546 12907 572
rect 12845 512 12859 546
rect 12893 512 12907 546
rect 12845 474 12907 512
rect 12845 440 12859 474
rect 12893 440 12907 474
rect 12845 402 12907 440
rect 13007 461 13041 797
rect 13007 411 13041 427
rect 13229 970 13237 988
rect 13229 954 13271 970
rect 13511 1004 13525 1038
rect 13559 1004 13573 1038
rect 14177 1038 14239 1076
rect 14349 1411 14735 1445
rect 14349 1343 14383 1377
rect 14349 1275 14383 1309
rect 14349 1207 14383 1241
rect 14349 1105 14383 1173
rect 14437 1343 14471 1359
rect 14437 1275 14471 1309
rect 14437 1207 14471 1241
rect 14437 1139 14471 1173
rect 14525 1343 14559 1377
rect 14525 1275 14559 1309
rect 14525 1207 14559 1241
rect 14525 1157 14559 1173
rect 14613 1343 14647 1359
rect 14613 1275 14647 1309
rect 14613 1207 14647 1241
rect 14613 1139 14647 1173
rect 14701 1343 14735 1377
rect 14701 1275 14735 1309
rect 14701 1207 14735 1241
rect 14701 1157 14735 1173
rect 14843 1436 14857 1470
rect 14891 1436 14905 1470
rect 14843 1398 14905 1436
rect 14843 1364 14857 1398
rect 14891 1364 14905 1398
rect 14843 1326 14905 1364
rect 14843 1292 14857 1326
rect 14891 1292 14905 1326
rect 14843 1254 14905 1292
rect 14843 1220 14857 1254
rect 14891 1220 14905 1254
rect 14843 1182 14905 1220
rect 14843 1148 14857 1182
rect 14891 1148 14905 1182
rect 14843 1110 14905 1148
rect 14437 1071 14743 1105
rect 14349 1055 14383 1071
rect 13511 966 13573 1004
rect 13229 905 13263 954
rect 13229 535 13263 871
rect 13511 932 13525 966
rect 13559 932 13573 966
rect 13511 868 13573 932
rect 13747 1004 13781 1020
rect 13229 461 13263 501
rect 13229 411 13263 427
rect 13511 546 13573 572
rect 13511 512 13525 546
rect 13559 512 13573 546
rect 13511 474 13573 512
rect 13511 440 13525 474
rect 13559 440 13573 474
rect 12845 368 12859 402
rect 12893 368 12907 402
rect 13511 402 13573 440
rect 13747 461 13781 945
rect 13747 411 13781 427
rect 14043 1004 14077 1020
rect 14043 683 14077 970
rect 14177 1004 14191 1038
rect 14225 1004 14239 1038
rect 14177 966 14239 1004
rect 14177 932 14191 966
rect 14225 932 14239 966
rect 14177 868 14239 932
rect 14339 1004 14373 1020
rect 14043 461 14077 649
rect 14043 411 14077 427
rect 14177 546 14239 572
rect 14177 512 14191 546
rect 14225 512 14239 546
rect 14177 474 14239 512
rect 14177 440 14191 474
rect 14225 440 14239 474
rect 12623 245 12657 342
rect 12845 330 12907 368
rect 12623 195 12657 211
rect 12720 289 12754 305
rect 12720 221 12754 255
rect 12526 151 12560 187
rect 12720 151 12754 187
rect 12560 117 12623 151
rect 12657 117 12720 151
rect 12526 101 12560 117
rect 12720 101 12754 117
rect 12845 296 12859 330
rect 12893 296 12907 330
rect 12845 258 12907 296
rect 12845 224 12859 258
rect 12893 224 12907 258
rect 12845 186 12907 224
rect 12845 152 12859 186
rect 12893 152 12907 186
rect 12845 114 12907 152
rect 12845 80 12859 114
rect 12893 80 12907 114
rect 12998 361 13032 377
rect 13192 361 13226 377
rect 13032 327 13095 361
rect 13129 327 13192 361
rect 12998 289 13032 327
rect 12998 221 13032 255
rect 13192 289 13226 327
rect 13386 361 13420 377
rect 13289 281 13323 297
rect 12998 151 13032 187
rect 12998 101 13032 117
rect 13095 236 13129 252
rect 12845 62 12907 80
rect 13095 62 13129 202
rect 13192 221 13226 255
rect 13288 247 13289 262
rect 13288 245 13323 247
rect 13322 231 13323 245
rect 13386 289 13420 327
rect 13288 195 13322 211
rect 13386 221 13420 255
rect 13192 151 13226 187
rect 13386 151 13420 187
rect 13226 117 13288 151
rect 13322 117 13386 151
rect 13192 101 13226 117
rect 13386 101 13420 117
rect 13511 368 13525 402
rect 13559 368 13573 402
rect 14177 402 14239 440
rect 14339 461 14373 970
rect 14339 411 14373 427
rect 14561 1004 14599 1020
rect 14561 970 14565 1004
rect 14561 954 14599 970
rect 14561 905 14595 954
rect 14561 461 14595 871
rect 14561 411 14595 427
rect 14709 831 14743 1071
rect 14843 1076 14857 1110
rect 14891 1076 14905 1110
rect 14843 1038 14905 1076
rect 14843 1004 14857 1038
rect 14891 1004 14905 1038
rect 14843 966 14905 1004
rect 14843 932 14857 966
rect 14891 932 14905 966
rect 14843 868 14905 932
rect 13511 330 13573 368
rect 13511 296 13525 330
rect 13559 296 13573 330
rect 13511 258 13573 296
rect 13511 224 13525 258
rect 13559 224 13573 258
rect 13511 186 13573 224
rect 13511 152 13525 186
rect 13559 152 13573 186
rect 13511 114 13573 152
rect 13511 80 13525 114
rect 13559 80 13573 114
rect 13664 361 13698 377
rect 13858 361 13892 377
rect 13698 327 13761 361
rect 13795 327 13858 361
rect 13664 289 13698 327
rect 13664 221 13698 255
rect 13858 289 13892 327
rect 14052 361 14086 377
rect 13664 151 13698 187
rect 13664 101 13698 117
rect 13761 236 13795 252
rect 13511 62 13573 80
rect 13761 62 13795 202
rect 13858 221 13892 255
rect 13955 281 13989 297
rect 13955 245 13989 247
rect 13955 195 13989 211
rect 14052 289 14086 327
rect 14052 221 14086 255
rect 13858 151 13892 187
rect 14052 151 14086 187
rect 13892 117 13955 151
rect 13989 117 14052 151
rect 13858 101 13892 117
rect 14052 101 14086 117
rect 14177 368 14191 402
rect 14225 368 14239 402
rect 14177 330 14239 368
rect 14177 296 14191 330
rect 14225 296 14239 330
rect 14177 258 14239 296
rect 14177 224 14191 258
rect 14225 224 14239 258
rect 14177 186 14239 224
rect 14177 152 14191 186
rect 14225 152 14239 186
rect 14177 114 14239 152
rect 14177 80 14191 114
rect 14225 80 14239 114
rect 14330 361 14364 377
rect 14524 361 14558 377
rect 14709 374 14743 797
rect 14364 327 14427 361
rect 14461 327 14524 361
rect 14330 289 14364 327
rect 14330 221 14364 255
rect 14524 289 14558 327
rect 14330 151 14364 187
rect 14330 101 14364 117
rect 14427 236 14461 252
rect 14177 62 14239 80
rect 14427 62 14461 202
rect 14524 221 14558 255
rect 14621 340 14743 374
rect 14843 546 14905 572
rect 14843 512 14857 546
rect 14891 512 14905 546
rect 14843 474 14905 512
rect 14843 440 14857 474
rect 14891 440 14905 474
rect 14843 402 14905 440
rect 14843 368 14857 402
rect 14891 368 14905 402
rect 14621 281 14655 340
rect 14843 330 14905 368
rect 14621 245 14655 247
rect 14621 195 14655 211
rect 14718 289 14752 306
rect 14718 221 14752 255
rect 14524 151 14558 187
rect 14718 151 14752 187
rect 14558 117 14621 151
rect 14655 117 14718 151
rect 14524 101 14558 117
rect 14718 101 14752 117
rect 14843 296 14857 330
rect 14891 296 14905 330
rect 14843 258 14905 296
rect 14843 224 14857 258
rect 14891 224 14905 258
rect 14843 186 14905 224
rect 14843 152 14857 186
rect 14891 152 14905 186
rect 14843 114 14905 152
rect 14843 80 14857 114
rect 14891 80 14905 114
rect 14843 62 14905 80
rect -31 47 13955 62
rect 13989 47 14905 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 343 47
rect 377 13 415 47
rect 449 13 513 47
rect 547 13 585 47
rect 619 13 657 47
rect 691 13 729 47
rect 763 13 801 47
rect 835 13 873 47
rect 907 13 1017 47
rect 1051 13 1089 47
rect 1123 13 1161 47
rect 1195 13 1233 47
rect 1267 13 1323 47
rect 1357 13 1395 47
rect 1429 13 1467 47
rect 1501 13 1539 47
rect 1573 13 1683 47
rect 1717 13 1755 47
rect 1789 13 1827 47
rect 1861 13 1899 47
rect 1933 13 1989 47
rect 2023 13 2061 47
rect 2095 13 2133 47
rect 2167 13 2205 47
rect 2239 13 2349 47
rect 2383 13 2421 47
rect 2455 13 2493 47
rect 2527 13 2565 47
rect 2599 13 2655 47
rect 2689 13 2727 47
rect 2761 13 2799 47
rect 2833 13 2871 47
rect 2905 13 3015 47
rect 3049 13 3087 47
rect 3121 13 3159 47
rect 3193 13 3231 47
rect 3265 13 3321 47
rect 3355 13 3393 47
rect 3427 13 3465 47
rect 3499 13 3537 47
rect 3571 13 3681 47
rect 3715 13 3753 47
rect 3787 13 3825 47
rect 3859 13 3897 47
rect 3931 13 3987 47
rect 4021 13 4059 47
rect 4093 13 4131 47
rect 4165 13 4203 47
rect 4237 13 4347 47
rect 4381 13 4419 47
rect 4453 13 4491 47
rect 4525 13 4563 47
rect 4597 13 4635 47
rect 4669 13 4707 47
rect 4741 13 4805 47
rect 4839 13 4877 47
rect 4911 13 4949 47
rect 4983 13 5021 47
rect 5055 13 5093 47
rect 5127 13 5165 47
rect 5199 13 5309 47
rect 5343 13 5381 47
rect 5415 13 5453 47
rect 5487 13 5525 47
rect 5559 13 5615 47
rect 5649 13 5687 47
rect 5721 13 5759 47
rect 5793 13 5831 47
rect 5865 13 5975 47
rect 6009 13 6047 47
rect 6081 13 6119 47
rect 6153 13 6191 47
rect 6225 13 6281 47
rect 6315 13 6353 47
rect 6387 13 6425 47
rect 6459 13 6497 47
rect 6531 13 6641 47
rect 6675 13 6713 47
rect 6747 13 6785 47
rect 6819 13 6857 47
rect 6891 13 6947 47
rect 6981 13 7019 47
rect 7053 13 7091 47
rect 7125 13 7163 47
rect 7197 13 7307 47
rect 7341 13 7379 47
rect 7413 13 7451 47
rect 7485 13 7523 47
rect 7557 13 7613 47
rect 7647 13 7685 47
rect 7719 13 7757 47
rect 7791 13 7829 47
rect 7863 13 7973 47
rect 8007 13 8045 47
rect 8079 13 8117 47
rect 8151 13 8189 47
rect 8223 13 8279 47
rect 8313 13 8351 47
rect 8385 13 8423 47
rect 8457 13 8495 47
rect 8529 13 8639 47
rect 8673 13 8711 47
rect 8745 13 8783 47
rect 8817 13 8855 47
rect 8889 13 8927 47
rect 8961 13 8999 47
rect 9033 13 9097 47
rect 9131 13 9169 47
rect 9203 13 9241 47
rect 9275 13 9313 47
rect 9347 13 9385 47
rect 9419 13 9457 47
rect 9491 13 9601 47
rect 9635 13 9673 47
rect 9707 13 9745 47
rect 9779 13 9817 47
rect 9851 13 9907 47
rect 9941 13 9979 47
rect 10013 13 10051 47
rect 10085 13 10123 47
rect 10157 13 10267 47
rect 10301 13 10339 47
rect 10373 13 10411 47
rect 10445 13 10483 47
rect 10517 13 10573 47
rect 10607 13 10645 47
rect 10679 13 10717 47
rect 10751 13 10789 47
rect 10823 13 10933 47
rect 10967 13 11005 47
rect 11039 13 11077 47
rect 11111 13 11149 47
rect 11183 13 11239 47
rect 11273 13 11311 47
rect 11345 13 11383 47
rect 11417 13 11455 47
rect 11489 13 11599 47
rect 11633 13 11671 47
rect 11705 13 11743 47
rect 11777 13 11815 47
rect 11849 13 11905 47
rect 11939 13 11977 47
rect 12011 13 12049 47
rect 12083 13 12121 47
rect 12155 13 12265 47
rect 12299 13 12337 47
rect 12371 13 12409 47
rect 12443 13 12481 47
rect 12515 13 12571 47
rect 12605 13 12643 47
rect 12677 13 12715 47
rect 12749 13 12787 47
rect 12821 13 12931 47
rect 12965 13 13003 47
rect 13037 13 13075 47
rect 13109 13 13147 47
rect 13181 13 13237 47
rect 13271 13 13309 47
rect 13343 13 13381 47
rect 13415 13 13453 47
rect 13487 13 13597 47
rect 13631 13 13669 47
rect 13703 13 13741 47
rect 13775 13 13813 47
rect 13847 13 13903 47
rect 13937 13 13975 47
rect 14009 13 14047 47
rect 14081 13 14119 47
rect 14153 13 14263 47
rect 14297 13 14335 47
rect 14369 13 14407 47
rect 14441 13 14479 47
rect 14513 13 14569 47
rect 14603 13 14641 47
rect 14675 13 14713 47
rect 14747 13 14785 47
rect 14819 13 14905 47
rect -31 0 14905 13
<< viali >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 343 1505 377 1539
rect 415 1505 449 1539
rect 513 1505 547 1539
rect 585 1505 619 1539
rect 657 1505 691 1539
rect 729 1505 763 1539
rect 801 1505 835 1539
rect 873 1505 907 1539
rect 1017 1505 1051 1539
rect 1089 1505 1123 1539
rect 1161 1505 1195 1539
rect 1233 1505 1267 1539
rect 1323 1505 1357 1539
rect 1395 1505 1429 1539
rect 1467 1505 1501 1539
rect 1539 1505 1573 1539
rect 1683 1505 1717 1539
rect 1755 1505 1789 1539
rect 1827 1505 1861 1539
rect 1899 1505 1933 1539
rect 1989 1505 2023 1539
rect 2061 1505 2095 1539
rect 2133 1505 2167 1539
rect 2205 1505 2239 1539
rect 2349 1505 2383 1539
rect 2421 1505 2455 1539
rect 2493 1505 2527 1539
rect 2565 1505 2599 1539
rect 2655 1505 2689 1539
rect 2727 1505 2761 1539
rect 2799 1505 2833 1539
rect 2871 1505 2905 1539
rect 3015 1505 3049 1539
rect 3087 1505 3121 1539
rect 3159 1505 3193 1539
rect 3231 1505 3265 1539
rect 3321 1505 3355 1539
rect 3393 1505 3427 1539
rect 3465 1505 3499 1539
rect 3537 1505 3571 1539
rect 3681 1505 3715 1539
rect 3753 1505 3787 1539
rect 3825 1505 3859 1539
rect 3897 1505 3931 1539
rect 3987 1505 4021 1539
rect 4059 1505 4093 1539
rect 4131 1505 4165 1539
rect 4203 1505 4237 1539
rect 4347 1505 4381 1539
rect 4419 1505 4453 1539
rect 4491 1505 4525 1539
rect 4563 1505 4597 1539
rect 4635 1505 4669 1539
rect 4707 1505 4741 1539
rect 4805 1505 4839 1539
rect 4877 1505 4911 1539
rect 4949 1505 4983 1539
rect 5021 1505 5055 1539
rect 5093 1505 5127 1539
rect 5165 1505 5199 1539
rect 5309 1505 5343 1539
rect 5381 1505 5415 1539
rect 5453 1505 5487 1539
rect 5525 1505 5559 1539
rect 5615 1505 5649 1539
rect 5687 1505 5721 1539
rect 5759 1505 5793 1539
rect 5831 1505 5865 1539
rect 5975 1505 6009 1539
rect 6047 1505 6081 1539
rect 6119 1505 6153 1539
rect 6191 1505 6225 1539
rect 6281 1505 6315 1539
rect 6353 1505 6387 1539
rect 6425 1505 6459 1539
rect 6497 1505 6531 1539
rect 6641 1505 6675 1539
rect 6713 1505 6747 1539
rect 6785 1505 6819 1539
rect 6857 1505 6891 1539
rect 6947 1505 6981 1539
rect 7019 1505 7053 1539
rect 7091 1505 7125 1539
rect 7163 1505 7197 1539
rect 7307 1505 7341 1539
rect 7379 1505 7413 1539
rect 7451 1505 7485 1539
rect 7523 1505 7557 1539
rect 7613 1505 7647 1539
rect 7685 1505 7719 1539
rect 7757 1505 7791 1539
rect 7829 1505 7863 1539
rect 7973 1505 8007 1539
rect 8045 1505 8079 1539
rect 8117 1505 8151 1539
rect 8189 1505 8223 1539
rect 8279 1505 8313 1539
rect 8351 1505 8385 1539
rect 8423 1505 8457 1539
rect 8495 1505 8529 1539
rect 8639 1505 8673 1539
rect 8711 1505 8745 1539
rect 8783 1505 8817 1539
rect 8855 1505 8889 1539
rect 8927 1505 8961 1539
rect 8999 1505 9033 1539
rect 9097 1505 9131 1539
rect 9169 1505 9203 1539
rect 9241 1505 9275 1539
rect 9313 1505 9347 1539
rect 9385 1505 9419 1539
rect 9457 1505 9491 1539
rect 9601 1505 9635 1539
rect 9673 1505 9707 1539
rect 9745 1505 9779 1539
rect 9817 1505 9851 1539
rect 9907 1505 9941 1539
rect 9979 1505 10013 1539
rect 10051 1505 10085 1539
rect 10123 1505 10157 1539
rect 10267 1505 10301 1539
rect 10339 1505 10373 1539
rect 10411 1505 10445 1539
rect 10483 1505 10517 1539
rect 10573 1505 10607 1539
rect 10645 1505 10679 1539
rect 10717 1505 10751 1539
rect 10789 1505 10823 1539
rect 10933 1505 10967 1539
rect 11005 1505 11039 1539
rect 11077 1505 11111 1539
rect 11149 1505 11183 1539
rect 11239 1505 11273 1539
rect 11311 1505 11345 1539
rect 11383 1505 11417 1539
rect 11455 1505 11489 1539
rect 11599 1505 11633 1539
rect 11671 1505 11705 1539
rect 11743 1505 11777 1539
rect 11815 1505 11849 1539
rect 11905 1505 11939 1539
rect 11977 1505 12011 1539
rect 12049 1505 12083 1539
rect 12121 1505 12155 1539
rect 12265 1505 12299 1539
rect 12337 1505 12371 1539
rect 12409 1505 12443 1539
rect 12481 1505 12515 1539
rect 12571 1505 12605 1539
rect 12643 1505 12677 1539
rect 12715 1505 12749 1539
rect 12787 1505 12821 1539
rect 12931 1505 12965 1539
rect 13003 1505 13037 1539
rect 13075 1505 13109 1539
rect 13147 1505 13181 1539
rect 13237 1505 13271 1539
rect 13309 1505 13343 1539
rect 13381 1505 13415 1539
rect 13453 1505 13487 1539
rect 13597 1505 13631 1539
rect 13669 1505 13703 1539
rect 13741 1505 13775 1539
rect 13813 1505 13847 1539
rect 13903 1505 13937 1539
rect 13975 1505 14009 1539
rect 14047 1505 14081 1539
rect 14119 1505 14153 1539
rect 14263 1505 14297 1539
rect 14335 1505 14369 1539
rect 14407 1505 14441 1539
rect 14479 1505 14513 1539
rect 14569 1505 14603 1539
rect 14641 1505 14675 1539
rect 14713 1505 14747 1539
rect 14785 1505 14819 1539
rect 205 871 239 905
rect 427 969 461 979
rect 427 945 461 969
rect 649 723 683 757
rect 797 797 831 831
rect 1167 797 1201 831
rect 1315 427 1349 461
rect 1463 723 1497 757
rect 1833 723 1867 757
rect 1981 871 2015 905
rect 2129 723 2163 757
rect 2499 723 2533 757
rect 2647 969 2653 979
rect 2653 969 2681 979
rect 2647 945 2681 969
rect 2795 871 2829 905
rect 3165 797 3199 831
rect 3313 649 3347 683
rect 3461 797 3495 831
rect 3831 797 3865 831
rect 3979 871 4013 905
rect 4497 871 4531 905
rect 4127 649 4161 683
rect 4719 969 4753 979
rect 4719 945 4753 969
rect 4941 723 4975 757
rect 5089 797 5123 831
rect 5459 797 5493 831
rect 5607 427 5641 461
rect 5755 723 5789 757
rect 6125 723 6159 757
rect 6273 871 6307 905
rect 6421 723 6455 757
rect 6791 723 6825 757
rect 6939 969 6945 979
rect 6945 969 6973 979
rect 6939 945 6973 969
rect 7087 871 7121 905
rect 7457 797 7491 831
rect 7605 501 7639 535
rect 7753 797 7787 831
rect 8123 797 8157 831
rect 8271 871 8305 905
rect 8789 871 8823 905
rect 8419 501 8453 535
rect 9011 969 9045 979
rect 9011 945 9045 969
rect 9233 723 9267 757
rect 9381 797 9415 831
rect 9751 797 9785 831
rect 9899 427 9933 461
rect 10047 723 10081 757
rect 10417 723 10451 757
rect 10565 871 10599 905
rect 10713 723 10747 757
rect 11083 723 11117 757
rect 11231 969 11237 979
rect 11237 969 11265 979
rect 11231 945 11265 969
rect 11379 871 11413 905
rect 11749 797 11783 831
rect 11897 797 11931 831
rect 12045 945 12079 979
rect 12415 969 12449 979
rect 12415 945 12449 969
rect 12563 871 12597 905
rect 13281 1071 13315 1105
rect 13681 1071 13715 1105
rect 13945 1071 13979 1105
rect 13007 970 13041 979
rect 13007 945 13041 970
rect 12711 797 12745 831
rect 13007 797 13041 831
rect 14349 1071 14383 1105
rect 13229 871 13263 905
rect 13747 970 13781 979
rect 13747 945 13781 970
rect 13229 501 13263 535
rect 14043 649 14077 683
rect 14043 427 14077 461
rect 13289 247 13323 281
rect 14339 427 14373 461
rect 14561 871 14595 905
rect 14709 797 14743 831
rect 13955 247 13989 281
rect 14621 247 14655 281
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 343 13 377 47
rect 415 13 449 47
rect 513 13 547 47
rect 585 13 619 47
rect 657 13 691 47
rect 729 13 763 47
rect 801 13 835 47
rect 873 13 907 47
rect 1017 13 1051 47
rect 1089 13 1123 47
rect 1161 13 1195 47
rect 1233 13 1267 47
rect 1323 13 1357 47
rect 1395 13 1429 47
rect 1467 13 1501 47
rect 1539 13 1573 47
rect 1683 13 1717 47
rect 1755 13 1789 47
rect 1827 13 1861 47
rect 1899 13 1933 47
rect 1989 13 2023 47
rect 2061 13 2095 47
rect 2133 13 2167 47
rect 2205 13 2239 47
rect 2349 13 2383 47
rect 2421 13 2455 47
rect 2493 13 2527 47
rect 2565 13 2599 47
rect 2655 13 2689 47
rect 2727 13 2761 47
rect 2799 13 2833 47
rect 2871 13 2905 47
rect 3015 13 3049 47
rect 3087 13 3121 47
rect 3159 13 3193 47
rect 3231 13 3265 47
rect 3321 13 3355 47
rect 3393 13 3427 47
rect 3465 13 3499 47
rect 3537 13 3571 47
rect 3681 13 3715 47
rect 3753 13 3787 47
rect 3825 13 3859 47
rect 3897 13 3931 47
rect 3987 13 4021 47
rect 4059 13 4093 47
rect 4131 13 4165 47
rect 4203 13 4237 47
rect 4347 13 4381 47
rect 4419 13 4453 47
rect 4491 13 4525 47
rect 4563 13 4597 47
rect 4635 13 4669 47
rect 4707 13 4741 47
rect 4805 13 4839 47
rect 4877 13 4911 47
rect 4949 13 4983 47
rect 5021 13 5055 47
rect 5093 13 5127 47
rect 5165 13 5199 47
rect 5309 13 5343 47
rect 5381 13 5415 47
rect 5453 13 5487 47
rect 5525 13 5559 47
rect 5615 13 5649 47
rect 5687 13 5721 47
rect 5759 13 5793 47
rect 5831 13 5865 47
rect 5975 13 6009 47
rect 6047 13 6081 47
rect 6119 13 6153 47
rect 6191 13 6225 47
rect 6281 13 6315 47
rect 6353 13 6387 47
rect 6425 13 6459 47
rect 6497 13 6531 47
rect 6641 13 6675 47
rect 6713 13 6747 47
rect 6785 13 6819 47
rect 6857 13 6891 47
rect 6947 13 6981 47
rect 7019 13 7053 47
rect 7091 13 7125 47
rect 7163 13 7197 47
rect 7307 13 7341 47
rect 7379 13 7413 47
rect 7451 13 7485 47
rect 7523 13 7557 47
rect 7613 13 7647 47
rect 7685 13 7719 47
rect 7757 13 7791 47
rect 7829 13 7863 47
rect 7973 13 8007 47
rect 8045 13 8079 47
rect 8117 13 8151 47
rect 8189 13 8223 47
rect 8279 13 8313 47
rect 8351 13 8385 47
rect 8423 13 8457 47
rect 8495 13 8529 47
rect 8639 13 8673 47
rect 8711 13 8745 47
rect 8783 13 8817 47
rect 8855 13 8889 47
rect 8927 13 8961 47
rect 8999 13 9033 47
rect 9097 13 9131 47
rect 9169 13 9203 47
rect 9241 13 9275 47
rect 9313 13 9347 47
rect 9385 13 9419 47
rect 9457 13 9491 47
rect 9601 13 9635 47
rect 9673 13 9707 47
rect 9745 13 9779 47
rect 9817 13 9851 47
rect 9907 13 9941 47
rect 9979 13 10013 47
rect 10051 13 10085 47
rect 10123 13 10157 47
rect 10267 13 10301 47
rect 10339 13 10373 47
rect 10411 13 10445 47
rect 10483 13 10517 47
rect 10573 13 10607 47
rect 10645 13 10679 47
rect 10717 13 10751 47
rect 10789 13 10823 47
rect 10933 13 10967 47
rect 11005 13 11039 47
rect 11077 13 11111 47
rect 11149 13 11183 47
rect 11239 13 11273 47
rect 11311 13 11345 47
rect 11383 13 11417 47
rect 11455 13 11489 47
rect 11599 13 11633 47
rect 11671 13 11705 47
rect 11743 13 11777 47
rect 11815 13 11849 47
rect 11905 13 11939 47
rect 11977 13 12011 47
rect 12049 13 12083 47
rect 12121 13 12155 47
rect 12265 13 12299 47
rect 12337 13 12371 47
rect 12409 13 12443 47
rect 12481 13 12515 47
rect 12571 13 12605 47
rect 12643 13 12677 47
rect 12715 13 12749 47
rect 12787 13 12821 47
rect 12931 13 12965 47
rect 13003 13 13037 47
rect 13075 13 13109 47
rect 13147 13 13181 47
rect 13237 13 13271 47
rect 13309 13 13343 47
rect 13381 13 13415 47
rect 13453 13 13487 47
rect 13597 13 13631 47
rect 13669 13 13703 47
rect 13741 13 13775 47
rect 13813 13 13847 47
rect 13903 13 13937 47
rect 13975 13 14009 47
rect 14047 13 14081 47
rect 14119 13 14153 47
rect 14263 13 14297 47
rect 14335 13 14369 47
rect 14407 13 14441 47
rect 14479 13 14513 47
rect 14569 13 14603 47
rect 14641 13 14675 47
rect 14713 13 14747 47
rect 14785 13 14819 47
<< metal1 >>
rect -31 1539 14905 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 343 1539
rect 377 1505 415 1539
rect 449 1505 513 1539
rect 547 1505 585 1539
rect 619 1505 657 1539
rect 691 1505 729 1539
rect 763 1505 801 1539
rect 835 1505 873 1539
rect 907 1505 1017 1539
rect 1051 1505 1089 1539
rect 1123 1505 1161 1539
rect 1195 1505 1233 1539
rect 1267 1505 1323 1539
rect 1357 1505 1395 1539
rect 1429 1505 1467 1539
rect 1501 1505 1539 1539
rect 1573 1505 1683 1539
rect 1717 1505 1755 1539
rect 1789 1505 1827 1539
rect 1861 1505 1899 1539
rect 1933 1505 1989 1539
rect 2023 1505 2061 1539
rect 2095 1505 2133 1539
rect 2167 1505 2205 1539
rect 2239 1505 2349 1539
rect 2383 1505 2421 1539
rect 2455 1505 2493 1539
rect 2527 1505 2565 1539
rect 2599 1505 2655 1539
rect 2689 1505 2727 1539
rect 2761 1505 2799 1539
rect 2833 1505 2871 1539
rect 2905 1505 3015 1539
rect 3049 1505 3087 1539
rect 3121 1505 3159 1539
rect 3193 1505 3231 1539
rect 3265 1505 3321 1539
rect 3355 1505 3393 1539
rect 3427 1505 3465 1539
rect 3499 1505 3537 1539
rect 3571 1505 3681 1539
rect 3715 1505 3753 1539
rect 3787 1505 3825 1539
rect 3859 1505 3897 1539
rect 3931 1505 3987 1539
rect 4021 1505 4059 1539
rect 4093 1505 4131 1539
rect 4165 1505 4203 1539
rect 4237 1505 4347 1539
rect 4381 1505 4419 1539
rect 4453 1505 4491 1539
rect 4525 1505 4563 1539
rect 4597 1505 4635 1539
rect 4669 1505 4707 1539
rect 4741 1505 4805 1539
rect 4839 1505 4877 1539
rect 4911 1505 4949 1539
rect 4983 1505 5021 1539
rect 5055 1505 5093 1539
rect 5127 1505 5165 1539
rect 5199 1505 5309 1539
rect 5343 1505 5381 1539
rect 5415 1505 5453 1539
rect 5487 1505 5525 1539
rect 5559 1505 5615 1539
rect 5649 1505 5687 1539
rect 5721 1505 5759 1539
rect 5793 1505 5831 1539
rect 5865 1505 5975 1539
rect 6009 1505 6047 1539
rect 6081 1505 6119 1539
rect 6153 1505 6191 1539
rect 6225 1505 6281 1539
rect 6315 1505 6353 1539
rect 6387 1505 6425 1539
rect 6459 1505 6497 1539
rect 6531 1505 6641 1539
rect 6675 1505 6713 1539
rect 6747 1505 6785 1539
rect 6819 1505 6857 1539
rect 6891 1505 6947 1539
rect 6981 1505 7019 1539
rect 7053 1505 7091 1539
rect 7125 1505 7163 1539
rect 7197 1505 7307 1539
rect 7341 1505 7379 1539
rect 7413 1505 7451 1539
rect 7485 1505 7523 1539
rect 7557 1505 7613 1539
rect 7647 1505 7685 1539
rect 7719 1505 7757 1539
rect 7791 1505 7829 1539
rect 7863 1505 7973 1539
rect 8007 1505 8045 1539
rect 8079 1505 8117 1539
rect 8151 1505 8189 1539
rect 8223 1505 8279 1539
rect 8313 1505 8351 1539
rect 8385 1505 8423 1539
rect 8457 1505 8495 1539
rect 8529 1505 8639 1539
rect 8673 1505 8711 1539
rect 8745 1505 8783 1539
rect 8817 1505 8855 1539
rect 8889 1505 8927 1539
rect 8961 1505 8999 1539
rect 9033 1505 9097 1539
rect 9131 1505 9169 1539
rect 9203 1505 9241 1539
rect 9275 1505 9313 1539
rect 9347 1505 9385 1539
rect 9419 1505 9457 1539
rect 9491 1505 9601 1539
rect 9635 1505 9673 1539
rect 9707 1505 9745 1539
rect 9779 1505 9817 1539
rect 9851 1505 9907 1539
rect 9941 1505 9979 1539
rect 10013 1505 10051 1539
rect 10085 1505 10123 1539
rect 10157 1505 10267 1539
rect 10301 1505 10339 1539
rect 10373 1505 10411 1539
rect 10445 1505 10483 1539
rect 10517 1505 10573 1539
rect 10607 1505 10645 1539
rect 10679 1505 10717 1539
rect 10751 1505 10789 1539
rect 10823 1505 10933 1539
rect 10967 1505 11005 1539
rect 11039 1505 11077 1539
rect 11111 1505 11149 1539
rect 11183 1505 11239 1539
rect 11273 1505 11311 1539
rect 11345 1505 11383 1539
rect 11417 1505 11455 1539
rect 11489 1505 11599 1539
rect 11633 1505 11671 1539
rect 11705 1505 11743 1539
rect 11777 1505 11815 1539
rect 11849 1505 11905 1539
rect 11939 1505 11977 1539
rect 12011 1505 12049 1539
rect 12083 1505 12121 1539
rect 12155 1505 12265 1539
rect 12299 1505 12337 1539
rect 12371 1505 12409 1539
rect 12443 1505 12481 1539
rect 12515 1505 12571 1539
rect 12605 1505 12643 1539
rect 12677 1505 12715 1539
rect 12749 1505 12787 1539
rect 12821 1505 12931 1539
rect 12965 1505 13003 1539
rect 13037 1505 13075 1539
rect 13109 1505 13147 1539
rect 13181 1505 13237 1539
rect 13271 1505 13309 1539
rect 13343 1505 13381 1539
rect 13415 1505 13453 1539
rect 13487 1505 13597 1539
rect 13631 1505 13669 1539
rect 13703 1505 13741 1539
rect 13775 1505 13813 1539
rect 13847 1505 13903 1539
rect 13937 1505 13975 1539
rect 14009 1505 14047 1539
rect 14081 1505 14119 1539
rect 14153 1505 14263 1539
rect 14297 1505 14335 1539
rect 14369 1505 14407 1539
rect 14441 1505 14479 1539
rect 14513 1505 14569 1539
rect 14603 1505 14641 1539
rect 14675 1505 14713 1539
rect 14747 1505 14785 1539
rect 14819 1505 14905 1539
rect -31 1492 14905 1505
rect 13275 1105 13321 1111
rect 13675 1105 13721 1111
rect 13939 1105 13985 1111
rect 14343 1105 14389 1111
rect 13269 1071 13281 1105
rect 13315 1071 13681 1105
rect 13715 1071 13727 1105
rect 13933 1071 13945 1105
rect 13979 1071 14349 1105
rect 14383 1071 14395 1105
rect 13275 1065 13321 1071
rect 13675 1065 13721 1071
rect 13939 1065 13985 1071
rect 14343 1065 14389 1071
rect 421 979 467 985
rect 2641 979 2687 985
rect 4713 979 4759 985
rect 6933 979 6979 985
rect 9005 979 9051 985
rect 11225 979 11271 985
rect 12039 979 12085 985
rect 12409 979 12455 985
rect 13001 979 13047 985
rect 13741 979 13787 985
rect 415 945 427 979
rect 461 945 2647 979
rect 2681 978 2693 979
rect 3349 978 4719 979
rect 2681 947 4719 978
rect 2681 945 2693 947
rect 3349 945 4719 947
rect 4753 945 6939 979
rect 6973 945 9011 979
rect 9045 945 11231 979
rect 11265 945 11277 979
rect 12033 945 12045 979
rect 12079 945 12415 979
rect 12449 945 12461 979
rect 12995 945 13007 979
rect 13041 945 13747 979
rect 13781 945 13793 979
rect 421 939 467 945
rect 2641 939 2687 945
rect 4713 939 4759 945
rect 6933 939 6979 945
rect 9005 939 9051 945
rect 11225 939 11271 945
rect 12039 939 12085 945
rect 12409 939 12455 945
rect 13001 939 13047 945
rect 13741 939 13787 945
rect 199 905 245 911
rect 1975 905 2021 911
rect 2789 905 2835 911
rect 3973 905 4019 911
rect 4491 905 4537 911
rect 6267 905 6313 911
rect 7081 905 7127 911
rect 8265 905 8311 911
rect 8783 905 8829 911
rect 10559 905 10605 911
rect 11373 905 11419 911
rect 12557 905 12603 911
rect 13223 905 13269 911
rect 14555 905 14601 911
rect 193 871 205 905
rect 239 871 1981 905
rect 2015 871 2795 905
rect 2829 871 3979 905
rect 4013 871 4025 905
rect 4485 871 4497 905
rect 4531 871 6273 905
rect 6307 871 7087 905
rect 7121 871 8271 905
rect 8305 871 8317 905
rect 8777 871 8789 905
rect 8823 871 10565 905
rect 10599 871 11379 905
rect 11413 871 12563 905
rect 12597 871 12609 905
rect 13217 871 13229 905
rect 13263 871 14561 905
rect 14595 871 14607 905
rect 199 865 245 871
rect 1975 865 2021 871
rect 2789 865 2835 871
rect 3973 865 4019 871
rect 4491 865 4537 871
rect 6267 865 6313 871
rect 7081 865 7127 871
rect 8265 865 8311 871
rect 8783 865 8829 871
rect 10559 865 10605 871
rect 11373 865 11419 871
rect 12557 865 12603 871
rect 13223 865 13269 871
rect 14555 865 14601 871
rect 791 831 837 837
rect 1161 831 1207 837
rect 3159 831 3205 837
rect 3455 831 3501 837
rect 3825 831 3871 837
rect 5083 831 5129 837
rect 5453 831 5499 837
rect 7451 831 7497 837
rect 7747 831 7793 837
rect 8117 831 8163 837
rect 9375 831 9421 837
rect 9745 831 9791 837
rect 11743 831 11789 837
rect 11891 831 11937 837
rect 12705 831 12751 837
rect 13001 831 13047 837
rect 14703 831 14749 837
rect 785 797 797 831
rect 831 797 1167 831
rect 1201 797 3165 831
rect 3199 797 3211 831
rect 3449 797 3461 831
rect 3495 797 3831 831
rect 3865 797 3877 831
rect 5077 797 5089 831
rect 5123 797 5459 831
rect 5493 797 7457 831
rect 7491 797 7503 831
rect 7741 797 7753 831
rect 7787 797 8123 831
rect 8157 797 8169 831
rect 9369 797 9381 831
rect 9415 797 9751 831
rect 9785 797 11749 831
rect 11783 797 11795 831
rect 11885 797 11897 831
rect 11931 797 12711 831
rect 12745 797 13007 831
rect 13041 797 13053 831
rect 14697 797 14709 831
rect 14743 797 14779 831
rect 791 791 837 797
rect 1161 791 1207 797
rect 3159 791 3205 797
rect 3455 791 3501 797
rect 3825 791 3871 797
rect 5083 791 5129 797
rect 5453 791 5499 797
rect 7451 791 7497 797
rect 7747 791 7793 797
rect 8117 791 8163 797
rect 9375 791 9421 797
rect 9745 791 9791 797
rect 11743 791 11789 797
rect 11891 791 11937 797
rect 12705 791 12751 797
rect 13001 791 13047 797
rect 14703 791 14749 797
rect 643 757 689 763
rect 1457 757 1503 763
rect 1827 757 1873 763
rect 2123 757 2169 763
rect 2493 757 2539 763
rect 4935 757 4981 763
rect 5749 757 5795 763
rect 6119 757 6165 763
rect 6415 757 6461 763
rect 6785 757 6831 763
rect 9227 757 9273 763
rect 10041 757 10087 763
rect 10411 757 10457 763
rect 10707 757 10753 763
rect 11077 757 11123 763
rect 637 723 649 757
rect 683 723 1463 757
rect 1497 723 1833 757
rect 1867 723 1879 757
rect 2117 723 2129 757
rect 2163 723 2499 757
rect 2533 723 2545 757
rect 4929 723 4941 757
rect 4975 723 5755 757
rect 5789 723 6125 757
rect 6159 723 6171 757
rect 6409 723 6421 757
rect 6455 723 6791 757
rect 6825 723 6837 757
rect 9221 723 9233 757
rect 9267 723 10047 757
rect 10081 723 10417 757
rect 10451 723 10463 757
rect 10701 723 10713 757
rect 10747 723 11083 757
rect 11117 723 11129 757
rect 643 717 689 723
rect 1457 717 1503 723
rect 1827 717 1873 723
rect 2123 717 2169 723
rect 2493 717 2539 723
rect 4935 717 4981 723
rect 5749 717 5795 723
rect 6119 717 6165 723
rect 6415 717 6461 723
rect 6785 717 6831 723
rect 9227 717 9273 723
rect 10041 717 10087 723
rect 10411 717 10457 723
rect 10707 717 10753 723
rect 11077 717 11123 723
rect 3307 683 3353 689
rect 4121 683 4167 689
rect 14037 683 14083 689
rect 3301 649 3313 683
rect 3347 649 4127 683
rect 4161 649 14043 683
rect 14077 649 14089 683
rect 3307 643 3353 649
rect 4121 643 4167 649
rect 14037 643 14083 649
rect 7599 535 7645 541
rect 8413 535 8459 541
rect 13223 535 13269 541
rect 7593 501 7605 535
rect 7639 501 8419 535
rect 8453 501 13229 535
rect 13263 501 13275 535
rect 7599 495 7645 501
rect 8413 495 8459 501
rect 13223 495 13269 501
rect 1309 461 1355 467
rect 5601 461 5647 467
rect 9893 461 9939 467
rect 14037 461 14083 467
rect 14333 461 14379 467
rect 1279 427 1315 461
rect 1349 427 5607 461
rect 5641 427 9899 461
rect 9933 427 9945 461
rect 14031 427 14043 461
rect 14077 427 14339 461
rect 14373 427 14385 461
rect 1309 421 1355 427
rect 5601 421 5647 427
rect 9893 421 9939 427
rect 14037 421 14083 427
rect 14333 421 14379 427
rect 13283 281 13329 287
rect 13949 281 13995 287
rect 14615 281 14661 287
rect 13277 247 13289 281
rect 13323 247 13955 281
rect 13989 247 14621 281
rect 14655 247 14667 281
rect 13283 241 13329 247
rect 13949 241 13995 247
rect 14615 241 14661 247
rect -31 47 14905 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 343 47
rect 377 13 415 47
rect 449 13 513 47
rect 547 13 585 47
rect 619 13 657 47
rect 691 13 729 47
rect 763 13 801 47
rect 835 13 873 47
rect 907 13 1017 47
rect 1051 13 1089 47
rect 1123 13 1161 47
rect 1195 13 1233 47
rect 1267 13 1323 47
rect 1357 13 1395 47
rect 1429 13 1467 47
rect 1501 13 1539 47
rect 1573 13 1683 47
rect 1717 13 1755 47
rect 1789 13 1827 47
rect 1861 13 1899 47
rect 1933 13 1989 47
rect 2023 13 2061 47
rect 2095 13 2133 47
rect 2167 13 2205 47
rect 2239 13 2349 47
rect 2383 13 2421 47
rect 2455 13 2493 47
rect 2527 13 2565 47
rect 2599 13 2655 47
rect 2689 13 2727 47
rect 2761 13 2799 47
rect 2833 13 2871 47
rect 2905 13 3015 47
rect 3049 13 3087 47
rect 3121 13 3159 47
rect 3193 13 3231 47
rect 3265 13 3321 47
rect 3355 13 3393 47
rect 3427 13 3465 47
rect 3499 13 3537 47
rect 3571 13 3681 47
rect 3715 13 3753 47
rect 3787 13 3825 47
rect 3859 13 3897 47
rect 3931 13 3987 47
rect 4021 13 4059 47
rect 4093 13 4131 47
rect 4165 13 4203 47
rect 4237 13 4347 47
rect 4381 13 4419 47
rect 4453 13 4491 47
rect 4525 13 4563 47
rect 4597 13 4635 47
rect 4669 13 4707 47
rect 4741 13 4805 47
rect 4839 13 4877 47
rect 4911 13 4949 47
rect 4983 13 5021 47
rect 5055 13 5093 47
rect 5127 13 5165 47
rect 5199 13 5309 47
rect 5343 13 5381 47
rect 5415 13 5453 47
rect 5487 13 5525 47
rect 5559 13 5615 47
rect 5649 13 5687 47
rect 5721 13 5759 47
rect 5793 13 5831 47
rect 5865 13 5975 47
rect 6009 13 6047 47
rect 6081 13 6119 47
rect 6153 13 6191 47
rect 6225 13 6281 47
rect 6315 13 6353 47
rect 6387 13 6425 47
rect 6459 13 6497 47
rect 6531 13 6641 47
rect 6675 13 6713 47
rect 6747 13 6785 47
rect 6819 13 6857 47
rect 6891 13 6947 47
rect 6981 13 7019 47
rect 7053 13 7091 47
rect 7125 13 7163 47
rect 7197 13 7307 47
rect 7341 13 7379 47
rect 7413 13 7451 47
rect 7485 13 7523 47
rect 7557 13 7613 47
rect 7647 13 7685 47
rect 7719 13 7757 47
rect 7791 13 7829 47
rect 7863 13 7973 47
rect 8007 13 8045 47
rect 8079 13 8117 47
rect 8151 13 8189 47
rect 8223 13 8279 47
rect 8313 13 8351 47
rect 8385 13 8423 47
rect 8457 13 8495 47
rect 8529 13 8639 47
rect 8673 13 8711 47
rect 8745 13 8783 47
rect 8817 13 8855 47
rect 8889 13 8927 47
rect 8961 13 8999 47
rect 9033 13 9097 47
rect 9131 13 9169 47
rect 9203 13 9241 47
rect 9275 13 9313 47
rect 9347 13 9385 47
rect 9419 13 9457 47
rect 9491 13 9601 47
rect 9635 13 9673 47
rect 9707 13 9745 47
rect 9779 13 9817 47
rect 9851 13 9907 47
rect 9941 13 9979 47
rect 10013 13 10051 47
rect 10085 13 10123 47
rect 10157 13 10267 47
rect 10301 13 10339 47
rect 10373 13 10411 47
rect 10445 13 10483 47
rect 10517 13 10573 47
rect 10607 13 10645 47
rect 10679 13 10717 47
rect 10751 13 10789 47
rect 10823 13 10933 47
rect 10967 13 11005 47
rect 11039 13 11077 47
rect 11111 13 11149 47
rect 11183 13 11239 47
rect 11273 13 11311 47
rect 11345 13 11383 47
rect 11417 13 11455 47
rect 11489 13 11599 47
rect 11633 13 11671 47
rect 11705 13 11743 47
rect 11777 13 11815 47
rect 11849 13 11905 47
rect 11939 13 11977 47
rect 12011 13 12049 47
rect 12083 13 12121 47
rect 12155 13 12265 47
rect 12299 13 12337 47
rect 12371 13 12409 47
rect 12443 13 12481 47
rect 12515 13 12571 47
rect 12605 13 12643 47
rect 12677 13 12715 47
rect 12749 13 12787 47
rect 12821 13 12931 47
rect 12965 13 13003 47
rect 13037 13 13075 47
rect 13109 13 13147 47
rect 13181 13 13237 47
rect 13271 13 13309 47
rect 13343 13 13381 47
rect 13415 13 13453 47
rect 13487 13 13597 47
rect 13631 13 13669 47
rect 13703 13 13741 47
rect 13775 13 13813 47
rect 13847 13 13903 47
rect 13937 13 13975 47
rect 14009 13 14047 47
rect 14081 13 14119 47
rect 14153 13 14263 47
rect 14297 13 14335 47
rect 14369 13 14407 47
rect 14441 13 14479 47
rect 14513 13 14569 47
rect 14603 13 14641 47
rect 14675 13 14713 47
rect 14747 13 14785 47
rect 14819 13 14905 47
rect -31 0 14905 13
<< labels >>
rlabel metal1 14709 797 14743 831 1 QN
port 1 n
rlabel metal1 1315 427 1349 461 1 D
port 2 n
rlabel metal1 427 945 461 979 1 CLK
port 3 n
rlabel metal1 72 1522 72 1522 1 VDD
port 4 n
rlabel metal1 72 30 72 30 1 VSS
port 5 n
<< end >>
