magic
tech sky130
magscale 1 2
timestamp 1645638725
<< nwell >>
rect 84 1264 508 1353
rect 84 941 507 1264
rect 84 759 508 941
<< psubdiff >>
rect 31 508 561 570
rect 31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 276 47
rect 310 13 353 47
rect 387 13 425 47
rect 459 13 497 47
rect 531 13 561 47
<< nsubdiff >>
rect 31 1283 55 1317
rect 89 1283 127 1317
rect 161 1283 199 1317
rect 233 1283 276 1317
rect 310 1283 353 1317
rect 387 1283 425 1317
rect 459 1283 497 1317
rect 531 1283 561 1317
rect 31 795 561 857
<< psubdiffcont >>
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 276 13 310 47
rect 353 13 387 47
rect 425 13 459 47
rect 497 13 531 47
<< nsubdiffcont >>
rect 55 1283 89 1317
rect 127 1283 161 1317
rect 199 1283 233 1317
rect 276 1283 310 1317
rect 353 1283 387 1317
rect 425 1283 459 1317
rect 497 1283 531 1317
<< poly >>
rect 147 418 255 448
rect 225 403 255 418
<< locali >>
rect 31 1317 561 1332
rect 31 1283 55 1317
rect 89 1283 127 1317
rect 161 1283 199 1317
rect 233 1283 276 1317
rect 310 1283 353 1317
rect 387 1283 425 1317
rect 459 1283 497 1317
rect 531 1283 561 1317
rect 31 1270 561 1283
rect 280 1269 314 1270
rect 192 961 226 1007
rect 368 961 402 1001
rect 192 927 402 961
rect 179 62 213 101
rect 372 62 406 101
rect 31 47 561 62
rect 31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 276 47
rect 310 13 353 47
rect 387 13 425 47
rect 459 13 497 47
rect 531 13 561 47
rect 31 0 561 13
<< viali >>
rect 55 1283 89 1317
rect 127 1283 161 1317
rect 199 1283 233 1317
rect 276 1283 310 1317
rect 353 1283 387 1317
rect 425 1283 459 1317
rect 497 1283 531 1317
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 276 13 310 47
rect 353 13 387 47
rect 425 13 459 47
rect 497 13 531 47
<< metal1 >>
rect 31 1317 561 1332
rect 31 1283 55 1317
rect 89 1283 127 1317
rect 161 1283 199 1317
rect 233 1283 276 1317
rect 310 1283 353 1317
rect 387 1283 425 1317
rect 459 1283 497 1317
rect 531 1283 561 1317
rect 31 1270 561 1283
rect 137 889 165 890
rect 131 456 165 889
rect 279 744 313 911
rect 280 675 314 744
rect 279 461 313 675
rect 276 427 313 461
rect 276 317 310 427
rect 31 47 561 62
rect 31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 276 47
rect 310 13 353 47
rect 387 13 425 47
rect 459 13 497 47
rect 531 13 561 47
rect 31 0 561 13
use pmos4  pmos4_0 pcells
timestamp 1645051079
transform 1 0 94 0 1 1228
box -36 -312 440 42
use poly_li1_contact_para  poly_li1_contact_para_0 pcells
timestamp 1645049503
transform 1 0 44 0 1 481
box 70 379 124 465
use diff_ring_side  diff_ring_side_1 pcells
timestamp 1645638419
transform 1 0 0 0 1 0
box -84 0 84 1353
use diff_ring_side  diff_ring_side_0
timestamp 1645638419
transform 1 0 592 0 1 0
box -84 0 84 1353
use li1_M1_contact_para_cent  li1_M1_contact_para_cent_0 pcells
timestamp 1645050557
transform 1 0 293 0 1 264
box -23 -33 23 53
use li1_M1_contact_perp_ext  li1_M1_contact_perp_ext_0 pcells
timestamp 1645050501
transform 1 0 296 0 1 944
box -23 -53 49 29
use nmos_top  nmos_top_0 pcells
timestamp 1645636714
transform -1 0 415 0 1 101
box -1 0 246 309
use poly_li1_contact_perp  poly_li1_contact_perp_0 pcells
timestamp 1645049645
transform -1 0 225 0 -1 896
box 44 399 110 481
<< labels >>
rlabel metal1 253 1325 253 1325 1 VDD
port 2 n
rlabel metal1 249 31 249 31 1 VSS
port 1 n
rlabel metal1 148 666 148 666 1 A
port 3 n
rlabel metal1 299 668 299 668 1 Y
port 4 n
<< end >>
