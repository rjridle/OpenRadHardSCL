magic
tech sky130A
magscale 1 2
timestamp 1651075983
<< nwell >>
rect 84 1554 363 1575
rect 31 1492 413 1554
rect 84 832 363 1492
<< pdiffc >>
rect 117 1106 151 1140
rect 205 1106 239 1140
rect 293 1106 327 1140
<< psubdiff >>
rect 17 510 427 572
rect 31 13 55 47
rect 89 13 127 47
rect 161 13 205 47
rect 239 13 283 47
rect 317 13 355 47
rect 389 13 413 47
<< nsubdiff >>
rect 31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 205 1539
rect 239 1505 283 1539
rect 317 1505 355 1539
rect 389 1505 413 1539
rect -31 868 475 930
<< psubdiffcont >>
rect 55 13 89 47
rect 127 13 161 47
rect 205 13 239 47
rect 283 13 317 47
rect 355 13 389 47
<< nsubdiffcont >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 205 1505 239 1539
rect 283 1505 317 1539
rect 355 1505 389 1539
<< poly >>
rect 155 409 185 441
<< locali >>
rect 31 1539 413 1554
rect 31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 205 1539
rect 239 1505 283 1539
rect 317 1505 355 1539
rect 389 1505 413 1539
rect 31 1492 413 1505
rect 117 1140 151 1157
rect 117 1062 151 1106
rect 205 1140 239 1157
rect 131 477 165 1003
rect 205 832 239 1106
rect 293 1140 327 1157
rect 293 1062 327 1106
rect 165 411 239 445
rect 205 262 239 411
rect 109 62 143 101
rect 205 62 239 117
rect 303 62 337 101
rect 31 47 413 62
rect 31 13 55 47
rect 89 13 127 47
rect 161 13 205 47
rect 239 13 283 47
rect 317 13 355 47
rect 389 13 413 47
rect 31 0 413 13
<< viali >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 205 1505 239 1539
rect 283 1505 317 1539
rect 355 1505 389 1539
rect 55 13 89 47
rect 127 13 161 47
rect 205 13 239 47
rect 283 13 317 47
rect 355 13 389 47
<< metal1 >>
rect -31 1539 475 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 205 1539
rect 239 1505 283 1539
rect 317 1505 355 1539
rect 389 1505 475 1539
rect -31 1492 475 1505
rect 205 797 239 831
rect -31 47 475 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 205 47
rect 239 13 283 47
rect 317 13 355 47
rect 389 13 475 47
rect -31 0 475 13
use nmos_top  nmos_top_0 pcells
timestamp 1648061425
transform -1 0 345 0 1 101
box 0 0 246 308
use pmos2  pmos2_0 pcells
timestamp 1648061063
transform 1 0 19 0 1 1450
box 52 -461 352 42
use diff_ring_side  diff_ring_side_1 pcells
timestamp 1648063806
transform 1 0 0 0 1 0
box -84 0 84 1575
use diff_ring_side  diff_ring_side_0
timestamp 1648063806
transform 1 0 444 0 1 0
box -84 0 84 1575
use poly_li1_contact  poly_li1_contact_1 pcells
timestamp 1648060378
transform 0 1 149 -1 0 445
box -32 -28 34 26
use li1_M1_contact  li1_M1_contact_0 pcells
timestamp 1648061256
transform -1 0 222 0 -1 814
box -53 -33 29 33
use poly_li1_contact  poly_li1_contact_0
timestamp 1648060378
transform 0 1 149 -1 0 987
box -32 -28 34 26
<< labels >>
rlabel metal1 205 797 239 831 1 Y
port 1 n
rlabel metal1 -31 1492 475 1554 1 VDD
rlabel metal1 -31 0 475 62 1 GND
<< end >>
