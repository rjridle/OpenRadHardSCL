* SPICE3 file created from TMRDFFRNQNX1.ext - technology: sky130A

.subckt TMRDFFRNQNX1 QN D CLK RN VDD GND
X0 VDD.t145 RN.t0 a_10507_187.t5 VDD.t144 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X1 GND a_10507_187.t7 a_10451_103.t0 GND sky130_fd_pr__nfet_01v8 ad=3.7611p pd=3.297u as=0p ps=0u w=0u l=0u
X2 a_14189_1050.t3 a_10637_1050.t7 VDD.t43 @�^a�U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X3 a_10959_989.t1 a_10637_1050.t8 VDD.t53 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X4 a_599_989.t3 D.t0 VDD.t3  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X5 a_16421_1051.t5 a_14511_989.t5 QN.t4 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X6 QN a_14511_989.t7 a_15652_101.t0 GND sky130_fd_pr__nfet_01v8 ad=5.373p pd=4.72u as=0p ps=0u w=0u l=0u
X7 a_5327_187.t6 CLK.t0 VDD.t151  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X8 VDD.t83 a_599_989.t7 a_2141_1050.t2 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X9 a_9331_989.t1 a_9009_1050.t7 VDD.t190  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X10 VDD.t99 CLK.t1 a_277_1050.t4 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X11 VDD.t51 a_5457_1050.t7 a_5779_989.t6  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X12 VDD.t6 a_5457_1050.t8 a_9009_1050.t0 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X13 VDD.t12 a_277_1050.t7 a_3829_1050.t6  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X14 VDD.t143 RN.t2 a_5779_989.t3 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X15 VDD.t70 a_9331_989.t5 a_9009_1050.t3  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X16 VDD.t81 CLK.t2 a_10507_187.t2 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X17 VDD.t188 CLK.t3 a_10637_1050.t6  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X18 a_9331_989.t4 a_5327_187.t7 VDD.t22 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X19 a_14189_1050.t5 RN.t3 VDD.t141  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X20 a_10959_989.t5 D.t2 VDD.t173 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X21 GND a_9331_989.t7 a_16318_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X22 a_599_989.t6 RN.t4 VDD.t139  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X23 a_3829_1050.t4 a_4151_989.t5 VDD.t103 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X24 VDD.t20 a_14511_989.t6 a_15757_1051.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X25 a_10637_1050.t5 a_10507_187.t8 VDD.t165 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X26 a_147_187.t6 CLK.t4 VDD.t194  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X27 a_4151_989.t1 a_3829_1050.t7 VDD.t32 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X28 GND a_5457_1050.t10 a_8823_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X29 a_9009_1050.t2 a_5457_1050.t9 VDD.t14  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X30 a_15757_1051.t3 a_9331_989.t6 VDD.t28 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X31 VDD.t204 a_14189_1050.t7 a_14511_989.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X32 VDD.t181 a_10959_989.t8 a_12501_1050.t1 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X33 GND a_5457_1050.t11 a_6233_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X34 VDD.t200 a_147_187.t9 a_2141_1050.t4  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X35 VDD.t169 a_599_989.t8 a_277_1050.t2 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X36 QN a_14511_989.t10 a_16984_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X37 VDD.t109 D.t4 a_5779_989.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X38 VDD.t137 RN.t6 a_9009_1050.t5 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X39 VDD.t167 a_2141_1050.t5 a_147_187.t4  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X40 VDD.t97 a_5327_187.t8 a_5457_1050.t6 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X41 VDD.t35 a_7321_1050.t5 a_5327_187.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X42 GND a_9009_1050.t9 a_9806_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X43 a_14189_1050.t1 a_14511_989.t8 VDD.t18 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X44 a_10959_989.t4 RN.t8 VDD.t135  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X45 a_147_187.t2 RN.t9 VDD.t133 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X46 GND a_5779_989.t8 a_7216_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X47 GND a_147_187.t12 a_91_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X48 GND a_7321_1050.t6 a_7861_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X49 a_4151_989.t3 a_147_187.t10 VDD.t74  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X50 a_7321_1050.t4 a_5327_187.t9 VDD.t1 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X51 QN.t6 a_4151_989.t6 a_16421_1051.t7  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X52 VDD.t38 a_10959_989.t9 a_10637_1050.t1 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X53 GND a_5327_187.t10 a_5271_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X54 a_15757_1051.t0 a_14511_989.t9 VDD.t47  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X55 VDD.t163 a_10507_187.t10 a_14511_989.t4 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X56 VDD.t161 a_10507_187.t11 a_12501_1050.t4  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X57 a_277_1050.t6 a_147_187.t11 VDD.t76 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X58 a_16421_1051.t1 a_4151_989.t7 a_15757_1051.t7  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X59 VDD.t196 a_9009_1050.t8 a_9331_989.t0 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X60 a_10507_187.t0 a_12501_1050.t5 VDD.t63  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X61 a_10507_187.t4 RN.t11 VDD.t131 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X62 a_10637_1050.t2 a_10959_989.t10 VDD.t65  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X63 a_7321_1050.t1 a_5779_989.t9 VDD.t153 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X64 VDD.t59 a_277_1050.t8 a_599_989.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X65 QN.t2 a_14511_989.t11 a_16421_1051.t4 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X66 VDD.t129 RN.t12 a_599_989.t5  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X67 VDD.t105 a_4151_989.t8 a_3829_1050.t3 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X68 GND a_12501_1050.t6 a_13041_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X69 QN a_4151_989.t10 a_16318_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X70 GND a_277_1050.t11 a_3643_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X71 VDD.t26 a_5779_989.t10 a_5457_1050.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X72 VDD.t127 RN.t14 a_5327_187.t4 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X73 a_16421_1051.t2 a_9331_989.t8 a_15757_1051.t5  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X74 a_2141_1050.t1 a_599_989.t10 VDD.t8 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X75 a_277_1050.t3 CLK.t7 VDD.t78  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X76 a_3829_1050.t5 a_277_1050.t9 VDD.t202 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X77 a_5779_989.t5 a_5457_1050.t12 VDD.t61  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X78 a_10507_187.t6 CLK.t8 VDD.t179 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X79 a_10637_1050.t0 CLK.t9 VDD.t10  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X80 VDD.t206 a_10637_1050.t10 a_14189_1050.t2 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X81 VDD.t87 a_10637_1050.t11 a_10959_989.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X82 GND a_3829_1050.t8 a_4626_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X83 VDD.t125 RN.t15 a_3829_1050.t1 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X84 VDD.t175 D.t6 a_599_989.t2  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X85 GND a_599_989.t12 a_2036_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X86 GND a_10637_1050.t12 a_14003_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X87 GND a_2141_1050.t7 a_2681_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X88 a_599_989.t0 a_277_1050.t10 VDD.t57 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X89 VDD.t45 CLK.t11 a_5457_1050.t4  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X90 VDD.t91 CLK.t12 a_5327_187.t2 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X91 a_2141_1050.t3 a_147_187.t13 VDD.t184  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X92 a_277_1050.t1 a_599_989.t11 VDD.t85 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X93 a_3829_1050.t0 RN.t16 VDD.t123  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X94 a_5779_989.t0 D.t7 VDD.t171 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X95 a_9009_1050.t4 RN.t17 VDD.t121  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X96 a_5327_187.t1 a_7321_1050.t7 VDD.t49 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X97 VDD.t89 a_5327_187.t12 a_9331_989.t3  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X98 GND a_9331_989.t11 a_15652_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X99 GND a_14189_1050.t8 a_14986_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X100 a_147_187.t3 a_2141_1050.t6 VDD.t107 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X101 a_5457_1050.t5 a_5327_187.t13 VDD.t95  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X102 VDD.t119 RN.t18 a_14189_1050.t4 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X103 VDD.t177 D.t8 a_10959_989.t6  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X104 VDD.t149 CLK.t14 a_147_187.t5 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X105 VDD.t93 a_5779_989.t11 a_7321_1050.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X106 VDD.t30 a_3829_1050.t9 a_4151_989.t0 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X107 VDD.t192 a_9331_989.t9 a_15757_1051.t2  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X108 GND a_277_1050.t12 a_1053_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X109 a_14511_989.t3 a_10507_187.t13 VDD.t159 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X110 a_12501_1050.t3 a_10507_187.t14 VDD.t157  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X111 a_9009_1050.t6 a_9331_989.t10 VDD.t198 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X112 a_5779_989.t2 RN.t21 VDD.t117  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X113 a_5457_1050.t3 CLK.t16 VDD.t147 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X114 a_15757_1051.t4 a_9331_989.t12 a_16421_1051.t6  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X115 VDD.t16 a_14511_989.t13 a_14189_1050.t0 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X116 GND a_4151_989.t13 a_16984_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X117 VDD.t115 RN.t23 a_147_187.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X118 VDD.t101 a_147_187.t14 a_4151_989.t2 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X119 VDD.t186 a_5327_187.t15 a_7321_1050.t3  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X120 a_16421_1051.t3 a_4151_989.t11 QN.t0 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X121 GND a_10637_1050.t9 a_11413_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X122 a_14511_989.t0 a_14189_1050.t9 VDD.t40  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X123 a_12501_1050.t0 a_10959_989.t12 VDD.t67 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X124 VDD.t113 RN.t25 a_10959_989.t3  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X125 a_5457_1050.t0 a_5779_989.t12 VDD.t24 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X126 a_5327_187.t3 RN.t26 VDD.t111  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X127 VDD.t55 a_147_187.t15 a_277_1050.t5 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X128 a_15757_1051.t6 a_4151_989.t12 a_16421_1051.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X129 GND a_10959_989.t7 a_12396_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X130 VDD.t155 a_10507_187.t15 a_10637_1050.t4 0ܪ{� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X131 VDD.t72 a_12501_1050.t7 a_10507_187.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
C0 CLK VDD 8.54fF
C1 D VDD 0.88fF
C2 RN VDD 2.66fF
C3 QN VDD 0.73fF
C4 CLK D 0.45fF
C5 CLK RN 1.13fF
C6 D RN 12.60fF
R0 RN.n17 RN.t15 479.223
R1 RN.n8 RN.t6 479.223
R2 RN.n0 RN.t18 479.223
R3 RN.n23 RN.t4 454.685
R4 RN.n20 RN.t9 454.685
R5 RN.n14 RN.t21 454.685
R6 RN.n11 RN.t26 454.685
R7 RN.n5 RN.t8 454.685
R8 RN.n2 RN.t11 454.685
R9 RN.n23 RN.t12 428.979
R10 RN.n20 RN.t23 428.979
R11 RN.n14 RN.t2 428.979
R12 RN.n11 RN.t14 428.979
R13 RN.n5 RN.t25 428.979
R14 RN.n2 RN.t0 428.979
R15 RN.n17 RN.t16 375.52
R16 RN.n8 RN.t17 375.52
R17 RN.n0 RN.t3 375.52
R18 RN.n24 RN.n23 254.865
R19 RN.n21 RN.n20 254.865
R20 RN.n15 RN.n14 254.865
R21 RN.n12 RN.n11 254.865
R22 RN.n6 RN.n5 254.865
R23 RN.n3 RN.n2 254.865
R24 RN.n18 RN.n17 252.188
R25 RN.n9 RN.n8 252.188
R26 RN.n1 RN.n0 252.188
R27 RN.n18 RN.t20 231.854
R28 RN.n9 RN.t7 231.854
R29 RN.n1 RN.t24 231.854
R30 RN.n24 RN.t19 228.106
R31 RN.n21 RN.t10 228.106
R32 RN.n15 RN.t5 228.106
R33 RN.n12 RN.t1 228.106
R34 RN.n6 RN.t22 228.106
R35 RN.n3 RN.t13 228.106
R36 RN.n10 RN.n7 10.293
R37 RN.n19 RN.n16 10.293
R38 RN.n4 RN.n1 7.325
R39 RN.n7 RN.n4 5.94
R40 RN.n16 RN.n13 5.94
R41 RN.n25 RN.n22 5.94
R42 RN.n4 RN.n3 4.65
R43 RN.n7 RN.n6 4.65
R44 RN.n10 RN.n9 4.65
R45 RN.n13 RN.n12 4.65
R46 RN.n16 RN.n15 4.65
R47 RN.n19 RN.n18 4.65
R48 RN.n22 RN.n21 4.65
R49 RN.n25 RN.n24 4.65
R50 RN.n13 RN.n10 2.675
R51 RN.n22 RN.n19 2.675
R52 RN.n25 RN 0.046
R53 a_10507_187.n10 a_10507_187.t15 512.525
R54 a_10507_187.n8 a_10507_187.t11 472.359
R55 a_10507_187.n6 a_10507_187.t10 472.359
R56 a_10507_187.n11 a_10507_187.t7 417.109
R57 a_10507_187.n8 a_10507_187.t14 384.527
R58 a_10507_187.n6 a_10507_187.t13 384.527
R59 a_10507_187.n10 a_10507_187.t8 371.139
R60 a_10507_187.n9 a_10507_187.t12 370.613
R61 a_10507_187.n7 a_10507_187.t9 370.613
R62 a_10507_187.n16 a_10507_187.n14 363.934
R63 a_10507_187.n11 a_10507_187.n10 179.837
R64 a_10507_187.n4 a_10507_187.n3 161.352
R65 a_10507_187.n9 a_10507_187.n8 127.096
R66 a_10507_187.n7 a_10507_187.n6 127.096
R67 a_10507_187.n14 a_10507_187.n5 123.481
R68 a_10507_187.n5 a_10507_187.n1 95.095
R69 a_10507_187.n4 a_10507_187.n2 95.095
R70 a_10507_187.n5 a_10507_187.n4 66.258
R71 a_10507_187.n16 a_10507_187.n15 30
R72 a_10507_187.n17 a_10507_187.n0 24.383
R73 a_10507_187.n17 a_10507_187.n16 23.684
R74 a_10507_187.n1 a_10507_187.t5 14.282
R75 a_10507_187.n1 a_10507_187.t4 14.282
R76 a_10507_187.n2 a_10507_187.t2 14.282
R77 a_10507_187.n2 a_10507_187.t6 14.282
R78 a_10507_187.n3 a_10507_187.t1 14.282
R79 a_10507_187.n3 a_10507_187.t0 14.282
R80 a_10507_187.n12 a_10507_187.n11 12.222
R81 a_10507_187.n13 a_10507_187.n7 10.046
R82 a_10507_187.n12 a_10507_187.n9 4.65
R83 a_10507_187.n14 a_10507_187.n13 4.65
R84 a_10507_187.n13 a_10507_187.n12 4.035
R85 VDD.n826 VDD.n815 144.705
R86 VDD.n901 VDD.n894 144.705
R87 VDD.n958 VDD.n951 144.705
R88 VDD.n1033 VDD.n1026 144.705
R89 VDD.n1108 VDD.n1101 144.705
R90 VDD.n1165 VDD.n1158 144.705
R91 VDD.n1240 VDD.n1233 144.705
R92 VDD.n1315 VDD.n1308 144.705
R93 VDD.n1372 VDD.n1365 144.705
R94 VDD.n656 VDD.n649 144.705
R95 VDD.n727 VDD.n720 144.705
R96 VDD.n599 VDD.n592 144.705
R97 VDD.n524 VDD.n517 144.705
R98 VDD.n449 VDD.n442 144.705
R99 VDD.n392 VDD.n385 144.705
R100 VDD.n317 VDD.n310 144.705
R101 VDD.n242 VDD.n235 144.705
R102 VDD.n185 VDD.n178 144.705
R103 VDD.n128 VDD.n121 144.705
R104 VDD.n75 VDD.n64 144.705
R105 VDD.n792 VDD.t169 143.754
R106 VDD.n868 VDD.t129 143.754
R107 VDD.n1000 VDD.t115 143.754
R108 VDD.n1075 VDD.t105 143.754
R109 VDD.n1207 VDD.t26 143.754
R110 VDD.n1282 VDD.t143 143.754
R111 VDD.n1414 VDD.t127 143.754
R112 VDD.n665 VDD.t70 143.754
R113 VDD.n533 VDD.t38 143.754
R114 VDD.n458 VDD.t113 143.754
R115 VDD.n326 VDD.t145 143.754
R116 VDD.n251 VDD.t16 143.754
R117 VDD.n926 VDD.t200 143.754
R118 VDD.n1133 VDD.t101 143.754
R119 VDD.n1340 VDD.t186 143.754
R120 VDD.n602 VDD.t89 143.754
R121 VDD.n395 VDD.t161 143.754
R122 VDD.n188 VDD.t163 143.754
R123 VDD.n153 VDD.t28 135.539
R124 VDD.n131 VDD.t20 135.539
R125 VDD.n757 VDD.t76 135.17
R126 VDD.n833 VDD.t57 135.17
R127 VDD.n904 VDD.t8 135.17
R128 VDD.n965 VDD.t107 135.17
R129 VDD.n1040 VDD.t202 135.17
R130 VDD.n1111 VDD.t32 135.17
R131 VDD.n1172 VDD.t95 135.17
R132 VDD.n1247 VDD.t61 135.17
R133 VDD.n1318 VDD.t153 135.17
R134 VDD.n1379 VDD.t49 135.17
R135 VDD.n695 VDD.t14 135.17
R136 VDD.n624 VDD.t190 135.17
R137 VDD.n563 VDD.t165 135.17
R138 VDD.n488 VDD.t53 135.17
R139 VDD.n417 VDD.t67 135.17
R140 VDD.n356 VDD.t63 135.17
R141 VDD.n281 VDD.t43 135.17
R142 VDD.n210 VDD.t40 135.17
R143 VDD.n141 VDD.n140 129.849
R144 VDD.n767 VDD.n766 129.472
R145 VDD.n783 VDD.n782 129.472
R146 VDD.n843 VDD.n842 129.472
R147 VDD.n859 VDD.n858 129.472
R148 VDD.n918 VDD.n917 129.472
R149 VDD.n975 VDD.n974 129.472
R150 VDD.n991 VDD.n990 129.472
R151 VDD.n1050 VDD.n1049 129.472
R152 VDD.n1066 VDD.n1065 129.472
R153 VDD.n1125 VDD.n1124 129.472
R154 VDD.n1182 VDD.n1181 129.472
R155 VDD.n1198 VDD.n1197 129.472
R156 VDD.n1257 VDD.n1256 129.472
R157 VDD.n1273 VDD.n1272 129.472
R158 VDD.n1332 VDD.n1331 129.472
R159 VDD.n1389 VDD.n1388 129.472
R160 VDD.n1405 VDD.n1404 129.472
R161 VDD.n686 VDD.n685 129.472
R162 VDD.n674 VDD.n673 129.472
R163 VDD.n612 VDD.n611 129.472
R164 VDD.n554 VDD.n553 129.472
R165 VDD.n542 VDD.n541 129.472
R166 VDD.n479 VDD.n478 129.472
R167 VDD.n467 VDD.n466 129.472
R168 VDD.n405 VDD.n404 129.472
R169 VDD.n347 VDD.n346 129.472
R170 VDD.n335 VDD.n334 129.472
R171 VDD.n272 VDD.n271 129.472
R172 VDD.n260 VDD.n259 129.472
R173 VDD.n198 VDD.n197 129.472
R174 VDD.n60 VDD.n59 92.5
R175 VDD.n58 VDD.n57 92.5
R176 VDD.n56 VDD.n55 92.5
R177 VDD.n54 VDD.n53 92.5
R178 VDD.n62 VDD.n61 92.5
R179 VDD.n117 VDD.n116 92.5
R180 VDD.n115 VDD.n114 92.5
R181 VDD.n113 VDD.n112 92.5
R182 VDD.n111 VDD.n110 92.5
R183 VDD.n119 VDD.n118 92.5
R184 VDD.n174 VDD.n173 92.5
R185 VDD.n172 VDD.n171 92.5
R186 VDD.n170 VDD.n169 92.5
R187 VDD.n168 VDD.n167 92.5
R188 VDD.n176 VDD.n175 92.5
R189 VDD.n231 VDD.n230 92.5
R190 VDD.n229 VDD.n228 92.5
R191 VDD.n227 VDD.n226 92.5
R192 VDD.n225 VDD.n224 92.5
R193 VDD.n233 VDD.n232 92.5
R194 VDD.n306 VDD.n305 92.5
R195 VDD.n304 VDD.n303 92.5
R196 VDD.n302 VDD.n301 92.5
R197 VDD.n300 VDD.n299 92.5
R198 VDD.n308 VDD.n307 92.5
R199 VDD.n381 VDD.n380 92.5
R200 VDD.n379 VDD.n378 92.5
R201 VDD.n377 VDD.n376 92.5
R202 VDD.n375 VDD.n374 92.5
R203 VDD.n383 VDD.n382 92.5
R204 VDD.n438 VDD.n437 92.5
R205 VDD.n436 VDD.n435 92.5
R206 VDD.n434 VDD.n433 92.5
R207 VDD.n432 VDD.n431 92.5
R208 VDD.n440 VDD.n439 92.5
R209 VDD.n513 VDD.n512 92.5
R210 VDD.n511 VDD.n510 92.5
R211 VDD.n509 VDD.n508 92.5
R212 VDD.n507 VDD.n506 92.5
R213 VDD.n515 VDD.n514 92.5
R214 VDD.n588 VDD.n587 92.5
R215 VDD.n586 VDD.n585 92.5
R216 VDD.n584 VDD.n583 92.5
R217 VDD.n582 VDD.n581 92.5
R218 VDD.n590 VDD.n589 92.5
R219 VDD.n645 VDD.n644 92.5
R220 VDD.n643 VDD.n642 92.5
R221 VDD.n641 VDD.n640 92.5
R222 VDD.n639 VDD.n638 92.5
R223 VDD.n647 VDD.n646 92.5
R224 VDD.n716 VDD.n715 92.5
R225 VDD.n714 VDD.n713 92.5
R226 VDD.n712 VDD.n711 92.5
R227 VDD.n710 VDD.n709 92.5
R228 VDD.n718 VDD.n717 92.5
R229 VDD.n1361 VDD.n1360 92.5
R230 VDD.n1359 VDD.n1358 92.5
R231 VDD.n1357 VDD.n1356 92.5
R232 VDD.n1355 VDD.n1354 92.5
R233 VDD.n1363 VDD.n1362 92.5
R234 VDD.n1304 VDD.n1303 92.5
R235 VDD.n1302 VDD.n1301 92.5
R236 VDD.n1300 VDD.n1299 92.5
R237 VDD.n1298 VDD.n1297 92.5
R238 VDD.n1306 VDD.n1305 92.5
R239 VDD.n1229 VDD.n1228 92.5
R240 VDD.n1227 VDD.n1226 92.5
R241 VDD.n1225 VDD.n1224 92.5
R242 VDD.n1223 VDD.n1222 92.5
R243 VDD.n1231 VDD.n1230 92.5
R244 VDD.n1154 VDD.n1153 92.5
R245 VDD.n1152 VDD.n1151 92.5
R246 VDD.n1150 VDD.n1149 92.5
R247 VDD.n1148 VDD.n1147 92.5
R248 VDD.n1156 VDD.n1155 92.5
R249 VDD.n1097 VDD.n1096 92.5
R250 VDD.n1095 VDD.n1094 92.5
R251 VDD.n1093 VDD.n1092 92.5
R252 VDD.n1091 VDD.n1090 92.5
R253 VDD.n1099 VDD.n1098 92.5
R254 VDD.n1022 VDD.n1021 92.5
R255 VDD.n1020 VDD.n1019 92.5
R256 VDD.n1018 VDD.n1017 92.5
R257 VDD.n1016 VDD.n1015 92.5
R258 VDD.n1024 VDD.n1023 92.5
R259 VDD.n947 VDD.n946 92.5
R260 VDD.n945 VDD.n944 92.5
R261 VDD.n943 VDD.n942 92.5
R262 VDD.n941 VDD.n940 92.5
R263 VDD.n949 VDD.n948 92.5
R264 VDD.n890 VDD.n889 92.5
R265 VDD.n888 VDD.n887 92.5
R266 VDD.n886 VDD.n885 92.5
R267 VDD.n884 VDD.n883 92.5
R268 VDD.n892 VDD.n891 92.5
R269 VDD.n811 VDD.n810 92.5
R270 VDD.n809 VDD.n808 92.5
R271 VDD.n807 VDD.n806 92.5
R272 VDD.n805 VDD.n804 92.5
R273 VDD.n813 VDD.n812 92.5
R274 VDD.n741 VDD.n740 92.5
R275 VDD.n739 VDD.n738 92.5
R276 VDD.n737 VDD.n736 92.5
R277 VDD.n735 VDD.n734 92.5
R278 VDD.n743 VDD.n742 92.5
R279 VDD.n14 VDD.n1 92.5
R280 VDD.n5 VDD.n4 92.5
R281 VDD.n7 VDD.n6 92.5
R282 VDD.n9 VDD.n8 92.5
R283 VDD.n11 VDD.n10 92.5
R284 VDD.n13 VDD.n12 92.5
R285 VDD.n21 VDD.n20 92.059
R286 VDD.n74 VDD.n73 92.059
R287 VDD.n127 VDD.n126 92.059
R288 VDD.n184 VDD.n183 92.059
R289 VDD.n241 VDD.n240 92.059
R290 VDD.n316 VDD.n315 92.059
R291 VDD.n391 VDD.n390 92.059
R292 VDD.n448 VDD.n447 92.059
R293 VDD.n523 VDD.n522 92.059
R294 VDD.n598 VDD.n597 92.059
R295 VDD.n655 VDD.n654 92.059
R296 VDD.n726 VDD.n725 92.059
R297 VDD.n1371 VDD.n1370 92.059
R298 VDD.n1314 VDD.n1313 92.059
R299 VDD.n1239 VDD.n1238 92.059
R300 VDD.n1164 VDD.n1163 92.059
R301 VDD.n1107 VDD.n1106 92.059
R302 VDD.n1032 VDD.n1031 92.059
R303 VDD.n957 VDD.n956 92.059
R304 VDD.n900 VDD.n899 92.059
R305 VDD.n825 VDD.n824 92.059
R306 VDD.n749 VDD.n748 92.059
R307 VDD.n20 VDD.n16 67.194
R308 VDD.n20 VDD.n17 67.194
R309 VDD.n20 VDD.n18 67.194
R310 VDD.n20 VDD.n19 67.194
R311 VDD.n733 VDD.n732 44.141
R312 VDD.n882 VDD.n881 44.141
R313 VDD.n939 VDD.n938 44.141
R314 VDD.n1014 VDD.n1013 44.141
R315 VDD.n1089 VDD.n1088 44.141
R316 VDD.n1146 VDD.n1145 44.141
R317 VDD.n1221 VDD.n1220 44.141
R318 VDD.n1296 VDD.n1295 44.141
R319 VDD.n1353 VDD.n1352 44.141
R320 VDD.n708 VDD.n707 44.141
R321 VDD.n637 VDD.n636 44.141
R322 VDD.n580 VDD.n579 44.141
R323 VDD.n505 VDD.n504 44.141
R324 VDD.n430 VDD.n429 44.141
R325 VDD.n373 VDD.n372 44.141
R326 VDD.n298 VDD.n297 44.141
R327 VDD.n223 VDD.n222 44.141
R328 VDD.n166 VDD.n165 44.141
R329 VDD.n109 VDD.n108 44.141
R330 VDD.n5 VDD.n3 44.141
R331 VDD.n881 VDD.n879 44.107
R332 VDD.n938 VDD.n936 44.107
R333 VDD.n1013 VDD.n1011 44.107
R334 VDD.n1088 VDD.n1086 44.107
R335 VDD.n1145 VDD.n1143 44.107
R336 VDD.n1220 VDD.n1218 44.107
R337 VDD.n1295 VDD.n1293 44.107
R338 VDD.n1352 VDD.n1350 44.107
R339 VDD.n707 VDD.n705 44.107
R340 VDD.n636 VDD.n634 44.107
R341 VDD.n579 VDD.n577 44.107
R342 VDD.n504 VDD.n502 44.107
R343 VDD.n429 VDD.n427 44.107
R344 VDD.n372 VDD.n370 44.107
R345 VDD.n297 VDD.n295 44.107
R346 VDD.n222 VDD.n220 44.107
R347 VDD.n165 VDD.n163 44.107
R348 VDD.n108 VDD.n106 44.107
R349 VDD.n732 VDD.n730 44.107
R350 VDD.n3 VDD.n2 44.107
R351 VDD.n20 VDD.n15 41.052
R352 VDD.n68 VDD.n66 39.742
R353 VDD.n68 VDD.n67 39.742
R354 VDD.n70 VDD.n69 39.742
R355 VDD.n123 VDD.n122 39.742
R356 VDD.n180 VDD.n179 39.742
R357 VDD.n237 VDD.n236 39.742
R358 VDD.n312 VDD.n311 39.742
R359 VDD.n387 VDD.n386 39.742
R360 VDD.n444 VDD.n443 39.742
R361 VDD.n519 VDD.n518 39.742
R362 VDD.n594 VDD.n593 39.742
R363 VDD.n651 VDD.n650 39.742
R364 VDD.n722 VDD.n721 39.742
R365 VDD.n1367 VDD.n1366 39.742
R366 VDD.n1310 VDD.n1309 39.742
R367 VDD.n1235 VDD.n1234 39.742
R368 VDD.n1160 VDD.n1159 39.742
R369 VDD.n1103 VDD.n1102 39.742
R370 VDD.n1028 VDD.n1027 39.742
R371 VDD.n953 VDD.n952 39.742
R372 VDD.n896 VDD.n895 39.742
R373 VDD.n745 VDD.n744 39.742
R374 VDD.n823 VDD.n820 39.742
R375 VDD.n823 VDD.n822 39.742
R376 VDD.n819 VDD.n818 39.742
R377 VDD.n108 VDD.n107 38
R378 VDD.n165 VDD.n164 38
R379 VDD.n222 VDD.n221 38
R380 VDD.n297 VDD.n296 38
R381 VDD.n372 VDD.n371 38
R382 VDD.n429 VDD.n428 38
R383 VDD.n504 VDD.n503 38
R384 VDD.n579 VDD.n578 38
R385 VDD.n636 VDD.n635 38
R386 VDD.n707 VDD.n706 38
R387 VDD.n1352 VDD.n1351 38
R388 VDD.n1295 VDD.n1294 38
R389 VDD.n1220 VDD.n1219 38
R390 VDD.n1145 VDD.n1144 38
R391 VDD.n1088 VDD.n1087 38
R392 VDD.n1013 VDD.n1012 38
R393 VDD.n938 VDD.n937 38
R394 VDD.n881 VDD.n880 38
R395 VDD.n732 VDD.n731 38
R396 VDD.n879 VDD.n878 36.774
R397 VDD.n936 VDD.n935 36.774
R398 VDD.n1011 VDD.n1010 36.774
R399 VDD.n1086 VDD.n1085 36.774
R400 VDD.n1143 VDD.n1142 36.774
R401 VDD.n1218 VDD.n1217 36.774
R402 VDD.n1293 VDD.n1292 36.774
R403 VDD.n1350 VDD.n1349 36.774
R404 VDD.n705 VDD.n704 36.774
R405 VDD.n634 VDD.n633 36.774
R406 VDD.n577 VDD.n576 36.774
R407 VDD.n502 VDD.n501 36.774
R408 VDD.n427 VDD.n426 36.774
R409 VDD.n370 VDD.n369 36.774
R410 VDD.n295 VDD.n294 36.774
R411 VDD.n220 VDD.n219 36.774
R412 VDD.n163 VDD.n162 36.774
R413 VDD.n106 VDD.n105 36.774
R414 VDD.n66 VDD.n65 36.774
R415 VDD.n822 VDD.n821 36.774
R416 VDD.n253 0ܪ{� 35.8
R417 VDD.n328 VDD.t144 35.8
R418 VDD.n460  35.8
R419 VDD.n535 0ܪ{� 35.8
R420 VDD.n667  35.8
R421 VDD.n1408 0ܪ{� 35.8
R422 VDD.n1276 0ܪ{� 35.8
R423 VDD.n1201  35.8
R424 VDD.n1069 0ܪ{� 35.8
R425 VDD.n994  35.8
R426 VDD.n862  35.8
R427 VDD.n786 0ܪ{� 35.8
R428 VDD.n277 �۪{� 33.243
R429 VDD.n352  33.243
R430 VDD.n484 0ܪ{� 33.243
R431 VDD.n559 0ܪ{� 33.243
R432 VDD.n691  33.243
R433 VDD.n1384 0ܪ{� 33.243
R434 VDD.n1252  33.243
R435 VDD.n1177  33.243
R436 VDD.n1045 0ܪ{� 33.243
R437 VDD.n970 0ܪ{� 33.243
R438 VDD.n838 0ܪ{� 33.243
R439 VDD.n762 0ܪ{� 33.243
R440 VDD.n1 VDD.n0 30.923
R441 VDD.n73 VDD.n71 26.38
R442 VDD.n73 VDD.n70 26.38
R443 VDD.n73 VDD.n68 26.38
R444 VDD.n73 VDD.n72 26.38
R445 VDD.n126 VDD.n124 26.38
R446 VDD.n126 VDD.n123 26.38
R447 VDD.n126 VDD.n125 26.38
R448 VDD.n183 VDD.n181 26.38
R449 VDD.n183 VDD.n180 26.38
R450 VDD.n183 VDD.n182 26.38
R451 VDD.n240 VDD.n238 26.38
R452 VDD.n240 VDD.n237 26.38
R453 VDD.n240 VDD.n239 26.38
R454 VDD.n315 VDD.n313 26.38
R455 VDD.n315 VDD.n312 26.38
R456 VDD.n315 VDD.n314 26.38
R457 VDD.n390 VDD.n388 26.38
R458 VDD.n390 VDD.n387 26.38
R459 VDD.n390 VDD.n389 26.38
R460 VDD.n447 VDD.n445 26.38
R461 VDD.n447 VDD.n444 26.38
R462 VDD.n447 VDD.n446 26.38
R463 VDD.n522 VDD.n520 26.38
R464 VDD.n522 VDD.n519 26.38
R465 VDD.n522 VDD.n521 26.38
R466 VDD.n597 VDD.n595 26.38
R467 VDD.n597 VDD.n594 26.38
R468 VDD.n597 VDD.n596 26.38
R469 VDD.n654 VDD.n652 26.38
R470 VDD.n654 VDD.n651 26.38
R471 VDD.n654 VDD.n653 26.38
R472 VDD.n725 VDD.n723 26.38
R473 VDD.n725 VDD.n722 26.38
R474 VDD.n725 VDD.n724 26.38
R475 VDD.n1370 VDD.n1368 26.38
R476 VDD.n1370 VDD.n1367 26.38
R477 VDD.n1370 VDD.n1369 26.38
R478 VDD.n1313 VDD.n1311 26.38
R479 VDD.n1313 VDD.n1310 26.38
R480 VDD.n1313 VDD.n1312 26.38
R481 VDD.n1238 VDD.n1236 26.38
R482 VDD.n1238 VDD.n1235 26.38
R483 VDD.n1238 VDD.n1237 26.38
R484 VDD.n1163 VDD.n1161 26.38
R485 VDD.n1163 VDD.n1160 26.38
R486 VDD.n1163 VDD.n1162 26.38
R487 VDD.n1106 VDD.n1104 26.38
R488 VDD.n1106 VDD.n1103 26.38
R489 VDD.n1106 VDD.n1105 26.38
R490 VDD.n1031 VDD.n1029 26.38
R491 VDD.n1031 VDD.n1028 26.38
R492 VDD.n1031 VDD.n1030 26.38
R493 VDD.n956 VDD.n954 26.38
R494 VDD.n956 VDD.n953 26.38
R495 VDD.n956 VDD.n955 26.38
R496 VDD.n899 VDD.n897 26.38
R497 VDD.n899 VDD.n896 26.38
R498 VDD.n899 VDD.n898 26.38
R499 VDD.n748 VDD.n746 26.38
R500 VDD.n748 VDD.n745 26.38
R501 VDD.n748 VDD.n747 26.38
R502 VDD.n824 VDD.n823 26.38
R503 VDD.n824 VDD.n819 26.38
R504 VDD.n824 VDD.n817 26.38
R505 VDD.n824 VDD.n816 26.38
R506 VDD.n751 VDD.n743 22.915
R507 VDD.n23 VDD.n14 22.915
R508 VDD.n28 0ܪ{� 20.457
R509 VDD.n93  20.457
R510 VDD.n136  20.457
R511 VDD.n193 0ܪ{� 20.457
R512 VDD.n400  20.457
R513 VDD.n607  20.457
R514 VDD.n1336  20.457
R515 VDD.n1129 0ܪ{� 20.457
R516 VDD.n922  20.457
R517 VDD.n39  17.9
R518 VDD.n82  17.9
R519 VDD.n149 0ܪ{� 17.9
R520 VDD.n206  17.9
R521 VDD.n413 0ܪ{� 17.9
R522 VDD.n620  17.9
R523 VDD.n1323 0ܪ{� 17.9
R524 VDD.n1116 0ܪ{� 17.9
R525 VDD.n909 0ܪ{� 17.9
R526 VDD.n257 0ܪ{� 15.343
R527 VDD.n332 0ܪ{� 15.343
R528 VDD.n464  15.343
R529 VDD.n539  15.343
R530 VDD.n671 0ܪ{� 15.343
R531 VDD.n1402  15.343
R532 VDD.n1270  15.343
R533 VDD.n1195 0ܪ{� 15.343
R534 VDD.n1063 0ܪ{� 15.343
R535 VDD.n988 0ܪ{� 15.343
R536 VDD.n856  15.343
R537 VDD.n780 0ܪ{� 15.343
R538 VDD.n743 VDD.n741 14.864
R539 VDD.n741 VDD.n739 14.864
R540 VDD.n739 VDD.n737 14.864
R541 VDD.n737 VDD.n735 14.864
R542 VDD.n735 VDD.n733 14.864
R543 VDD.n892 VDD.n890 14.864
R544 VDD.n890 VDD.n888 14.864
R545 VDD.n888 VDD.n886 14.864
R546 VDD.n886 VDD.n884 14.864
R547 VDD.n884 VDD.n882 14.864
R548 VDD.n949 VDD.n947 14.864
R549 VDD.n947 VDD.n945 14.864
R550 VDD.n945 VDD.n943 14.864
R551 VDD.n943 VDD.n941 14.864
R552 VDD.n941 VDD.n939 14.864
R553 VDD.n1024 VDD.n1022 14.864
R554 VDD.n1022 VDD.n1020 14.864
R555 VDD.n1020 VDD.n1018 14.864
R556 VDD.n1018 VDD.n1016 14.864
R557 VDD.n1016 VDD.n1014 14.864
R558 VDD.n1099 VDD.n1097 14.864
R559 VDD.n1097 VDD.n1095 14.864
R560 VDD.n1095 VDD.n1093 14.864
R561 VDD.n1093 VDD.n1091 14.864
R562 VDD.n1091 VDD.n1089 14.864
R563 VDD.n1156 VDD.n1154 14.864
R564 VDD.n1154 VDD.n1152 14.864
R565 VDD.n1152 VDD.n1150 14.864
R566 VDD.n1150 VDD.n1148 14.864
R567 VDD.n1148 VDD.n1146 14.864
R568 VDD.n1231 VDD.n1229 14.864
R569 VDD.n1229 VDD.n1227 14.864
R570 VDD.n1227 VDD.n1225 14.864
R571 VDD.n1225 VDD.n1223 14.864
R572 VDD.n1223 VDD.n1221 14.864
R573 VDD.n1306 VDD.n1304 14.864
R574 VDD.n1304 VDD.n1302 14.864
R575 VDD.n1302 VDD.n1300 14.864
R576 VDD.n1300 VDD.n1298 14.864
R577 VDD.n1298 VDD.n1296 14.864
R578 VDD.n1363 VDD.n1361 14.864
R579 VDD.n1361 VDD.n1359 14.864
R580 VDD.n1359 VDD.n1357 14.864
R581 VDD.n1357 VDD.n1355 14.864
R582 VDD.n1355 VDD.n1353 14.864
R583 VDD.n718 VDD.n716 14.864
R584 VDD.n716 VDD.n714 14.864
R585 VDD.n714 VDD.n712 14.864
R586 VDD.n712 VDD.n710 14.864
R587 VDD.n710 VDD.n708 14.864
R588 VDD.n647 VDD.n645 14.864
R589 VDD.n645 VDD.n643 14.864
R590 VDD.n643 VDD.n641 14.864
R591 VDD.n641 VDD.n639 14.864
R592 VDD.n639 VDD.n637 14.864
R593 VDD.n590 VDD.n588 14.864
R594 VDD.n588 VDD.n586 14.864
R595 VDD.n586 VDD.n584 14.864
R596 VDD.n584 VDD.n582 14.864
R597 VDD.n582 VDD.n580 14.864
R598 VDD.n515 VDD.n513 14.864
R599 VDD.n513 VDD.n511 14.864
R600 VDD.n511 VDD.n509 14.864
R601 VDD.n509 VDD.n507 14.864
R602 VDD.n507 VDD.n505 14.864
R603 VDD.n440 VDD.n438 14.864
R604 VDD.n438 VDD.n436 14.864
R605 VDD.n436 VDD.n434 14.864
R606 VDD.n434 VDD.n432 14.864
R607 VDD.n432 VDD.n430 14.864
R608 VDD.n383 VDD.n381 14.864
R609 VDD.n381 VDD.n379 14.864
R610 VDD.n379 VDD.n377 14.864
R611 VDD.n377 VDD.n375 14.864
R612 VDD.n375 VDD.n373 14.864
R613 VDD.n308 VDD.n306 14.864
R614 VDD.n306 VDD.n304 14.864
R615 VDD.n304 VDD.n302 14.864
R616 VDD.n302 VDD.n300 14.864
R617 VDD.n300 VDD.n298 14.864
R618 VDD.n233 VDD.n231 14.864
R619 VDD.n231 VDD.n229 14.864
R620 VDD.n229 VDD.n227 14.864
R621 VDD.n227 VDD.n225 14.864
R622 VDD.n225 VDD.n223 14.864
R623 VDD.n176 VDD.n174 14.864
R624 VDD.n174 VDD.n172 14.864
R625 VDD.n172 VDD.n170 14.864
R626 VDD.n170 VDD.n168 14.864
R627 VDD.n168 VDD.n166 14.864
R628 VDD.n119 VDD.n117 14.864
R629 VDD.n117 VDD.n115 14.864
R630 VDD.n115 VDD.n113 14.864
R631 VDD.n113 VDD.n111 14.864
R632 VDD.n111 VDD.n109 14.864
R633 VDD.n62 VDD.n60 14.864
R634 VDD.n60 VDD.n58 14.864
R635 VDD.n58 VDD.n56 14.864
R636 VDD.n56 VDD.n54 14.864
R637 VDD.n54 VDD.n52 14.864
R638 VDD.n52 VDD.n51 14.864
R639 VDD.n813 VDD.n811 14.864
R640 VDD.n811 VDD.n809 14.864
R641 VDD.n809 VDD.n807 14.864
R642 VDD.n807 VDD.n805 14.864
R643 VDD.n805 VDD.n803 14.864
R644 VDD.n803 VDD.n802 14.864
R645 VDD.n14 VDD.n13 14.864
R646 VDD.n13 VDD.n11 14.864
R647 VDD.n11 VDD.n9 14.864
R648 VDD.n9 VDD.n7 14.864
R649 VDD.n7 VDD.n5 14.864
R650 VDD.n76 VDD.n63 14.864
R651 VDD.n129 VDD.n120 14.864
R652 VDD.n186 VDD.n177 14.864
R653 VDD.n243 VDD.n234 14.864
R654 VDD.n318 VDD.n309 14.864
R655 VDD.n393 VDD.n384 14.864
R656 VDD.n450 VDD.n441 14.864
R657 VDD.n525 VDD.n516 14.864
R658 VDD.n600 VDD.n591 14.864
R659 VDD.n657 VDD.n648 14.864
R660 VDD.n728 VDD.n719 14.864
R661 VDD.n1373 VDD.n1364 14.864
R662 VDD.n1316 VDD.n1307 14.864
R663 VDD.n1241 VDD.n1232 14.864
R664 VDD.n1166 VDD.n1157 14.864
R665 VDD.n1109 VDD.n1100 14.864
R666 VDD.n1034 VDD.n1025 14.864
R667 VDD.n959 VDD.n950 14.864
R668 VDD.n902 VDD.n893 14.864
R669 VDD.n827 VDD.n814 14.864
R670 VDD.n766 VDD.t78 14.282
R671 VDD.n766 VDD.t55 14.282
R672 VDD.n782 VDD.t85 14.282
R673 VDD.n782 VDD.t99 14.282
R674 VDD.n842 VDD.t3 14.282
R675 VDD.n842 VDD.t59 14.282
R676 VDD.n858 VDD.t139 14.282
R677 VDD.n858 VDD.t175 14.282
R678 VDD.n917 VDD.t184 14.282
R679 VDD.n917 VDD.t83 14.282
R680 VDD.n974 VDD.t194 14.282
R681 VDD.n974 VDD.t167 14.282
R682 VDD.n990 VDD.t133 14.282
R683 VDD.n990 VDD.t149 14.282
R684 VDD.n1049 VDD.t123 14.282
R685 VDD.n1049 VDD.t12 14.282
R686 VDD.n1065 VDD.t103 14.282
R687 VDD.n1065 VDD.t125 14.282
R688 VDD.n1124 VDD.t74 14.282
R689 VDD.n1124 VDD.t30 14.282
R690 VDD.n1181 VDD.t147 14.282
R691 VDD.n1181 VDD.t97 14.282
R692 VDD.n1197 VDD.t24 14.282
R693 VDD.n1197 VDD.t45 14.282
R694 VDD.n1256 VDD.t171 14.282
R695 VDD.n1256 VDD.t51 14.282
R696 VDD.n1272 VDD.t117 14.282
R697 VDD.n1272 VDD.t109 14.282
R698 VDD.n1331 VDD.t1 14.282
R699 VDD.n1331 VDD.t93 14.282
R700 VDD.n1388 VDD.t151 14.282
R701 VDD.n1388 VDD.t35 14.282
R702 VDD.n1404 VDD.t111 14.282
R703 VDD.n1404 VDD.t91 14.282
R704 VDD.n685 VDD.t121 14.282
R705 VDD.n685 VDD.t6 14.282
R706 VDD.n673 VDD.t198 14.282
R707 VDD.n673 VDD.t137 14.282
R708 VDD.n611 VDD.t22 14.282
R709 VDD.n611 VDD.t196 14.282
R710 VDD.n553 VDD.t10 14.282
R711 VDD.n553 VDD.t155 14.282
R712 VDD.n541 VDD.t65 14.282
R713 VDD.n541 VDD.t188 14.282
R714 VDD.n478 VDD.t173 14.282
R715 VDD.n478 VDD.t87 14.282
R716 VDD.n466 VDD.t135 14.282
R717 VDD.n466 VDD.t177 14.282
R718 VDD.n404 VDD.t157 14.282
R719 VDD.n404 VDD.t181 14.282
R720 VDD.n346 VDD.t179 14.282
R721 VDD.n346 VDD.t72 14.282
R722 VDD.n334 VDD.t131 14.282
R723 VDD.n334 VDD.t81 14.282
R724 VDD.n271 VDD.t141 14.282
R725 VDD.n271 VDD.t206 14.282
R726 VDD.n259 VDD.t18 14.282
R727 VDD.n259 VDD.t119 14.282
R728 VDD.n197 VDD.t159 14.282
R729 VDD.n197 VDD.t204 14.282
R730 VDD.n140 VDD.t47 14.282
R731 VDD.n140 VDD.t192 14.282
R732 VDD.n273 0ܪ{� 12.786
R733 VDD.n348  12.786
R734 VDD.n480  12.786
R735 VDD.n555 0ܪ{� 12.786
R736 VDD.n687 0ܪ{� 12.786
R737 VDD.n1390  12.786
R738 VDD.n1258  12.786
R739 VDD.n1183 0ܪ{� 12.786
R740 VDD.n1051  12.786
R741 VDD.n976  12.786
R742 VDD.n844  12.786
R743 VDD.n768 0ܪ{� 12.786
R744 VDD.n143 VDD.n141 9.083
R745 VDD.n200 VDD.n198 9.083
R746 VDD.n407 VDD.n405 9.083
R747 VDD.n614 VDD.n612 9.083
R748 VDD.n1334 VDD.n1332 9.083
R749 VDD.n1127 VDD.n1125 9.083
R750 VDD.n920 VDD.n918 9.083
R751 VDD.n23 VDD.n22 8.855
R752 VDD.n22 VDD.n21 8.855
R753 VDD.n26 VDD.n25 8.855
R754 VDD.n25 VDD.n24 8.855
R755 VDD.n30 VDD.n29 8.855
R756 VDD.n29 VDD.n28 8.855
R757 VDD.n33 VDD.n32 8.855
R758 VDD.n32 0ܪ{� 8.855
R759 VDD.n37 VDD.n36 8.855
R760 VDD.n36 VDD.n35 8.855
R761 VDD.n41 VDD.n40 8.855
R762 VDD.n40 VDD.n39 8.855
R763 VDD.n45 VDD.n44 8.855
R764 VDD.n44 VDD.n43 8.855
R765 VDD.n49 VDD.n48 8.855
R766 VDD.n48 VDD.n47 8.855
R767 VDD.n76 VDD.n75 8.855
R768 VDD.n75 VDD.n74 8.855
R769 VDD.n80 VDD.n79 8.855
R770 VDD.n79 VDD.n78 8.855
R771 VDD.n84 VDD.n83 8.855
R772 VDD.n83 VDD.n82 8.855
R773 VDD.n88 VDD.n87 8.855
R774 VDD.n87 VDD.n86 8.855
R775 VDD.n91 VDD.n90 8.855
R776 VDD.n90  8.855
R777 VDD.n95 VDD.n94 8.855
R778 VDD.n94 VDD.n93 8.855
R779 VDD.n99 VDD.n98 8.855
R780 VDD.n98 VDD.n97 8.855
R781 VDD.n103 VDD.n102 8.855
R782 VDD.n102 VDD.n101 8.855
R783 VDD.n129 VDD.n128 8.855
R784 VDD.n128 VDD.n127 8.855
R785 VDD.n134 VDD.n133 8.855
R786 VDD.n133 VDD.n132 8.855
R787 VDD.n138 VDD.n137 8.855
R788 VDD.n137 VDD.n136 8.855
R789 VDD.n143 VDD.n142 8.855
R790 VDD.n142  8.855
R791 VDD.n147 VDD.n146 8.855
R792 VDD.n146 VDD.n145 8.855
R793 VDD.n151 VDD.n150 8.855
R794 VDD.n150 VDD.n149 8.855
R795 VDD.n156 VDD.n155 8.855
R796 VDD.n155 VDD.n154 8.855
R797 VDD.n160 VDD.n159 8.855
R798 VDD.n159 VDD.n158 8.855
R799 VDD.n186 VDD.n185 8.855
R800 VDD.n185 VDD.n184 8.855
R801 VDD.n191 VDD.n190 8.855
R802 VDD.n190 VDD.n189 8.855
R803 VDD.n195 VDD.n194 8.855
R804 VDD.n194 VDD.n193 8.855
R805 VDD.n200 VDD.n199 8.855
R806 VDD.n199 0ܪ{� 8.855
R807 VDD.n204 VDD.n203 8.855
R808 VDD.n203 VDD.n202 8.855
R809 VDD.n208 VDD.n207 8.855
R810 VDD.n207 VDD.n206 8.855
R811 VDD.n213 VDD.n212 8.855
R812 VDD.n212 VDD.n211 8.855
R813 VDD.n217 VDD.n216 8.855
R814 VDD.n216 VDD.n215 8.855
R815 VDD.n243 VDD.n242 8.855
R816 VDD.n242 VDD.n241 8.855
R817 VDD.n247 VDD.n246 8.855
R818 VDD.n246 VDD.n245 8.855
R819 VDD.n251 VDD.n250 8.855
R820 VDD.n250 VDD.n249 8.855
R821 VDD.n255 VDD.n254 8.855
R822 VDD.n254 VDD.n253 8.855
R823 VDD.n261 VDD.n258 8.855
R824 VDD.n258 VDD.n257 8.855
R825 VDD.n265 VDD.n264 8.855
R826 VDD.n264 VDD.n263 8.855
R827 VDD.n269 VDD.n268 8.855
R828 VDD.n268 VDD.n267 8.855
R829 VDD.n275 VDD.n274 8.855
R830 VDD.n274 VDD.n273 8.855
R831 VDD.n279 VDD.n278 8.855
R832 VDD.n278 VDD.n277 8.855
R833 VDD.n284 VDD.n283 8.855
R834 VDD.n283 VDD.n282 8.855
R835 VDD.n288 VDD.n287 8.855
R836 VDD.n287 VDD.n286 8.855
R837 VDD.n292 VDD.n291 8.855
R838 VDD.n291 VDD.n290 8.855
R839 VDD.n318 VDD.n317 8.855
R840 VDD.n317 VDD.n316 8.855
R841 VDD.n322 VDD.n321 8.855
R842 VDD.n321 VDD.n320 8.855
R843 VDD.n326 VDD.n325 8.855
R844 VDD.n325 VDD.n324 8.855
R845 VDD.n330 VDD.n329 8.855
R846 VDD.n329 VDD.n328 8.855
R847 VDD.n336 VDD.n333 8.855
R848 VDD.n333 VDD.n332 8.855
R849 VDD.n340 VDD.n339 8.855
R850 VDD.n339 VDD.n338 8.855
R851 VDD.n344 VDD.n343 8.855
R852 VDD.n343 VDD.n342 8.855
R853 VDD.n350 VDD.n349 8.855
R854 VDD.n349 VDD.n348 8.855
R855 VDD.n354 VDD.n353 8.855
R856 VDD.n353 VDD.n352 8.855
R857 VDD.n359 VDD.n358 8.855
R858 VDD.n358 VDD.n357 8.855
R859 VDD.n363 VDD.n362 8.855
R860 VDD.n362 VDD.n361 8.855
R861 VDD.n367 VDD.n366 8.855
R862 VDD.n366 VDD.n365 8.855
R863 VDD.n393 VDD.n392 8.855
R864 VDD.n392 VDD.n391 8.855
R865 VDD.n398 VDD.n397 8.855
R866 VDD.n397 VDD.n396 8.855
R867 VDD.n402 VDD.n401 8.855
R868 VDD.n401 VDD.n400 8.855
R869 VDD.n407 VDD.n406 8.855
R870 VDD.n406  8.855
R871 VDD.n411 VDD.n410 8.855
R872 VDD.n410 VDD.n409 8.855
R873 VDD.n415 VDD.n414 8.855
R874 VDD.n414 VDD.n413 8.855
R875 VDD.n420 VDD.n419 8.855
R876 VDD.n419 VDD.n418 8.855
R877 VDD.n424 VDD.n423 8.855
R878 VDD.n423 VDD.n422 8.855
R879 VDD.n450 VDD.n449 8.855
R880 VDD.n449 VDD.n448 8.855
R881 VDD.n454 VDD.n453 8.855
R882 VDD.n453 VDD.n452 8.855
R883 VDD.n458 VDD.n457 8.855
R884 VDD.n457 VDD.n456 8.855
R885 VDD.n462 VDD.n461 8.855
R886 VDD.n461 VDD.n460 8.855
R887 VDD.n468 VDD.n465 8.855
R888 VDD.n465 VDD.n464 8.855
R889 VDD.n472 VDD.n471 8.855
R890 VDD.n471 VDD.n470 8.855
R891 VDD.n476 VDD.n475 8.855
R892 VDD.n475 VDD.n474 8.855
R893 VDD.n482 VDD.n481 8.855
R894 VDD.n481 VDD.n480 8.855
R895 VDD.n486 VDD.n485 8.855
R896 VDD.n485 VDD.n484 8.855
R897 VDD.n491 VDD.n490 8.855
R898 VDD.n490 VDD.n489 8.855
R899 VDD.n495 VDD.n494 8.855
R900 VDD.n494 VDD.n493 8.855
R901 VDD.n499 VDD.n498 8.855
R902 VDD.n498 VDD.n497 8.855
R903 VDD.n525 VDD.n524 8.855
R904 VDD.n524 VDD.n523 8.855
R905 VDD.n529 VDD.n528 8.855
R906 VDD.n528 VDD.n527 8.855
R907 VDD.n533 VDD.n532 8.855
R908 VDD.n532 VDD.n531 8.855
R909 VDD.n537 VDD.n536 8.855
R910 VDD.n536 VDD.n535 8.855
R911 VDD.n543 VDD.n540 8.855
R912 VDD.n540 VDD.n539 8.855
R913 VDD.n547 VDD.n546 8.855
R914 VDD.n546 VDD.n545 8.855
R915 VDD.n551 VDD.n550 8.855
R916 VDD.n550 VDD.n549 8.855
R917 VDD.n557 VDD.n556 8.855
R918 VDD.n556 VDD.n555 8.855
R919 VDD.n561 VDD.n560 8.855
R920 VDD.n560 VDD.n559 8.855
R921 VDD.n566 VDD.n565 8.855
R922 VDD.n565 VDD.n564 8.855
R923 VDD.n570 VDD.n569 8.855
R924 VDD.n569 VDD.n568 8.855
R925 VDD.n574 VDD.n573 8.855
R926 VDD.n573 VDD.n572 8.855
R927 VDD.n600 VDD.n599 8.855
R928 VDD.n599 VDD.n598 8.855
R929 VDD.n605 VDD.n604 8.855
R930 VDD.n604 VDD.n603 8.855
R931 VDD.n609 VDD.n608 8.855
R932 VDD.n608 VDD.n607 8.855
R933 VDD.n614 VDD.n613 8.855
R934 VDD.n613 0ܪ{� 8.855
R935 VDD.n618 VDD.n617 8.855
R936 VDD.n617 VDD.n616 8.855
R937 VDD.n622 VDD.n621 8.855
R938 VDD.n621 VDD.n620 8.855
R939 VDD.n627 VDD.n626 8.855
R940 VDD.n626 VDD.n625 8.855
R941 VDD.n631 VDD.n630 8.855
R942 VDD.n630 VDD.n629 8.855
R943 VDD.n657 VDD.n656 8.855
R944 VDD.n656 VDD.n655 8.855
R945 VDD.n661 VDD.n660 8.855
R946 VDD.n660 VDD.n659 8.855
R947 VDD.n665 VDD.n664 8.855
R948 VDD.n664 VDD.n663 8.855
R949 VDD.n669 VDD.n668 8.855
R950 VDD.n668 VDD.n667 8.855
R951 VDD.n675 VDD.n672 8.855
R952 VDD.n672 VDD.n671 8.855
R953 VDD.n679 VDD.n678 8.855
R954 VDD.n678 VDD.n677 8.855
R955 VDD.n683 VDD.n682 8.855
R956 VDD.n682 VDD.n681 8.855
R957 VDD.n689 VDD.n688 8.855
R958 VDD.n688 VDD.n687 8.855
R959 VDD.n693 VDD.n692 8.855
R960 VDD.n692 VDD.n691 8.855
R961 VDD.n698 VDD.n697 8.855
R962 VDD.n697 VDD.n696 8.855
R963 VDD.n702 VDD.n701 8.855
R964 VDD.n701 VDD.n700 8.855
R965 VDD.n728 VDD.n727 8.855
R966 VDD.n727 VDD.n726 8.855
R967 VDD.n1422 VDD.n1421 8.855
R968 VDD.n1421 VDD.n1420 8.855
R969 VDD.n1418 VDD.n1417 8.855
R970 VDD.n1417 VDD.n1416 8.855
R971 VDD.n1414 VDD.n1413 8.855
R972 VDD.n1413 VDD.n1412 8.855
R973 VDD.n1410 VDD.n1409 8.855
R974 VDD.n1409 VDD.n1408 8.855
R975 VDD.n1406 VDD.n1403 8.855
R976 VDD.n1403 VDD.n1402 8.855
R977 VDD.n1400 VDD.n1399 8.855
R978 VDD.n1399 VDD.n1398 8.855
R979 VDD.n1396 VDD.n1395 8.855
R980 VDD.n1395 VDD.n1394 8.855
R981 VDD.n1392 VDD.n1391 8.855
R982 VDD.n1391 VDD.n1390 8.855
R983 VDD.n1386 VDD.n1385 8.855
R984 VDD.n1385 VDD.n1384 8.855
R985 VDD.n1382 VDD.n1381 8.855
R986 VDD.n1381 VDD.n1380 8.855
R987 VDD.n1377 VDD.n1376 8.855
R988 VDD.n1376 VDD.n1375 8.855
R989 VDD.n1373 VDD.n1372 8.855
R990 VDD.n1372 VDD.n1371 8.855
R991 VDD.n1347 VDD.n1346 8.855
R992 VDD.n1346 VDD.n1345 8.855
R993 VDD.n1343 VDD.n1342 8.855
R994 VDD.n1342 VDD.n1341 8.855
R995 VDD.n1338 VDD.n1337 8.855
R996 VDD.n1337 VDD.n1336 8.855
R997 VDD.n1334 VDD.n1333 8.855
R998 VDD.n1333 0ܪ{� 8.855
R999 VDD.n1329 VDD.n1328 8.855
R1000 VDD.n1328 VDD.n1327 8.855
R1001 VDD.n1325 VDD.n1324 8.855
R1002 VDD.n1324 VDD.n1323 8.855
R1003 VDD.n1321 VDD.n1320 8.855
R1004 VDD.n1320 VDD.n1319 8.855
R1005 VDD.n1316 VDD.n1315 8.855
R1006 VDD.n1315 VDD.n1314 8.855
R1007 VDD.n1290 VDD.n1289 8.855
R1008 VDD.n1289 VDD.n1288 8.855
R1009 VDD.n1286 VDD.n1285 8.855
R1010 VDD.n1285 VDD.n1284 8.855
R1011 VDD.n1282 VDD.n1281 8.855
R1012 VDD.n1281 VDD.n1280 8.855
R1013 VDD.n1278 VDD.n1277 8.855
R1014 VDD.n1277 VDD.n1276 8.855
R1015 VDD.n1274 VDD.n1271 8.855
R1016 VDD.n1271 VDD.n1270 8.855
R1017 VDD.n1268 VDD.n1267 8.855
R1018 VDD.n1267 VDD.n1266 8.855
R1019 VDD.n1264 VDD.n1263 8.855
R1020 VDD.n1263 VDD.n1262 8.855
R1021 VDD.n1260 VDD.n1259 8.855
R1022 VDD.n1259 VDD.n1258 8.855
R1023 VDD.n1254 VDD.n1253 8.855
R1024 VDD.n1253 VDD.n1252 8.855
R1025 VDD.n1250 VDD.n1249 8.855
R1026 VDD.n1249 VDD.n1248 8.855
R1027 VDD.n1245 VDD.n1244 8.855
R1028 VDD.n1244 VDD.n1243 8.855
R1029 VDD.n1241 VDD.n1240 8.855
R1030 VDD.n1240 VDD.n1239 8.855
R1031 VDD.n1215 VDD.n1214 8.855
R1032 VDD.n1214 VDD.n1213 8.855
R1033 VDD.n1211 VDD.n1210 8.855
R1034 VDD.n1210 VDD.n1209 8.855
R1035 VDD.n1207 VDD.n1206 8.855
R1036 VDD.n1206 VDD.n1205 8.855
R1037 VDD.n1203 VDD.n1202 8.855
R1038 VDD.n1202 VDD.n1201 8.855
R1039 VDD.n1199 VDD.n1196 8.855
R1040 VDD.n1196 VDD.n1195 8.855
R1041 VDD.n1193 VDD.n1192 8.855
R1042 VDD.n1192 VDD.n1191 8.855
R1043 VDD.n1189 VDD.n1188 8.855
R1044 VDD.n1188 VDD.n1187 8.855
R1045 VDD.n1185 VDD.n1184 8.855
R1046 VDD.n1184 VDD.n1183 8.855
R1047 VDD.n1179 VDD.n1178 8.855
R1048 VDD.n1178 VDD.n1177 8.855
R1049 VDD.n1175 VDD.n1174 8.855
R1050 VDD.n1174 VDD.n1173 8.855
R1051 VDD.n1170 VDD.n1169 8.855
R1052 VDD.n1169 VDD.n1168 8.855
R1053 VDD.n1166 VDD.n1165 8.855
R1054 VDD.n1165 VDD.n1164 8.855
R1055 VDD.n1140 VDD.n1139 8.855
R1056 VDD.n1139 VDD.n1138 8.855
R1057 VDD.n1136 VDD.n1135 8.855
R1058 VDD.n1135 VDD.n1134 8.855
R1059 VDD.n1131 VDD.n1130 8.855
R1060 VDD.n1130 VDD.n1129 8.855
R1061 VDD.n1127 VDD.n1126 8.855
R1062 VDD.n1126  8.855
R1063 VDD.n1122 VDD.n1121 8.855
R1064 VDD.n1121 VDD.n1120 8.855
R1065 VDD.n1118 VDD.n1117 8.855
R1066 VDD.n1117 VDD.n1116 8.855
R1067 VDD.n1114 VDD.n1113 8.855
R1068 VDD.n1113 VDD.n1112 8.855
R1069 VDD.n1109 VDD.n1108 8.855
R1070 VDD.n1108 VDD.n1107 8.855
R1071 VDD.n1083 VDD.n1082 8.855
R1072 VDD.n1082 VDD.n1081 8.855
R1073 VDD.n1079 VDD.n1078 8.855
R1074 VDD.n1078 VDD.n1077 8.855
R1075 VDD.n1075 VDD.n1074 8.855
R1076 VDD.n1074 VDD.n1073 8.855
R1077 VDD.n1071 VDD.n1070 8.855
R1078 VDD.n1070 VDD.n1069 8.855
R1079 VDD.n1067 VDD.n1064 8.855
R1080 VDD.n1064 VDD.n1063 8.855
R1081 VDD.n1061 VDD.n1060 8.855
R1082 VDD.n1060 VDD.n1059 8.855
R1083 VDD.n1057 VDD.n1056 8.855
R1084 VDD.n1056 VDD.n1055 8.855
R1085 VDD.n1053 VDD.n1052 8.855
R1086 VDD.n1052 VDD.n1051 8.855
R1087 VDD.n1047 VDD.n1046 8.855
R1088 VDD.n1046 VDD.n1045 8.855
R1089 VDD.n1043 VDD.n1042 8.855
R1090 VDD.n1042 VDD.n1041 8.855
R1091 VDD.n1038 VDD.n1037 8.855
R1092 VDD.n1037 VDD.n1036 8.855
R1093 VDD.n1034 VDD.n1033 8.855
R1094 VDD.n1033 VDD.n1032 8.855
R1095 VDD.n1008 VDD.n1007 8.855
R1096 VDD.n1007 VDD.n1006 8.855
R1097 VDD.n1004 VDD.n1003 8.855
R1098 VDD.n1003 VDD.n1002 8.855
R1099 VDD.n1000 VDD.n999 8.855
R1100 VDD.n999 VDD.n998 8.855
R1101 VDD.n996 VDD.n995 8.855
R1102 VDD.n995 VDD.n994 8.855
R1103 VDD.n992 VDD.n989 8.855
R1104 VDD.n989 VDD.n988 8.855
R1105 VDD.n986 VDD.n985 8.855
R1106 VDD.n985 VDD.n984 8.855
R1107 VDD.n982 VDD.n981 8.855
R1108 VDD.n981 VDD.n980 8.855
R1109 VDD.n978 VDD.n977 8.855
R1110 VDD.n977 VDD.n976 8.855
R1111 VDD.n972 VDD.n971 8.855
R1112 VDD.n971 VDD.n970 8.855
R1113 VDD.n968 VDD.n967 8.855
R1114 VDD.n967 VDD.n966 8.855
R1115 VDD.n963 VDD.n962 8.855
R1116 VDD.n962 VDD.n961 8.855
R1117 VDD.n959 VDD.n958 8.855
R1118 VDD.n958 VDD.n957 8.855
R1119 VDD.n933 VDD.n932 8.855
R1120 VDD.n932 VDD.n931 8.855
R1121 VDD.n929 VDD.n928 8.855
R1122 VDD.n928 VDD.n927 8.855
R1123 VDD.n924 VDD.n923 8.855
R1124 VDD.n923 VDD.n922 8.855
R1125 VDD.n920 VDD.n919 8.855
R1126 VDD.n919  8.855
R1127 VDD.n915 VDD.n914 8.855
R1128 VDD.n914 VDD.n913 8.855
R1129 VDD.n911 VDD.n910 8.855
R1130 VDD.n910 VDD.n909 8.855
R1131 VDD.n907 VDD.n906 8.855
R1132 VDD.n906 VDD.n905 8.855
R1133 VDD.n902 VDD.n901 8.855
R1134 VDD.n901 VDD.n900 8.855
R1135 VDD.n876 VDD.n875 8.855
R1136 VDD.n875 VDD.n874 8.855
R1137 VDD.n872 VDD.n871 8.855
R1138 VDD.n871 VDD.n870 8.855
R1139 VDD.n868 VDD.n867 8.855
R1140 VDD.n867 VDD.n866 8.855
R1141 VDD.n864 VDD.n863 8.855
R1142 VDD.n863 VDD.n862 8.855
R1143 VDD.n860 VDD.n857 8.855
R1144 VDD.n857 VDD.n856 8.855
R1145 VDD.n854 VDD.n853 8.855
R1146 VDD.n853 VDD.n852 8.855
R1147 VDD.n850 VDD.n849 8.855
R1148 VDD.n849 VDD.n848 8.855
R1149 VDD.n846 VDD.n845 8.855
R1150 VDD.n845 VDD.n844 8.855
R1151 VDD.n840 VDD.n839 8.855
R1152 VDD.n839 VDD.n838 8.855
R1153 VDD.n836 VDD.n835 8.855
R1154 VDD.n835 VDD.n834 8.855
R1155 VDD.n831 VDD.n830 8.855
R1156 VDD.n830 VDD.n829 8.855
R1157 VDD.n827 VDD.n826 8.855
R1158 VDD.n826 VDD.n825 8.855
R1159 VDD.n800 VDD.n799 8.855
R1160 VDD.n799 VDD.n798 8.855
R1161 VDD.n796 VDD.n795 8.855
R1162 VDD.n795 VDD.n794 8.855
R1163 VDD.n792 VDD.n791 8.855
R1164 VDD.n791 VDD.n790 8.855
R1165 VDD.n788 VDD.n787 8.855
R1166 VDD.n787 VDD.n786 8.855
R1167 VDD.n784 VDD.n781 8.855
R1168 VDD.n781 VDD.n780 8.855
R1169 VDD.n778 VDD.n777 8.855
R1170 VDD.n777 VDD.n776 8.855
R1171 VDD.n774 VDD.n773 8.855
R1172 VDD.n773 VDD.n772 8.855
R1173 VDD.n770 VDD.n769 8.855
R1174 VDD.n769 VDD.n768 8.855
R1175 VDD.n764 VDD.n763 8.855
R1176 VDD.n763 VDD.n762 8.855
R1177 VDD.n760 VDD.n759 8.855
R1178 VDD.n759 VDD.n758 8.855
R1179 VDD.n755 VDD.n754 8.855
R1180 VDD.n754 VDD.n753 8.855
R1181 VDD.n751 VDD.n750 8.855
R1182 VDD.n750 VDD.n749 8.855
R1183 VDD.n893 VDD.n892 8.051
R1184 VDD.n950 VDD.n949 8.051
R1185 VDD.n1025 VDD.n1024 8.051
R1186 VDD.n1100 VDD.n1099 8.051
R1187 VDD.n1157 VDD.n1156 8.051
R1188 VDD.n1232 VDD.n1231 8.051
R1189 VDD.n1307 VDD.n1306 8.051
R1190 VDD.n1364 VDD.n1363 8.051
R1191 VDD.n719 VDD.n718 8.051
R1192 VDD.n648 VDD.n647 8.051
R1193 VDD.n591 VDD.n590 8.051
R1194 VDD.n516 VDD.n515 8.051
R1195 VDD.n441 VDD.n440 8.051
R1196 VDD.n384 VDD.n383 8.051
R1197 VDD.n309 VDD.n308 8.051
R1198 VDD.n234 VDD.n233 8.051
R1199 VDD.n177 VDD.n176 8.051
R1200 VDD.n120 VDD.n119 8.051
R1201 VDD.n63 VDD.n62 8.051
R1202 VDD.n814 VDD.n813 8.051
R1203 VDD.n267  7.671
R1204 VDD.n342 0ܪ{� 7.671
R1205 VDD.n474 0ܪ{� 7.671
R1206 VDD.n549  7.671
R1207 VDD.n681  7.671
R1208 VDD.n1394  7.671
R1209 VDD.n1262 0ܪ{� 7.671
R1210 VDD.n1187 0ܪ{� 7.671
R1211 VDD.n1055  7.671
R1212 VDD.n980  7.671
R1213 VDD.n848  7.671
R1214 VDD.n772  7.671
R1215 VDD.n275 VDD.n272 7.019
R1216 VDD.n350 VDD.n347 7.019
R1217 VDD.n482 VDD.n479 7.019
R1218 VDD.n557 VDD.n554 7.019
R1219 VDD.n689 VDD.n686 7.019
R1220 VDD.n1392 VDD.n1389 7.019
R1221 VDD.n1260 VDD.n1257 7.019
R1222 VDD.n1185 VDD.n1182 7.019
R1223 VDD.n1053 VDD.n1050 7.019
R1224 VDD.n978 VDD.n975 7.019
R1225 VDD.n846 VDD.n843 7.019
R1226 VDD.n770 VDD.n767 7.019
R1227 VDD.n261 VDD.n260 6.606
R1228 VDD.n336 VDD.n335 6.606
R1229 VDD.n468 VDD.n467 6.606
R1230 VDD.n543 VDD.n542 6.606
R1231 VDD.n675 VDD.n674 6.606
R1232 VDD.n1406 VDD.n1405 6.606
R1233 VDD.n1274 VDD.n1273 6.606
R1234 VDD.n1199 VDD.n1198 6.606
R1235 VDD.n1067 VDD.n1066 6.606
R1236 VDD.n992 VDD.n991 6.606
R1237 VDD.n860 VDD.n859 6.606
R1238 VDD.n784 VDD.n783 6.606
R1239 VDD.n263 0ܪ{� 5.114
R1240 VDD.n338 0ܪ{� 5.114
R1241 VDD.n470  5.114
R1242 VDD.n545  5.114
R1243 VDD.n677 0ܪ{� 5.114
R1244 VDD.n1398 0ܪ{� 5.114
R1245 VDD.n1266  5.114
R1246 VDD.n1191  5.114
R1247 VDD.n1059 0ܪ{� 5.114
R1248 VDD.n984 0ܪ{� 5.114
R1249 VDD.n852  5.114
R1250 VDD.n776 0ܪ{� 5.114
R1251 VDD.n31 VDD.n30 4.65
R1252 VDD.n34 VDD.n33 4.65
R1253 VDD.n38 VDD.n37 4.65
R1254 VDD.n42 VDD.n41 4.65
R1255 VDD.n46 VDD.n45 4.65
R1256 VDD.n50 VDD.n49 4.65
R1257 VDD.n77 VDD.n76 4.65
R1258 VDD.n81 VDD.n80 4.65
R1259 VDD.n85 VDD.n84 4.65
R1260 VDD.n89 VDD.n88 4.65
R1261 VDD.n92 VDD.n91 4.65
R1262 VDD.n96 VDD.n95 4.65
R1263 VDD.n100 VDD.n99 4.65
R1264 VDD.n104 VDD.n103 4.65
R1265 VDD.n130 VDD.n129 4.65
R1266 VDD.n135 VDD.n134 4.65
R1267 VDD.n139 VDD.n138 4.65
R1268 VDD.n144 VDD.n143 4.65
R1269 VDD.n148 VDD.n147 4.65
R1270 VDD.n152 VDD.n151 4.65
R1271 VDD.n157 VDD.n156 4.65
R1272 VDD.n161 VDD.n160 4.65
R1273 VDD.n187 VDD.n186 4.65
R1274 VDD.n192 VDD.n191 4.65
R1275 VDD.n196 VDD.n195 4.65
R1276 VDD.n201 VDD.n200 4.65
R1277 VDD.n205 VDD.n204 4.65
R1278 VDD.n209 VDD.n208 4.65
R1279 VDD.n214 VDD.n213 4.65
R1280 VDD.n218 VDD.n217 4.65
R1281 VDD.n244 VDD.n243 4.65
R1282 VDD.n248 VDD.n247 4.65
R1283 VDD.n252 VDD.n251 4.65
R1284 VDD.n256 VDD.n255 4.65
R1285 VDD.n262 VDD.n261 4.65
R1286 VDD.n266 VDD.n265 4.65
R1287 VDD.n270 VDD.n269 4.65
R1288 VDD.n276 VDD.n275 4.65
R1289 VDD.n280 VDD.n279 4.65
R1290 VDD.n285 VDD.n284 4.65
R1291 VDD.n289 VDD.n288 4.65
R1292 VDD.n293 VDD.n292 4.65
R1293 VDD.n319 VDD.n318 4.65
R1294 VDD.n323 VDD.n322 4.65
R1295 VDD.n327 VDD.n326 4.65
R1296 VDD.n331 VDD.n330 4.65
R1297 VDD.n337 VDD.n336 4.65
R1298 VDD.n341 VDD.n340 4.65
R1299 VDD.n345 VDD.n344 4.65
R1300 VDD.n351 VDD.n350 4.65
R1301 VDD.n355 VDD.n354 4.65
R1302 VDD.n360 VDD.n359 4.65
R1303 VDD.n364 VDD.n363 4.65
R1304 VDD.n368 VDD.n367 4.65
R1305 VDD.n394 VDD.n393 4.65
R1306 VDD.n399 VDD.n398 4.65
R1307 VDD.n403 VDD.n402 4.65
R1308 VDD.n408 VDD.n407 4.65
R1309 VDD.n412 VDD.n411 4.65
R1310 VDD.n416 VDD.n415 4.65
R1311 VDD.n421 VDD.n420 4.65
R1312 VDD.n425 VDD.n424 4.65
R1313 VDD.n451 VDD.n450 4.65
R1314 VDD.n455 VDD.n454 4.65
R1315 VDD.n459 VDD.n458 4.65
R1316 VDD.n463 VDD.n462 4.65
R1317 VDD.n469 VDD.n468 4.65
R1318 VDD.n473 VDD.n472 4.65
R1319 VDD.n477 VDD.n476 4.65
R1320 VDD.n483 VDD.n482 4.65
R1321 VDD.n487 VDD.n486 4.65
R1322 VDD.n492 VDD.n491 4.65
R1323 VDD.n496 VDD.n495 4.65
R1324 VDD.n500 VDD.n499 4.65
R1325 VDD.n526 VDD.n525 4.65
R1326 VDD.n530 VDD.n529 4.65
R1327 VDD.n534 VDD.n533 4.65
R1328 VDD.n538 VDD.n537 4.65
R1329 VDD.n544 VDD.n543 4.65
R1330 VDD.n548 VDD.n547 4.65
R1331 VDD.n552 VDD.n551 4.65
R1332 VDD.n558 VDD.n557 4.65
R1333 VDD.n562 VDD.n561 4.65
R1334 VDD.n567 VDD.n566 4.65
R1335 VDD.n571 VDD.n570 4.65
R1336 VDD.n575 VDD.n574 4.65
R1337 VDD.n601 VDD.n600 4.65
R1338 VDD.n606 VDD.n605 4.65
R1339 VDD.n610 VDD.n609 4.65
R1340 VDD.n615 VDD.n614 4.65
R1341 VDD.n619 VDD.n618 4.65
R1342 VDD.n623 VDD.n622 4.65
R1343 VDD.n628 VDD.n627 4.65
R1344 VDD.n632 VDD.n631 4.65
R1345 VDD.n658 VDD.n657 4.65
R1346 VDD.n662 VDD.n661 4.65
R1347 VDD.n666 VDD.n665 4.65
R1348 VDD.n670 VDD.n669 4.65
R1349 VDD.n676 VDD.n675 4.65
R1350 VDD.n680 VDD.n679 4.65
R1351 VDD.n684 VDD.n683 4.65
R1352 VDD.n690 VDD.n689 4.65
R1353 VDD.n694 VDD.n693 4.65
R1354 VDD.n699 VDD.n698 4.65
R1355 VDD.n703 VDD.n702 4.65
R1356 VDD.n729 VDD.n728 4.65
R1357 VDD.n1423 VDD.n1422 4.65
R1358 VDD.n1419 VDD.n1418 4.65
R1359 VDD.n1415 VDD.n1414 4.65
R1360 VDD.n1411 VDD.n1410 4.65
R1361 VDD.n1407 VDD.n1406 4.65
R1362 VDD.n1401 VDD.n1400 4.65
R1363 VDD.n1397 VDD.n1396 4.65
R1364 VDD.n1393 VDD.n1392 4.65
R1365 VDD.n1387 VDD.n1386 4.65
R1366 VDD.n1383 VDD.n1382 4.65
R1367 VDD.n1378 VDD.n1377 4.65
R1368 VDD.n1374 VDD.n1373 4.65
R1369 VDD.n1348 VDD.n1347 4.65
R1370 VDD.n1344 VDD.n1343 4.65
R1371 VDD.n1339 VDD.n1338 4.65
R1372 VDD.n1335 VDD.n1334 4.65
R1373 VDD.n1330 VDD.n1329 4.65
R1374 VDD.n1326 VDD.n1325 4.65
R1375 VDD.n1322 VDD.n1321 4.65
R1376 VDD.n1317 VDD.n1316 4.65
R1377 VDD.n1291 VDD.n1290 4.65
R1378 VDD.n1287 VDD.n1286 4.65
R1379 VDD.n1283 VDD.n1282 4.65
R1380 VDD.n1279 VDD.n1278 4.65
R1381 VDD.n1275 VDD.n1274 4.65
R1382 VDD.n1269 VDD.n1268 4.65
R1383 VDD.n1265 VDD.n1264 4.65
R1384 VDD.n1261 VDD.n1260 4.65
R1385 VDD.n1255 VDD.n1254 4.65
R1386 VDD.n1251 VDD.n1250 4.65
R1387 VDD.n1246 VDD.n1245 4.65
R1388 VDD.n1242 VDD.n1241 4.65
R1389 VDD.n1216 VDD.n1215 4.65
R1390 VDD.n1212 VDD.n1211 4.65
R1391 VDD.n1208 VDD.n1207 4.65
R1392 VDD.n1204 VDD.n1203 4.65
R1393 VDD.n1200 VDD.n1199 4.65
R1394 VDD.n1194 VDD.n1193 4.65
R1395 VDD.n1190 VDD.n1189 4.65
R1396 VDD.n1186 VDD.n1185 4.65
R1397 VDD.n1180 VDD.n1179 4.65
R1398 VDD.n1176 VDD.n1175 4.65
R1399 VDD.n1171 VDD.n1170 4.65
R1400 VDD.n1167 VDD.n1166 4.65
R1401 VDD.n1141 VDD.n1140 4.65
R1402 VDD.n1137 VDD.n1136 4.65
R1403 VDD.n1132 VDD.n1131 4.65
R1404 VDD.n1128 VDD.n1127 4.65
R1405 VDD.n1123 VDD.n1122 4.65
R1406 VDD.n1119 VDD.n1118 4.65
R1407 VDD.n1115 VDD.n1114 4.65
R1408 VDD.n1110 VDD.n1109 4.65
R1409 VDD.n1084 VDD.n1083 4.65
R1410 VDD.n1080 VDD.n1079 4.65
R1411 VDD.n1076 VDD.n1075 4.65
R1412 VDD.n1072 VDD.n1071 4.65
R1413 VDD.n1068 VDD.n1067 4.65
R1414 VDD.n1062 VDD.n1061 4.65
R1415 VDD.n1058 VDD.n1057 4.65
R1416 VDD.n1054 VDD.n1053 4.65
R1417 VDD.n1048 VDD.n1047 4.65
R1418 VDD.n1044 VDD.n1043 4.65
R1419 VDD.n1039 VDD.n1038 4.65
R1420 VDD.n1035 VDD.n1034 4.65
R1421 VDD.n1009 VDD.n1008 4.65
R1422 VDD.n1005 VDD.n1004 4.65
R1423 VDD.n1001 VDD.n1000 4.65
R1424 VDD.n997 VDD.n996 4.65
R1425 VDD.n993 VDD.n992 4.65
R1426 VDD.n987 VDD.n986 4.65
R1427 VDD.n983 VDD.n982 4.65
R1428 VDD.n979 VDD.n978 4.65
R1429 VDD.n973 VDD.n972 4.65
R1430 VDD.n969 VDD.n968 4.65
R1431 VDD.n964 VDD.n963 4.65
R1432 VDD.n960 VDD.n959 4.65
R1433 VDD.n934 VDD.n933 4.65
R1434 VDD.n930 VDD.n929 4.65
R1435 VDD.n925 VDD.n924 4.65
R1436 VDD.n921 VDD.n920 4.65
R1437 VDD.n916 VDD.n915 4.65
R1438 VDD.n912 VDD.n911 4.65
R1439 VDD.n908 VDD.n907 4.65
R1440 VDD.n903 VDD.n902 4.65
R1441 VDD.n877 VDD.n876 4.65
R1442 VDD.n873 VDD.n872 4.65
R1443 VDD.n869 VDD.n868 4.65
R1444 VDD.n865 VDD.n864 4.65
R1445 VDD.n861 VDD.n860 4.65
R1446 VDD.n855 VDD.n854 4.65
R1447 VDD.n851 VDD.n850 4.65
R1448 VDD.n847 VDD.n846 4.65
R1449 VDD.n841 VDD.n840 4.65
R1450 VDD.n837 VDD.n836 4.65
R1451 VDD.n832 VDD.n831 4.65
R1452 VDD.n828 VDD.n827 4.65
R1453 VDD.n801 VDD.n800 4.65
R1454 VDD.n797 VDD.n796 4.65
R1455 VDD.n793 VDD.n792 4.65
R1456 VDD.n789 VDD.n788 4.65
R1457 VDD.n785 VDD.n784 4.65
R1458 VDD.n779 VDD.n778 4.65
R1459 VDD.n775 VDD.n774 4.65
R1460 VDD.n771 VDD.n770 4.65
R1461 VDD.n765 VDD.n764 4.65
R1462 VDD.n761 VDD.n760 4.65
R1463 VDD.n756 VDD.n755 4.65
R1464 VDD.n752 VDD.n751 4.65
R1465 VDD.n27 VDD.n23 2.933
R1466 VDD.n156 VDD.n153 2.89
R1467 VDD.n213 VDD.n210 2.89
R1468 VDD.n420 VDD.n417 2.89
R1469 VDD.n627 VDD.n624 2.89
R1470 VDD.n1321 VDD.n1318 2.89
R1471 VDD.n1114 VDD.n1111 2.89
R1472 VDD.n907 VDD.n904 2.89
R1473 VDD.n27 VDD.n26 2.844
R1474 VDD.n35 0ܪ{� 2.557
R1475 VDD.n86  2.557
R1476 VDD.n145  2.557
R1477 VDD.n202  2.557
R1478 VDD.n409 0ܪ{� 2.557
R1479 VDD.n616 0ܪ{� 2.557
R1480 VDD.n1327  2.557
R1481 VDD.n1120 0ܪ{� 2.557
R1482 VDD.n913 0ܪ{� 2.557
R1483 VDD.n134 VDD.n131 2.477
R1484 VDD.n191 VDD.n188 2.477
R1485 VDD.n398 VDD.n395 2.477
R1486 VDD.n605 VDD.n602 2.477
R1487 VDD.n1343 VDD.n1340 2.477
R1488 VDD.n1136 VDD.n1133 2.477
R1489 VDD.n929 VDD.n926 2.477
R1490 VDD.n31 VDD.n27 1.063
R1491 VDD.n284 VDD.n281 0.412
R1492 VDD.n359 VDD.n356 0.412
R1493 VDD.n491 VDD.n488 0.412
R1494 VDD.n566 VDD.n563 0.412
R1495 VDD.n698 VDD.n695 0.412
R1496 VDD.n1382 VDD.n1379 0.412
R1497 VDD.n1250 VDD.n1247 0.412
R1498 VDD.n1175 VDD.n1172 0.412
R1499 VDD.n1043 VDD.n1040 0.412
R1500 VDD.n968 VDD.n965 0.412
R1501 VDD.n836 VDD.n833 0.412
R1502 VDD.n760 VDD.n757 0.412
R1503 VDD.n77 VDD.n50 0.29
R1504 VDD.n130 VDD.n104 0.29
R1505 VDD.n187 VDD.n161 0.29
R1506 VDD.n244 VDD.n218 0.29
R1507 VDD.n319 VDD.n293 0.29
R1508 VDD.n394 VDD.n368 0.29
R1509 VDD.n451 VDD.n425 0.29
R1510 VDD.n526 VDD.n500 0.29
R1511 VDD.n601 VDD.n575 0.29
R1512 VDD.n658 VDD.n632 0.29
R1513 VDD.n1374 VDD.n1348 0.29
R1514 VDD.n1317 VDD.n1291 0.29
R1515 VDD.n1242 VDD.n1216 0.29
R1516 VDD.n1167 VDD.n1141 0.29
R1517 VDD.n1110 VDD.n1084 0.29
R1518 VDD.n1035 VDD.n1009 0.29
R1519 VDD.n960 VDD.n934 0.29
R1520 VDD.n903 VDD.n877 0.29
R1521 VDD.n828 VDD.n801 0.29
R1522 VDD VDD.n1423 0.219
R1523 VDD.n752 VDD 0.207
R1524 VDD.n270 VDD.n266 0.197
R1525 VDD.n345 VDD.n341 0.197
R1526 VDD.n477 VDD.n473 0.197
R1527 VDD.n552 VDD.n548 0.197
R1528 VDD.n684 VDD.n680 0.197
R1529 VDD.n1401 VDD.n1397 0.197
R1530 VDD.n1269 VDD.n1265 0.197
R1531 VDD.n1194 VDD.n1190 0.197
R1532 VDD.n1062 VDD.n1058 0.197
R1533 VDD.n987 VDD.n983 0.197
R1534 VDD.n855 VDD.n851 0.197
R1535 VDD.n779 VDD.n775 0.197
R1536 VDD.n38 VDD.n34 0.181
R1537 VDD.n92 VDD.n89 0.181
R1538 VDD.n148 VDD.n144 0.181
R1539 VDD.n205 VDD.n201 0.181
R1540 VDD.n412 VDD.n408 0.181
R1541 VDD.n619 VDD.n615 0.181
R1542 VDD.n1335 VDD.n1330 0.181
R1543 VDD.n1128 VDD.n1123 0.181
R1544 VDD.n921 VDD.n916 0.181
R1545 VDD.n34 VDD.n31 0.145
R1546 VDD.n42 VDD.n38 0.145
R1547 VDD.n46 VDD.n42 0.145
R1548 VDD.n50 VDD.n46 0.145
R1549 VDD.n81 VDD.n77 0.145
R1550 VDD.n85 VDD.n81 0.145
R1551 VDD.n89 VDD.n85 0.145
R1552 VDD.n96 VDD.n92 0.145
R1553 VDD.n100 VDD.n96 0.145
R1554 VDD.n104 VDD.n100 0.145
R1555 VDD.n135 VDD.n130 0.145
R1556 VDD.n139 VDD.n135 0.145
R1557 VDD.n144 VDD.n139 0.145
R1558 VDD.n152 VDD.n148 0.145
R1559 VDD.n157 VDD.n152 0.145
R1560 VDD.n161 VDD.n157 0.145
R1561 VDD.n192 VDD.n187 0.145
R1562 VDD.n196 VDD.n192 0.145
R1563 VDD.n201 VDD.n196 0.145
R1564 VDD.n209 VDD.n205 0.145
R1565 VDD.n214 VDD.n209 0.145
R1566 VDD.n218 VDD.n214 0.145
R1567 VDD.n248 VDD.n244 0.145
R1568 VDD.n252 VDD.n248 0.145
R1569 VDD.n256 VDD.n252 0.145
R1570 VDD.n262 VDD.n256 0.145
R1571 VDD.n266 VDD.n262 0.145
R1572 VDD.n276 VDD.n270 0.145
R1573 VDD.n280 VDD.n276 0.145
R1574 VDD.n285 VDD.n280 0.145
R1575 VDD.n289 VDD.n285 0.145
R1576 VDD.n293 VDD.n289 0.145
R1577 VDD.n323 VDD.n319 0.145
R1578 VDD.n327 VDD.n323 0.145
R1579 VDD.n331 VDD.n327 0.145
R1580 VDD.n337 VDD.n331 0.145
R1581 VDD.n341 VDD.n337 0.145
R1582 VDD.n351 VDD.n345 0.145
R1583 VDD.n355 VDD.n351 0.145
R1584 VDD.n360 VDD.n355 0.145
R1585 VDD.n364 VDD.n360 0.145
R1586 VDD.n368 VDD.n364 0.145
R1587 VDD.n399 VDD.n394 0.145
R1588 VDD.n403 VDD.n399 0.145
R1589 VDD.n408 VDD.n403 0.145
R1590 VDD.n416 VDD.n412 0.145
R1591 VDD.n421 VDD.n416 0.145
R1592 VDD.n425 VDD.n421 0.145
R1593 VDD.n455 VDD.n451 0.145
R1594 VDD.n459 VDD.n455 0.145
R1595 VDD.n463 VDD.n459 0.145
R1596 VDD.n469 VDD.n463 0.145
R1597 VDD.n473 VDD.n469 0.145
R1598 VDD.n483 VDD.n477 0.145
R1599 VDD.n487 VDD.n483 0.145
R1600 VDD.n492 VDD.n487 0.145
R1601 VDD.n496 VDD.n492 0.145
R1602 VDD.n500 VDD.n496 0.145
R1603 VDD.n530 VDD.n526 0.145
R1604 VDD.n534 VDD.n530 0.145
R1605 VDD.n538 VDD.n534 0.145
R1606 VDD.n544 VDD.n538 0.145
R1607 VDD.n548 VDD.n544 0.145
R1608 VDD.n558 VDD.n552 0.145
R1609 VDD.n562 VDD.n558 0.145
R1610 VDD.n567 VDD.n562 0.145
R1611 VDD.n571 VDD.n567 0.145
R1612 VDD.n575 VDD.n571 0.145
R1613 VDD.n606 VDD.n601 0.145
R1614 VDD.n610 VDD.n606 0.145
R1615 VDD.n615 VDD.n610 0.145
R1616 VDD.n623 VDD.n619 0.145
R1617 VDD.n628 VDD.n623 0.145
R1618 VDD.n632 VDD.n628 0.145
R1619 VDD.n662 VDD.n658 0.145
R1620 VDD.n666 VDD.n662 0.145
R1621 VDD.n670 VDD.n666 0.145
R1622 VDD.n676 VDD.n670 0.145
R1623 VDD.n680 VDD.n676 0.145
R1624 VDD.n690 VDD.n684 0.145
R1625 VDD.n694 VDD.n690 0.145
R1626 VDD.n699 VDD.n694 0.145
R1627 VDD.n703 VDD.n699 0.145
R1628 VDD.n729 VDD.n703 0.145
R1629 VDD.n1423 VDD.n1419 0.145
R1630 VDD.n1419 VDD.n1415 0.145
R1631 VDD.n1415 VDD.n1411 0.145
R1632 VDD.n1411 VDD.n1407 0.145
R1633 VDD.n1407 VDD.n1401 0.145
R1634 VDD.n1397 VDD.n1393 0.145
R1635 VDD.n1393 VDD.n1387 0.145
R1636 VDD.n1387 VDD.n1383 0.145
R1637 VDD.n1383 VDD.n1378 0.145
R1638 VDD.n1378 VDD.n1374 0.145
R1639 VDD.n1348 VDD.n1344 0.145
R1640 VDD.n1344 VDD.n1339 0.145
R1641 VDD.n1339 VDD.n1335 0.145
R1642 VDD.n1330 VDD.n1326 0.145
R1643 VDD.n1326 VDD.n1322 0.145
R1644 VDD.n1322 VDD.n1317 0.145
R1645 VDD.n1291 VDD.n1287 0.145
R1646 VDD.n1287 VDD.n1283 0.145
R1647 VDD.n1283 VDD.n1279 0.145
R1648 VDD.n1279 VDD.n1275 0.145
R1649 VDD.n1275 VDD.n1269 0.145
R1650 VDD.n1265 VDD.n1261 0.145
R1651 VDD.n1261 VDD.n1255 0.145
R1652 VDD.n1255 VDD.n1251 0.145
R1653 VDD.n1251 VDD.n1246 0.145
R1654 VDD.n1246 VDD.n1242 0.145
R1655 VDD.n1216 VDD.n1212 0.145
R1656 VDD.n1212 VDD.n1208 0.145
R1657 VDD.n1208 VDD.n1204 0.145
R1658 VDD.n1204 VDD.n1200 0.145
R1659 VDD.n1200 VDD.n1194 0.145
R1660 VDD.n1190 VDD.n1186 0.145
R1661 VDD.n1186 VDD.n1180 0.145
R1662 VDD.n1180 VDD.n1176 0.145
R1663 VDD.n1176 VDD.n1171 0.145
R1664 VDD.n1171 VDD.n1167 0.145
R1665 VDD.n1141 VDD.n1137 0.145
R1666 VDD.n1137 VDD.n1132 0.145
R1667 VDD.n1132 VDD.n1128 0.145
R1668 VDD.n1123 VDD.n1119 0.145
R1669 VDD.n1119 VDD.n1115 0.145
R1670 VDD.n1115 VDD.n1110 0.145
R1671 VDD.n1084 VDD.n1080 0.145
R1672 VDD.n1080 VDD.n1076 0.145
R1673 VDD.n1076 VDD.n1072 0.145
R1674 VDD.n1072 VDD.n1068 0.145
R1675 VDD.n1068 VDD.n1062 0.145
R1676 VDD.n1058 VDD.n1054 0.145
R1677 VDD.n1054 VDD.n1048 0.145
R1678 VDD.n1048 VDD.n1044 0.145
R1679 VDD.n1044 VDD.n1039 0.145
R1680 VDD.n1039 VDD.n1035 0.145
R1681 VDD.n1009 VDD.n1005 0.145
R1682 VDD.n1005 VDD.n1001 0.145
R1683 VDD.n1001 VDD.n997 0.145
R1684 VDD.n997 VDD.n993 0.145
R1685 VDD.n993 VDD.n987 0.145
R1686 VDD.n983 VDD.n979 0.145
R1687 VDD.n979 VDD.n973 0.145
R1688 VDD.n973 VDD.n969 0.145
R1689 VDD.n969 VDD.n964 0.145
R1690 VDD.n964 VDD.n960 0.145
R1691 VDD.n934 VDD.n930 0.145
R1692 VDD.n930 VDD.n925 0.145
R1693 VDD.n925 VDD.n921 0.145
R1694 VDD.n916 VDD.n912 0.145
R1695 VDD.n912 VDD.n908 0.145
R1696 VDD.n908 VDD.n903 0.145
R1697 VDD.n877 VDD.n873 0.145
R1698 VDD.n873 VDD.n869 0.145
R1699 VDD.n869 VDD.n865 0.145
R1700 VDD.n865 VDD.n861 0.145
R1701 VDD.n861 VDD.n855 0.145
R1702 VDD.n851 VDD.n847 0.145
R1703 VDD.n847 VDD.n841 0.145
R1704 VDD.n841 VDD.n837 0.145
R1705 VDD.n837 VDD.n832 0.145
R1706 VDD.n832 VDD.n828 0.145
R1707 VDD.n801 VDD.n797 0.145
R1708 VDD.n797 VDD.n793 0.145
R1709 VDD.n793 VDD.n789 0.145
R1710 VDD.n789 VDD.n785 0.145
R1711 VDD.n785 VDD.n779 0.145
R1712 VDD.n775 VDD.n771 0.145
R1713 VDD.n771 VDD.n765 0.145
R1714 VDD.n765 VDD.n761 0.145
R1715 VDD.n761 VDD.n756 0.145
R1716 VDD.n756 VDD.n752 0.145
R1717 VDD VDD.n729 0.07
R1718 a_10637_1050.n4 a_10637_1050.t11 512.525
R1719 a_10637_1050.n2 a_10637_1050.t10 512.525
R1720 a_10637_1050.n5 a_10637_1050.t9 389.251
R1721 a_10637_1050.n3 a_10637_1050.t12 389.251
R1722 a_10637_1050.n4 a_10637_1050.t8 371.139
R1723 a_10637_1050.n2 a_10637_1050.t7 371.139
R1724 a_10637_1050.n8 a_10637_1050.n7 357.814
R1725 a_10637_1050.n5 a_10637_1050.n4 207.695
R1726 a_10637_1050.n3 a_10637_1050.n2 207.695
R1727 a_10637_1050.n11 a_10637_1050.n10 161.352
R1728 a_10637_1050.n9 a_10637_1050.n8 151.34
R1729 a_10637_1050.n9 a_10637_1050.n1 95.095
R1730 a_10637_1050.n10 a_10637_1050.n0 95.095
R1731 a_10637_1050.n10 a_10637_1050.n9 66.258
R1732 a_10637_1050.n1 a_10637_1050.t1 14.282
R1733 a_10637_1050.n1 a_10637_1050.t2 14.282
R1734 a_10637_1050.n0 a_10637_1050.t6 14.282
R1735 a_10637_1050.n0 a_10637_1050.t0 14.282
R1736 a_10637_1050.n11 a_10637_1050.t4 14.282
R1737 a_10637_1050.t5 a_10637_1050.n11 14.282
R1738 a_10637_1050.n6 a_10637_1050.n3 14.126
R1739 a_10637_1050.n8 a_10637_1050.n6 5.965
R1740 a_10637_1050.n6 a_10637_1050.n5 4.65
R1741 a_14189_1050.n2 a_14189_1050.t7 480.392
R1742 a_14189_1050.n2 a_14189_1050.t9 403.272
R1743 a_14189_1050.n3 a_14189_1050.t8 385.063
R1744 a_14189_1050.n5 a_14189_1050.n4 357.814
R1745 a_14189_1050.n8 a_14189_1050.n7 161.352
R1746 a_14189_1050.n6 a_14189_1050.n5 151.34
R1747 a_14189_1050.n3 a_14189_1050.n2 143.429
R1748 a_14189_1050.n6 a_14189_1050.n1 95.095
R1749 a_14189_1050.n7 a_14189_1050.n0 95.095
R1750 a_14189_1050.n7 a_14189_1050.n6 66.258
R1751 a_14189_1050.n1 a_14189_1050.t0 14.282
R1752 a_14189_1050.n1 a_14189_1050.t1 14.282
R1753 a_14189_1050.n0 a_14189_1050.t4 14.282
R1754 a_14189_1050.n0 a_14189_1050.t5 14.282
R1755 a_14189_1050.n8 a_14189_1050.t2 14.282
R1756 a_14189_1050.t3 a_14189_1050.n8 14.282
R1757 a_14189_1050.n5 a_14189_1050.n3 10.615
R1758 a_10959_989.n2 a_10959_989.t8 480.392
R1759 a_10959_989.n4 a_10959_989.t10 454.685
R1760 a_10959_989.n4 a_10959_989.t9 428.979
R1761 a_10959_989.n2 a_10959_989.t12 403.272
R1762 a_10959_989.n3 a_10959_989.t7 357.204
R1763 a_10959_989.n5 a_10959_989.t11 311.683
R1764 a_10959_989.n11 a_10959_989.n10 308.216
R1765 a_10959_989.n12 a_10959_989.n11 179.199
R1766 a_10959_989.n5 a_10959_989.n4 171.288
R1767 a_10959_989.n3 a_10959_989.n2 171.288
R1768 a_10959_989.n14 a_10959_989.n13 161.352
R1769 a_10959_989.n12 a_10959_989.n1 95.095
R1770 a_10959_989.n13 a_10959_989.n0 95.095
R1771 a_10959_989.n13 a_10959_989.n12 66.258
R1772 a_10959_989.n10 a_10959_989.n9 30
R1773 a_10959_989.n8 a_10959_989.n7 24.383
R1774 a_10959_989.n10 a_10959_989.n8 23.684
R1775 a_10959_989.n1 a_10959_989.t3 14.282
R1776 a_10959_989.n1 a_10959_989.t4 14.282
R1777 a_10959_989.n0 a_10959_989.t6 14.282
R1778 a_10959_989.n0 a_10959_989.t5 14.282
R1779 a_10959_989.n14 a_10959_989.t0 14.282
R1780 a_10959_989.t1 a_10959_989.n14 14.282
R1781 a_10959_989.n6 a_10959_989.n5 8.685
R1782 a_10959_989.n6 a_10959_989.n3 5.965
R1783 a_10959_989.n11 a_10959_989.n6 4.65
R1784 D.n5 D.t6 479.223
R1785 D.n2 D.t4 479.223
R1786 D.n0 D.t8 479.223
R1787 D.n5 D.t0 375.52
R1788 D.n2 D.t7 375.52
R1789 D.n0 D.t2 375.52
R1790 D.n6 D.n5 280.047
R1791 D.n3 D.n2 280.047
R1792 D.n1 D.n0 280.047
R1793 D.n6 D.t1 136.76
R1794 D.n3 D.t5 136.76
R1795 D.n1 D.t3 136.76
R1796 D.n4 D.n1 23.649
R1797 D.n7 D.n4 18.999
R1798 D.n4 D.n3 4.65
R1799 D.n7 D.n6 4.65
R1800 D.n7 D 0.046
R1801 a_599_989.n1 a_599_989.t7 480.392
R1802 a_599_989.n3 a_599_989.t11 454.685
R1803 a_599_989.n3 a_599_989.t8 428.979
R1804 a_599_989.n1 a_599_989.t10 403.272
R1805 a_599_989.n2 a_599_989.t12 357.204
R1806 a_599_989.n4 a_599_989.t9 311.683
R1807 a_599_989.n10 a_599_989.n9 308.216
R1808 a_599_989.n11 a_599_989.n10 179.199
R1809 a_599_989.n4 a_599_989.n3 171.288
R1810 a_599_989.n2 a_599_989.n1 171.288
R1811 a_599_989.n13 a_599_989.n12 161.352
R1812 a_599_989.n11 a_599_989.n0 95.095
R1813 a_599_989.n14 a_599_989.n13 95.094
R1814 a_599_989.n13 a_599_989.n11 66.258
R1815 a_599_989.n9 a_599_989.n8 30
R1816 a_599_989.n7 a_599_989.n6 24.383
R1817 a_599_989.n9 a_599_989.n7 23.684
R1818 a_599_989.n0 a_599_989.t5 14.282
R1819 a_599_989.n0 a_599_989.t6 14.282
R1820 a_599_989.n12 a_599_989.t1 14.282
R1821 a_599_989.n12 a_599_989.t0 14.282
R1822 a_599_989.n14 a_599_989.t2 14.282
R1823 a_599_989.t3 a_599_989.n14 14.282
R1824 a_599_989.n5 a_599_989.n4 8.685
R1825 a_599_989.n5 a_599_989.n2 5.965
R1826 a_599_989.n10 a_599_989.n5 4.65
R1827 a_11413_103.t0 a_11413_103.n0 117.777
R1828 a_11413_103.n2 a_11413_103.n1 66.629
R1829 a_11413_103.t0 a_11413_103.n8 59.616
R1830 a_11413_103.n5 a_11413_103.n3 54.496
R1831 a_11413_103.n5 a_11413_103.n4 54.496
R1832 a_11413_103.t0 a_11413_103.n2 20.262
R1833 a_11413_103.n7 a_11413_103.n5 7.859
R1834 a_11413_103.t0 a_11413_103.n7 3.034
R1835 a_11413_103.n7 a_11413_103.n6 0.443
R1836 GND.n30 GND.n29 237.558
R1837 GND.n449 GND.n448 237.558
R1838 GND.n494 GND.n493 237.558
R1839 GND.n527 GND.n526 237.558
R1840 GND.n571 GND.n570 237.558
R1841 GND.n613 GND.n612 237.558
R1842 GND.n646 GND.n645 237.558
R1843 GND.n690 GND.n689 237.558
R1844 GND.n732 GND.n731 237.558
R1845 GND.n764 GND.n763 237.558
R1846 GND.n364 GND.n363 237.558
R1847 GND.n402 GND.n401 237.558
R1848 GND.n334 GND.n333 237.558
R1849 GND.n289 GND.n288 237.558
R1850 GND.n245 GND.n244 237.558
R1851 GND.n212 GND.n211 237.558
R1852 GND.n170 GND.n169 237.558
R1853 GND.n125 GND.n124 237.558
R1854 GND.n92 GND.n91 237.558
R1855 GND.n60 GND.n59 237.558
R1856 GND.n27 GND.n26 210.82
R1857 GND.n57 GND.n56 210.82
R1858 GND.n451 GND.n450 210.82
R1859 GND.n496 GND.n495 210.82
R1860 GND.n529 GND.n528 210.82
R1861 GND.n573 GND.n572 210.82
R1862 GND.n615 GND.n614 210.82
R1863 GND.n648 GND.n647 210.82
R1864 GND.n692 GND.n691 210.82
R1865 GND.n734 GND.n733 210.82
R1866 GND.n766 GND.n765 210.82
R1867 GND.n404 GND.n403 210.82
R1868 GND.n361 GND.n360 210.82
R1869 GND.n331 GND.n330 210.82
R1870 GND.n286 GND.n285 210.82
R1871 GND.n242 GND.n241 210.82
R1872 GND.n209 GND.n208 210.82
R1873 GND.n167 GND.n166 210.82
R1874 GND.n122 GND.n121 210.82
R1875 GND.n89 GND.n88 210.82
R1876 GND.n199 GND.n198 173.365
R1877 GND.n701 GND.n700 173.365
R1878 GND.n582 GND.n581 173.365
R1879 GND.n46 GND.n45 172.612
R1880 GND.n350 GND.n349 172.612
R1881 GND.n276 GND.n275 167.358
R1882 GND.n395 GND.n394 167.358
R1883 GND.n777 GND.n776 167.358
R1884 GND.n659 GND.n658 167.358
R1885 GND.n540 GND.n539 167.358
R1886 GND.n418 GND.n417 167.358
R1887 GND.n78 GND.n77 166.605
R1888 GND.n744 GND.n743 166.605
R1889 GND.n16 GND.n15 166.605
R1890 GND.n157 GND.n156 152.358
R1891 GND.n321 GND.n320 152.358
R1892 GND.n463 GND.n462 152.358
R1893 GND.n111 GND.n110 151.605
R1894 GND.n231 GND.n230 151.605
R1895 GND.n626 GND.n625 151.605
R1896 GND.n507 GND.n506 151.605
R1897 GND.n110 GND.n109 28.421
R1898 GND.n156 GND.n155 28.421
R1899 GND.n230 GND.n229 28.421
R1900 GND.n320 GND.n319 28.421
R1901 GND.n625 GND.n624 28.421
R1902 GND.n506 GND.n505 28.421
R1903 GND.n462 GND.n461 28.421
R1904 GND.n110 GND.n108 25.263
R1905 GND.n156 GND.n154 25.263
R1906 GND.n230 GND.n228 25.263
R1907 GND.n320 GND.n318 25.263
R1908 GND.n625 GND.n623 25.263
R1909 GND.n506 GND.n504 25.263
R1910 GND.n462 GND.n460 25.263
R1911 GND.n108 GND.n107 24.383
R1912 GND.n154 GND.n153 24.383
R1913 GND.n228 GND.n227 24.383
R1914 GND.n318 GND.n317 24.383
R1915 GND.n623 GND.n622 24.383
R1916 GND.n504 GND.n503 24.383
R1917 GND.n460 GND.n459 24.383
R1918 GND.n77 GND.n75 23.03
R1919 GND.n275 GND.n273 23.03
R1920 GND.n394 GND.n392 23.03
R1921 GND.n776 GND.n774 23.03
R1922 GND.n743 GND.n741 23.03
R1923 GND.n658 GND.n656 23.03
R1924 GND.n539 GND.n537 23.03
R1925 GND.n417 GND.n415 23.03
R1926 GND.n15 GND.n13 23.03
R1927 GND.n28 GND.n27 18.953
R1928 GND.n58 GND.n57 18.953
R1929 GND.n452 GND.n451 18.953
R1930 GND.n497 GND.n496 18.953
R1931 GND.n530 GND.n529 18.953
R1932 GND.n574 GND.n573 18.953
R1933 GND.n616 GND.n615 18.953
R1934 GND.n649 GND.n648 18.953
R1935 GND.n693 GND.n692 18.953
R1936 GND.n735 GND.n734 18.953
R1937 GND.n767 GND.n766 18.953
R1938 GND.n405 GND.n404 18.953
R1939 GND.n362 GND.n361 18.953
R1940 GND.n332 GND.n331 18.953
R1941 GND.n287 GND.n286 18.953
R1942 GND.n243 GND.n242 18.953
R1943 GND.n210 GND.n209 18.953
R1944 GND.n168 GND.n167 18.953
R1945 GND.n123 GND.n122 18.953
R1946 GND.n90 GND.n89 18.953
R1947 GND.n31 GND.n28 14.864
R1948 GND.n61 GND.n58 14.864
R1949 GND.n93 GND.n90 14.864
R1950 GND.n126 GND.n123 14.864
R1951 GND.n171 GND.n168 14.864
R1952 GND.n213 GND.n210 14.864
R1953 GND.n246 GND.n243 14.864
R1954 GND.n290 GND.n287 14.864
R1955 GND.n335 GND.n332 14.864
R1956 GND.n365 GND.n362 14.864
R1957 GND.n406 GND.n405 14.864
R1958 GND.n768 GND.n767 14.864
R1959 GND.n736 GND.n735 14.864
R1960 GND.n694 GND.n693 14.864
R1961 GND.n650 GND.n649 14.864
R1962 GND.n617 GND.n616 14.864
R1963 GND.n575 GND.n574 14.864
R1964 GND.n531 GND.n530 14.864
R1965 GND.n498 GND.n497 14.864
R1966 GND.n453 GND.n452 14.864
R1967 GND.n412 GND.n411 9.154
R1968 GND.n419 GND.n414 9.154
R1969 GND.n422 GND.n421 9.154
R1970 GND.n425 GND.n424 9.154
R1971 GND.n428 GND.n427 9.154
R1972 GND.n431 GND.n430 9.154
R1973 GND.n434 GND.n433 9.154
R1974 GND.n437 GND.n436 9.154
R1975 GND.n440 GND.n439 9.154
R1976 GND.n443 GND.n442 9.154
R1977 GND.n446 GND.n445 9.154
R1978 GND.n453 GND.n449 9.154
R1979 GND.n456 GND.n455 9.154
R1980 GND.n464 GND.n458 9.154
R1981 GND.n467 GND.n466 9.154
R1982 GND.n470 GND.n469 9.154
R1983 GND.n473 GND.n472 9.154
R1984 GND.n476 GND.n475 9.154
R1985 GND.n479 GND.n478 9.154
R1986 GND.n482 GND.n481 9.154
R1987 GND.n485 GND.n484 9.154
R1988 GND.n488 GND.n487 9.154
R1989 GND.n491 GND.n490 9.154
R1990 GND.n498 GND.n494 9.154
R1991 GND.n501 GND.n500 9.154
R1992 GND.n509 GND.n508 9.154
R1993 GND.n512 GND.n511 9.154
R1994 GND.n515 GND.n514 9.154
R1995 GND.n518 GND.n517 9.154
R1996 GND.n521 GND.n520 9.154
R1997 GND.n524 GND.n523 9.154
R1998 GND.n531 GND.n527 9.154
R1999 GND.n534 GND.n533 9.154
R2000 GND.n541 GND.n536 9.154
R2001 GND.n544 GND.n543 9.154
R2002 GND.n547 GND.n546 9.154
R2003 GND.n550 GND.n549 9.154
R2004 GND.n553 GND.n552 9.154
R2005 GND.n556 GND.n555 9.154
R2006 GND.n559 GND.n558 9.154
R2007 GND.n562 GND.n561 9.154
R2008 GND.n565 GND.n564 9.154
R2009 GND.n568 GND.n567 9.154
R2010 GND.n575 GND.n571 9.154
R2011 GND.n578 GND.n577 9.154
R2012 GND.n583 GND.n580 9.154
R2013 GND.n586 GND.n585 9.154
R2014 GND.n589 GND.n588 9.154
R2015 GND.n592 GND.n591 9.154
R2016 GND.n595 GND.n594 9.154
R2017 GND.n598 GND.n597 9.154
R2018 GND.n601 GND.n600 9.154
R2019 GND.n604 GND.n603 9.154
R2020 GND.n607 GND.n606 9.154
R2021 GND.n610 GND.n609 9.154
R2022 GND.n617 GND.n613 9.154
R2023 GND.n620 GND.n619 9.154
R2024 GND.n628 GND.n627 9.154
R2025 GND.n631 GND.n630 9.154
R2026 GND.n634 GND.n633 9.154
R2027 GND.n637 GND.n636 9.154
R2028 GND.n640 GND.n639 9.154
R2029 GND.n643 GND.n642 9.154
R2030 GND.n650 GND.n646 9.154
R2031 GND.n653 GND.n652 9.154
R2032 GND.n660 GND.n655 9.154
R2033 GND.n663 GND.n662 9.154
R2034 GND.n666 GND.n665 9.154
R2035 GND.n669 GND.n668 9.154
R2036 GND.n672 GND.n671 9.154
R2037 GND.n675 GND.n674 9.154
R2038 GND.n678 GND.n677 9.154
R2039 GND.n681 GND.n680 9.154
R2040 GND.n684 GND.n683 9.154
R2041 GND.n687 GND.n686 9.154
R2042 GND.n694 GND.n690 9.154
R2043 GND.n697 GND.n696 9.154
R2044 GND.n702 GND.n699 9.154
R2045 GND.n705 GND.n704 9.154
R2046 GND.n708 GND.n707 9.154
R2047 GND.n711 GND.n710 9.154
R2048 GND.n714 GND.n713 9.154
R2049 GND.n717 GND.n716 9.154
R2050 GND.n720 GND.n719 9.154
R2051 GND.n723 GND.n722 9.154
R2052 GND.n726 GND.n725 9.154
R2053 GND.n729 GND.n728 9.154
R2054 GND.n736 GND.n732 9.154
R2055 GND.n739 GND.n738 9.154
R2056 GND.n746 GND.n745 9.154
R2057 GND.n749 GND.n748 9.154
R2058 GND.n752 GND.n751 9.154
R2059 GND.n755 GND.n754 9.154
R2060 GND.n758 GND.n757 9.154
R2061 GND.n761 GND.n760 9.154
R2062 GND.n768 GND.n764 9.154
R2063 GND.n771 GND.n770 9.154
R2064 GND.n778 GND.n773 9.154
R2065 GND.n781 GND.n780 9.154
R2066 GND.n784 GND.n783 9.154
R2067 GND.n787 GND.n786 9.154
R2068 GND.n790 GND.n789 9.154
R2069 GND.n793 GND.n792 9.154
R2070 GND.n796 GND.n795 9.154
R2071 GND.n799 GND.n798 9.154
R2072 GND.n802 GND.n801 9.154
R2073 GND.n805 GND.n804 9.154
R2074 GND.n406 GND.n402 9.154
R2075 GND.n399 GND.n398 9.154
R2076 GND.n396 GND.n391 9.154
R2077 GND.n389 GND.n388 9.154
R2078 GND.n386 GND.n385 9.154
R2079 GND.n383 GND.n382 9.154
R2080 GND.n380 GND.n379 9.154
R2081 GND.n377 GND.n376 9.154
R2082 GND.n374 GND.n373 9.154
R2083 GND.n371 GND.n370 9.154
R2084 GND.n368 GND.n367 9.154
R2085 GND.n365 GND.n364 9.154
R2086 GND.n358 GND.n357 9.154
R2087 GND.n355 GND.n354 9.154
R2088 GND.n352 GND.n351 9.154
R2089 GND.n347 GND.n346 9.154
R2090 GND.n344 GND.n343 9.154
R2091 GND.n341 GND.n340 9.154
R2092 GND.n338 GND.n337 9.154
R2093 GND.n335 GND.n334 9.154
R2094 GND.n328 GND.n327 9.154
R2095 GND.n325 GND.n324 9.154
R2096 GND.n322 GND.n316 9.154
R2097 GND.n314 GND.n313 9.154
R2098 GND.n311 GND.n310 9.154
R2099 GND.n308 GND.n307 9.154
R2100 GND.n305 GND.n304 9.154
R2101 GND.n302 GND.n301 9.154
R2102 GND.n299 GND.n298 9.154
R2103 GND.n296 GND.n295 9.154
R2104 GND.n293 GND.n292 9.154
R2105 GND.n290 GND.n289 9.154
R2106 GND.n283 GND.n282 9.154
R2107 GND.n280 GND.n279 9.154
R2108 GND.n277 GND.n272 9.154
R2109 GND.n270 GND.n269 9.154
R2110 GND.n267 GND.n266 9.154
R2111 GND.n264 GND.n263 9.154
R2112 GND.n261 GND.n260 9.154
R2113 GND.n258 GND.n257 9.154
R2114 GND.n255 GND.n254 9.154
R2115 GND.n252 GND.n251 9.154
R2116 GND.n249 GND.n248 9.154
R2117 GND.n246 GND.n245 9.154
R2118 GND.n239 GND.n238 9.154
R2119 GND.n236 GND.n235 9.154
R2120 GND.n233 GND.n232 9.154
R2121 GND.n225 GND.n224 9.154
R2122 GND.n222 GND.n221 9.154
R2123 GND.n219 GND.n218 9.154
R2124 GND.n216 GND.n215 9.154
R2125 GND.n213 GND.n212 9.154
R2126 GND.n206 GND.n205 9.154
R2127 GND.n203 GND.n202 9.154
R2128 GND.n200 GND.n197 9.154
R2129 GND.n195 GND.n194 9.154
R2130 GND.n192 GND.n191 9.154
R2131 GND.n189 GND.n188 9.154
R2132 GND.n186 GND.n185 9.154
R2133 GND.n183 GND.n182 9.154
R2134 GND.n180 GND.n179 9.154
R2135 GND.n177 GND.n176 9.154
R2136 GND.n174 GND.n173 9.154
R2137 GND.n171 GND.n170 9.154
R2138 GND.n164 GND.n163 9.154
R2139 GND.n161 GND.n160 9.154
R2140 GND.n158 GND.n152 9.154
R2141 GND.n150 GND.n149 9.154
R2142 GND.n147 GND.n146 9.154
R2143 GND.n144 GND.n143 9.154
R2144 GND.n141 GND.n140 9.154
R2145 GND.n138 GND.n137 9.154
R2146 GND.n135 GND.n134 9.154
R2147 GND.n132 GND.n131 9.154
R2148 GND.n129 GND.n128 9.154
R2149 GND.n126 GND.n125 9.154
R2150 GND.n119 GND.n118 9.154
R2151 GND.n116 GND.n115 9.154
R2152 GND.n113 GND.n112 9.154
R2153 GND.n105 GND.n104 9.154
R2154 GND.n102 GND.n101 9.154
R2155 GND.n99 GND.n98 9.154
R2156 GND.n96 GND.n95 9.154
R2157 GND.n93 GND.n92 9.154
R2158 GND.n86 GND.n85 9.154
R2159 GND.n83 GND.n82 9.154
R2160 GND.n80 GND.n79 9.154
R2161 GND.n73 GND.n72 9.154
R2162 GND.n70 GND.n69 9.154
R2163 GND.n67 GND.n66 9.154
R2164 GND.n64 GND.n63 9.154
R2165 GND.n61 GND.n60 9.154
R2166 GND.n54 GND.n53 9.154
R2167 GND.n51 GND.n50 9.154
R2168 GND.n48 GND.n47 9.154
R2169 GND.n43 GND.n42 9.154
R2170 GND.n40 GND.n39 9.154
R2171 GND.n1 GND.n0 9.154
R2172 GND.n5 GND.n4 9.154
R2173 GND.n8 GND.n7 9.154
R2174 GND.n11 GND.n10 9.154
R2175 GND.n18 GND.n17 9.154
R2176 GND.n21 GND.n20 9.154
R2177 GND.n24 GND.n23 9.154
R2178 GND.n31 GND.n30 9.154
R2179 GND.n34 GND.n33 9.154
R2180 GND.n37 GND.n36 9.154
R2181 GND.n77 GND.n76 8.128
R2182 GND.n275 GND.n274 8.128
R2183 GND.n394 GND.n393 8.128
R2184 GND.n776 GND.n775 8.128
R2185 GND.n743 GND.n742 8.128
R2186 GND.n658 GND.n657 8.128
R2187 GND.n539 GND.n538 8.128
R2188 GND.n417 GND.n416 8.128
R2189 GND.n15 GND.n14 8.128
R2190 GND.n410 GND.n409 4.65
R2191 GND.n41 GND.n40 4.65
R2192 GND.n44 GND.n43 4.65
R2193 GND.n49 GND.n48 4.65
R2194 GND.n52 GND.n51 4.65
R2195 GND.n55 GND.n54 4.65
R2196 GND.n62 GND.n61 4.65
R2197 GND.n65 GND.n64 4.65
R2198 GND.n68 GND.n67 4.65
R2199 GND.n71 GND.n70 4.65
R2200 GND.n74 GND.n73 4.65
R2201 GND.n81 GND.n80 4.65
R2202 GND.n84 GND.n83 4.65
R2203 GND.n87 GND.n86 4.65
R2204 GND.n94 GND.n93 4.65
R2205 GND.n97 GND.n96 4.65
R2206 GND.n100 GND.n99 4.65
R2207 GND.n103 GND.n102 4.65
R2208 GND.n106 GND.n105 4.65
R2209 GND.n114 GND.n113 4.65
R2210 GND.n117 GND.n116 4.65
R2211 GND.n120 GND.n119 4.65
R2212 GND.n127 GND.n126 4.65
R2213 GND.n130 GND.n129 4.65
R2214 GND.n133 GND.n132 4.65
R2215 GND.n136 GND.n135 4.65
R2216 GND.n139 GND.n138 4.65
R2217 GND.n142 GND.n141 4.65
R2218 GND.n145 GND.n144 4.65
R2219 GND.n148 GND.n147 4.65
R2220 GND.n151 GND.n150 4.65
R2221 GND.n159 GND.n158 4.65
R2222 GND.n162 GND.n161 4.65
R2223 GND.n165 GND.n164 4.65
R2224 GND.n172 GND.n171 4.65
R2225 GND.n175 GND.n174 4.65
R2226 GND.n178 GND.n177 4.65
R2227 GND.n181 GND.n180 4.65
R2228 GND.n184 GND.n183 4.65
R2229 GND.n187 GND.n186 4.65
R2230 GND.n190 GND.n189 4.65
R2231 GND.n193 GND.n192 4.65
R2232 GND.n196 GND.n195 4.65
R2233 GND.n201 GND.n200 4.65
R2234 GND.n204 GND.n203 4.65
R2235 GND.n207 GND.n206 4.65
R2236 GND.n214 GND.n213 4.65
R2237 GND.n217 GND.n216 4.65
R2238 GND.n220 GND.n219 4.65
R2239 GND.n223 GND.n222 4.65
R2240 GND.n226 GND.n225 4.65
R2241 GND.n234 GND.n233 4.65
R2242 GND.n237 GND.n236 4.65
R2243 GND.n240 GND.n239 4.65
R2244 GND.n247 GND.n246 4.65
R2245 GND.n250 GND.n249 4.65
R2246 GND.n253 GND.n252 4.65
R2247 GND.n256 GND.n255 4.65
R2248 GND.n259 GND.n258 4.65
R2249 GND.n262 GND.n261 4.65
R2250 GND.n265 GND.n264 4.65
R2251 GND.n268 GND.n267 4.65
R2252 GND.n271 GND.n270 4.65
R2253 GND.n278 GND.n277 4.65
R2254 GND.n281 GND.n280 4.65
R2255 GND.n284 GND.n283 4.65
R2256 GND.n291 GND.n290 4.65
R2257 GND.n294 GND.n293 4.65
R2258 GND.n297 GND.n296 4.65
R2259 GND.n300 GND.n299 4.65
R2260 GND.n303 GND.n302 4.65
R2261 GND.n306 GND.n305 4.65
R2262 GND.n309 GND.n308 4.65
R2263 GND.n312 GND.n311 4.65
R2264 GND.n315 GND.n314 4.65
R2265 GND.n323 GND.n322 4.65
R2266 GND.n326 GND.n325 4.65
R2267 GND.n329 GND.n328 4.65
R2268 GND.n336 GND.n335 4.65
R2269 GND.n339 GND.n338 4.65
R2270 GND.n342 GND.n341 4.65
R2271 GND.n345 GND.n344 4.65
R2272 GND.n348 GND.n347 4.65
R2273 GND.n353 GND.n352 4.65
R2274 GND.n356 GND.n355 4.65
R2275 GND.n359 GND.n358 4.65
R2276 GND.n366 GND.n365 4.65
R2277 GND.n369 GND.n368 4.65
R2278 GND.n372 GND.n371 4.65
R2279 GND.n375 GND.n374 4.65
R2280 GND.n378 GND.n377 4.65
R2281 GND.n381 GND.n380 4.65
R2282 GND.n384 GND.n383 4.65
R2283 GND.n387 GND.n386 4.65
R2284 GND.n390 GND.n389 4.65
R2285 GND.n397 GND.n396 4.65
R2286 GND.n400 GND.n399 4.65
R2287 GND.n407 GND.n406 4.65
R2288 GND.n806 GND.n805 4.65
R2289 GND.n803 GND.n802 4.65
R2290 GND.n800 GND.n799 4.65
R2291 GND.n797 GND.n796 4.65
R2292 GND.n794 GND.n793 4.65
R2293 GND.n791 GND.n790 4.65
R2294 GND.n788 GND.n787 4.65
R2295 GND.n785 GND.n784 4.65
R2296 GND.n782 GND.n781 4.65
R2297 GND.n779 GND.n778 4.65
R2298 GND.n772 GND.n771 4.65
R2299 GND.n769 GND.n768 4.65
R2300 GND.n762 GND.n761 4.65
R2301 GND.n759 GND.n758 4.65
R2302 GND.n756 GND.n755 4.65
R2303 GND.n753 GND.n752 4.65
R2304 GND.n750 GND.n749 4.65
R2305 GND.n747 GND.n746 4.65
R2306 GND.n740 GND.n739 4.65
R2307 GND.n737 GND.n736 4.65
R2308 GND.n730 GND.n729 4.65
R2309 GND.n727 GND.n726 4.65
R2310 GND.n724 GND.n723 4.65
R2311 GND.n721 GND.n720 4.65
R2312 GND.n718 GND.n717 4.65
R2313 GND.n715 GND.n714 4.65
R2314 GND.n712 GND.n711 4.65
R2315 GND.n709 GND.n708 4.65
R2316 GND.n706 GND.n705 4.65
R2317 GND.n703 GND.n702 4.65
R2318 GND.n698 GND.n697 4.65
R2319 GND.n695 GND.n694 4.65
R2320 GND.n688 GND.n687 4.65
R2321 GND.n685 GND.n684 4.65
R2322 GND.n682 GND.n681 4.65
R2323 GND.n679 GND.n678 4.65
R2324 GND.n676 GND.n675 4.65
R2325 GND.n673 GND.n672 4.65
R2326 GND.n670 GND.n669 4.65
R2327 GND.n667 GND.n666 4.65
R2328 GND.n664 GND.n663 4.65
R2329 GND.n661 GND.n660 4.65
R2330 GND.n654 GND.n653 4.65
R2331 GND.n651 GND.n650 4.65
R2332 GND.n644 GND.n643 4.65
R2333 GND.n641 GND.n640 4.65
R2334 GND.n638 GND.n637 4.65
R2335 GND.n635 GND.n634 4.65
R2336 GND.n632 GND.n631 4.65
R2337 GND.n629 GND.n628 4.65
R2338 GND.n621 GND.n620 4.65
R2339 GND.n618 GND.n617 4.65
R2340 GND.n611 GND.n610 4.65
R2341 GND.n608 GND.n607 4.65
R2342 GND.n605 GND.n604 4.65
R2343 GND.n602 GND.n601 4.65
R2344 GND.n599 GND.n598 4.65
R2345 GND.n596 GND.n595 4.65
R2346 GND.n593 GND.n592 4.65
R2347 GND.n590 GND.n589 4.65
R2348 GND.n587 GND.n586 4.65
R2349 GND.n584 GND.n583 4.65
R2350 GND.n579 GND.n578 4.65
R2351 GND.n576 GND.n575 4.65
R2352 GND.n569 GND.n568 4.65
R2353 GND.n566 GND.n565 4.65
R2354 GND.n563 GND.n562 4.65
R2355 GND.n560 GND.n559 4.65
R2356 GND.n557 GND.n556 4.65
R2357 GND.n554 GND.n553 4.65
R2358 GND.n551 GND.n550 4.65
R2359 GND.n548 GND.n547 4.65
R2360 GND.n545 GND.n544 4.65
R2361 GND.n542 GND.n541 4.65
R2362 GND.n535 GND.n534 4.65
R2363 GND.n532 GND.n531 4.65
R2364 GND.n525 GND.n524 4.65
R2365 GND.n522 GND.n521 4.65
R2366 GND.n519 GND.n518 4.65
R2367 GND.n516 GND.n515 4.65
R2368 GND.n513 GND.n512 4.65
R2369 GND.n510 GND.n509 4.65
R2370 GND.n502 GND.n501 4.65
R2371 GND.n499 GND.n498 4.65
R2372 GND.n492 GND.n491 4.65
R2373 GND.n489 GND.n488 4.65
R2374 GND.n486 GND.n485 4.65
R2375 GND.n483 GND.n482 4.65
R2376 GND.n480 GND.n479 4.65
R2377 GND.n477 GND.n476 4.65
R2378 GND.n474 GND.n473 4.65
R2379 GND.n471 GND.n470 4.65
R2380 GND.n468 GND.n467 4.65
R2381 GND.n465 GND.n464 4.65
R2382 GND.n457 GND.n456 4.65
R2383 GND.n454 GND.n453 4.65
R2384 GND.n447 GND.n446 4.65
R2385 GND.n444 GND.n443 4.65
R2386 GND.n441 GND.n440 4.65
R2387 GND.n438 GND.n437 4.65
R2388 GND.n435 GND.n434 4.65
R2389 GND.n432 GND.n431 4.65
R2390 GND.n429 GND.n428 4.65
R2391 GND.n426 GND.n425 4.65
R2392 GND.n423 GND.n422 4.65
R2393 GND.n420 GND.n419 4.65
R2394 GND.n413 GND.n412 4.65
R2395 GND.n6 GND.n5 4.65
R2396 GND.n9 GND.n8 4.65
R2397 GND.n12 GND.n11 4.65
R2398 GND.n19 GND.n18 4.65
R2399 GND.n22 GND.n21 4.65
R2400 GND.n25 GND.n24 4.65
R2401 GND.n32 GND.n31 4.65
R2402 GND.n35 GND.n34 4.65
R2403 GND.n38 GND.n37 4.65
R2404 GND.n18 GND.n16 4.129
R2405 GND.n48 GND.n46 4.129
R2406 GND.n80 GND.n78 4.129
R2407 GND.n113 GND.n111 4.129
R2408 GND.n233 GND.n231 4.129
R2409 GND.n352 GND.n350 4.129
R2410 GND.n746 GND.n744 4.129
R2411 GND.n628 GND.n626 4.129
R2412 GND.n509 GND.n507 4.129
R2413 GND.n3 GND.n2 3.408
R2414 GND.n3 GND.n1 2.844
R2415 GND.n6 GND.n3 1.063
R2416 GND.n409 GND.n408 0.474
R2417 GND.n32 GND.n25 0.29
R2418 GND.n62 GND.n55 0.29
R2419 GND.n94 GND.n87 0.29
R2420 GND.n127 GND.n120 0.29
R2421 GND.n172 GND.n165 0.29
R2422 GND.n214 GND.n207 0.29
R2423 GND.n247 GND.n240 0.29
R2424 GND.n291 GND.n284 0.29
R2425 GND.n336 GND.n329 0.29
R2426 GND.n366 GND.n359 0.29
R2427 GND.n769 GND.n762 0.29
R2428 GND.n737 GND.n730 0.29
R2429 GND.n695 GND.n688 0.29
R2430 GND.n651 GND.n644 0.29
R2431 GND.n618 GND.n611 0.29
R2432 GND.n576 GND.n569 0.29
R2433 GND.n532 GND.n525 0.29
R2434 GND.n499 GND.n492 0.29
R2435 GND.n454 GND.n447 0.29
R2436 GND GND.n806 0.219
R2437 GND.n410 GND 0.207
R2438 GND.n158 GND.n157 0.206
R2439 GND.n200 GND.n199 0.206
R2440 GND.n277 GND.n276 0.206
R2441 GND.n322 GND.n321 0.206
R2442 GND.n396 GND.n395 0.206
R2443 GND.n778 GND.n777 0.206
R2444 GND.n702 GND.n701 0.206
R2445 GND.n660 GND.n659 0.206
R2446 GND.n583 GND.n582 0.206
R2447 GND.n541 GND.n540 0.206
R2448 GND.n464 GND.n463 0.206
R2449 GND.n419 GND.n418 0.206
R2450 GND.n145 GND.n142 0.197
R2451 GND.n190 GND.n187 0.197
R2452 GND.n265 GND.n262 0.197
R2453 GND.n309 GND.n306 0.197
R2454 GND.n384 GND.n381 0.197
R2455 GND.n791 GND.n788 0.197
R2456 GND.n715 GND.n712 0.197
R2457 GND.n673 GND.n670 0.197
R2458 GND.n596 GND.n593 0.197
R2459 GND.n554 GND.n551 0.197
R2460 GND.n477 GND.n474 0.197
R2461 GND.n432 GND.n429 0.197
R2462 GND.n12 GND.n9 0.181
R2463 GND.n44 GND.n41 0.181
R2464 GND.n74 GND.n71 0.181
R2465 GND.n106 GND.n103 0.181
R2466 GND.n226 GND.n223 0.181
R2467 GND.n348 GND.n345 0.181
R2468 GND.n753 GND.n750 0.181
R2469 GND.n635 GND.n632 0.181
R2470 GND.n516 GND.n513 0.181
R2471 GND.n9 GND.n6 0.145
R2472 GND.n19 GND.n12 0.145
R2473 GND.n22 GND.n19 0.145
R2474 GND.n25 GND.n22 0.145
R2475 GND.n35 GND.n32 0.145
R2476 GND.n38 GND.n35 0.145
R2477 GND.n41 GND.n38 0.145
R2478 GND.n49 GND.n44 0.145
R2479 GND.n52 GND.n49 0.145
R2480 GND.n55 GND.n52 0.145
R2481 GND.n65 GND.n62 0.145
R2482 GND.n68 GND.n65 0.145
R2483 GND.n71 GND.n68 0.145
R2484 GND.n81 GND.n74 0.145
R2485 GND.n84 GND.n81 0.145
R2486 GND.n87 GND.n84 0.145
R2487 GND.n97 GND.n94 0.145
R2488 GND.n100 GND.n97 0.145
R2489 GND.n103 GND.n100 0.145
R2490 GND.n114 GND.n106 0.145
R2491 GND.n117 GND.n114 0.145
R2492 GND.n120 GND.n117 0.145
R2493 GND.n130 GND.n127 0.145
R2494 GND.n133 GND.n130 0.145
R2495 GND.n136 GND.n133 0.145
R2496 GND.n139 GND.n136 0.145
R2497 GND.n142 GND.n139 0.145
R2498 GND.n148 GND.n145 0.145
R2499 GND.n151 GND.n148 0.145
R2500 GND.n159 GND.n151 0.145
R2501 GND.n162 GND.n159 0.145
R2502 GND.n165 GND.n162 0.145
R2503 GND.n175 GND.n172 0.145
R2504 GND.n178 GND.n175 0.145
R2505 GND.n181 GND.n178 0.145
R2506 GND.n184 GND.n181 0.145
R2507 GND.n187 GND.n184 0.145
R2508 GND.n193 GND.n190 0.145
R2509 GND.n196 GND.n193 0.145
R2510 GND.n201 GND.n196 0.145
R2511 GND.n204 GND.n201 0.145
R2512 GND.n207 GND.n204 0.145
R2513 GND.n217 GND.n214 0.145
R2514 GND.n220 GND.n217 0.145
R2515 GND.n223 GND.n220 0.145
R2516 GND.n234 GND.n226 0.145
R2517 GND.n237 GND.n234 0.145
R2518 GND.n240 GND.n237 0.145
R2519 GND.n250 GND.n247 0.145
R2520 GND.n253 GND.n250 0.145
R2521 GND.n256 GND.n253 0.145
R2522 GND.n259 GND.n256 0.145
R2523 GND.n262 GND.n259 0.145
R2524 GND.n268 GND.n265 0.145
R2525 GND.n271 GND.n268 0.145
R2526 GND.n278 GND.n271 0.145
R2527 GND.n281 GND.n278 0.145
R2528 GND.n284 GND.n281 0.145
R2529 GND.n294 GND.n291 0.145
R2530 GND.n297 GND.n294 0.145
R2531 GND.n300 GND.n297 0.145
R2532 GND.n303 GND.n300 0.145
R2533 GND.n306 GND.n303 0.145
R2534 GND.n312 GND.n309 0.145
R2535 GND.n315 GND.n312 0.145
R2536 GND.n323 GND.n315 0.145
R2537 GND.n326 GND.n323 0.145
R2538 GND.n329 GND.n326 0.145
R2539 GND.n339 GND.n336 0.145
R2540 GND.n342 GND.n339 0.145
R2541 GND.n345 GND.n342 0.145
R2542 GND.n353 GND.n348 0.145
R2543 GND.n356 GND.n353 0.145
R2544 GND.n359 GND.n356 0.145
R2545 GND.n369 GND.n366 0.145
R2546 GND.n372 GND.n369 0.145
R2547 GND.n375 GND.n372 0.145
R2548 GND.n378 GND.n375 0.145
R2549 GND.n381 GND.n378 0.145
R2550 GND.n387 GND.n384 0.145
R2551 GND.n390 GND.n387 0.145
R2552 GND.n397 GND.n390 0.145
R2553 GND.n400 GND.n397 0.145
R2554 GND.n407 GND.n400 0.145
R2555 GND.n806 GND.n803 0.145
R2556 GND.n803 GND.n800 0.145
R2557 GND.n800 GND.n797 0.145
R2558 GND.n797 GND.n794 0.145
R2559 GND.n794 GND.n791 0.145
R2560 GND.n788 GND.n785 0.145
R2561 GND.n785 GND.n782 0.145
R2562 GND.n782 GND.n779 0.145
R2563 GND.n779 GND.n772 0.145
R2564 GND.n772 GND.n769 0.145
R2565 GND.n762 GND.n759 0.145
R2566 GND.n759 GND.n756 0.145
R2567 GND.n756 GND.n753 0.145
R2568 GND.n750 GND.n747 0.145
R2569 GND.n747 GND.n740 0.145
R2570 GND.n740 GND.n737 0.145
R2571 GND.n730 GND.n727 0.145
R2572 GND.n727 GND.n724 0.145
R2573 GND.n724 GND.n721 0.145
R2574 GND.n721 GND.n718 0.145
R2575 GND.n718 GND.n715 0.145
R2576 GND.n712 GND.n709 0.145
R2577 GND.n709 GND.n706 0.145
R2578 GND.n706 GND.n703 0.145
R2579 GND.n703 GND.n698 0.145
R2580 GND.n698 GND.n695 0.145
R2581 GND.n688 GND.n685 0.145
R2582 GND.n685 GND.n682 0.145
R2583 GND.n682 GND.n679 0.145
R2584 GND.n679 GND.n676 0.145
R2585 GND.n676 GND.n673 0.145
R2586 GND.n670 GND.n667 0.145
R2587 GND.n667 GND.n664 0.145
R2588 GND.n664 GND.n661 0.145
R2589 GND.n661 GND.n654 0.145
R2590 GND.n654 GND.n651 0.145
R2591 GND.n644 GND.n641 0.145
R2592 GND.n641 GND.n638 0.145
R2593 GND.n638 GND.n635 0.145
R2594 GND.n632 GND.n629 0.145
R2595 GND.n629 GND.n621 0.145
R2596 GND.n621 GND.n618 0.145
R2597 GND.n611 GND.n608 0.145
R2598 GND.n608 GND.n605 0.145
R2599 GND.n605 GND.n602 0.145
R2600 GND.n602 GND.n599 0.145
R2601 GND.n599 GND.n596 0.145
R2602 GND.n593 GND.n590 0.145
R2603 GND.n590 GND.n587 0.145
R2604 GND.n587 GND.n584 0.145
R2605 GND.n584 GND.n579 0.145
R2606 GND.n579 GND.n576 0.145
R2607 GND.n569 GND.n566 0.145
R2608 GND.n566 GND.n563 0.145
R2609 GND.n563 GND.n560 0.145
R2610 GND.n560 GND.n557 0.145
R2611 GND.n557 GND.n554 0.145
R2612 GND.n551 GND.n548 0.145
R2613 GND.n548 GND.n545 0.145
R2614 GND.n545 GND.n542 0.145
R2615 GND.n542 GND.n535 0.145
R2616 GND.n535 GND.n532 0.145
R2617 GND.n525 GND.n522 0.145
R2618 GND.n522 GND.n519 0.145
R2619 GND.n519 GND.n516 0.145
R2620 GND.n513 GND.n510 0.145
R2621 GND.n510 GND.n502 0.145
R2622 GND.n502 GND.n499 0.145
R2623 GND.n492 GND.n489 0.145
R2624 GND.n489 GND.n486 0.145
R2625 GND.n486 GND.n483 0.145
R2626 GND.n483 GND.n480 0.145
R2627 GND.n480 GND.n477 0.145
R2628 GND.n474 GND.n471 0.145
R2629 GND.n471 GND.n468 0.145
R2630 GND.n468 GND.n465 0.145
R2631 GND.n465 GND.n457 0.145
R2632 GND.n457 GND.n454 0.145
R2633 GND.n447 GND.n444 0.145
R2634 GND.n444 GND.n441 0.145
R2635 GND.n441 GND.n438 0.145
R2636 GND.n438 GND.n435 0.145
R2637 GND.n435 GND.n432 0.145
R2638 GND.n429 GND.n426 0.145
R2639 GND.n426 GND.n423 0.145
R2640 GND.n423 GND.n420 0.145
R2641 GND.n420 GND.n413 0.145
R2642 GND.n413 GND.n410 0.145
R2643 GND GND.n407 0.07
R2644 a_14511_989.n2 a_14511_989.t5 475.572
R2645 a_14511_989.n1 a_14511_989.t6 469.145
R2646 a_14511_989.n6 a_14511_989.t8 454.685
R2647 a_14511_989.n6 a_14511_989.t13 428.979
R2648 a_14511_989.n2 a_14511_989.t11 384.527
R2649 a_14511_989.n1 a_14511_989.t9 384.527
R2650 a_14511_989.n3 a_14511_989.t10 370.613
R2651 a_14511_989.n5 a_14511_989.t7 314.896
R2652 a_14511_989.n7 a_14511_989.t12 311.683
R2653 a_14511_989.n13 a_14511_989.n12 305.581
R2654 a_14511_989.n7 a_14511_989.n6 171.288
R2655 a_14511_989.n14 a_14511_989.n13 159.999
R2656 a_14511_989.n15 a_14511_989.n14 157.963
R2657 a_14511_989.n3 a_14511_989.n2 128.028
R2658 a_14511_989.n4 a_14511_989.n1 126.97
R2659 a_14511_989.n14 a_14511_989.n0 91.706
R2660 a_14511_989.n5 a_14511_989.n4 55.717
R2661 a_14511_989.n12 a_14511_989.n11 30
R2662 a_14511_989.n10 a_14511_989.n9 24.383
R2663 a_14511_989.n12 a_14511_989.n10 23.684
R2664 a_14511_989.n0 a_14511_989.t4 14.282
R2665 a_14511_989.n0 a_14511_989.t3 14.282
R2666 a_14511_989.t1 a_14511_989.n15 14.282
R2667 a_14511_989.n15 a_14511_989.t0 14.282
R2668 a_14511_989.n4 a_14511_989.n3 14.151
R2669 a_14511_989.n8 a_14511_989.n7 7.597
R2670 a_14511_989.n8 a_14511_989.n5 6.509
R2671 a_14511_989.n13 a_14511_989.n8 4.65
R2672 QN.n15 QN.n14 227.387
R2673 QN.n2 QN.n1 165.613
R2674 QN.n15 QN.n2 132.893
R2675 QN.n10 QN.n5 126.225
R2676 QN.n10 QN.n9 112.771
R2677 QN.n14 QN.n13 106.052
R2678 QN.n2 QN.n0 99.355
R2679 QN.n13 QN.n11 80.526
R2680 QN.n9 QN.n8 30
R2681 QN.n13 QN.n12 30
R2682 QN.n7 QN.n6 24.383
R2683 QN.n9 QN.n7 23.684
R2684 QN.n5 QN.n4 22.578
R2685 QN.n0 QN.t4 14.282
R2686 QN.n0 QN.t2 14.282
R2687 QN.n1 QN.t0 14.282
R2688 QN.n1 QN.t6 14.282
R2689 QN.n5 QN.n3 8.58
R2690 QN.n14 QN.n10 7.053
R2691 QN.n16 QN.n15 4.65
R2692 QN.n16 QN 0.046
R2693 a_16421_1051.t5 a_16421_1051.n5 179.898
R2694 a_16421_1051.n3 a_16421_1051.n2 165.613
R2695 a_16421_1051.n3 a_16421_1051.n1 142.653
R2696 a_16421_1051.n5 a_16421_1051.n4 106.183
R2697 a_16421_1051.n5 a_16421_1051.n0 99.355
R2698 a_16421_1051.n4 a_16421_1051.n3 82.665
R2699 a_16421_1051.n4 a_16421_1051.t7 73.712
R2700 a_16421_1051.n1 a_16421_1051.t0 14.282
R2701 a_16421_1051.n1 a_16421_1051.t1 14.282
R2702 a_16421_1051.n2 a_16421_1051.t6 14.282
R2703 a_16421_1051.n2 a_16421_1051.t2 14.282
R2704 a_16421_1051.n0 a_16421_1051.t4 14.282
R2705 a_16421_1051.n0 a_16421_1051.t3 14.282
R2706 a_8142_210.n12 a_8142_210.n10 171.558
R2707 a_8142_210.n7 a_8142_210.n6 117.622
R2708 a_8142_210.n5 a_8142_210.n4 92.5
R2709 a_8142_210.n9 a_8142_210.n8 92.5
R2710 a_8142_210.n10 a_8142_210.t1 75.764
R2711 a_8142_210.n5 a_8142_210.n3 65.02
R2712 a_8142_210.n13 a_8142_210.n0 49.6
R2713 a_8142_210.n7 a_8142_210.n5 36.517
R2714 a_8142_210.n3 a_8142_210.n2 35.865
R2715 a_8142_210.n12 a_8142_210.n11 27.2
R2716 a_8142_210.n13 a_8142_210.n12 22.4
R2717 a_8142_210.n9 a_8142_210.n7 19.952
R2718 a_8142_210.t1 a_8142_210.n1 7.04
R2719 a_8142_210.n10 a_8142_210.n9 1.505
R2720 a_5327_187.n4 a_5327_187.t8 512.525
R2721 a_5327_187.n2 a_5327_187.t15 472.359
R2722 a_5327_187.n0 a_5327_187.t12 472.359
R2723 a_5327_187.n5 a_5327_187.t10 417.109
R2724 a_5327_187.n2 a_5327_187.t9 384.527
R2725 a_5327_187.n0 a_5327_187.t7 384.527
R2726 a_5327_187.n11 a_5327_187.n10 379.457
R2727 a_5327_187.n4 a_5327_187.t13 371.139
R2728 a_5327_187.n3 a_5327_187.t14 370.613
R2729 a_5327_187.n1 a_5327_187.t11 370.613
R2730 a_5327_187.n5 a_5327_187.n4 179.837
R2731 a_5327_187.n14 a_5327_187.n13 161.352
R2732 a_5327_187.n3 a_5327_187.n2 127.096
R2733 a_5327_187.n1 a_5327_187.n0 127.096
R2734 a_5327_187.n15 a_5327_187.n11 123.481
R2735 a_5327_187.n14 a_5327_187.n12 95.095
R2736 a_5327_187.n16 a_5327_187.n15 95.094
R2737 a_5327_187.n15 a_5327_187.n14 66.258
R2738 a_5327_187.n10 a_5327_187.n9 22.578
R2739 a_5327_187.n12 a_5327_187.t2 14.282
R2740 a_5327_187.n12 a_5327_187.t6 14.282
R2741 a_5327_187.n13 a_5327_187.t0 14.282
R2742 a_5327_187.n13 a_5327_187.t1 14.282
R2743 a_5327_187.t4 a_5327_187.n16 14.282
R2744 a_5327_187.n16 a_5327_187.t3 14.282
R2745 a_5327_187.n6 a_5327_187.n5 12.222
R2746 a_5327_187.n7 a_5327_187.n1 10.046
R2747 a_5327_187.n10 a_5327_187.n8 8.58
R2748 a_5327_187.n6 a_5327_187.n3 4.65
R2749 a_5327_187.n11 a_5327_187.n7 4.65
R2750 a_5327_187.n7 a_5327_187.n6 4.035
R2751 CLK.n14 CLK.t1 459.505
R2752 CLK.n11 CLK.t14 459.505
R2753 CLK.n8 CLK.t11 459.505
R2754 CLK.n5 CLK.t12 459.505
R2755 CLK.n2 CLK.t3 459.505
R2756 CLK.n0 CLK.t2 459.505
R2757 CLK.n15 CLK.t10 399.181
R2758 CLK.n12 CLK.t17 399.181
R2759 CLK.n9 CLK.t13 399.181
R2760 CLK.n6 CLK.t6 399.181
R2761 CLK.n3 CLK.t5 399.181
R2762 CLK.n1 CLK.t15 399.181
R2763 CLK.n14 CLK.t7 384.527
R2764 CLK.n11 CLK.t4 384.527
R2765 CLK.n8 CLK.t16 384.527
R2766 CLK.n5 CLK.t0 384.527
R2767 CLK.n2 CLK.t9 384.527
R2768 CLK.n0 CLK.t8 384.527
R2769 CLK.n15 CLK.n14 33.832
R2770 CLK.n1 CLK.n0 33.832
R2771 CLK.n3 CLK.n2 33.832
R2772 CLK.n6 CLK.n5 33.832
R2773 CLK.n9 CLK.n8 33.832
R2774 CLK.n12 CLK.n11 33.832
R2775 CLK.n4 CLK.n1 11.555
R2776 CLK.n7 CLK.n4 9.476
R2777 CLK.n10 CLK.n7 9.476
R2778 CLK.n13 CLK.n10 9.476
R2779 CLK.n16 CLK.n13 9.476
R2780 CLK.n4 CLK.n3 2.079
R2781 CLK.n7 CLK.n6 2.079
R2782 CLK.n10 CLK.n9 2.079
R2783 CLK.n13 CLK.n12 2.079
R2784 CLK.n16 CLK.n15 2.079
R2785 CLK.n16 CLK 0.046
R2786 a_2141_1050.n1 a_2141_1050.t5 512.525
R2787 a_2141_1050.n1 a_2141_1050.t6 371.139
R2788 a_2141_1050.n2 a_2141_1050.t7 361.392
R2789 a_2141_1050.n4 a_2141_1050.n3 327.32
R2790 a_2141_1050.n2 a_2141_1050.n1 235.554
R2791 a_2141_1050.n5 a_2141_1050.n4 159.999
R2792 a_2141_1050.n6 a_2141_1050.n5 157.963
R2793 a_2141_1050.n5 a_2141_1050.n0 91.706
R2794 a_2141_1050.n0 a_2141_1050.t4 14.282
R2795 a_2141_1050.n0 a_2141_1050.t3 14.282
R2796 a_2141_1050.t2 a_2141_1050.n6 14.282
R2797 a_2141_1050.n6 a_2141_1050.t1 14.282
R2798 a_2141_1050.n4 a_2141_1050.n2 10.615
R2799 a_9009_1050.n1 a_9009_1050.t8 480.392
R2800 a_9009_1050.n1 a_9009_1050.t7 403.272
R2801 a_9009_1050.n2 a_9009_1050.t9 385.063
R2802 a_9009_1050.n4 a_9009_1050.n3 357.814
R2803 a_9009_1050.n7 a_9009_1050.n6 161.352
R2804 a_9009_1050.n5 a_9009_1050.n4 151.34
R2805 a_9009_1050.n2 a_9009_1050.n1 143.429
R2806 a_9009_1050.n5 a_9009_1050.n0 95.095
R2807 a_9009_1050.n8 a_9009_1050.n7 95.094
R2808 a_9009_1050.n7 a_9009_1050.n5 66.258
R2809 a_9009_1050.n0 a_9009_1050.t3 14.282
R2810 a_9009_1050.n0 a_9009_1050.t6 14.282
R2811 a_9009_1050.n6 a_9009_1050.t0 14.282
R2812 a_9009_1050.n6 a_9009_1050.t2 14.282
R2813 a_9009_1050.t5 a_9009_1050.n8 14.282
R2814 a_9009_1050.n8 a_9009_1050.t4 14.282
R2815 a_9009_1050.n4 a_9009_1050.n2 10.615
R2816 a_9331_989.n3 a_9331_989.t9 512.525
R2817 a_9331_989.n1 a_9331_989.t12 477.179
R2818 a_9331_989.n6 a_9331_989.t10 454.685
R2819 a_9331_989.n2 a_9331_989.t7 440.954
R2820 a_9331_989.n6 a_9331_989.t5 428.979
R2821 a_9331_989.n1 a_9331_989.t8 406.485
R2822 a_9331_989.n3 a_9331_989.t6 371.139
R2823 a_9331_989.n5 a_9331_989.t11 322.918
R2824 a_9331_989.n7 a_9331_989.t13 283.824
R2825 a_9331_989.n13 a_9331_989.n12 277.722
R2826 a_9331_989.n7 a_9331_989.n6 199.147
R2827 a_9331_989.n14 a_9331_989.n13 187.858
R2828 a_9331_989.n15 a_9331_989.n14 157.963
R2829 a_9331_989.n5 a_9331_989.n4 111.608
R2830 a_9331_989.n14 a_9331_989.n0 91.706
R2831 a_9331_989.n4 a_9331_989.n3 77.972
R2832 a_9331_989.n12 a_9331_989.n11 30
R2833 a_9331_989.n8 a_9331_989.n5 24.737
R2834 a_9331_989.n10 a_9331_989.n9 24.383
R2835 a_9331_989.n12 a_9331_989.n10 23.684
R2836 a_9331_989.n2 a_9331_989.n1 21.4
R2837 a_9331_989.n0 a_9331_989.t3 14.282
R2838 a_9331_989.n0 a_9331_989.t4 14.282
R2839 a_9331_989.n15 a_9331_989.t0 14.282
R2840 a_9331_989.t1 a_9331_989.n15 14.282
R2841 a_9331_989.n8 a_9331_989.n7 7.597
R2842 a_9331_989.n4 a_9331_989.n2 6.833
R2843 a_9331_989.n13 a_9331_989.n8 4.65
R2844 a_147_187.n4 a_147_187.t15 512.525
R2845 a_147_187.n2 a_147_187.t9 472.359
R2846 a_147_187.n0 a_147_187.t14 472.359
R2847 a_147_187.n5 a_147_187.t12 417.109
R2848 a_147_187.n2 a_147_187.t13 384.527
R2849 a_147_187.n0 a_147_187.t10 384.527
R2850 a_147_187.n4 a_147_187.t11 371.139
R2851 a_147_187.n3 a_147_187.t8 370.613
R2852 a_147_187.n1 a_147_187.t7 370.613
R2853 a_147_187.n12 a_147_187.n11 363.934
R2854 a_147_187.n5 a_147_187.n4 179.837
R2855 a_147_187.n15 a_147_187.n14 161.352
R2856 a_147_187.n3 a_147_187.n2 127.096
R2857 a_147_187.n1 a_147_187.n0 127.096
R2858 a_147_187.n16 a_147_187.n12 123.481
R2859 a_147_187.n15 a_147_187.n13 95.095
R2860 a_147_187.n17 a_147_187.n16 95.094
R2861 a_147_187.n16 a_147_187.n15 66.258
R2862 a_147_187.n11 a_147_187.n10 30
R2863 a_147_187.n9 a_147_187.n8 24.383
R2864 a_147_187.n11 a_147_187.n9 23.684
R2865 a_147_187.n13 a_147_187.t5 14.282
R2866 a_147_187.n13 a_147_187.t6 14.282
R2867 a_147_187.n14 a_147_187.t4 14.282
R2868 a_147_187.n14 a_147_187.t3 14.282
R2869 a_147_187.n17 a_147_187.t1 14.282
R2870 a_147_187.t2 a_147_187.n17 14.282
R2871 a_147_187.n6 a_147_187.n5 12.222
R2872 a_147_187.n7 a_147_187.n1 10.046
R2873 a_147_187.n6 a_147_187.n3 4.65
R2874 a_147_187.n12 a_147_187.n7 4.65
R2875 a_147_187.n7 a_147_187.n6 4.035
R2876 a_4626_101.n5 a_4626_101.n4 62.817
R2877 a_4626_101.n2 a_4626_101.n0 41.528
R2878 a_4626_101.n5 a_4626_101.n3 26.202
R2879 a_4626_101.t0 a_4626_101.n5 19.737
R2880 a_4626_101.t0 a_4626_101.n6 8.137
R2881 a_4626_101.n2 a_4626_101.n1 3.644
R2882 a_4626_101.t0 a_4626_101.n2 1.093
R2883 a_4151_989.n1 a_4151_989.t11 512.525
R2884 a_4151_989.n0 a_4151_989.t7 512.525
R2885 a_4151_989.n5 a_4151_989.t5 454.685
R2886 a_4151_989.n5 a_4151_989.t8 428.979
R2887 a_4151_989.n1 a_4151_989.t6 371.139
R2888 a_4151_989.n0 a_4151_989.t12 371.139
R2889 a_4151_989.n2 a_4151_989.n1 343.521
R2890 a_4151_989.n4 a_4151_989.n0 287.803
R2891 a_4151_989.n9 a_4151_989.n8 271.602
R2892 a_4151_989.n6 a_4151_989.t9 244.718
R2893 a_4151_989.n6 a_4151_989.n5 227.006
R2894 a_4151_989.n11 a_4151_989.n9 215.717
R2895 a_4151_989.n2 a_4151_989.t13 172.106
R2896 a_4151_989.n3 a_4151_989.t10 165.68
R2897 a_4151_989.n11 a_4151_989.n10 157.964
R2898 a_4151_989.n12 a_4151_989.n11 91.705
R2899 a_4151_989.n4 a_4151_989.n3 55.717
R2900 a_4151_989.n7 a_4151_989.n4 47.59
R2901 a_4151_989.n10 a_4151_989.t0 14.282
R2902 a_4151_989.n10 a_4151_989.t1 14.282
R2903 a_4151_989.n12 a_4151_989.t2 14.282
R2904 a_4151_989.t3 a_4151_989.n12 14.282
R2905 a_4151_989.n3 a_4151_989.n2 10.343
R2906 a_4151_989.n7 a_4151_989.n6 7.597
R2907 a_4151_989.n9 a_4151_989.n7 4.65
R2908 a_1053_103.n5 a_1053_103.n4 66.708
R2909 a_1053_103.n2 a_1053_103.n0 32.662
R2910 a_1053_103.n5 a_1053_103.n3 19.496
R2911 a_1053_103.t0 a_1053_103.n5 13.756
R2912 a_1053_103.t0 a_1053_103.n2 3.034
R2913 a_1053_103.n2 a_1053_103.n1 0.443
R2914 a_1334_210.n10 a_1334_210.n8 171.558
R2915 a_1334_210.n8 a_1334_210.t1 75.764
R2916 a_1334_210.n11 a_1334_210.n0 49.6
R2917 a_1334_210.n3 a_1334_210.n2 27.476
R2918 a_1334_210.n10 a_1334_210.n9 27.2
R2919 a_1334_210.n11 a_1334_210.n10 22.4
R2920 a_1334_210.t1 a_1334_210.n5 20.241
R2921 a_1334_210.n7 a_1334_210.n6 19.952
R2922 a_1334_210.t1 a_1334_210.n3 13.984
R2923 a_1334_210.n5 a_1334_210.n4 13.494
R2924 a_1334_210.t1 a_1334_210.n1 7.04
R2925 a_1334_210.n8 a_1334_210.n7 1.505
R2926 a_277_1050.n2 a_277_1050.t8 512.525
R2927 a_277_1050.n0 a_277_1050.t7 512.525
R2928 a_277_1050.n3 a_277_1050.t12 389.251
R2929 a_277_1050.n1 a_277_1050.t11 389.251
R2930 a_277_1050.n2 a_277_1050.t10 371.139
R2931 a_277_1050.n0 a_277_1050.t9 371.139
R2932 a_277_1050.n9 a_277_1050.n8 336.075
R2933 a_277_1050.n3 a_277_1050.n2 207.695
R2934 a_277_1050.n1 a_277_1050.n0 207.695
R2935 a_277_1050.n12 a_277_1050.n11 161.352
R2936 a_277_1050.n13 a_277_1050.n9 151.34
R2937 a_277_1050.n12 a_277_1050.n10 95.095
R2938 a_277_1050.n14 a_277_1050.n13 95.094
R2939 a_277_1050.n13 a_277_1050.n12 66.258
R2940 a_277_1050.n8 a_277_1050.n7 30
R2941 a_277_1050.n6 a_277_1050.n5 24.383
R2942 a_277_1050.n8 a_277_1050.n6 23.684
R2943 a_277_1050.n10 a_277_1050.t4 14.282
R2944 a_277_1050.n10 a_277_1050.t3 14.282
R2945 a_277_1050.n11 a_277_1050.t5 14.282
R2946 a_277_1050.n11 a_277_1050.t6 14.282
R2947 a_277_1050.t2 a_277_1050.n14 14.282
R2948 a_277_1050.n14 a_277_1050.t1 14.282
R2949 a_277_1050.n4 a_277_1050.n1 14.126
R2950 a_277_1050.n9 a_277_1050.n4 5.965
R2951 a_277_1050.n4 a_277_1050.n3 4.65
R2952 a_5457_1050.n3 a_5457_1050.t7 512.525
R2953 a_5457_1050.n1 a_5457_1050.t8 512.525
R2954 a_5457_1050.n4 a_5457_1050.t11 389.251
R2955 a_5457_1050.n2 a_5457_1050.t10 389.251
R2956 a_5457_1050.n3 a_5457_1050.t12 371.139
R2957 a_5457_1050.n1 a_5457_1050.t9 371.139
R2958 a_5457_1050.n7 a_5457_1050.n6 357.814
R2959 a_5457_1050.n4 a_5457_1050.n3 207.695
R2960 a_5457_1050.n2 a_5457_1050.n1 207.695
R2961 a_5457_1050.n10 a_5457_1050.n9 161.352
R2962 a_5457_1050.n8 a_5457_1050.n7 151.34
R2963 a_5457_1050.n8 a_5457_1050.n0 95.095
R2964 a_5457_1050.n11 a_5457_1050.n10 95.094
R2965 a_5457_1050.n10 a_5457_1050.n8 66.258
R2966 a_5457_1050.n0 a_5457_1050.t1 14.282
R2967 a_5457_1050.n0 a_5457_1050.t0 14.282
R2968 a_5457_1050.n9 a_5457_1050.t6 14.282
R2969 a_5457_1050.n9 a_5457_1050.t5 14.282
R2970 a_5457_1050.t4 a_5457_1050.n11 14.282
R2971 a_5457_1050.n11 a_5457_1050.t3 14.282
R2972 a_5457_1050.n5 a_5457_1050.n2 14.126
R2973 a_5457_1050.n7 a_5457_1050.n5 5.965
R2974 a_5457_1050.n5 a_5457_1050.n4 4.65
R2975 a_5779_989.n1 a_5779_989.t11 480.392
R2976 a_5779_989.n3 a_5779_989.t12 454.685
R2977 a_5779_989.n3 a_5779_989.t10 428.979
R2978 a_5779_989.n1 a_5779_989.t9 403.272
R2979 a_5779_989.n2 a_5779_989.t8 357.204
R2980 a_5779_989.n4 a_5779_989.t7 311.683
R2981 a_5779_989.n10 a_5779_989.n9 308.216
R2982 a_5779_989.n11 a_5779_989.n10 179.199
R2983 a_5779_989.n4 a_5779_989.n3 171.288
R2984 a_5779_989.n2 a_5779_989.n1 171.288
R2985 a_5779_989.n13 a_5779_989.n12 161.352
R2986 a_5779_989.n11 a_5779_989.n0 95.095
R2987 a_5779_989.n14 a_5779_989.n13 95.094
R2988 a_5779_989.n13 a_5779_989.n11 66.258
R2989 a_5779_989.n9 a_5779_989.n8 30
R2990 a_5779_989.n7 a_5779_989.n6 24.383
R2991 a_5779_989.n9 a_5779_989.n7 23.684
R2992 a_5779_989.n0 a_5779_989.t3 14.282
R2993 a_5779_989.n0 a_5779_989.t2 14.282
R2994 a_5779_989.n12 a_5779_989.t6 14.282
R2995 a_5779_989.n12 a_5779_989.t5 14.282
R2996 a_5779_989.t1 a_5779_989.n14 14.282
R2997 a_5779_989.n14 a_5779_989.t0 14.282
R2998 a_5779_989.n5 a_5779_989.n4 8.685
R2999 a_5779_989.n5 a_5779_989.n2 5.965
R3000 a_5779_989.n10 a_5779_989.n5 4.65
R3001 a_12396_101.n5 a_12396_101.n4 62.817
R3002 a_12396_101.n2 a_12396_101.n0 41.528
R3003 a_12396_101.n5 a_12396_101.n3 26.202
R3004 a_12396_101.t0 a_12396_101.n5 19.737
R3005 a_12396_101.t0 a_12396_101.n6 8.137
R3006 a_12396_101.n2 a_12396_101.n1 3.644
R3007 a_12396_101.t0 a_12396_101.n2 1.093
R3008 a_3829_1050.n1 a_3829_1050.t9 480.392
R3009 a_3829_1050.n1 a_3829_1050.t7 403.272
R3010 a_3829_1050.n2 a_3829_1050.t8 385.063
R3011 a_3829_1050.n7 a_3829_1050.n6 336.075
R3012 a_3829_1050.n10 a_3829_1050.n9 161.352
R3013 a_3829_1050.n8 a_3829_1050.n7 151.34
R3014 a_3829_1050.n2 a_3829_1050.n1 143.429
R3015 a_3829_1050.n8 a_3829_1050.n0 95.095
R3016 a_3829_1050.n11 a_3829_1050.n10 95.094
R3017 a_3829_1050.n10 a_3829_1050.n8 66.258
R3018 a_3829_1050.n6 a_3829_1050.n5 30
R3019 a_3829_1050.n4 a_3829_1050.n3 24.383
R3020 a_3829_1050.n6 a_3829_1050.n4 23.684
R3021 a_3829_1050.n0 a_3829_1050.t3 14.282
R3022 a_3829_1050.n0 a_3829_1050.t4 14.282
R3023 a_3829_1050.n9 a_3829_1050.t6 14.282
R3024 a_3829_1050.n9 a_3829_1050.t5 14.282
R3025 a_3829_1050.t1 a_3829_1050.n11 14.282
R3026 a_3829_1050.n11 a_3829_1050.t0 14.282
R3027 a_3829_1050.n7 a_3829_1050.n2 10.615
R3028 a_2036_101.n11 a_2036_101.n10 68.43
R3029 a_2036_101.n3 a_2036_101.n2 62.817
R3030 a_2036_101.n7 a_2036_101.n6 38.626
R3031 a_2036_101.n6 a_2036_101.n5 35.955
R3032 a_2036_101.n3 a_2036_101.n1 26.202
R3033 a_2036_101.t0 a_2036_101.n3 19.737
R3034 a_2036_101.t1 a_2036_101.n8 8.137
R3035 a_2036_101.t0 a_2036_101.n4 7.273
R3036 a_2036_101.t0 a_2036_101.n0 6.109
R3037 a_2036_101.t1 a_2036_101.n7 4.864
R3038 a_2036_101.t0 a_2036_101.n12 2.074
R3039 a_2036_101.n12 a_2036_101.t1 0.937
R3040 a_2036_101.t1 a_2036_101.n11 0.763
R3041 a_2036_101.n11 a_2036_101.n9 0.185
R3042 a_10451_103.n5 a_10451_103.n4 66.708
R3043 a_10451_103.n2 a_10451_103.n0 32.662
R3044 a_10451_103.n5 a_10451_103.n3 19.496
R3045 a_10451_103.t0 a_10451_103.n5 13.756
R3046 a_10451_103.t0 a_10451_103.n2 3.034
R3047 a_10451_103.n2 a_10451_103.n1 0.443
R3048 a_15757_1051.n2 a_15757_1051.t6 179.895
R3049 a_15757_1051.n4 a_15757_1051.n0 157.021
R3050 a_15757_1051.n5 a_15757_1051.n4 124.954
R3051 a_15757_1051.n3 a_15757_1051.n2 106.183
R3052 a_15757_1051.n2 a_15757_1051.n1 99.355
R3053 a_15757_1051.n4 a_15757_1051.n3 82.65
R3054 a_15757_1051.n3 a_15757_1051.t5 73.712
R3055 a_15757_1051.n1 a_15757_1051.t7 14.282
R3056 a_15757_1051.n1 a_15757_1051.t4 14.282
R3057 a_15757_1051.n0 a_15757_1051.t2 14.282
R3058 a_15757_1051.n0 a_15757_1051.t3 14.282
R3059 a_15757_1051.t1 a_15757_1051.n5 14.282
R3060 a_15757_1051.n5 a_15757_1051.t0 14.282
R3061 a_15652_101.n4 a_15652_101.n2 41.528
R3062 a_15652_101.n1 a_15652_101.n0 33.123
R3063 a_15652_101.t0 a_15652_101.n1 10.642
R3064 a_15652_101.n6 a_15652_101.n5 7.966
R3065 a_15652_101.n4 a_15652_101.n3 3.644
R3066 a_15652_101.t0 a_15652_101.n4 1.093
R3067 a_15652_101.t0 a_15652_101.n6 0.088
R3068 a_6514_210.n10 a_6514_210.n8 171.558
R3069 a_6514_210.n8 a_6514_210.t1 75.764
R3070 a_6514_210.n3 a_6514_210.n2 27.476
R3071 a_6514_210.n10 a_6514_210.n9 27.2
R3072 a_6514_210.n11 a_6514_210.n0 23.498
R3073 a_6514_210.n11 a_6514_210.n10 22.4
R3074 a_6514_210.t1 a_6514_210.n5 20.241
R3075 a_6514_210.n7 a_6514_210.n6 19.952
R3076 a_6514_210.t1 a_6514_210.n3 13.984
R3077 a_6514_210.n5 a_6514_210.n4 13.494
R3078 a_6514_210.t1 a_6514_210.n1 7.04
R3079 a_6514_210.n8 a_6514_210.n7 1.505
R3080 a_11694_210.n10 a_11694_210.n8 171.558
R3081 a_11694_210.n8 a_11694_210.t1 75.764
R3082 a_11694_210.n11 a_11694_210.n0 49.6
R3083 a_11694_210.n3 a_11694_210.n2 27.476
R3084 a_11694_210.n10 a_11694_210.n9 27.2
R3085 a_11694_210.n11 a_11694_210.n10 22.4
R3086 a_11694_210.t1 a_11694_210.n5 20.241
R3087 a_11694_210.n7 a_11694_210.n6 19.952
R3088 a_11694_210.t1 a_11694_210.n3 13.984
R3089 a_11694_210.n5 a_11694_210.n4 13.494
R3090 a_11694_210.t1 a_11694_210.n1 7.04
R3091 a_11694_210.n8 a_11694_210.n7 1.505
R3092 a_14986_101.n11 a_14986_101.n10 68.43
R3093 a_14986_101.n3 a_14986_101.n2 62.817
R3094 a_14986_101.n7 a_14986_101.n6 38.626
R3095 a_14986_101.n6 a_14986_101.n5 35.955
R3096 a_14986_101.n3 a_14986_101.n1 26.202
R3097 a_14986_101.t0 a_14986_101.n3 19.737
R3098 a_14986_101.t1 a_14986_101.n8 8.137
R3099 a_14986_101.t0 a_14986_101.n4 7.273
R3100 a_14986_101.t0 a_14986_101.n0 6.109
R3101 a_14986_101.t1 a_14986_101.n7 4.864
R3102 a_14986_101.t0 a_14986_101.n12 2.074
R3103 a_14986_101.n12 a_14986_101.t1 0.937
R3104 a_14986_101.t1 a_14986_101.n11 0.763
R3105 a_14986_101.n11 a_14986_101.n9 0.185
R3106 a_12501_1050.n1 a_12501_1050.t7 512.525
R3107 a_12501_1050.n1 a_12501_1050.t5 371.139
R3108 a_12501_1050.n2 a_12501_1050.t6 361.392
R3109 a_12501_1050.n4 a_12501_1050.n3 327.32
R3110 a_12501_1050.n2 a_12501_1050.n1 235.554
R3111 a_12501_1050.n5 a_12501_1050.n4 159.999
R3112 a_12501_1050.n6 a_12501_1050.n5 157.963
R3113 a_12501_1050.n5 a_12501_1050.n0 91.706
R3114 a_12501_1050.n0 a_12501_1050.t4 14.282
R3115 a_12501_1050.n0 a_12501_1050.t3 14.282
R3116 a_12501_1050.t1 a_12501_1050.n6 14.282
R3117 a_12501_1050.n6 a_12501_1050.t0 14.282
R3118 a_12501_1050.n4 a_12501_1050.n2 10.615
R3119 a_7321_1050.n1 a_7321_1050.t5 512.525
R3120 a_7321_1050.n1 a_7321_1050.t7 371.139
R3121 a_7321_1050.n2 a_7321_1050.t6 361.392
R3122 a_7321_1050.n7 a_7321_1050.n6 305.581
R3123 a_7321_1050.n2 a_7321_1050.n1 235.554
R3124 a_7321_1050.n8 a_7321_1050.n7 159.999
R3125 a_7321_1050.n9 a_7321_1050.n8 157.963
R3126 a_7321_1050.n8 a_7321_1050.n0 91.706
R3127 a_7321_1050.n6 a_7321_1050.n5 30
R3128 a_7321_1050.n4 a_7321_1050.n3 24.383
R3129 a_7321_1050.n6 a_7321_1050.n4 23.684
R3130 a_7321_1050.n0 a_7321_1050.t3 14.282
R3131 a_7321_1050.n0 a_7321_1050.t4 14.282
R3132 a_7321_1050.n9 a_7321_1050.t0 14.282
R3133 a_7321_1050.t1 a_7321_1050.n9 14.282
R3134 a_7321_1050.n7 a_7321_1050.n2 10.615
R3135 a_8823_103.t0 a_8823_103.n7 59.616
R3136 a_8823_103.n4 a_8823_103.n2 54.496
R3137 a_8823_103.n4 a_8823_103.n3 54.496
R3138 a_8823_103.n1 a_8823_103.n0 24.679
R3139 a_8823_103.n6 a_8823_103.n4 7.859
R3140 a_8823_103.t0 a_8823_103.n1 7.505
R3141 a_8823_103.t0 a_8823_103.n6 3.034
R3142 a_8823_103.n6 a_8823_103.n5 0.443
R3143 a_9104_210.n10 a_9104_210.n8 171.558
R3144 a_9104_210.n8 a_9104_210.t1 75.764
R3145 a_9104_210.n11 a_9104_210.n0 49.6
R3146 a_9104_210.n3 a_9104_210.n2 27.476
R3147 a_9104_210.n10 a_9104_210.n9 27.2
R3148 a_9104_210.n11 a_9104_210.n10 22.4
R3149 a_9104_210.t1 a_9104_210.n5 20.241
R3150 a_9104_210.n7 a_9104_210.n6 19.952
R3151 a_9104_210.t1 a_9104_210.n3 13.984
R3152 a_9104_210.n5 a_9104_210.n4 13.494
R3153 a_9104_210.t1 a_9104_210.n1 7.04
R3154 a_9104_210.n8 a_9104_210.n7 1.505
R3155 a_16318_101.n2 a_16318_101.n0 42.755
R3156 a_16318_101.n2 a_16318_101.n1 2.198
R3157 a_16318_101.t0 a_16318_101.n2 0.106
R3158 a_372_210.n9 a_372_210.n7 171.558
R3159 a_372_210.t0 a_372_210.n9 75.765
R3160 a_372_210.n3 a_372_210.n1 74.827
R3161 a_372_210.n3 a_372_210.n2 27.476
R3162 a_372_210.n7 a_372_210.n6 27.2
R3163 a_372_210.n5 a_372_210.n4 23.498
R3164 a_372_210.n7 a_372_210.n5 22.4
R3165 a_372_210.t0 a_372_210.n11 20.241
R3166 a_372_210.t0 a_372_210.n3 13.984
R3167 a_372_210.n11 a_372_210.n10 13.494
R3168 a_372_210.t0 a_372_210.n0 8.137
R3169 a_372_210.n9 a_372_210.n8 1.505
R3170 a_10732_210.n8 a_10732_210.n6 185.173
R3171 a_10732_210.t0 a_10732_210.n8 75.765
R3172 a_10732_210.n3 a_10732_210.n1 74.827
R3173 a_10732_210.n3 a_10732_210.n2 27.476
R3174 a_10732_210.n6 a_10732_210.n5 22.349
R3175 a_10732_210.t0 a_10732_210.n10 20.241
R3176 a_10732_210.t0 a_10732_210.n3 13.984
R3177 a_10732_210.n10 a_10732_210.n9 13.494
R3178 a_10732_210.n6 a_10732_210.n4 8.443
R3179 a_10732_210.t0 a_10732_210.n0 8.137
R3180 a_10732_210.n8 a_10732_210.n7 1.505
R3181 a_6233_103.t0 a_6233_103.n7 59.616
R3182 a_6233_103.n4 a_6233_103.n2 54.496
R3183 a_6233_103.n4 a_6233_103.n3 54.496
R3184 a_6233_103.n1 a_6233_103.n0 24.679
R3185 a_6233_103.t0 a_6233_103.n1 7.505
R3186 a_6233_103.n6 a_6233_103.n5 2.455
R3187 a_6233_103.n6 a_6233_103.n4 0.636
R3188 a_6233_103.t0 a_6233_103.n6 0.246
R3189 a_5552_210.n9 a_5552_210.n7 171.558
R3190 a_5552_210.t0 a_5552_210.n9 75.765
R3191 a_5552_210.n3 a_5552_210.n1 74.827
R3192 a_5552_210.n3 a_5552_210.n2 27.476
R3193 a_5552_210.n7 a_5552_210.n6 27.2
R3194 a_5552_210.n5 a_5552_210.n4 23.498
R3195 a_5552_210.n7 a_5552_210.n5 22.4
R3196 a_5552_210.t0 a_5552_210.n11 20.241
R3197 a_5552_210.t0 a_5552_210.n3 13.984
R3198 a_5552_210.n11 a_5552_210.n10 13.494
R3199 a_5552_210.t0 a_5552_210.n0 8.137
R3200 a_5552_210.n9 a_5552_210.n8 1.505
R3201 a_16984_101.n3 a_16984_101.n1 42.788
R3202 a_16984_101.t0 a_16984_101.n0 8.137
R3203 a_16984_101.n3 a_16984_101.n2 4.665
R3204 a_16984_101.t0 a_16984_101.n3 0.06
R3205 a_2962_210.n9 a_2962_210.n7 171.558
R3206 a_2962_210.t0 a_2962_210.n9 75.765
R3207 a_2962_210.n3 a_2962_210.n1 74.827
R3208 a_2962_210.n3 a_2962_210.n2 27.476
R3209 a_2962_210.n7 a_2962_210.n6 27.2
R3210 a_2962_210.n5 a_2962_210.n4 23.498
R3211 a_2962_210.n7 a_2962_210.n5 22.4
R3212 a_2962_210.t0 a_2962_210.n11 20.241
R3213 a_2962_210.t0 a_2962_210.n3 13.984
R3214 a_2962_210.n11 a_2962_210.n10 13.494
R3215 a_2962_210.t0 a_2962_210.n0 8.137
R3216 a_2962_210.n9 a_2962_210.n8 1.505
R3217 a_7861_103.n5 a_7861_103.n4 66.708
R3218 a_7861_103.n2 a_7861_103.n0 25.439
R3219 a_7861_103.n5 a_7861_103.n3 19.496
R3220 a_7861_103.t0 a_7861_103.n5 13.756
R3221 a_7861_103.n2 a_7861_103.n1 2.455
R3222 a_7861_103.t0 a_7861_103.n2 0.246
R3223 a_9806_101.n11 a_9806_101.n10 68.43
R3224 a_9806_101.n3 a_9806_101.n2 62.817
R3225 a_9806_101.n7 a_9806_101.n6 38.626
R3226 a_9806_101.n6 a_9806_101.n5 35.955
R3227 a_9806_101.n3 a_9806_101.n1 26.202
R3228 a_9806_101.t0 a_9806_101.n3 19.737
R3229 a_9806_101.t1 a_9806_101.n8 8.137
R3230 a_9806_101.t0 a_9806_101.n4 7.273
R3231 a_9806_101.t0 a_9806_101.n0 6.109
R3232 a_9806_101.t1 a_9806_101.n7 4.864
R3233 a_9806_101.t0 a_9806_101.n12 2.074
R3234 a_9806_101.n12 a_9806_101.t1 0.937
R3235 a_9806_101.t1 a_9806_101.n11 0.763
R3236 a_9806_101.n11 a_9806_101.n9 0.185
R3237 a_7216_101.n11 a_7216_101.n10 68.43
R3238 a_7216_101.n3 a_7216_101.n2 62.817
R3239 a_7216_101.n7 a_7216_101.n6 38.626
R3240 a_7216_101.n6 a_7216_101.n5 35.955
R3241 a_7216_101.n3 a_7216_101.n1 26.202
R3242 a_7216_101.t0 a_7216_101.n3 19.737
R3243 a_7216_101.t1 a_7216_101.n8 8.137
R3244 a_7216_101.t0 a_7216_101.n4 7.273
R3245 a_7216_101.t0 a_7216_101.n0 6.109
R3246 a_7216_101.t1 a_7216_101.n7 4.864
R3247 a_7216_101.t0 a_7216_101.n12 2.074
R3248 a_7216_101.n12 a_7216_101.t1 0.937
R3249 a_7216_101.t1 a_7216_101.n11 0.763
R3250 a_7216_101.n11 a_7216_101.n9 0.185
R3251 a_91_103.t0 a_91_103.n7 59.616
R3252 a_91_103.n4 a_91_103.n2 54.496
R3253 a_91_103.n4 a_91_103.n3 54.496
R3254 a_91_103.n1 a_91_103.n0 24.679
R3255 a_91_103.t0 a_91_103.n1 7.505
R3256 a_91_103.n6 a_91_103.n5 2.455
R3257 a_91_103.n6 a_91_103.n4 0.636
R3258 a_91_103.t0 a_91_103.n6 0.246
R3259 a_5271_103.t0 a_5271_103.n7 59.616
R3260 a_5271_103.n4 a_5271_103.n2 54.496
R3261 a_5271_103.n4 a_5271_103.n3 54.496
R3262 a_5271_103.n1 a_5271_103.n0 24.679
R3263 a_5271_103.t0 a_5271_103.n1 7.505
R3264 a_5271_103.n6 a_5271_103.n5 2.455
R3265 a_5271_103.n6 a_5271_103.n4 0.636
R3266 a_5271_103.t0 a_5271_103.n6 0.246
R3267 a_3924_210.n10 a_3924_210.n8 171.558
R3268 a_3924_210.n8 a_3924_210.t1 75.764
R3269 a_3924_210.n3 a_3924_210.n2 27.476
R3270 a_3924_210.n10 a_3924_210.n9 27.2
R3271 a_3924_210.n11 a_3924_210.n0 23.498
R3272 a_3924_210.n11 a_3924_210.n10 22.4
R3273 a_3924_210.t1 a_3924_210.n5 20.241
R3274 a_3924_210.n7 a_3924_210.n6 19.952
R3275 a_3924_210.t1 a_3924_210.n3 13.984
R3276 a_3924_210.n5 a_3924_210.n4 13.494
R3277 a_3924_210.t1 a_3924_210.n1 7.04
R3278 a_3924_210.n8 a_3924_210.n7 1.505
R3279 a_13322_210.n9 a_13322_210.n7 171.558
R3280 a_13322_210.t0 a_13322_210.n9 75.765
R3281 a_13322_210.n3 a_13322_210.n1 74.827
R3282 a_13322_210.n3 a_13322_210.n2 27.476
R3283 a_13322_210.n7 a_13322_210.n6 27.2
R3284 a_13322_210.n5 a_13322_210.n4 23.498
R3285 a_13322_210.n7 a_13322_210.n5 22.4
R3286 a_13322_210.t0 a_13322_210.n11 20.241
R3287 a_13322_210.t0 a_13322_210.n3 13.984
R3288 a_13322_210.n11 a_13322_210.n10 13.494
R3289 a_13322_210.t0 a_13322_210.n0 8.137
R3290 a_13322_210.n9 a_13322_210.n8 1.505
R3291 a_14284_210.n10 a_14284_210.n8 171.558
R3292 a_14284_210.n8 a_14284_210.t1 75.764
R3293 a_14284_210.n3 a_14284_210.n2 27.476
R3294 a_14284_210.n10 a_14284_210.n9 27.2
R3295 a_14284_210.n11 a_14284_210.n0 23.498
R3296 a_14284_210.n11 a_14284_210.n10 22.4
R3297 a_14284_210.t1 a_14284_210.n5 20.241
R3298 a_14284_210.n7 a_14284_210.n6 19.952
R3299 a_14284_210.t1 a_14284_210.n3 13.984
R3300 a_14284_210.n5 a_14284_210.n4 13.494
R3301 a_14284_210.t1 a_14284_210.n1 7.04
R3302 a_14284_210.n8 a_14284_210.n7 1.505
R3303 a_13041_103.n5 a_13041_103.n4 66.708
R3304 a_13041_103.n2 a_13041_103.n0 25.439
R3305 a_13041_103.n5 a_13041_103.n3 19.496
R3306 a_13041_103.t0 a_13041_103.n5 13.756
R3307 a_13041_103.n2 a_13041_103.n1 2.455
R3308 a_13041_103.t0 a_13041_103.n2 0.246
R3309 a_3643_103.t0 a_3643_103.n7 59.616
R3310 a_3643_103.n4 a_3643_103.n2 54.496
R3311 a_3643_103.n4 a_3643_103.n3 54.496
R3312 a_3643_103.n1 a_3643_103.n0 24.679
R3313 a_3643_103.t0 a_3643_103.n1 7.505
R3314 a_3643_103.n6 a_3643_103.n5 2.455
R3315 a_3643_103.n6 a_3643_103.n4 0.636
R3316 a_3643_103.t0 a_3643_103.n6 0.246
R3317 a_14003_103.n5 a_14003_103.n4 66.708
R3318 a_14003_103.n2 a_14003_103.n0 25.439
R3319 a_14003_103.n5 a_14003_103.n3 19.496
R3320 a_14003_103.t0 a_14003_103.n5 13.756
R3321 a_14003_103.n2 a_14003_103.n1 2.455
R3322 a_14003_103.t0 a_14003_103.n2 0.246
R3323 a_2681_103.n5 a_2681_103.n4 66.708
R3324 a_2681_103.n2 a_2681_103.n0 25.439
R3325 a_2681_103.n5 a_2681_103.n3 19.496
R3326 a_2681_103.t0 a_2681_103.n5 13.756
R3327 a_2681_103.n2 a_2681_103.n1 2.455
R3328 a_2681_103.t0 a_2681_103.n2 0.246
C7 RN GND 7.36fF
C8 VDD GND 28.70fF
C9 a_2681_103.n0 GND 0.11fF
C10 a_2681_103.n1 GND 0.04fF
C11 a_2681_103.n2 GND 0.03fF
C12 a_2681_103.n3 GND 0.07fF
C13 a_2681_103.n4 GND 0.08fF
C14 a_2681_103.n5 GND 0.03fF
C15 a_14003_103.n0 GND 0.11fF
C16 a_14003_103.n1 GND 0.04fF
C17 a_14003_103.n2 GND 0.03fF
C18 a_14003_103.n3 GND 0.07fF
C19 a_14003_103.n4 GND 0.08fF
C20 a_14003_103.n5 GND 0.03fF
C21 a_3643_103.n0 GND 0.08fF
C22 a_3643_103.n1 GND 0.07fF
C23 a_3643_103.n2 GND 0.04fF
C24 a_3643_103.n3 GND 0.06fF
C25 a_3643_103.n4 GND 0.03fF
C26 a_3643_103.n5 GND 0.04fF
C27 a_3643_103.n7 GND 0.08fF
C28 a_13041_103.n0 GND 0.11fF
C29 a_13041_103.n1 GND 0.04fF
C30 a_13041_103.n2 GND 0.03fF
C31 a_13041_103.n3 GND 0.07fF
C32 a_13041_103.n4 GND 0.08fF
C33 a_13041_103.n5 GND 0.03fF
C34 a_14284_210.n0 GND 0.02fF
C35 a_14284_210.n1 GND 0.09fF
C36 a_14284_210.n2 GND 0.12fF
C37 a_14284_210.n3 GND 0.08fF
C38 a_14284_210.n4 GND 0.08fF
C39 a_14284_210.n5 GND 0.02fF
C40 a_14284_210.t1 GND 0.29fF
C41 a_14284_210.n6 GND 0.09fF
C42 a_14284_210.n7 GND 0.02fF
C43 a_14284_210.n8 GND 0.13fF
C44 a_14284_210.n9 GND 0.02fF
C45 a_14284_210.n10 GND 0.03fF
C46 a_14284_210.n11 GND 0.03fF
C47 a_13322_210.n0 GND 0.07fF
C48 a_13322_210.n1 GND 0.09fF
C49 a_13322_210.n2 GND 0.12fF
C50 a_13322_210.n3 GND 0.08fF
C51 a_13322_210.n4 GND 0.02fF
C52 a_13322_210.n5 GND 0.03fF
C53 a_13322_210.n6 GND 0.02fF
C54 a_13322_210.n7 GND 0.03fF
C55 a_13322_210.n8 GND 0.02fF
C56 a_13322_210.n9 GND 0.13fF
C57 a_13322_210.n10 GND 0.08fF
C58 a_13322_210.n11 GND 0.02fF
C59 a_13322_210.t0 GND 0.31fF
C60 a_3924_210.n0 GND 0.02fF
C61 a_3924_210.n1 GND 0.09fF
C62 a_3924_210.n2 GND 0.12fF
C63 a_3924_210.n3 GND 0.08fF
C64 a_3924_210.n4 GND 0.08fF
C65 a_3924_210.n5 GND 0.02fF
C66 a_3924_210.t1 GND 0.29fF
C67 a_3924_210.n6 GND 0.09fF
C68 a_3924_210.n7 GND 0.02fF
C69 a_3924_210.n8 GND 0.13fF
C70 a_3924_210.n9 GND 0.02fF
C71 a_3924_210.n10 GND 0.03fF
C72 a_3924_210.n11 GND 0.03fF
C73 a_5271_103.n0 GND 0.08fF
C74 a_5271_103.n1 GND 0.07fF
C75 a_5271_103.n2 GND 0.04fF
C76 a_5271_103.n3 GND 0.06fF
C77 a_5271_103.n4 GND 0.03fF
C78 a_5271_103.n5 GND 0.04fF
C79 a_5271_103.n7 GND 0.08fF
C80 a_91_103.n0 GND 0.08fF
C81 a_91_103.n1 GND 0.07fF
C82 a_91_103.n2 GND 0.04fF
C83 a_91_103.n3 GND 0.06fF
C84 a_91_103.n4 GND 0.03fF
C85 a_91_103.n5 GND 0.03fF
C86 a_91_103.n7 GND 0.08fF
C87 a_7216_101.n0 GND 0.02fF
C88 a_7216_101.n1 GND 0.09fF
C89 a_7216_101.n2 GND 0.08fF
C90 a_7216_101.n3 GND 0.03fF
C91 a_7216_101.n4 GND 0.01fF
C92 a_7216_101.n5 GND 0.04fF
C93 a_7216_101.n6 GND 0.04fF
C94 a_7216_101.n7 GND 0.02fF
C95 a_7216_101.n8 GND 0.05fF
C96 a_7216_101.n9 GND 0.15fF
C97 a_7216_101.n10 GND 0.08fF
C98 a_7216_101.n11 GND 0.08fF
C99 a_7216_101.t1 GND 0.23fF
C100 a_7216_101.n12 GND 0.01fF
C101 a_9806_101.n0 GND 0.02fF
C102 a_9806_101.n1 GND 0.09fF
C103 a_9806_101.n2 GND 0.08fF
C104 a_9806_101.n3 GND 0.03fF
C105 a_9806_101.n4 GND 0.01fF
C106 a_9806_101.n5 GND 0.04fF
C107 a_9806_101.n6 GND 0.04fF
C108 a_9806_101.n7 GND 0.02fF
C109 a_9806_101.n8 GND 0.05fF
C110 a_9806_101.n9 GND 0.15fF
C111 a_9806_101.n10 GND 0.08fF
C112 a_9806_101.n11 GND 0.08fF
C113 a_9806_101.t1 GND 0.23fF
C114 a_9806_101.n12 GND 0.01fF
C115 a_7861_103.n0 GND 0.11fF
C116 a_7861_103.n1 GND 0.04fF
C117 a_7861_103.n2 GND 0.03fF
C118 a_7861_103.n3 GND 0.07fF
C119 a_7861_103.n4 GND 0.08fF
C120 a_7861_103.n5 GND 0.03fF
C121 a_2962_210.n0 GND 0.07fF
C122 a_2962_210.n1 GND 0.09fF
C123 a_2962_210.n2 GND 0.12fF
C124 a_2962_210.n3 GND 0.08fF
C125 a_2962_210.n4 GND 0.02fF
C126 a_2962_210.n5 GND 0.03fF
C127 a_2962_210.n6 GND 0.02fF
C128 a_2962_210.n7 GND 0.03fF
C129 a_2962_210.n8 GND 0.02fF
C130 a_2962_210.n9 GND 0.13fF
C131 a_2962_210.n10 GND 0.08fF
C132 a_2962_210.n11 GND 0.02fF
C133 a_2962_210.t0 GND 0.31fF
C134 a_16984_101.n0 GND 0.05fF
C135 a_16984_101.n1 GND 0.13fF
C136 a_16984_101.n2 GND 0.04fF
C137 a_16984_101.n3 GND 0.18fF
C138 a_5552_210.n0 GND 0.07fF
C139 a_5552_210.n1 GND 0.09fF
C140 a_5552_210.n2 GND 0.12fF
C141 a_5552_210.n3 GND 0.08fF
C142 a_5552_210.n4 GND 0.02fF
C143 a_5552_210.n5 GND 0.03fF
C144 a_5552_210.n6 GND 0.02fF
C145 a_5552_210.n7 GND 0.03fF
C146 a_5552_210.n8 GND 0.02fF
C147 a_5552_210.n9 GND 0.13fF
C148 a_5552_210.n10 GND 0.08fF
C149 a_5552_210.n11 GND 0.02fF
C150 a_5552_210.t0 GND 0.31fF
C151 a_6233_103.n0 GND 0.08fF
C152 a_6233_103.n1 GND 0.07fF
C153 a_6233_103.n2 GND 0.04fF
C154 a_6233_103.n3 GND 0.06fF
C155 a_6233_103.n4 GND 0.03fF
C156 a_6233_103.n5 GND 0.04fF
C157 a_6233_103.n7 GND 0.08fF
C158 a_10732_210.n0 GND 0.07fF
C159 a_10732_210.n1 GND 0.09fF
C160 a_10732_210.n2 GND 0.12fF
C161 a_10732_210.n3 GND 0.08fF
C162 a_10732_210.n4 GND 0.02fF
C163 a_10732_210.n5 GND 0.03fF
C164 a_10732_210.n6 GND 0.05fF
C165 a_10732_210.n7 GND 0.02fF
C166 a_10732_210.n8 GND 0.14fF
C167 a_10732_210.n9 GND 0.08fF
C168 a_10732_210.n10 GND 0.02fF
C169 a_10732_210.t0 GND 0.31fF
C170 a_372_210.n0 GND 0.07fF
C171 a_372_210.n1 GND 0.09fF
C172 a_372_210.n2 GND 0.12fF
C173 a_372_210.n3 GND 0.08fF
C174 a_372_210.n4 GND 0.02fF
C175 a_372_210.n5 GND 0.03fF
C176 a_372_210.n6 GND 0.02fF
C177 a_372_210.n7 GND 0.03fF
C178 a_372_210.n8 GND 0.02fF
C179 a_372_210.n9 GND 0.13fF
C180 a_372_210.n10 GND 0.08fF
C181 a_372_210.n11 GND 0.02fF
C182 a_372_210.t0 GND 0.31fF
C183 a_16318_101.n0 GND 0.13fF
C184 a_16318_101.n1 GND 0.14fF
C185 a_16318_101.n2 GND 0.14fF
C186 a_9104_210.n0 GND 0.02fF
C187 a_9104_210.n1 GND 0.09fF
C188 a_9104_210.n2 GND 0.12fF
C189 a_9104_210.n3 GND 0.08fF
C190 a_9104_210.n4 GND 0.08fF
C191 a_9104_210.n5 GND 0.02fF
C192 a_9104_210.t1 GND 0.29fF
C193 a_9104_210.n6 GND 0.09fF
C194 a_9104_210.n7 GND 0.02fF
C195 a_9104_210.n8 GND 0.13fF
C196 a_9104_210.n9 GND 0.02fF
C197 a_9104_210.n10 GND 0.03fF
C198 a_9104_210.n11 GND 0.02fF
C199 a_8823_103.n0 GND 0.08fF
C200 a_8823_103.n1 GND 0.07fF
C201 a_8823_103.n2 GND 0.04fF
C202 a_8823_103.n3 GND 0.06fF
C203 a_8823_103.n4 GND 0.11fF
C204 a_8823_103.n5 GND 0.04fF
C205 a_8823_103.n7 GND 0.08fF
C206 a_7321_1050.n0 GND 0.39fF
C207 a_7321_1050.n1 GND 0.33fF
C208 a_7321_1050.n2 GND 0.67fF
C209 a_7321_1050.n3 GND 0.04fF
C210 a_7321_1050.n4 GND 0.06fF
C211 a_7321_1050.n5 GND 0.03fF
C212 a_7321_1050.n6 GND 0.23fF
C213 a_7321_1050.n7 GND 0.69fF
C214 a_7321_1050.n8 GND 0.59fF
C215 a_7321_1050.n9 GND 0.51fF
C216 a_12501_1050.n0 GND 0.42fF
C217 a_12501_1050.n1 GND 0.36fF
C218 a_12501_1050.n2 GND 0.72fF
C219 a_12501_1050.n3 GND 0.37fF
C220 a_12501_1050.n4 GND 0.76fF
C221 a_12501_1050.n5 GND 0.64fF
C222 a_12501_1050.n6 GND 0.54fF
C223 a_14986_101.n0 GND 0.02fF
C224 a_14986_101.n1 GND 0.09fF
C225 a_14986_101.n2 GND 0.08fF
C226 a_14986_101.n3 GND 0.03fF
C227 a_14986_101.n4 GND 0.01fF
C228 a_14986_101.n5 GND 0.04fF
C229 a_14986_101.n6 GND 0.04fF
C230 a_14986_101.n7 GND 0.02fF
C231 a_14986_101.n8 GND 0.05fF
C232 a_14986_101.n9 GND 0.15fF
C233 a_14986_101.n10 GND 0.08fF
C234 a_14986_101.n11 GND 0.08fF
C235 a_14986_101.t1 GND 0.23fF
C236 a_14986_101.n12 GND 0.01fF
C237 a_11694_210.n0 GND 0.02fF
C238 a_11694_210.n1 GND 0.09fF
C239 a_11694_210.n2 GND 0.12fF
C240 a_11694_210.n3 GND 0.08fF
C241 a_11694_210.n4 GND 0.08fF
C242 a_11694_210.n5 GND 0.02fF
C243 a_11694_210.t1 GND 0.29fF
C244 a_11694_210.n6 GND 0.09fF
C245 a_11694_210.n7 GND 0.02fF
C246 a_11694_210.n8 GND 0.13fF
C247 a_11694_210.n9 GND 0.02fF
C248 a_11694_210.n10 GND 0.03fF
C249 a_11694_210.n11 GND 0.02fF
C250 a_6514_210.n0 GND 0.02fF
C251 a_6514_210.n1 GND 0.09fF
C252 a_6514_210.n2 GND 0.12fF
C253 a_6514_210.n3 GND 0.08fF
C254 a_6514_210.n4 GND 0.08fF
C255 a_6514_210.n5 GND 0.02fF
C256 a_6514_210.t1 GND 0.29fF
C257 a_6514_210.n6 GND 0.09fF
C258 a_6514_210.n7 GND 0.02fF
C259 a_6514_210.n8 GND 0.13fF
C260 a_6514_210.n9 GND 0.02fF
C261 a_6514_210.n10 GND 0.03fF
C262 a_6514_210.n11 GND 0.03fF
C263 a_15652_101.n0 GND 0.09fF
C264 a_15652_101.n1 GND 0.07fF
C265 a_15652_101.n2 GND 0.11fF
C266 a_15652_101.n3 GND 0.02fF
C267 a_15652_101.n4 GND 0.02fF
C268 a_15652_101.n5 GND 0.06fF
C269 a_15652_101.n6 GND 0.21fF
C270 a_15757_1051.n0 GND 0.43fF
C271 a_15757_1051.n1 GND 0.32fF
C272 a_15757_1051.n2 GND 0.52fF
C273 a_15757_1051.n3 GND 0.30fF
C274 a_15757_1051.n4 GND 0.80fF
C275 a_15757_1051.n5 GND 0.36fF
C276 a_10451_103.n0 GND 0.13fF
C277 a_10451_103.n1 GND 0.04fF
C278 a_10451_103.n2 GND 0.09fF
C279 a_10451_103.n3 GND 0.07fF
C280 a_10451_103.n4 GND 0.08fF
C281 a_10451_103.n5 GND 0.03fF
C282 a_2036_101.n0 GND 0.02fF
C283 a_2036_101.n1 GND 0.09fF
C284 a_2036_101.n2 GND 0.08fF
C285 a_2036_101.n3 GND 0.03fF
C286 a_2036_101.n4 GND 0.01fF
C287 a_2036_101.n5 GND 0.04fF
C288 a_2036_101.n6 GND 0.04fF
C289 a_2036_101.n7 GND 0.02fF
C290 a_2036_101.n8 GND 0.05fF
C291 a_2036_101.n9 GND 0.15fF
C292 a_2036_101.n10 GND 0.08fF
C293 a_2036_101.n11 GND 0.08fF
C294 a_2036_101.t1 GND 0.23fF
C295 a_2036_101.n12 GND 0.01fF
C296 a_3829_1050.n0 GND 0.35fF
C297 a_3829_1050.n1 GND 0.28fF
C298 a_3829_1050.n2 GND 0.55fF
C299 a_3829_1050.n3 GND 0.04fF
C300 a_3829_1050.n4 GND 0.05fF
C301 a_3829_1050.n5 GND 0.03fF
C302 a_3829_1050.n6 GND 0.23fF
C303 a_3829_1050.n7 GND 0.63fF
C304 a_3829_1050.n8 GND 0.38fF
C305 a_3829_1050.n9 GND 0.45fF
C306 a_3829_1050.n10 GND 0.43fF
C307 a_3829_1050.n11 GND 0.35fF
C308 a_12396_101.n0 GND 0.08fF
C309 a_12396_101.n1 GND 0.02fF
C310 a_12396_101.n2 GND 0.02fF
C311 a_12396_101.n3 GND 0.09fF
C312 a_12396_101.n4 GND 0.08fF
C313 a_12396_101.n5 GND 0.03fF
C314 a_12396_101.n6 GND 0.05fF
C315 a_5779_989.n0 GND 0.46fF
C316 a_5779_989.n1 GND 0.39fF
C317 a_5779_989.n2 GND 0.56fF
C318 a_5779_989.n3 GND 0.39fF
C319 a_5779_989.t7 GND 0.63fF
C320 a_5779_989.n4 GND 0.75fF
C321 a_5779_989.n5 GND 1.19fF
C322 a_5779_989.n6 GND 0.05fF
C323 a_5779_989.n7 GND 0.06fF
C324 a_5779_989.n8 GND 0.04fF
C325 a_5779_989.n9 GND 0.27fF
C326 a_5779_989.n10 GND 0.62fF
C327 a_5779_989.n11 GND 0.53fF
C328 a_5779_989.n12 GND 0.59fF
C329 a_5779_989.n13 GND 0.56fF
C330 a_5779_989.n14 GND 0.46fF
C331 a_5457_1050.n0 GND 0.60fF
C332 a_5457_1050.n1 GND 0.47fF
C333 a_5457_1050.n2 GND 1.86fF
C334 a_5457_1050.n3 GND 0.47fF
C335 a_5457_1050.n4 GND 0.74fF
C336 a_5457_1050.n5 GND 2.64fF
C337 a_5457_1050.n6 GND 0.57fF
C338 a_5457_1050.n7 GND 0.90fF
C339 a_5457_1050.n8 GND 0.65fF
C340 a_5457_1050.n9 GND 0.77fF
C341 a_5457_1050.n10 GND 0.73fF
C342 a_5457_1050.n11 GND 0.60fF
C343 a_277_1050.n0 GND 0.43fF
C344 a_277_1050.n1 GND 1.71fF
C345 a_277_1050.n2 GND 0.43fF
C346 a_277_1050.n3 GND 0.68fF
C347 a_277_1050.n4 GND 2.43fF
C348 a_277_1050.n5 GND 0.06fF
C349 a_277_1050.n6 GND 0.08fF
C350 a_277_1050.n7 GND 0.05fF
C351 a_277_1050.n8 GND 0.36fF
C352 a_277_1050.n9 GND 0.80fF
C353 a_277_1050.n10 GND 0.56fF
C354 a_277_1050.n11 GND 0.71fF
C355 a_277_1050.n12 GND 0.67fF
C356 a_277_1050.n13 GND 0.59fF
C357 a_277_1050.n14 GND 0.56fF
C358 a_1334_210.n0 GND 0.02fF
C359 a_1334_210.n1 GND 0.09fF
C360 a_1334_210.n2 GND 0.12fF
C361 a_1334_210.n3 GND 0.08fF
C362 a_1334_210.n4 GND 0.08fF
C363 a_1334_210.n5 GND 0.02fF
C364 a_1334_210.t1 GND 0.29fF
C365 a_1334_210.n6 GND 0.09fF
C366 a_1334_210.n7 GND 0.02fF
C367 a_1334_210.n8 GND 0.13fF
C368 a_1334_210.n9 GND 0.02fF
C369 a_1334_210.n10 GND 0.03fF
C370 a_1334_210.n11 GND 0.02fF
C371 a_1053_103.n0 GND 0.13fF
C372 a_1053_103.n1 GND 0.04fF
C373 a_1053_103.n2 GND 0.09fF
C374 a_1053_103.n3 GND 0.07fF
C375 a_1053_103.n4 GND 0.08fF
C376 a_1053_103.n5 GND 0.03fF
C377 a_4151_989.n0 GND 0.86fF
C378 a_4151_989.n1 GND 0.98fF
C379 a_4151_989.n2 GND 1.36fF
C380 a_4151_989.n3 GND 0.74fF
C381 a_4151_989.n4 GND 10.33fF
C382 a_4151_989.n5 GND 0.85fF
C383 a_4151_989.t9 GND 1.09fF
C384 a_4151_989.n6 GND 1.19fF
C385 a_4151_989.n7 GND 12.86fF
C386 a_4151_989.n8 GND 0.62fF
C387 a_4151_989.n9 GND 1.14fF
C388 a_4151_989.n10 GND 1.10fF
C389 a_4151_989.n11 GND 1.43fF
C390 a_4151_989.n12 GND 0.86fF
C391 a_4626_101.n0 GND 0.08fF
C392 a_4626_101.n1 GND 0.02fF
C393 a_4626_101.n2 GND 0.02fF
C394 a_4626_101.n3 GND 0.09fF
C395 a_4626_101.n4 GND 0.08fF
C396 a_4626_101.n5 GND 0.03fF
C397 a_4626_101.n6 GND 0.05fF
C398 a_147_187.n0 GND 0.46fF
C399 a_147_187.t7 GND 0.95fF
C400 a_147_187.n1 GND 1.20fF
C401 a_147_187.n2 GND 0.46fF
C402 a_147_187.t8 GND 0.95fF
C403 a_147_187.n3 GND 0.64fF
C404 a_147_187.n4 GND 0.47fF
C405 a_147_187.n5 GND 1.67fF
C406 a_147_187.n6 GND 2.70fF
C407 a_147_187.n7 GND 2.24fF
C408 a_147_187.n8 GND 0.07fF
C409 a_147_187.n9 GND 0.09fF
C410 a_147_187.n10 GND 0.06fF
C411 a_147_187.n11 GND 0.47fF
C412 a_147_187.n12 GND 0.87fF
C413 a_147_187.n13 GND 0.65fF
C414 a_147_187.n14 GND 0.82fF
C415 a_147_187.n15 GND 0.78fF
C416 a_147_187.n16 GND 0.64fF
C417 a_147_187.n17 GND 0.65fF
C418 a_9331_989.n0 GND 0.76fF
C419 a_9331_989.n1 GND 0.49fF
C420 a_9331_989.n2 GND 1.52fF
C421 a_9331_989.n3 GND 0.48fF
C422 a_9331_989.n4 GND 1.10fF
C423 a_9331_989.n5 GND 4.30fF
C424 a_9331_989.n6 GND 0.70fF
C425 a_9331_989.t13 GND 1.00fF
C426 a_9331_989.n7 GND 1.08fF
C427 a_9331_989.n8 GND 6.33fF
C428 a_9331_989.n9 GND 0.08fF
C429 a_9331_989.n10 GND 0.11fF
C430 a_9331_989.n11 GND 0.07fF
C431 a_9331_989.n12 GND 0.38fF
C432 a_9331_989.n13 GND 0.98fF
C433 a_9331_989.n14 GND 1.20fF
C434 a_9331_989.n15 GND 0.97fF
C435 a_9009_1050.n0 GND 0.37fF
C436 a_9009_1050.n1 GND 0.29fF
C437 a_9009_1050.n2 GND 0.58fF
C438 a_9009_1050.n3 GND 0.35fF
C439 a_9009_1050.n4 GND 0.68fF
C440 a_9009_1050.n5 GND 0.40fF
C441 a_9009_1050.n6 GND 0.47fF
C442 a_9009_1050.n7 GND 0.45fF
C443 a_9009_1050.n8 GND 0.37fF
C444 a_2141_1050.n0 GND 0.38fF
C445 a_2141_1050.n1 GND 0.32fF
C446 a_2141_1050.n2 GND 0.64fF
C447 a_2141_1050.n3 GND 0.33fF
C448 a_2141_1050.n4 GND 0.68fF
C449 a_2141_1050.n5 GND 0.57fF
C450 a_2141_1050.n6 GND 0.48fF
C451 a_5327_187.n0 GND 0.49fF
C452 a_5327_187.t11 GND 1.03fF
C453 a_5327_187.n1 GND 1.30fF
C454 a_5327_187.n2 GND 0.49fF
C455 a_5327_187.t14 GND 1.03fF
C456 a_5327_187.n3 GND 0.69fF
C457 a_5327_187.n4 GND 0.51fF
C458 a_5327_187.n5 GND 1.81fF
C459 a_5327_187.n6 GND 2.92fF
C460 a_5327_187.n7 GND 2.42fF
C461 a_5327_187.n8 GND 0.08fF
C462 a_5327_187.n9 GND 0.10fF
C463 a_5327_187.n10 GND 0.54fF
C464 a_5327_187.n11 GND 0.96fF
C465 a_5327_187.n12 GND 0.70fF
C466 a_5327_187.n13 GND 0.89fF
C467 a_5327_187.n14 GND 0.84fF
C468 a_5327_187.n15 GND 0.69fF
C469 a_5327_187.n16 GND 0.70fF
C470 a_8142_210.n0 GND 0.02fF
C471 a_8142_210.n1 GND 0.09fF
C472 a_8142_210.t1 GND 0.23fF
C473 a_8142_210.n2 GND 0.10fF
C474 a_8142_210.n3 GND 0.07fF
C475 a_8142_210.n4 GND 0.04fF
C476 a_8142_210.n5 GND 0.08fF
C477 a_8142_210.n6 GND 0.09fF
C478 a_8142_210.n7 GND 0.04fF
C479 a_8142_210.n8 GND 0.02fF
C480 a_8142_210.n9 GND 0.01fF
C481 a_8142_210.n10 GND 0.13fF
C482 a_8142_210.n11 GND 0.02fF
C483 a_8142_210.n12 GND 0.03fF
C484 a_8142_210.n13 GND 0.02fF
C485 a_16421_1051.n0 GND 0.28fF
C486 a_16421_1051.n1 GND 0.28fF
C487 a_16421_1051.n2 GND 0.36fF
C488 a_16421_1051.n3 GND 0.69fF
C489 a_16421_1051.n4 GND 0.27fF
C490 a_16421_1051.n5 GND 0.45fF
C491 QN.n0 GND 0.30fF
C492 QN.n1 GND 0.38fF
C493 QN.n2 GND 0.46fF
C494 QN.n3 GND 0.04fF
C495 QN.n4 GND 0.05fF
C496 QN.n5 GND 0.06fF
C497 QN.n6 GND 0.04fF
C498 QN.n7 GND 0.05fF
C499 QN.n8 GND 0.03fF
C500 QN.n9 GND 0.04fF
C501 QN.n10 GND 1.07fF
C502 QN.n11 GND 0.06fF
C503 QN.n12 GND 0.03fF
C504 QN.n13 GND 0.06fF
C505 QN.n14 GND 0.37fF
C506 QN.n15 GND 0.35fF
C507 QN.n16 GND 0.01fF
C508 a_14511_989.n0 GND 0.41fF
C509 a_14511_989.n1 GND 0.29fF
C510 a_14511_989.n2 GND 0.31fF
C511 a_14511_989.n3 GND 1.06fF
C512 a_14511_989.n4 GND 0.73fF
C513 a_14511_989.n5 GND 0.41fF
C514 a_14511_989.n6 GND 0.35fF
C515 a_14511_989.t12 GND 0.56fF
C516 a_14511_989.n7 GND 0.59fF
C517 a_14511_989.n8 GND 1.00fF
C518 a_14511_989.n9 GND 0.04fF
C519 a_14511_989.n10 GND 0.06fF
C520 a_14511_989.n11 GND 0.04fF
C521 a_14511_989.n12 GND 0.24fF
C522 a_14511_989.n13 GND 0.53fF
C523 a_14511_989.n14 GND 0.62fF
C524 a_14511_989.n15 GND 0.53fF
C525 a_11413_103.n0 GND 0.03fF
C526 a_11413_103.n1 GND 0.09fF
C527 a_11413_103.n2 GND 0.08fF
C528 a_11413_103.n3 GND 0.04fF
C529 a_11413_103.n4 GND 0.05fF
C530 a_11413_103.n5 GND 0.11fF
C531 a_11413_103.n6 GND 0.04fF
C532 a_11413_103.n8 GND 0.08fF
C533 a_599_989.n0 GND 0.41fF
C534 a_599_989.n1 GND 0.34fF
C535 a_599_989.n2 GND 0.49fF
C536 a_599_989.n3 GND 0.34fF
C537 a_599_989.t9 GND 0.56fF
C538 a_599_989.n4 GND 0.66fF
C539 a_599_989.n5 GND 1.06fF
C540 a_599_989.n6 GND 0.04fF
C541 a_599_989.n7 GND 0.06fF
C542 a_599_989.n8 GND 0.04fF
C543 a_599_989.n9 GND 0.24fF
C544 a_599_989.n10 GND 0.55fF
C545 a_599_989.n11 GND 0.47fF
C546 a_599_989.n12 GND 0.52fF
C547 a_599_989.n13 GND 0.49fF
C548 a_599_989.n14 GND 0.41fF
C549 a_10959_989.n0 GND 0.54fF
C550 a_10959_989.n1 GND 0.54fF
C551 a_10959_989.n2 GND 0.45fF
C552 a_10959_989.n3 GND 0.65fF
C553 a_10959_989.n4 GND 0.45fF
C554 a_10959_989.t11 GND 0.73fF
C555 a_10959_989.n5 GND 0.87fF
C556 a_10959_989.n6 GND 1.38fF
C557 a_10959_989.n7 GND 0.06fF
C558 a_10959_989.n8 GND 0.07fF
C559 a_10959_989.n9 GND 0.05fF
C560 a_10959_989.n10 GND 0.31fF
C561 a_10959_989.n11 GND 0.72fF
C562 a_10959_989.n12 GND 0.62fF
C563 a_10959_989.n13 GND 0.65fF
C564 a_10959_989.n14 GND 0.68fF
C565 a_14189_1050.n0 GND 0.37fF
C566 a_14189_1050.n1 GND 0.37fF
C567 a_14189_1050.n2 GND 0.29fF
C568 a_14189_1050.n3 GND 0.58fF
C569 a_14189_1050.n4 GND 0.35fF
C570 a_14189_1050.n5 GND 0.68fF
C571 a_14189_1050.n6 GND 0.39fF
C572 a_14189_1050.n7 GND 0.44fF
C573 a_14189_1050.n8 GND 0.47fF
C574 a_10637_1050.n0 GND 0.63fF
C575 a_10637_1050.n1 GND 0.63fF
C576 a_10637_1050.n2 GND 0.49fF
C577 a_10637_1050.n3 GND 1.93fF
C578 a_10637_1050.n4 GND 0.49fF
C579 a_10637_1050.n5 GND 0.77fF
C580 a_10637_1050.n6 GND 2.74fF
C581 a_10637_1050.n7 GND 0.59fF
C582 a_10637_1050.n8 GND 0.93fF
C583 a_10637_1050.n9 GND 0.67fF
C584 a_10637_1050.n10 GND 0.75fF
C585 a_10637_1050.n11 GND 0.80fF
C586 VDD.n1 GND 0.03fF
C587 VDD.n2 GND 0.14fF
C588 VDD.n3 GND 0.03fF
C589 VDD.n4 GND 0.02fF
C590 VDD.n5 GND 0.06fF
C591 VDD.n6 GND 0.02fF
C592 VDD.n7 GND 0.02fF
C593 VDD.n8 GND 0.02fF
C594 VDD.n9 GND 0.02fF
C595 VDD.n10 GND 0.02fF
C596 VDD.n11 GND 0.02fF
C597 VDD.n12 GND 0.02fF
C598 VDD.n13 GND 0.02fF
C599 VDD.n14 GND 0.04fF
C600 VDD.n15 GND 0.01fF
C601 VDD.n20 GND 0.48fF
C602 VDD.n21 GND 0.29fF
C603 VDD.n22 GND 0.02fF
C604 VDD.n23 GND 0.04fF
C605 VDD.n24 GND 0.26fF
C606 VDD.n25 GND 0.01fF
C607 VDD.n26 GND 0.02fF
C608 VDD.n27 GND 0.01fF
C609 VDD.n28 GND 0.18fF
C610 VDD.n29 GND 0.01fF
C611 VDD.n30 GND 0.02fF
C612 VDD.n31 GND 0.08fF
C613 VDD.n32 GND 0.01fF
C614 VDD.n33 GND 0.03fF
C615 VDD.n34 GND 0.03fF
C616 VDD.n35 GND 0.15fF
C617 VDD.n36 GND 0.01fF
C618 VDD.n37 GND 0.03fF
C619 VDD.n38 GND 0.03fF
C620 VDD.n39 GND 0.17fF
C621 VDD.n40 GND 0.01fF
C622 VDD.n41 GND 0.02fF
C623 VDD.n42 GND 0.02fF
C624 VDD.n43 GND 0.26fF
C625 VDD.n44 GND 0.01fF
C626 VDD.n45 GND 0.02fF
C627 VDD.n46 GND 0.02fF
C628 VDD.n47 GND 0.29fF
C629 VDD.n48 GND 0.01fF
C630 VDD.n49 GND 0.02fF
C631 VDD.n50 GND 0.04fF
C632 VDD.n51 GND 0.06fF
C633 VDD.n52 GND 0.02fF
C634 VDD.n53 GND 0.02fF
C635 VDD.n54 GND 0.02fF
C636 VDD.n55 GND 0.02fF
C637 VDD.n56 GND 0.02fF
C638 VDD.n57 GND 0.02fF
C639 VDD.n58 GND 0.02fF
C640 VDD.n59 GND 0.02fF
C641 VDD.n60 GND 0.02fF
C642 VDD.n61 GND 0.02fF
C643 VDD.n62 GND 0.02fF
C644 VDD.n63 GND 0.03fF
C645 VDD.n64 GND 0.02fF
C646 VDD.n65 GND 0.23fF
C647 VDD.n66 GND 0.02fF
C648 VDD.n67 GND 0.02fF
C649 VDD.n69 GND 0.02fF
C650 VDD.n73 GND 0.29fF
C651 VDD.n74 GND 0.29fF
C652 VDD.n75 GND 0.01fF
C653 VDD.n76 GND 0.02fF
C654 VDD.n77 GND 0.04fF
C655 VDD.n78 GND 0.26fF
C656 VDD.n79 GND 0.01fF
C657 VDD.n80 GND 0.02fF
C658 VDD.n81 GND 0.02fF
C659 VDD.n82 GND 0.17fF
C660 VDD.n83 GND 0.01fF
C661 VDD.n84 GND 0.02fF
C662 VDD.n85 GND 0.02fF
C663 VDD.n86 GND 0.15fF
C664 VDD.n87 GND 0.01fF
C665 VDD.n88 GND 0.03fF
C666 VDD.n89 GND 0.03fF
C667 VDD.n90 GND 0.01fF
C668 VDD.n91 GND 0.03fF
C669 VDD.n92 GND 0.03fF
C670 VDD.n93 GND 0.18fF
C671 VDD.n94 GND 0.01fF
C672 VDD.n95 GND 0.02fF
C673 VDD.n96 GND 0.02fF
C674 VDD.n97 GND 0.26fF
C675 VDD.n98 GND 0.01fF
C676 VDD.n99 GND 0.02fF
C677 VDD.n100 GND 0.02fF
C678 VDD.n101 GND 0.29fF
C679 VDD.n102 GND 0.01fF
C680 VDD.n103 GND 0.02fF
C681 VDD.n104 GND 0.04fF
C682 VDD.n105 GND 0.23fF
C683 VDD.n106 GND 0.02fF
C684 VDD.n107 GND 0.02fF
C685 VDD.n108 GND 0.02fF
C686 VDD.n109 GND 0.06fF
C687 VDD.n110 GND 0.02fF
C688 VDD.n111 GND 0.02fF
C689 VDD.n112 GND 0.02fF
C690 VDD.n113 GND 0.02fF
C691 VDD.n114 GND 0.02fF
C692 VDD.n115 GND 0.02fF
C693 VDD.n116 GND 0.02fF
C694 VDD.n117 GND 0.02fF
C695 VDD.n118 GND 0.02fF
C696 VDD.n119 GND 0.02fF
C697 VDD.n120 GND 0.03fF
C698 VDD.n121 GND 0.02fF
C699 VDD.n122 GND 0.02fF
C700 VDD.n126 GND 0.29fF
C701 VDD.n127 GND 0.29fF
C702 VDD.n128 GND 0.01fF
C703 VDD.n129 GND 0.02fF
C704 VDD.n130 GND 0.04fF
C705 VDD.n131 GND 0.07fF
C706 VDD.n132 GND 0.26fF
C707 VDD.n133 GND 0.01fF
C708 VDD.n134 GND 0.01fF
C709 VDD.n135 GND 0.02fF
C710 VDD.n136 GND 0.18fF
C711 VDD.n137 GND 0.01fF
C712 VDD.n138 GND 0.02fF
C713 VDD.n139 GND 0.02fF
C714 VDD.n140 GND 0.09fF
C715 VDD.n141 GND 0.05fF
C716 VDD.n142 GND 0.01fF
C717 VDD.n143 GND 0.02fF
C718 VDD.n144 GND 0.03fF
C719 VDD.n145 GND 0.15fF
C720 VDD.n146 GND 0.01fF
C721 VDD.n147 GND 0.02fF
C722 VDD.n148 GND 0.03fF
C723 VDD.n149 GND 0.17fF
C724 VDD.n150 GND 0.01fF
C725 VDD.n151 GND 0.02fF
C726 VDD.n152 GND 0.02fF
C727 VDD.n153 GND 0.07fF
C728 VDD.n154 GND 0.26fF
C729 VDD.n155 GND 0.01fF
C730 VDD.n156 GND 0.01fF
C731 VDD.n157 GND 0.02fF
C732 VDD.n158 GND 0.29fF
C733 VDD.n159 GND 0.01fF
C734 VDD.n160 GND 0.02fF
C735 VDD.n161 GND 0.04fF
C736 VDD.n162 GND 0.23fF
C737 VDD.n163 GND 0.02fF
C738 VDD.n164 GND 0.02fF
C739 VDD.n165 GND 0.02fF
C740 VDD.n166 GND 0.06fF
C741 VDD.n167 GND 0.02fF
C742 VDD.n168 GND 0.02fF
C743 VDD.n169 GND 0.02fF
C744 VDD.n170 GND 0.02fF
C745 VDD.n171 GND 0.02fF
C746 VDD.n172 GND 0.02fF
C747 VDD.n173 GND 0.02fF
C748 VDD.n174 GND 0.02fF
C749 VDD.n175 GND 0.02fF
C750 VDD.n176 GND 0.02fF
C751 VDD.n177 GND 0.03fF
C752 VDD.n178 GND 0.02fF
C753 VDD.n179 GND 0.02fF
C754 VDD.n183 GND 0.29fF
C755 VDD.n184 GND 0.29fF
C756 VDD.n185 GND 0.01fF
C757 VDD.n186 GND 0.02fF
C758 VDD.n187 GND 0.04fF
C759 VDD.n188 GND 0.06fF
C760 VDD.n189 GND 0.26fF
C761 VDD.n190 GND 0.01fF
C762 VDD.n191 GND 0.01fF
C763 VDD.n192 GND 0.02fF
C764 VDD.n193 GND 0.18fF
C765 VDD.n194 GND 0.01fF
C766 VDD.n195 GND 0.02fF
C767 VDD.n196 GND 0.02fF
C768 VDD.n197 GND 0.09fF
C769 VDD.n198 GND 0.05fF
C770 VDD.n199 GND 0.01fF
C771 VDD.n200 GND 0.02fF
C772 VDD.n201 GND 0.03fF
C773 VDD.n202 GND 0.15fF
C774 VDD.n203 GND 0.01fF
C775 VDD.n204 GND 0.02fF
C776 VDD.n205 GND 0.03fF
C777 VDD.n206 GND 0.17fF
C778 VDD.n207 GND 0.01fF
C779 VDD.n208 GND 0.02fF
C780 VDD.n209 GND 0.02fF
C781 VDD.n210 GND 0.07fF
C782 VDD.n211 GND 0.26fF
C783 VDD.n212 GND 0.01fF
C784 VDD.n213 GND 0.01fF
C785 VDD.n214 GND 0.02fF
C786 VDD.n215 GND 0.29fF
C787 VDD.n216 GND 0.01fF
C788 VDD.n217 GND 0.02fF
C789 VDD.n218 GND 0.04fF
C790 VDD.n219 GND 0.28fF
C791 VDD.n220 GND 0.02fF
C792 VDD.n221 GND 0.02fF
C793 VDD.n222 GND 0.02fF
C794 VDD.n223 GND 0.06fF
C795 VDD.n224 GND 0.02fF
C796 VDD.n225 GND 0.02fF
C797 VDD.n226 GND 0.02fF
C798 VDD.n227 GND 0.02fF
C799 VDD.n228 GND 0.02fF
C800 VDD.n229 GND 0.02fF
C801 VDD.n230 GND 0.02fF
C802 VDD.n231 GND 0.02fF
C803 VDD.n232 GND 0.02fF
C804 VDD.n233 GND 0.02fF
C805 VDD.n234 GND 0.03fF
C806 VDD.n235 GND 0.02fF
C807 VDD.n236 GND 0.02fF
C808 VDD.n240 GND 0.29fF
C809 VDD.n241 GND 0.29fF
C810 VDD.n242 GND 0.01fF
C811 VDD.n243 GND 0.02fF
C812 VDD.n244 GND 0.04fF
C813 VDD.n245 GND 0.29fF
C814 VDD.n246 GND 0.01fF
C815 VDD.n247 GND 0.02fF
C816 VDD.n248 GND 0.02fF
C817 VDD.n249 GND 0.23fF
C818 VDD.n250 GND 0.01fF
C819 VDD.n251 GND 0.07fF
C820 VDD.n252 GND 0.02fF
C821 VDD.n253 GND 0.18fF
C822 VDD.n254 GND 0.01fF
C823 VDD.n255 GND 0.02fF
C824 VDD.n256 GND 0.02fF
C825 VDD.n257 GND 0.17fF
C826 VDD.n258 GND 0.01fF
C827 VDD.n259 GND 0.09fF
C828 VDD.n260 GND 0.05fF
C829 VDD.n261 GND 0.02fF
C830 VDD.n262 GND 0.02fF
C831 VDD.n263 GND 0.15fF
C832 VDD.n264 GND 0.02fF
C833 VDD.n265 GND 0.02fF
C834 VDD.n266 GND 0.03fF
C835 VDD.n267 GND 0.16fF
C836 VDD.n268 GND 0.02fF
C837 VDD.n269 GND 0.02fF
C838 VDD.n270 GND 0.03fF
C839 VDD.n271 GND 0.09fF
C840 VDD.n272 GND 0.05fF
C841 VDD.n273 GND 0.16fF
C842 VDD.n274 GND 0.01fF
C843 VDD.n275 GND 0.02fF
C844 VDD.n276 GND 0.02fF
C845 VDD.n277 GND 0.18fF
C846 VDD.n278 GND 0.01fF
C847 VDD.n279 GND 0.02fF
C848 VDD.n280 GND 0.02fF
C849 VDD.n281 GND 0.07fF
C850 VDD.n282 GND 0.24fF
C851 VDD.n283 GND 0.01fF
C852 VDD.n284 GND 0.01fF
C853 VDD.n285 GND 0.02fF
C854 VDD.n286 GND 0.29fF
C855 VDD.n287 GND 0.01fF
C856 VDD.n288 GND 0.02fF
C857 VDD.n289 GND 0.02fF
C858 VDD.n290 GND 0.29fF
C859 VDD.n291 GND 0.01fF
C860 VDD.n292 GND 0.02fF
C861 VDD.n293 GND 0.04fF
C862 VDD.n294 GND 0.33fF
C863 VDD.n295 GND 0.02fF
C864 VDD.n296 GND 0.02fF
C865 VDD.n297 GND 0.02fF
C866 VDD.n298 GND 0.06fF
C867 VDD.n299 GND 0.02fF
C868 VDD.n300 GND 0.02fF
C869 VDD.n301 GND 0.02fF
C870 VDD.n302 GND 0.02fF
C871 VDD.n303 GND 0.02fF
C872 VDD.n304 GND 0.02fF
C873 VDD.n305 GND 0.02fF
C874 VDD.n306 GND 0.02fF
C875 VDD.n307 GND 0.02fF
C876 VDD.n308 GND 0.02fF
C877 VDD.n309 GND 0.03fF
C878 VDD.n310 GND 0.02fF
C879 VDD.n311 GND 0.02fF
C880 VDD.n315 GND 0.29fF
C881 VDD.n316 GND 0.29fF
C882 VDD.n317 GND 0.01fF
C883 VDD.n318 GND 0.02fF
C884 VDD.n319 GND 0.04fF
C885 VDD.n320 GND 0.29fF
C886 VDD.n321 GND 0.01fF
C887 VDD.n322 GND 0.02fF
C888 VDD.n323 GND 0.02fF
C889 VDD.n324 GND 0.23fF
C890 VDD.n325 GND 0.01fF
C891 VDD.n326 GND 0.07fF
C892 VDD.n327 GND 0.02fF
C893 VDD.n328 GND 0.18fF
C894 VDD.n329 GND 0.01fF
C895 VDD.n330 GND 0.02fF
C896 VDD.n331 GND 0.02fF
C897 VDD.n332 GND 0.17fF
C898 VDD.n333 GND 0.01fF
C899 VDD.n334 GND 0.09fF
C900 VDD.n335 GND 0.05fF
C901 VDD.n336 GND 0.02fF
C902 VDD.n337 GND 0.02fF
C903 VDD.n338 GND 0.15fF
C904 VDD.n339 GND 0.02fF
C905 VDD.n340 GND 0.02fF
C906 VDD.n341 GND 0.03fF
C907 VDD.n342 GND 0.16fF
C908 VDD.n343 GND 0.02fF
C909 VDD.n344 GND 0.02fF
C910 VDD.n345 GND 0.03fF
C911 VDD.n346 GND 0.09fF
C912 VDD.n347 GND 0.05fF
C913 VDD.n348 GND 0.16fF
C914 VDD.n349 GND 0.01fF
C915 VDD.n350 GND 0.02fF
C916 VDD.n351 GND 0.02fF
C917 VDD.n352 GND 0.18fF
C918 VDD.n353 GND 0.01fF
C919 VDD.n354 GND 0.02fF
C920 VDD.n355 GND 0.02fF
C921 VDD.n356 GND 0.07fF
C922 VDD.n357 GND 0.24fF
C923 VDD.n358 GND 0.01fF
C924 VDD.n359 GND 0.01fF
C925 VDD.n360 GND 0.02fF
C926 VDD.n361 GND 0.29fF
C927 VDD.n362 GND 0.01fF
C928 VDD.n363 GND 0.02fF
C929 VDD.n364 GND 0.02fF
C930 VDD.n365 GND 0.29fF
C931 VDD.n366 GND 0.01fF
C932 VDD.n367 GND 0.02fF
C933 VDD.n368 GND 0.04fF
C934 VDD.n369 GND 0.28fF
C935 VDD.n370 GND 0.02fF
C936 VDD.n371 GND 0.02fF
C937 VDD.n372 GND 0.02fF
C938 VDD.n373 GND 0.06fF
C939 VDD.n374 GND 0.02fF
C940 VDD.n375 GND 0.02fF
C941 VDD.n376 GND 0.02fF
C942 VDD.n377 GND 0.02fF
C943 VDD.n378 GND 0.02fF
C944 VDD.n379 GND 0.02fF
C945 VDD.n380 GND 0.02fF
C946 VDD.n381 GND 0.02fF
C947 VDD.n382 GND 0.02fF
C948 VDD.n383 GND 0.02fF
C949 VDD.n384 GND 0.03fF
C950 VDD.n385 GND 0.02fF
C951 VDD.n386 GND 0.02fF
C952 VDD.n390 GND 0.29fF
C953 VDD.n391 GND 0.29fF
C954 VDD.n392 GND 0.01fF
C955 VDD.n393 GND 0.02fF
C956 VDD.n394 GND 0.04fF
C957 VDD.n395 GND 0.06fF
C958 VDD.n396 GND 0.26fF
C959 VDD.n397 GND 0.01fF
C960 VDD.n398 GND 0.01fF
C961 VDD.n399 GND 0.02fF
C962 VDD.n400 GND 0.18fF
C963 VDD.n401 GND 0.01fF
C964 VDD.n402 GND 0.02fF
C965 VDD.n403 GND 0.02fF
C966 VDD.n404 GND 0.09fF
C967 VDD.n405 GND 0.05fF
C968 VDD.n406 GND 0.01fF
C969 VDD.n407 GND 0.02fF
C970 VDD.n408 GND 0.03fF
C971 VDD.n409 GND 0.15fF
C972 VDD.n410 GND 0.01fF
C973 VDD.n411 GND 0.02fF
C974 VDD.n412 GND 0.03fF
C975 VDD.n413 GND 0.17fF
C976 VDD.n414 GND 0.01fF
C977 VDD.n415 GND 0.02fF
C978 VDD.n416 GND 0.02fF
C979 VDD.n417 GND 0.07fF
C980 VDD.n418 GND 0.26fF
C981 VDD.n419 GND 0.01fF
C982 VDD.n420 GND 0.01fF
C983 VDD.n421 GND 0.02fF
C984 VDD.n422 GND 0.29fF
C985 VDD.n423 GND 0.01fF
C986 VDD.n424 GND 0.02fF
C987 VDD.n425 GND 0.04fF
C988 VDD.n426 GND 0.28fF
C989 VDD.n427 GND 0.02fF
C990 VDD.n428 GND 0.02fF
C991 VDD.n429 GND 0.02fF
C992 VDD.n430 GND 0.06fF
C993 VDD.n431 GND 0.02fF
C994 VDD.n432 GND 0.02fF
C995 VDD.n433 GND 0.02fF
C996 VDD.n434 GND 0.02fF
C997 VDD.n435 GND 0.02fF
C998 VDD.n436 GND 0.02fF
C999 VDD.n437 GND 0.02fF
C1000 VDD.n438 GND 0.02fF
C1001 VDD.n439 GND 0.02fF
C1002 VDD.n440 GND 0.02fF
C1003 VDD.n441 GND 0.03fF
C1004 VDD.n442 GND 0.02fF
C1005 VDD.n443 GND 0.02fF
C1006 VDD.n447 GND 0.29fF
C1007 VDD.n448 GND 0.29fF
C1008 VDD.n449 GND 0.01fF
C1009 VDD.n450 GND 0.02fF
C1010 VDD.n451 GND 0.04fF
C1011 VDD.n452 GND 0.29fF
C1012 VDD.n453 GND 0.01fF
C1013 VDD.n454 GND 0.02fF
C1014 VDD.n455 GND 0.02fF
C1015 VDD.n456 GND 0.23fF
C1016 VDD.n457 GND 0.01fF
C1017 VDD.n458 GND 0.07fF
C1018 VDD.n459 GND 0.02fF
C1019 VDD.n460 GND 0.18fF
C1020 VDD.n461 GND 0.01fF
C1021 VDD.n462 GND 0.02fF
C1022 VDD.n463 GND 0.02fF
C1023 VDD.n464 GND 0.17fF
C1024 VDD.n465 GND 0.01fF
C1025 VDD.n466 GND 0.09fF
C1026 VDD.n467 GND 0.05fF
C1027 VDD.n468 GND 0.02fF
C1028 VDD.n469 GND 0.02fF
C1029 VDD.n470 GND 0.15fF
C1030 VDD.n471 GND 0.02fF
C1031 VDD.n472 GND 0.02fF
C1032 VDD.n473 GND 0.03fF
C1033 VDD.n474 GND 0.16fF
C1034 VDD.n475 GND 0.02fF
C1035 VDD.n476 GND 0.02fF
C1036 VDD.n477 GND 0.03fF
C1037 VDD.n478 GND 0.09fF
C1038 VDD.n479 GND 0.05fF
C1039 VDD.n480 GND 0.16fF
C1040 VDD.n481 GND 0.01fF
C1041 VDD.n482 GND 0.02fF
C1042 VDD.n483 GND 0.02fF
C1043 VDD.n484 GND 0.18fF
C1044 VDD.n485 GND 0.01fF
C1045 VDD.n486 GND 0.02fF
C1046 VDD.n487 GND 0.02fF
C1047 VDD.n488 GND 0.07fF
C1048 VDD.n489 GND 0.24fF
C1049 VDD.n490 GND 0.01fF
C1050 VDD.n491 GND 0.01fF
C1051 VDD.n492 GND 0.02fF
C1052 VDD.n493 GND 0.29fF
C1053 VDD.n494 GND 0.01fF
C1054 VDD.n495 GND 0.02fF
C1055 VDD.n496 GND 0.02fF
C1056 VDD.n497 GND 0.29fF
C1057 VDD.n498 GND 0.01fF
C1058 VDD.n499 GND 0.02fF
C1059 VDD.n500 GND 0.04fF
C1060 VDD.n501 GND 0.33fF
C1061 VDD.n502 GND 0.02fF
C1062 VDD.n503 GND 0.02fF
C1063 VDD.n504 GND 0.02fF
C1064 VDD.n505 GND 0.06fF
C1065 VDD.n506 GND 0.02fF
C1066 VDD.n507 GND 0.02fF
C1067 VDD.n508 GND 0.02fF
C1068 VDD.n509 GND 0.02fF
C1069 VDD.n510 GND 0.02fF
C1070 VDD.n511 GND 0.02fF
C1071 VDD.n512 GND 0.02fF
C1072 VDD.n513 GND 0.02fF
C1073 VDD.n514 GND 0.02fF
C1074 VDD.n515 GND 0.02fF
C1075 VDD.n516 GND 0.03fF
C1076 VDD.n517 GND 0.02fF
C1077 VDD.n518 GND 0.02fF
C1078 VDD.n522 GND 0.29fF
C1079 VDD.n523 GND 0.29fF
C1080 VDD.n524 GND 0.01fF
C1081 VDD.n525 GND 0.02fF
C1082 VDD.n526 GND 0.04fF
C1083 VDD.n527 GND 0.29fF
C1084 VDD.n528 GND 0.01fF
C1085 VDD.n529 GND 0.02fF
C1086 VDD.n530 GND 0.02fF
C1087 VDD.n531 GND 0.23fF
C1088 VDD.n532 GND 0.01fF
C1089 VDD.n533 GND 0.07fF
C1090 VDD.n534 GND 0.02fF
C1091 VDD.n535 GND 0.18fF
C1092 VDD.n536 GND 0.01fF
C1093 VDD.n537 GND 0.02fF
C1094 VDD.n538 GND 0.02fF
C1095 VDD.n539 GND 0.17fF
C1096 VDD.n540 GND 0.01fF
C1097 VDD.n541 GND 0.09fF
C1098 VDD.n542 GND 0.05fF
C1099 VDD.n543 GND 0.02fF
C1100 VDD.n544 GND 0.02fF
C1101 VDD.n545 GND 0.15fF
C1102 VDD.n546 GND 0.02fF
C1103 VDD.n547 GND 0.02fF
C1104 VDD.n548 GND 0.03fF
C1105 VDD.n549 GND 0.16fF
C1106 VDD.n550 GND 0.02fF
C1107 VDD.n551 GND 0.02fF
C1108 VDD.n552 GND 0.03fF
C1109 VDD.n553 GND 0.09fF
C1110 VDD.n554 GND 0.05fF
C1111 VDD.n555 GND 0.16fF
C1112 VDD.n556 GND 0.01fF
C1113 VDD.n557 GND 0.02fF
C1114 VDD.n558 GND 0.02fF
C1115 VDD.n559 GND 0.18fF
C1116 VDD.n560 GND 0.01fF
C1117 VDD.n561 GND 0.02fF
C1118 VDD.n562 GND 0.02fF
C1119 VDD.n563 GND 0.07fF
C1120 VDD.n564 GND 0.24fF
C1121 VDD.n565 GND 0.01fF
C1122 VDD.n566 GND 0.01fF
C1123 VDD.n567 GND 0.02fF
C1124 VDD.n568 GND 0.29fF
C1125 VDD.n569 GND 0.01fF
C1126 VDD.n570 GND 0.02fF
C1127 VDD.n571 GND 0.02fF
C1128 VDD.n572 GND 0.29fF
C1129 VDD.n573 GND 0.01fF
C1130 VDD.n574 GND 0.02fF
C1131 VDD.n575 GND 0.04fF
C1132 VDD.n576 GND 0.28fF
C1133 VDD.n577 GND 0.02fF
C1134 VDD.n578 GND 0.02fF
C1135 VDD.n579 GND 0.02fF
C1136 VDD.n580 GND 0.06fF
C1137 VDD.n581 GND 0.02fF
C1138 VDD.n582 GND 0.02fF
C1139 VDD.n583 GND 0.02fF
C1140 VDD.n584 GND 0.02fF
C1141 VDD.n585 GND 0.02fF
C1142 VDD.n586 GND 0.02fF
C1143 VDD.n587 GND 0.02fF
C1144 VDD.n588 GND 0.02fF
C1145 VDD.n589 GND 0.02fF
C1146 VDD.n590 GND 0.02fF
C1147 VDD.n591 GND 0.03fF
C1148 VDD.n592 GND 0.02fF
C1149 VDD.n593 GND 0.02fF
C1150 VDD.n597 GND 0.29fF
C1151 VDD.n598 GND 0.29fF
C1152 VDD.n599 GND 0.01fF
C1153 VDD.n600 GND 0.02fF
C1154 VDD.n601 GND 0.04fF
C1155 VDD.n602 GND 0.06fF
C1156 VDD.n603 GND 0.26fF
C1157 VDD.n604 GND 0.01fF
C1158 VDD.n605 GND 0.01fF
C1159 VDD.n606 GND 0.02fF
C1160 VDD.n607 GND 0.18fF
C1161 VDD.n608 GND 0.01fF
C1162 VDD.n609 GND 0.02fF
C1163 VDD.n610 GND 0.02fF
C1164 VDD.n611 GND 0.09fF
C1165 VDD.n612 GND 0.05fF
C1166 VDD.n613 GND 0.01fF
C1167 VDD.n614 GND 0.02fF
C1168 VDD.n615 GND 0.03fF
C1169 VDD.n616 GND 0.15fF
C1170 VDD.n617 GND 0.01fF
C1171 VDD.n618 GND 0.02fF
C1172 VDD.n619 GND 0.03fF
C1173 VDD.n620 GND 0.17fF
C1174 VDD.n621 GND 0.01fF
C1175 VDD.n622 GND 0.02fF
C1176 VDD.n623 GND 0.02fF
C1177 VDD.n624 GND 0.07fF
C1178 VDD.n625 GND 0.26fF
C1179 VDD.n626 GND 0.01fF
C1180 VDD.n627 GND 0.01fF
C1181 VDD.n628 GND 0.02fF
C1182 VDD.n629 GND 0.29fF
C1183 VDD.n630 GND 0.01fF
C1184 VDD.n631 GND 0.02fF
C1185 VDD.n632 GND 0.04fF
C1186 VDD.n633 GND 0.28fF
C1187 VDD.n634 GND 0.02fF
C1188 VDD.n635 GND 0.02fF
C1189 VDD.n636 GND 0.02fF
C1190 VDD.n637 GND 0.06fF
C1191 VDD.n638 GND 0.02fF
C1192 VDD.n639 GND 0.02fF
C1193 VDD.n640 GND 0.02fF
C1194 VDD.n641 GND 0.02fF
C1195 VDD.n642 GND 0.02fF
C1196 VDD.n643 GND 0.02fF
C1197 VDD.n644 GND 0.02fF
C1198 VDD.n645 GND 0.02fF
C1199 VDD.n646 GND 0.02fF
C1200 VDD.n647 GND 0.02fF
C1201 VDD.n648 GND 0.03fF
C1202 VDD.n649 GND 0.02fF
C1203 VDD.n650 GND 0.02fF
C1204 VDD.n654 GND 0.29fF
C1205 VDD.n655 GND 0.29fF
C1206 VDD.n656 GND 0.01fF
C1207 VDD.n657 GND 0.02fF
C1208 VDD.n658 GND 0.04fF
C1209 VDD.n659 GND 0.29fF
C1210 VDD.n660 GND 0.01fF
C1211 VDD.n661 GND 0.02fF
C1212 VDD.n662 GND 0.02fF
C1213 VDD.n663 GND 0.23fF
C1214 VDD.n664 GND 0.01fF
C1215 VDD.n665 GND 0.07fF
C1216 VDD.n666 GND 0.02fF
C1217 VDD.n667 GND 0.18fF
C1218 VDD.n668 GND 0.01fF
C1219 VDD.n669 GND 0.02fF
C1220 VDD.n670 GND 0.02fF
C1221 VDD.n671 GND 0.17fF
C1222 VDD.n672 GND 0.01fF
C1223 VDD.n673 GND 0.09fF
C1224 VDD.n674 GND 0.05fF
C1225 VDD.n675 GND 0.02fF
C1226 VDD.n676 GND 0.02fF
C1227 VDD.n677 GND 0.15fF
C1228 VDD.n678 GND 0.02fF
C1229 VDD.n679 GND 0.02fF
C1230 VDD.n680 GND 0.03fF
C1231 VDD.n681 GND 0.16fF
C1232 VDD.n682 GND 0.02fF
C1233 VDD.n683 GND 0.02fF
C1234 VDD.n684 GND 0.03fF
C1235 VDD.n685 GND 0.09fF
C1236 VDD.n686 GND 0.05fF
C1237 VDD.n687 GND 0.16fF
C1238 VDD.n688 GND 0.01fF
C1239 VDD.n689 GND 0.02fF
C1240 VDD.n690 GND 0.02fF
C1241 VDD.n691 GND 0.18fF
C1242 VDD.n692 GND 0.01fF
C1243 VDD.n693 GND 0.02fF
C1244 VDD.n694 GND 0.02fF
C1245 VDD.n695 GND 0.07fF
C1246 VDD.n696 GND 0.24fF
C1247 VDD.n697 GND 0.01fF
C1248 VDD.n698 GND 0.01fF
C1249 VDD.n699 GND 0.02fF
C1250 VDD.n700 GND 0.29fF
C1251 VDD.n701 GND 0.01fF
C1252 VDD.n702 GND 0.02fF
C1253 VDD.n703 GND 0.02fF
C1254 VDD.n704 GND 0.33fF
C1255 VDD.n705 GND 0.02fF
C1256 VDD.n706 GND 0.02fF
C1257 VDD.n707 GND 0.02fF
C1258 VDD.n708 GND 0.06fF
C1259 VDD.n709 GND 0.02fF
C1260 VDD.n710 GND 0.02fF
C1261 VDD.n711 GND 0.02fF
C1262 VDD.n712 GND 0.02fF
C1263 VDD.n713 GND 0.02fF
C1264 VDD.n714 GND 0.02fF
C1265 VDD.n715 GND 0.02fF
C1266 VDD.n716 GND 0.02fF
C1267 VDD.n717 GND 0.02fF
C1268 VDD.n718 GND 0.02fF
C1269 VDD.n719 GND 0.03fF
C1270 VDD.n720 GND 0.02fF
C1271 VDD.n721 GND 0.02fF
C1272 VDD.n725 GND 0.29fF
C1273 VDD.n726 GND 0.29fF
C1274 VDD.n727 GND 0.01fF
C1275 VDD.n728 GND 0.02fF
C1276 VDD.n729 GND 0.02fF
C1277 VDD.n730 GND 0.19fF
C1278 VDD.n731 GND 0.02fF
C1279 VDD.n732 GND 0.02fF
C1280 VDD.n733 GND 0.06fF
C1281 VDD.n734 GND 0.02fF
C1282 VDD.n735 GND 0.02fF
C1283 VDD.n736 GND 0.02fF
C1284 VDD.n737 GND 0.02fF
C1285 VDD.n738 GND 0.02fF
C1286 VDD.n739 GND 0.02fF
C1287 VDD.n740 GND 0.02fF
C1288 VDD.n741 GND 0.02fF
C1289 VDD.n742 GND 0.03fF
C1290 VDD.n743 GND 0.04fF
C1291 VDD.n744 GND 0.02fF
C1292 VDD.n748 GND 0.48fF
C1293 VDD.n749 GND 0.29fF
C1294 VDD.n750 GND 0.02fF
C1295 VDD.n751 GND 0.03fF
C1296 VDD.n752 GND 0.03fF
C1297 VDD.n753 GND 0.29fF
C1298 VDD.n754 GND 0.01fF
C1299 VDD.n755 GND 0.02fF
C1300 VDD.n756 GND 0.02fF
C1301 VDD.n757 GND 0.07fF
C1302 VDD.n758 GND 0.24fF
C1303 VDD.n759 GND 0.01fF
C1304 VDD.n760 GND 0.01fF
C1305 VDD.n761 GND 0.02fF
C1306 VDD.n762 GND 0.18fF
C1307 VDD.n763 GND 0.01fF
C1308 VDD.n764 GND 0.02fF
C1309 VDD.n765 GND 0.02fF
C1310 VDD.n766 GND 0.09fF
C1311 VDD.n767 GND 0.05fF
C1312 VDD.n768 GND 0.16fF
C1313 VDD.n769 GND 0.01fF
C1314 VDD.n770 GND 0.02fF
C1315 VDD.n771 GND 0.02fF
C1316 VDD.n772 GND 0.16fF
C1317 VDD.n773 GND 0.02fF
C1318 VDD.n774 GND 0.02fF
C1319 VDD.n775 GND 0.03fF
C1320 VDD.n776 GND 0.15fF
C1321 VDD.n777 GND 0.02fF
C1322 VDD.n778 GND 0.02fF
C1323 VDD.n779 GND 0.03fF
C1324 VDD.n780 GND 0.17fF
C1325 VDD.n781 GND 0.01fF
C1326 VDD.n782 GND 0.09fF
C1327 VDD.n783 GND 0.05fF
C1328 VDD.n784 GND 0.02fF
C1329 VDD.n785 GND 0.02fF
C1330 VDD.n786 GND 0.18fF
C1331 VDD.n787 GND 0.01fF
C1332 VDD.n788 GND 0.02fF
C1333 VDD.n789 GND 0.02fF
C1334 VDD.n790 GND 0.23fF
C1335 VDD.n791 GND 0.01fF
C1336 VDD.n792 GND 0.07fF
C1337 VDD.n793 GND 0.02fF
C1338 VDD.n794 GND 0.29fF
C1339 VDD.n795 GND 0.01fF
C1340 VDD.n796 GND 0.02fF
C1341 VDD.n797 GND 0.02fF
C1342 VDD.n798 GND 0.29fF
C1343 VDD.n799 GND 0.01fF
C1344 VDD.n800 GND 0.02fF
C1345 VDD.n801 GND 0.04fF
C1346 VDD.n802 GND 0.06fF
C1347 VDD.n803 GND 0.02fF
C1348 VDD.n804 GND 0.02fF
C1349 VDD.n805 GND 0.02fF
C1350 VDD.n806 GND 0.02fF
C1351 VDD.n807 GND 0.02fF
C1352 VDD.n808 GND 0.02fF
C1353 VDD.n809 GND 0.02fF
C1354 VDD.n810 GND 0.02fF
C1355 VDD.n811 GND 0.02fF
C1356 VDD.n812 GND 0.02fF
C1357 VDD.n813 GND 0.02fF
C1358 VDD.n814 GND 0.03fF
C1359 VDD.n815 GND 0.02fF
C1360 VDD.n818 GND 0.02fF
C1361 VDD.n820 GND 0.02fF
C1362 VDD.n821 GND 0.33fF
C1363 VDD.n822 GND 0.02fF
C1364 VDD.n824 GND 0.29fF
C1365 VDD.n825 GND 0.29fF
C1366 VDD.n826 GND 0.01fF
C1367 VDD.n827 GND 0.02fF
C1368 VDD.n828 GND 0.04fF
C1369 VDD.n829 GND 0.29fF
C1370 VDD.n830 GND 0.01fF
C1371 VDD.n831 GND 0.02fF
C1372 VDD.n832 GND 0.02fF
C1373 VDD.n833 GND 0.07fF
C1374 VDD.n834 GND 0.24fF
C1375 VDD.n835 GND 0.01fF
C1376 VDD.n836 GND 0.01fF
C1377 VDD.n837 GND 0.02fF
C1378 VDD.n838 GND 0.18fF
C1379 VDD.n839 GND 0.01fF
C1380 VDD.n840 GND 0.02fF
C1381 VDD.n841 GND 0.02fF
C1382 VDD.n842 GND 0.09fF
C1383 VDD.n843 GND 0.05fF
C1384 VDD.n844 GND 0.16fF
C1385 VDD.n845 GND 0.01fF
C1386 VDD.n846 GND 0.02fF
C1387 VDD.n847 GND 0.02fF
C1388 VDD.n848 GND 0.16fF
C1389 VDD.n849 GND 0.02fF
C1390 VDD.n850 GND 0.02fF
C1391 VDD.n851 GND 0.03fF
C1392 VDD.n852 GND 0.15fF
C1393 VDD.n853 GND 0.02fF
C1394 VDD.n854 GND 0.02fF
C1395 VDD.n855 GND 0.03fF
C1396 VDD.n856 GND 0.17fF
C1397 VDD.n857 GND 0.01fF
C1398 VDD.n858 GND 0.09fF
C1399 VDD.n859 GND 0.05fF
C1400 VDD.n860 GND 0.02fF
C1401 VDD.n861 GND 0.02fF
C1402 VDD.n862 GND 0.18fF
C1403 VDD.n863 GND 0.01fF
C1404 VDD.n864 GND 0.02fF
C1405 VDD.n865 GND 0.02fF
C1406 VDD.n866 GND 0.23fF
C1407 VDD.n867 GND 0.01fF
C1408 VDD.n868 GND 0.07fF
C1409 VDD.n869 GND 0.02fF
C1410 VDD.n870 GND 0.29fF
C1411 VDD.n871 GND 0.01fF
C1412 VDD.n872 GND 0.02fF
C1413 VDD.n873 GND 0.02fF
C1414 VDD.n874 GND 0.29fF
C1415 VDD.n875 GND 0.01fF
C1416 VDD.n876 GND 0.02fF
C1417 VDD.n877 GND 0.04fF
C1418 VDD.n878 GND 0.28fF
C1419 VDD.n879 GND 0.02fF
C1420 VDD.n880 GND 0.02fF
C1421 VDD.n881 GND 0.02fF
C1422 VDD.n882 GND 0.06fF
C1423 VDD.n883 GND 0.02fF
C1424 VDD.n884 GND 0.02fF
C1425 VDD.n885 GND 0.02fF
C1426 VDD.n886 GND 0.02fF
C1427 VDD.n887 GND 0.02fF
C1428 VDD.n888 GND 0.02fF
C1429 VDD.n889 GND 0.02fF
C1430 VDD.n890 GND 0.02fF
C1431 VDD.n891 GND 0.02fF
C1432 VDD.n892 GND 0.02fF
C1433 VDD.n893 GND 0.03fF
C1434 VDD.n894 GND 0.02fF
C1435 VDD.n895 GND 0.02fF
C1436 VDD.n899 GND 0.29fF
C1437 VDD.n900 GND 0.29fF
C1438 VDD.n901 GND 0.01fF
C1439 VDD.n902 GND 0.02fF
C1440 VDD.n903 GND 0.04fF
C1441 VDD.n904 GND 0.07fF
C1442 VDD.n905 GND 0.26fF
C1443 VDD.n906 GND 0.01fF
C1444 VDD.n907 GND 0.01fF
C1445 VDD.n908 GND 0.02fF
C1446 VDD.n909 GND 0.17fF
C1447 VDD.n910 GND 0.01fF
C1448 VDD.n911 GND 0.02fF
C1449 VDD.n912 GND 0.02fF
C1450 VDD.n913 GND 0.15fF
C1451 VDD.n914 GND 0.01fF
C1452 VDD.n915 GND 0.02fF
C1453 VDD.n916 GND 0.03fF
C1454 VDD.n917 GND 0.09fF
C1455 VDD.n918 GND 0.05fF
C1456 VDD.n919 GND 0.01fF
C1457 VDD.n920 GND 0.02fF
C1458 VDD.n921 GND 0.03fF
C1459 VDD.n922 GND 0.18fF
C1460 VDD.n923 GND 0.01fF
C1461 VDD.n924 GND 0.02fF
C1462 VDD.n925 GND 0.02fF
C1463 VDD.n926 GND 0.06fF
C1464 VDD.n927 GND 0.26fF
C1465 VDD.n928 GND 0.01fF
C1466 VDD.n929 GND 0.01fF
C1467 VDD.n930 GND 0.02fF
C1468 VDD.n931 GND 0.29fF
C1469 VDD.n932 GND 0.01fF
C1470 VDD.n933 GND 0.02fF
C1471 VDD.n934 GND 0.04fF
C1472 VDD.n935 GND 0.28fF
C1473 VDD.n936 GND 0.02fF
C1474 VDD.n937 GND 0.02fF
C1475 VDD.n938 GND 0.02fF
C1476 VDD.n939 GND 0.06fF
C1477 VDD.n940 GND 0.02fF
C1478 VDD.n941 GND 0.02fF
C1479 VDD.n942 GND 0.02fF
C1480 VDD.n943 GND 0.02fF
C1481 VDD.n944 GND 0.02fF
C1482 VDD.n945 GND 0.02fF
C1483 VDD.n946 GND 0.02fF
C1484 VDD.n947 GND 0.02fF
C1485 VDD.n948 GND 0.02fF
C1486 VDD.n949 GND 0.02fF
C1487 VDD.n950 GND 0.03fF
C1488 VDD.n951 GND 0.02fF
C1489 VDD.n952 GND 0.02fF
C1490 VDD.n956 GND 0.29fF
C1491 VDD.n957 GND 0.29fF
C1492 VDD.n958 GND 0.01fF
C1493 VDD.n959 GND 0.02fF
C1494 VDD.n960 GND 0.04fF
C1495 VDD.n961 GND 0.29fF
C1496 VDD.n962 GND 0.01fF
C1497 VDD.n963 GND 0.02fF
C1498 VDD.n964 GND 0.02fF
C1499 VDD.n965 GND 0.07fF
C1500 VDD.n966 GND 0.24fF
C1501 VDD.n967 GND 0.01fF
C1502 VDD.n968 GND 0.01fF
C1503 VDD.n969 GND 0.02fF
C1504 VDD.n970 GND 0.18fF
C1505 VDD.n971 GND 0.01fF
C1506 VDD.n972 GND 0.02fF
C1507 VDD.n973 GND 0.02fF
C1508 VDD.n974 GND 0.09fF
C1509 VDD.n975 GND 0.05fF
C1510 VDD.n976 GND 0.16fF
C1511 VDD.n977 GND 0.01fF
C1512 VDD.n978 GND 0.02fF
C1513 VDD.n979 GND 0.02fF
C1514 VDD.n980 GND 0.16fF
C1515 VDD.n981 GND 0.02fF
C1516 VDD.n982 GND 0.02fF
C1517 VDD.n983 GND 0.03fF
C1518 VDD.n984 GND 0.15fF
C1519 VDD.n985 GND 0.02fF
C1520 VDD.n986 GND 0.02fF
C1521 VDD.n987 GND 0.03fF
C1522 VDD.n988 GND 0.17fF
C1523 VDD.n989 GND 0.01fF
C1524 VDD.n990 GND 0.09fF
C1525 VDD.n991 GND 0.05fF
C1526 VDD.n992 GND 0.02fF
C1527 VDD.n993 GND 0.02fF
C1528 VDD.n994 GND 0.18fF
C1529 VDD.n995 GND 0.01fF
C1530 VDD.n996 GND 0.02fF
C1531 VDD.n997 GND 0.02fF
C1532 VDD.n998 GND 0.23fF
C1533 VDD.n999 GND 0.01fF
C1534 VDD.n1000 GND 0.07fF
C1535 VDD.n1001 GND 0.02fF
C1536 VDD.n1002 GND 0.29fF
C1537 VDD.n1003 GND 0.01fF
C1538 VDD.n1004 GND 0.02fF
C1539 VDD.n1005 GND 0.02fF
C1540 VDD.n1006 GND 0.29fF
C1541 VDD.n1007 GND 0.01fF
C1542 VDD.n1008 GND 0.02fF
C1543 VDD.n1009 GND 0.04fF
C1544 VDD.n1010 GND 0.33fF
C1545 VDD.n1011 GND 0.02fF
C1546 VDD.n1012 GND 0.02fF
C1547 VDD.n1013 GND 0.02fF
C1548 VDD.n1014 GND 0.06fF
C1549 VDD.n1015 GND 0.02fF
C1550 VDD.n1016 GND 0.02fF
C1551 VDD.n1017 GND 0.02fF
C1552 VDD.n1018 GND 0.02fF
C1553 VDD.n1019 GND 0.02fF
C1554 VDD.n1020 GND 0.02fF
C1555 VDD.n1021 GND 0.02fF
C1556 VDD.n1022 GND 0.02fF
C1557 VDD.n1023 GND 0.02fF
C1558 VDD.n1024 GND 0.02fF
C1559 VDD.n1025 GND 0.03fF
C1560 VDD.n1026 GND 0.02fF
C1561 VDD.n1027 GND 0.02fF
C1562 VDD.n1031 GND 0.29fF
C1563 VDD.n1032 GND 0.29fF
C1564 VDD.n1033 GND 0.01fF
C1565 VDD.n1034 GND 0.02fF
C1566 VDD.n1035 GND 0.04fF
C1567 VDD.n1036 GND 0.29fF
C1568 VDD.n1037 GND 0.01fF
C1569 VDD.n1038 GND 0.02fF
C1570 VDD.n1039 GND 0.02fF
C1571 VDD.n1040 GND 0.07fF
C1572 VDD.n1041 GND 0.24fF
C1573 VDD.n1042 GND 0.01fF
C1574 VDD.n1043 GND 0.01fF
C1575 VDD.n1044 GND 0.02fF
C1576 VDD.n1045 GND 0.18fF
C1577 VDD.n1046 GND 0.01fF
C1578 VDD.n1047 GND 0.02fF
C1579 VDD.n1048 GND 0.02fF
C1580 VDD.n1049 GND 0.09fF
C1581 VDD.n1050 GND 0.05fF
C1582 VDD.n1051 GND 0.16fF
C1583 VDD.n1052 GND 0.01fF
C1584 VDD.n1053 GND 0.02fF
C1585 VDD.n1054 GND 0.02fF
C1586 VDD.n1055 GND 0.16fF
C1587 VDD.n1056 GND 0.02fF
C1588 VDD.n1057 GND 0.02fF
C1589 VDD.n1058 GND 0.03fF
C1590 VDD.n1059 GND 0.15fF
C1591 VDD.n1060 GND 0.02fF
C1592 VDD.n1061 GND 0.02fF
C1593 VDD.n1062 GND 0.03fF
C1594 VDD.n1063 GND 0.17fF
C1595 VDD.n1064 GND 0.01fF
C1596 VDD.n1065 GND 0.09fF
C1597 VDD.n1066 GND 0.05fF
C1598 VDD.n1067 GND 0.02fF
C1599 VDD.n1068 GND 0.02fF
C1600 VDD.n1069 GND 0.18fF
C1601 VDD.n1070 GND 0.01fF
C1602 VDD.n1071 GND 0.02fF
C1603 VDD.n1072 GND 0.02fF
C1604 VDD.n1073 GND 0.23fF
C1605 VDD.n1074 GND 0.01fF
C1606 VDD.n1075 GND 0.07fF
C1607 VDD.n1076 GND 0.02fF
C1608 VDD.n1077 GND 0.29fF
C1609 VDD.n1078 GND 0.01fF
C1610 VDD.n1079 GND 0.02fF
C1611 VDD.n1080 GND 0.02fF
C1612 VDD.n1081 GND 0.29fF
C1613 VDD.n1082 GND 0.01fF
C1614 VDD.n1083 GND 0.02fF
C1615 VDD.n1084 GND 0.04fF
C1616 VDD.n1085 GND 0.28fF
C1617 VDD.n1086 GND 0.02fF
C1618 VDD.n1087 GND 0.02fF
C1619 VDD.n1088 GND 0.02fF
C1620 VDD.n1089 GND 0.06fF
C1621 VDD.n1090 GND 0.02fF
C1622 VDD.n1091 GND 0.02fF
C1623 VDD.n1092 GND 0.02fF
C1624 VDD.n1093 GND 0.02fF
C1625 VDD.n1094 GND 0.02fF
C1626 VDD.n1095 GND 0.02fF
C1627 VDD.n1096 GND 0.02fF
C1628 VDD.n1097 GND 0.02fF
C1629 VDD.n1098 GND 0.02fF
C1630 VDD.n1099 GND 0.02fF
C1631 VDD.n1100 GND 0.03fF
C1632 VDD.n1101 GND 0.02fF
C1633 VDD.n1102 GND 0.02fF
C1634 VDD.n1106 GND 0.29fF
C1635 VDD.n1107 GND 0.29fF
C1636 VDD.n1108 GND 0.01fF
C1637 VDD.n1109 GND 0.02fF
C1638 VDD.n1110 GND 0.04fF
C1639 VDD.n1111 GND 0.07fF
C1640 VDD.n1112 GND 0.26fF
C1641 VDD.n1113 GND 0.01fF
C1642 VDD.n1114 GND 0.01fF
C1643 VDD.n1115 GND 0.02fF
C1644 VDD.n1116 GND 0.17fF
C1645 VDD.n1117 GND 0.01fF
C1646 VDD.n1118 GND 0.02fF
C1647 VDD.n1119 GND 0.02fF
C1648 VDD.n1120 GND 0.15fF
C1649 VDD.n1121 GND 0.01fF
C1650 VDD.n1122 GND 0.02fF
C1651 VDD.n1123 GND 0.03fF
C1652 VDD.n1124 GND 0.09fF
C1653 VDD.n1125 GND 0.05fF
C1654 VDD.n1126 GND 0.01fF
C1655 VDD.n1127 GND 0.02fF
C1656 VDD.n1128 GND 0.03fF
C1657 VDD.n1129 GND 0.18fF
C1658 VDD.n1130 GND 0.01fF
C1659 VDD.n1131 GND 0.02fF
C1660 VDD.n1132 GND 0.02fF
C1661 VDD.n1133 GND 0.06fF
C1662 VDD.n1134 GND 0.26fF
C1663 VDD.n1135 GND 0.01fF
C1664 VDD.n1136 GND 0.01fF
C1665 VDD.n1137 GND 0.02fF
C1666 VDD.n1138 GND 0.29fF
C1667 VDD.n1139 GND 0.01fF
C1668 VDD.n1140 GND 0.02fF
C1669 VDD.n1141 GND 0.04fF
C1670 VDD.n1142 GND 0.28fF
C1671 VDD.n1143 GND 0.02fF
C1672 VDD.n1144 GND 0.02fF
C1673 VDD.n1145 GND 0.02fF
C1674 VDD.n1146 GND 0.06fF
C1675 VDD.n1147 GND 0.02fF
C1676 VDD.n1148 GND 0.02fF
C1677 VDD.n1149 GND 0.02fF
C1678 VDD.n1150 GND 0.02fF
C1679 VDD.n1151 GND 0.02fF
C1680 VDD.n1152 GND 0.02fF
C1681 VDD.n1153 GND 0.02fF
C1682 VDD.n1154 GND 0.02fF
C1683 VDD.n1155 GND 0.02fF
C1684 VDD.n1156 GND 0.02fF
C1685 VDD.n1157 GND 0.03fF
C1686 VDD.n1158 GND 0.02fF
C1687 VDD.n1159 GND 0.02fF
C1688 VDD.n1163 GND 0.29fF
C1689 VDD.n1164 GND 0.29fF
C1690 VDD.n1165 GND 0.01fF
C1691 VDD.n1166 GND 0.02fF
C1692 VDD.n1167 GND 0.04fF
C1693 VDD.n1168 GND 0.29fF
C1694 VDD.n1169 GND 0.01fF
C1695 VDD.n1170 GND 0.02fF
C1696 VDD.n1171 GND 0.02fF
C1697 VDD.n1172 GND 0.07fF
C1698 VDD.n1173 GND 0.24fF
C1699 VDD.n1174 GND 0.01fF
C1700 VDD.n1175 GND 0.01fF
C1701 VDD.n1176 GND 0.02fF
C1702 VDD.n1177 GND 0.18fF
C1703 VDD.n1178 GND 0.01fF
C1704 VDD.n1179 GND 0.02fF
C1705 VDD.n1180 GND 0.02fF
C1706 VDD.n1181 GND 0.09fF
C1707 VDD.n1182 GND 0.05fF
C1708 VDD.n1183 GND 0.16fF
C1709 VDD.n1184 GND 0.01fF
C1710 VDD.n1185 GND 0.02fF
C1711 VDD.n1186 GND 0.02fF
C1712 VDD.n1187 GND 0.16fF
C1713 VDD.n1188 GND 0.02fF
C1714 VDD.n1189 GND 0.02fF
C1715 VDD.n1190 GND 0.03fF
C1716 VDD.n1191 GND 0.15fF
C1717 VDD.n1192 GND 0.02fF
C1718 VDD.n1193 GND 0.02fF
C1719 VDD.n1194 GND 0.03fF
C1720 VDD.n1195 GND 0.17fF
C1721 VDD.n1196 GND 0.01fF
C1722 VDD.n1197 GND 0.09fF
C1723 VDD.n1198 GND 0.05fF
C1724 VDD.n1199 GND 0.02fF
C1725 VDD.n1200 GND 0.02fF
C1726 VDD.n1201 GND 0.18fF
C1727 VDD.n1202 GND 0.01fF
C1728 VDD.n1203 GND 0.02fF
C1729 VDD.n1204 GND 0.02fF
C1730 VDD.n1205 GND 0.23fF
C1731 VDD.n1206 GND 0.01fF
C1732 VDD.n1207 GND 0.07fF
C1733 VDD.n1208 GND 0.02fF
C1734 VDD.n1209 GND 0.29fF
C1735 VDD.n1210 GND 0.01fF
C1736 VDD.n1211 GND 0.02fF
C1737 VDD.n1212 GND 0.02fF
C1738 VDD.n1213 GND 0.29fF
C1739 VDD.n1214 GND 0.01fF
C1740 VDD.n1215 GND 0.02fF
C1741 VDD.n1216 GND 0.04fF
C1742 VDD.n1217 GND 0.33fF
C1743 VDD.n1218 GND 0.02fF
C1744 VDD.n1219 GND 0.02fF
C1745 VDD.n1220 GND 0.02fF
C1746 VDD.n1221 GND 0.06fF
C1747 VDD.n1222 GND 0.02fF
C1748 VDD.n1223 GND 0.02fF
C1749 VDD.n1224 GND 0.02fF
C1750 VDD.n1225 GND 0.02fF
C1751 VDD.n1226 GND 0.02fF
C1752 VDD.n1227 GND 0.02fF
C1753 VDD.n1228 GND 0.02fF
C1754 VDD.n1229 GND 0.02fF
C1755 VDD.n1230 GND 0.02fF
C1756 VDD.n1231 GND 0.02fF
C1757 VDD.n1232 GND 0.03fF
C1758 VDD.n1233 GND 0.02fF
C1759 VDD.n1234 GND 0.02fF
C1760 VDD.n1238 GND 0.29fF
C1761 VDD.n1239 GND 0.29fF
C1762 VDD.n1240 GND 0.01fF
C1763 VDD.n1241 GND 0.02fF
C1764 VDD.n1242 GND 0.04fF
C1765 VDD.n1243 GND 0.29fF
C1766 VDD.n1244 GND 0.01fF
C1767 VDD.n1245 GND 0.02fF
C1768 VDD.n1246 GND 0.02fF
C1769 VDD.n1247 GND 0.07fF
C1770 VDD.n1248 GND 0.24fF
C1771 VDD.n1249 GND 0.01fF
C1772 VDD.n1250 GND 0.01fF
C1773 VDD.n1251 GND 0.02fF
C1774 VDD.n1252 GND 0.18fF
C1775 VDD.n1253 GND 0.01fF
C1776 VDD.n1254 GND 0.02fF
C1777 VDD.n1255 GND 0.02fF
C1778 VDD.n1256 GND 0.09fF
C1779 VDD.n1257 GND 0.05fF
C1780 VDD.n1258 GND 0.16fF
C1781 VDD.n1259 GND 0.01fF
C1782 VDD.n1260 GND 0.02fF
C1783 VDD.n1261 GND 0.02fF
C1784 VDD.n1262 GND 0.16fF
C1785 VDD.n1263 GND 0.02fF
C1786 VDD.n1264 GND 0.02fF
C1787 VDD.n1265 GND 0.03fF
C1788 VDD.n1266 GND 0.15fF
C1789 VDD.n1267 GND 0.02fF
C1790 VDD.n1268 GND 0.02fF
C1791 VDD.n1269 GND 0.03fF
C1792 VDD.n1270 GND 0.17fF
C1793 VDD.n1271 GND 0.01fF
C1794 VDD.n1272 GND 0.09fF
C1795 VDD.n1273 GND 0.05fF
C1796 VDD.n1274 GND 0.02fF
C1797 VDD.n1275 GND 0.02fF
C1798 VDD.n1276 GND 0.18fF
C1799 VDD.n1277 GND 0.01fF
C1800 VDD.n1278 GND 0.02fF
C1801 VDD.n1279 GND 0.02fF
C1802 VDD.n1280 GND 0.23fF
C1803 VDD.n1281 GND 0.01fF
C1804 VDD.n1282 GND 0.07fF
C1805 VDD.n1283 GND 0.02fF
C1806 VDD.n1284 GND 0.29fF
C1807 VDD.n1285 GND 0.01fF
C1808 VDD.n1286 GND 0.02fF
C1809 VDD.n1287 GND 0.02fF
C1810 VDD.n1288 GND 0.29fF
C1811 VDD.n1289 GND 0.01fF
C1812 VDD.n1290 GND 0.02fF
C1813 VDD.n1291 GND 0.04fF
C1814 VDD.n1292 GND 0.28fF
C1815 VDD.n1293 GND 0.02fF
C1816 VDD.n1294 GND 0.02fF
C1817 VDD.n1295 GND 0.02fF
C1818 VDD.n1296 GND 0.06fF
C1819 VDD.n1297 GND 0.02fF
C1820 VDD.n1298 GND 0.02fF
C1821 VDD.n1299 GND 0.02fF
C1822 VDD.n1300 GND 0.02fF
C1823 VDD.n1301 GND 0.02fF
C1824 VDD.n1302 GND 0.02fF
C1825 VDD.n1303 GND 0.02fF
C1826 VDD.n1304 GND 0.02fF
C1827 VDD.n1305 GND 0.02fF
C1828 VDD.n1306 GND 0.02fF
C1829 VDD.n1307 GND 0.03fF
C1830 VDD.n1308 GND 0.02fF
C1831 VDD.n1309 GND 0.02fF
C1832 VDD.n1313 GND 0.29fF
C1833 VDD.n1314 GND 0.29fF
C1834 VDD.n1315 GND 0.01fF
C1835 VDD.n1316 GND 0.02fF
C1836 VDD.n1317 GND 0.04fF
C1837 VDD.n1318 GND 0.07fF
C1838 VDD.n1319 GND 0.26fF
C1839 VDD.n1320 GND 0.01fF
C1840 VDD.n1321 GND 0.01fF
C1841 VDD.n1322 GND 0.02fF
C1842 VDD.n1323 GND 0.17fF
C1843 VDD.n1324