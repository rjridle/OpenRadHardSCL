* SPICE3 file created from HA.ext - technology: sky130A

.subckt HA SUM COUT A B VDD GND
X0 VDD.t31 A.t0 a_217_1050.t3 �w˶U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X1 GND a_1917_990.t3 a_2332_101.t0 GND sky130_fd_pr__nfet_01v8 ad=3.9597p pd=2.901u as=0p ps=0u w=0u l=0u
X2 COUT.t2 a_217_1050.t5 VDD.t19 �t�˶U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X3 a_1295_209.t2 A.t1 VDD.t29 ��*̶U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X4 VDD.t11 B.t1 a_217_1050.t1 P�*̶U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X5 GND A.t2 a_112_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X6 SUM.t3 a_1295_209.t3 a_2351_1051.t3  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X7 VDD.t13 B.t3 a_1917_990.t2 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X8 SUM a_1295_209.t4 a_2332_101.t1 GND sky130_fd_pr__nfet_01v8 ad=3.582p pd=3.14u as=0p ps=0u w=0u l=0u
X9 a_1685_1051.t1 a_1917_990.t4 SUM.t0  ,��r sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X10 a_217_1050.t4 A.t3 VDD.t27 VDD.t26 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X11 SUM.t1 a_1917_990.t5 a_1685_1051.t0  ,��r sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X12 GND A.t6 a_1666_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X13 a_217_1050.t0 B.t4 VDD.t7 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X14 VDD.t17 a_217_1050.t7 COUT.t1  ,��r sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X15 VDD.t25 A.t4 a_1685_1051.t3 �+��r sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X16 VDD.t23 A.t5 a_1295_209.t1  ,��r sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X17 a_2351_1051.t1 B.t5 VDD.t5 �+��r sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X18 a_1917_990.t1 B.t6 VDD.t15  ,��r sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X19 a_2351_1051.t2 a_1295_209.t5 SUM.t5 �+��r sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X20 a_1685_1051.t2 A.t8 VDD.t21  ,��r sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X21 VDD.t3 B.t8 a_2351_1051.t0 �+��r sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X22 SUM B.t0 a_1666_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X23 COUT a_217_1050.t6 GND.t3 GND sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=0p ps=0u w=0u l=0u
C0 B SUM 0.89fF
C1 VDD B 2.34fF
C2 COUT B 0.07fF
C3 VDD SUM 1.04fF
C4 A B 1.08fF
C5 VDD COUT 1.10fF
C6 A SUM 0.08fF
C7 A VDD 2.56fF
C8 A COUT 0.12fF
R0 A.n2 A.t5 512.525
R1 A.n5 A.t0 480.392
R2 A.n0 A.t8 480.392
R3 A.n6 A.t2 412.921
R4 A.n1 A.t6 412.921
R5 A.n5 A.t3 403.272
R6 A.n0 A.t4 403.272
R7 A.n2 A.t1 371.139
R8 A.n3 A.t7 366.428
R9 A.n3 A.n2 163.771
R10 A.n1 A.n0 115.947
R11 A.n6 A.n5 115.571
R12 A.n4 A.n1 6.509
R13 A.n4 A.n3 4.65
R14 A.n7 A.n6 4.65
R15 A.n7 A.n4 3.763
R16 A.n7 A 0.046
R17 a_217_1050.n3 a_217_1050.t7 512.525
R18 a_217_1050.n3 a_217_1050.t5 371.139
R19 a_217_1050.n7 a_217_1050.n5 284.244
R20 a_217_1050.n4 a_217_1050.t6 282.852
R21 a_217_1050.n4 a_217_1050.n3 247.347
R22 a_217_1050.n5 a_217_1050.n2 187.858
R23 a_217_1050.n2 a_217_1050.n1 157.964
R24 a_217_1050.n2 a_217_1050.n0 91.706
R25 a_217_1050.n7 a_217_1050.n6 15.218
R26 a_217_1050.n0 a_217_1050.t1 14.282
R27 a_217_1050.n0 a_217_1050.t0 14.282
R28 a_217_1050.n1 a_217_1050.t3 14.282
R29 a_217_1050.n1 a_217_1050.t4 14.282
R30 a_217_1050.n8 a_217_1050.n7 12.014
R31 a_217_1050.n5 a_217_1050.n4 10.343
R32 VDD.n140 VDD.n139 173.148
R33 VDD.n85 VDD.n84 173.148
R34 VDD.n227 VDD.n216 144.705
R35 VDD.n255 VDD.n248 144.705
R36 VDD.n121 VDD.n114 144.705
R37 VDD.n315 VDD.n308 144.705
R38 VDD.n66 VDD.n55 144.705
R39 VDD.n194 VDD.t11 143.754
R40 VDD.n172 VDD.t27 135.17
R41 VDD.n232 VDD.t19 135.17
R42 VDD.n239 VDD.t17 135.17
R43 VDD.n274 VDD.t29 135.17
R44 VDD.n283 VDD.t23 135.17
R45 VDD.n35 VDD.t15 135.17
R46 VDD.n24 VDD.t13 135.17
R47 VDD.n186 VDD.n185 129.472
R48 VDD.n51 VDD.n50 92.5
R49 VDD.n49 VDD.n48 92.5
R50 VDD.n47 VDD.n46 92.5
R51 VDD.n45 VDD.n44 92.5
R52 VDD.n53 VDD.n52 92.5
R53 VDD.n110 VDD.n109 92.5
R54 VDD.n108 VDD.n107 92.5
R55 VDD.n106 VDD.n105 92.5
R56 VDD.n104 VDD.n103 92.5
R57 VDD.n112 VDD.n111 92.5
R58 VDD.n304 VDD.n303 92.5
R59 VDD.n302 VDD.n301 92.5
R60 VDD.n300 VDD.n299 92.5
R61 VDD.n298 VDD.n297 92.5
R62 VDD.n306 VDD.n305 92.5
R63 VDD.n268 VDD.n267 92.5
R64 VDD.n266 VDD.n265 92.5
R65 VDD.n264 VDD.n263 92.5
R66 VDD.n262 VDD.n261 92.5
R67 VDD.n270 VDD.n269 92.5
R68 VDD.n212 VDD.n211 92.5
R69 VDD.n210 VDD.n209 92.5
R70 VDD.n208 VDD.n207 92.5
R71 VDD.n206 VDD.n205 92.5
R72 VDD.n214 VDD.n213 92.5
R73 VDD.n160 VDD.n159 92.5
R74 VDD.n158 VDD.n157 92.5
R75 VDD.n156 VDD.n155 92.5
R76 VDD.n154 VDD.n153 92.5
R77 VDD.n162 VDD.n161 92.5
R78 VDD.n14 VDD.n1 92.5
R79 VDD.n5 VDD.n4 92.5
R80 VDD.n7 VDD.n6 92.5
R81 VDD.n9 VDD.n8 92.5
R82 VDD.n11 VDD.n10 92.5
R83 VDD.n13 VDD.n12 92.5
R84 VDD.n21 VDD.n20 92.059
R85 VDD.n65 VDD.n64 92.059
R86 VDD.n120 VDD.n119 92.059
R87 VDD.n314 VDD.n313 92.059
R88 VDD.n254 VDD.n253 92.059
R89 VDD.n226 VDD.n225 92.059
R90 VDD.n168 VDD.n167 92.059
R91 VDD.n20 VDD.n16 67.194
R92 VDD.n20 VDD.n17 67.194
R93 VDD.n20 VDD.n18 67.194
R94 VDD.n20 VDD.n19 67.194
R95 VDD.n152 VDD.n151 44.141
R96 VDD.n260 VDD.n259 44.141
R97 VDD.n296 VDD.n295 44.141
R98 VDD.n102 VDD.n101 44.141
R99 VDD.n5 VDD.n3 44.141
R100 VDD.n259 VDD.n257 44.107
R101 VDD.n295 VDD.n293 44.107
R102 VDD.n101 VDD.n99 44.107
R103 VDD.n151 VDD.n149 44.107
R104 VDD.n3 VDD.n2 44.107
R105 VDD.n25 VDD.t12 43.472
R106 VDD.n33  ,��r 43.472
R107 VDD.n284  ,��r 43.472
R108 VDD.n275 ��*̶U 43.472
R109 VDD.n240  ,��r 43.472
R110 VDD.n230 �t�˶U 43.472
R111 VDD.n20 VDD.n15 41.052
R112 VDD.n59 VDD.n57 39.742
R113 VDD.n59 VDD.n58 39.742
R114 VDD.n61 VDD.n60 39.742
R115 VDD.n116 VDD.n115 39.742
R116 VDD.n310 VDD.n309 39.742
R117 VDD.n250 VDD.n249 39.742
R118 VDD.n164 VDD.n163 39.742
R119 VDD.n224 VDD.n221 39.742
R120 VDD.n224 VDD.n223 39.742
R121 VDD.n220 VDD.n219 39.742
R122 VDD.n101 VDD.n100 38
R123 VDD.n295 VDD.n294 38
R124 VDD.n259 VDD.n258 38
R125 VDD.n151 VDD.n150 38
R126 VDD.n257 VDD.n256 36.774
R127 VDD.n293 VDD.n292 36.774
R128 VDD.n99 VDD.n98 36.774
R129 VDD.n57 VDD.n56 36.774
R130 VDD.n223 VDD.n222 36.774
R131 VDD.n1 VDD.n0 30.923
R132 VDD.n64 VDD.n62 26.38
R133 VDD.n64 VDD.n61 26.38
R134 VDD.n64 VDD.n59 26.38
R135 VDD.n64 VDD.n63 26.38
R136 VDD.n119 VDD.n117 26.38
R137 VDD.n119 VDD.n116 26.38
R138 VDD.n119 VDD.n118 26.38
R139 VDD.n313 VDD.n311 26.38
R140 VDD.n313 VDD.n310 26.38
R141 VDD.n313 VDD.n312 26.38
R142 VDD.n253 VDD.n251 26.38
R143 VDD.n253 VDD.n250 26.38
R144 VDD.n253 VDD.n252 26.38
R145 VDD.n167 VDD.n165 26.38
R146 VDD.n167 VDD.n164 26.38
R147 VDD.n167 VDD.n166 26.38
R148 VDD.n225 VDD.n224 26.38
R149 VDD.n225 VDD.n220 26.38
R150 VDD.n225 VDD.n218 26.38
R151 VDD.n225 VDD.n217 26.38
R152 VDD.n170 VDD.n162 22.915
R153 VDD.n23 VDD.n14 22.915
R154 VDD.n73 �+��r 20.457
R155 VDD.n128  ,��r 20.457
R156 VDD.n190 P�*̶U 20.457
R157 VDD.n86 �+��r 17.9
R158 VDD.n141 �+��r 17.9
R159 VDD.n177 VDD.t26 17.9
R160 VDD.n162 VDD.n160 14.864
R161 VDD.n160 VDD.n158 14.864
R162 VDD.n158 VDD.n156 14.864
R163 VDD.n156 VDD.n154 14.864
R164 VDD.n154 VDD.n152 14.864
R165 VDD.n270 VDD.n268 14.864
R166 VDD.n268 VDD.n266 14.864
R167 VDD.n266 VDD.n264 14.864
R168 VDD.n264 VDD.n262 14.864
R169 VDD.n262 VDD.n260 14.864
R170 VDD.n306 VDD.n304 14.864
R171 VDD.n304 VDD.n302 14.864
R172 VDD.n302 VDD.n300 14.864
R173 VDD.n300 VDD.n298 14.864
R174 VDD.n298 VDD.n296 14.864
R175 VDD.n112 VDD.n110 14.864
R176 VDD.n110 VDD.n108 14.864
R177 VDD.n108 VDD.n106 14.864
R178 VDD.n106 VDD.n104 14.864
R179 VDD.n104 VDD.n102 14.864
R180 VDD.n53 VDD.n51 14.864
R181 VDD.n51 VDD.n49 14.864
R182 VDD.n49 VDD.n47 14.864
R183 VDD.n47 VDD.n45 14.864
R184 VDD.n45 VDD.n43 14.864
R185 VDD.n43 VDD.n42 14.864
R186 VDD.n214 VDD.n212 14.864
R187 VDD.n212 VDD.n210 14.864
R188 VDD.n210 VDD.n208 14.864
R189 VDD.n208 VDD.n206 14.864
R190 VDD.n206 VDD.n204 14.864
R191 VDD.n204 VDD.n203 14.864
R192 VDD.n14 VDD.n13 14.864
R193 VDD.n13 VDD.n11 14.864
R194 VDD.n11 VDD.n9 14.864
R195 VDD.n9 VDD.n7 14.864
R196 VDD.n7 VDD.n5 14.864
R197 VDD.n67 VDD.n54 14.864
R198 VDD.n122 VDD.n113 14.864
R199 VDD.n316 VDD.n307 14.864
R200 VDD.n272 VDD.n271 14.864
R201 VDD.n228 VDD.n215 14.864
R202 VDD.n185 VDD.t7 14.282
R203 VDD.n185 VDD.t31 14.282
R204 VDD.n139 VDD.t21 14.282
R205 VDD.n139 VDD.t25 14.282
R206 VDD.n84 VDD.t5 14.282
R207 VDD.n84 VDD.t3 14.282
R208 VDD.n188 VDD.n186 9.083
R209 VDD.n23 VDD.n22 8.855
R210 VDD.n22 VDD.n21 8.855
R211 VDD.n27 VDD.n26 8.855
R212 VDD.n26 VDD.n25 8.855
R213 VDD.n31 VDD.n30 8.855
R214 VDD.n30 VDD.n29 8.855
R215 VDD.n36 VDD.n34 8.855
R216 VDD.n34 VDD.n33 8.855
R217 VDD.n40 VDD.n39 8.855
R218 VDD.n39 VDD.n38 8.855
R219 VDD.n67 VDD.n66 8.855
R220 VDD.n66 VDD.n65 8.855
R221 VDD.n71 VDD.n70 8.855
R222 VDD.n70 VDD.n69 8.855
R223 VDD.n75 VDD.n74 8.855
R224 VDD.n74 VDD.n73 8.855
R225 VDD.n78 VDD.n77 8.855
R226 VDD.n77 ��\̶U 8.855
R227 VDD.n82 VDD.n81 8.855
R228 VDD.n81 VDD.n80 8.855
R229 VDD.n88 VDD.n87 8.855
R230 VDD.n87 VDD.n86 8.855
R231 VDD.n92 VDD.n91 8.855
R232 VDD.n91 VDD.n90 8.855
R233 VDD.n96 VDD.n95 8.855
R234 VDD.n95 VDD.n94 8.855
R235 VDD.n122 VDD.n121 8.855
R236 VDD.n121 VDD.n120 8.855
R237 VDD.n126 VDD.n125 8.855
R238 VDD.n125 VDD.n124 8.855
R239 VDD.n130 VDD.n129 8.855
R240 VDD.n129 VDD.n128 8.855
R241 VDD.n133 VDD.n132 8.855
R242 VDD.n132  ,��r 8.855
R243 VDD.n137 VDD.n136 8.855
R244 VDD.n136 VDD.n135 8.855
R245 VDD.n143 VDD.n142 8.855
R246 VDD.n142 VDD.n141 8.855
R247 VDD.n147 VDD.n146 8.855
R248 VDD.n146 VDD.n145 8.855
R249 VDD.n316 VDD.n315 8.855
R250 VDD.n315 VDD.n314 8.855
R251 VDD.n290 VDD.n289 8.855
R252 VDD.n289 VDD.n288 8.855
R253 VDD.n286 VDD.n285 8.855
R254 VDD.n285 VDD.n284 8.855
R255 VDD.n281 VDD.n280 8.855
R256 VDD.n280 VDD.n279 8.855
R257 VDD.n277 VDD.n276 8.855
R258 VDD.n276 VDD.n275 8.855
R259 VDD.n272 VDD.n255 8.855
R260 VDD.n255 VDD.n254 8.855
R261 VDD.n246 VDD.n245 8.855
R262 VDD.n245 VDD.n244 8.855
R263 VDD.n242 VDD.n241 8.855
R264 VDD.n241 VDD.n240 8.855
R265 VDD.n237 VDD.n236 8.855
R266 VDD.n236 VDD.n235 8.855
R267 VDD.n233 VDD.n231 8.855
R268 VDD.n231 VDD.n230 8.855
R269 VDD.n228 VDD.n227 8.855
R270 VDD.n227 VDD.n226 8.855
R271 VDD.n201 VDD.n200 8.855
R272 VDD.n200 VDD.n199 8.855
R273 VDD.n197 VDD.n196 8.855
R274 VDD.n196 VDD.n195 8.855
R275 VDD.n192 VDD.n191 8.855
R276 VDD.n191 VDD.n190 8.855
R277 VDD.n188 VDD.n187 8.855
R278 VDD.n187 VDD.t6 8.855
R279 VDD.n183 VDD.n182 8.855
R280 VDD.n182 VDD.n181 8.855
R281 VDD.n179 VDD.n178 8.855
R282 VDD.n178 VDD.n177 8.855
R283 VDD.n175 VDD.n174 8.855
R284 VDD.n174 VDD.n173 8.855
R285 VDD.n170 VDD.n169 8.855
R286 VDD.n169 VDD.n168 8.855
R287 VDD.n271 VDD.n270 8.051
R288 VDD.n307 VDD.n306 8.051
R289 VDD.n113 VDD.n112 8.051
R290 VDD.n54 VDD.n53 8.051
R291 VDD.n215 VDD.n214 8.051
R292 VDD.n88 VDD.n85 6.193
R293 VDD.n143 VDD.n140 6.193
R294 VDD.n28 VDD.n23 4.795
R295 VDD.n28 VDD.n27 4.65
R296 VDD.n32 VDD.n31 4.65
R297 VDD.n37 VDD.n36 4.65
R298 VDD.n41 VDD.n40 4.65
R299 VDD.n68 VDD.n67 4.65
R300 VDD.n72 VDD.n71 4.65
R301 VDD.n76 VDD.n75 4.65
R302 VDD.n79 VDD.n78 4.65
R303 VDD.n83 VDD.n82 4.65
R304 VDD.n89 VDD.n88 4.65
R305 VDD.n93 VDD.n92 4.65
R306 VDD.n97 VDD.n96 4.65
R307 VDD.n123 VDD.n122 4.65
R308 VDD.n127 VDD.n126 4.65
R309 VDD.n131 VDD.n130 4.65
R310 VDD.n134 VDD.n133 4.65
R311 VDD.n138 VDD.n137 4.65
R312 VDD.n144 VDD.n143 4.65
R313 VDD.n148 VDD.n147 4.65
R314 VDD.n317 VDD.n316 4.65
R315 VDD.n291 VDD.n290 4.65
R316 VDD.n287 VDD.n286 4.65
R317 VDD.n282 VDD.n281 4.65
R318 VDD.n278 VDD.n277 4.65
R319 VDD.n273 VDD.n272 4.65
R320 VDD.n247 VDD.n246 4.65
R321 VDD.n243 VDD.n242 4.65
R322 VDD.n238 VDD.n237 4.65
R323 VDD.n234 VDD.n233 4.65
R324 VDD.n229 VDD.n228 4.65
R325 VDD.n202 VDD.n201 4.65
R326 VDD.n198 VDD.n197 4.65
R327 VDD.n193 VDD.n192 4.65
R328 VDD.n189 VDD.n188 4.65
R329 VDD.n184 VDD.n183 4.65
R330 VDD.n180 VDD.n179 4.65
R331 VDD.n176 VDD.n175 4.65
R332 VDD.n171 VDD.n170 4.65
R333 VDD.n175 VDD.n172 2.89
R334 VDD.n80 �+��r 2.557
R335 VDD.n135  ,��r 2.557
R336 VDD.n181 �w˶U 2.557
R337 VDD.n197 VDD.n194 2.477
R338 VDD.n27 VDD.n24 2.064
R339 VDD.n36 VDD.n35 2.064
R340 VDD.n286 VDD.n283 2.064
R341 VDD.n277 VDD.n274 2.064
R342 VDD.n242 VDD.n239 2.064
R343 VDD.n233 VDD.n232 2.064
R344 VDD.n68 VDD.n41 0.29
R345 VDD.n123 VDD.n97 0.29
R346 VDD.n317 VDD.n291 0.29
R347 VDD.n273 VDD.n247 0.29
R348 VDD.n229 VDD.n202 0.29
R349 VDD.n171 VDD 0.207
R350 VDD.n83 VDD.n79 0.181
R351 VDD.n138 VDD.n134 0.181
R352 VDD.n189 VDD.n184 0.181
R353 VDD.n32 VDD.n28 0.157
R354 VDD.n37 VDD.n32 0.157
R355 VDD.n287 VDD.n282 0.157
R356 VDD.n282 VDD.n278 0.157
R357 VDD.n243 VDD.n238 0.157
R358 VDD.n238 VDD.n234 0.157
R359 VDD.n41 VDD.n37 0.145
R360 VDD.n72 VDD.n68 0.145
R361 VDD.n76 VDD.n72 0.145
R362 VDD.n79 VDD.n76 0.145
R363 VDD.n89 VDD.n83 0.145
R364 VDD.n93 VDD.n89 0.145
R365 VDD.n97 VDD.n93 0.145
R366 VDD.n127 VDD.n123 0.145
R367 VDD.n131 VDD.n127 0.145
R368 VDD.n134 VDD.n131 0.145
R369 VDD.n144 VDD.n138 0.145
R370 VDD.n148 VDD.n144 0.145
R371 VDD.n291 VDD.n287 0.145
R372 VDD.n278 VDD.n273 0.145
R373 VDD.n247 VDD.n243 0.145
R374 VDD.n234 VDD.n229 0.145
R375 VDD.n202 VDD.n198 0.145
R376 VDD.n198 VDD.n193 0.145
R377 VDD.n193 VDD.n189 0.145
R378 VDD.n184 VDD.n180 0.145
R379 VDD.n180 VDD.n176 0.145
R380 VDD.n176 VDD.n171 0.145
R381 VDD VDD.n317 0.078
R382 VDD VDD.n148 0.066
R383 COUT.n5 COUT.n0 299.141
R384 COUT.n5 COUT.n4 244.592
R385 COUT.n4 COUT.n3 30
R386 COUT.n2 COUT.n1 24.383
R387 COUT.n4 COUT.n2 23.684
R388 COUT.n0 COUT.t1 14.282
R389 COUT.n0 COUT.t2 14.282
R390 COUT.n6 COUT.n5 4.65
R391 COUT.n6 COUT 0.046
R392 a_1295_209.n0 a_1295_209.t3 477.179
R393 a_1295_209.n0 a_1295_209.t5 406.485
R394 a_1295_209.n1 a_1295_209.t4 341.566
R395 a_1295_209.n6 a_1295_209.n5 272.451
R396 a_1295_209.n7 a_1295_209.n6 271.281
R397 a_1295_209.n1 a_1295_209.n0 199.524
R398 a_1295_209.n5 a_1295_209.n4 30
R399 a_1295_209.n3 a_1295_209.n2 24.383
R400 a_1295_209.n5 a_1295_209.n3 23.684
R401 a_1295_209.n7 a_1295_209.t1 14.282
R402 a_1295_209.t2 a_1295_209.n7 14.282
R403 a_1295_209.n6 a_1295_209.n1 13.879
R404 B.n0 B.t6 512.525
R405 B.n3 B.t5 480.392
R406 B.n5 B.t1 472.359
R407 B.n3 B.t8 403.272
R408 B.n5 B.t4 384.527
R409 B.n0 B.t3 371.139
R410 B.n6 B.t7 314.896
R411 B.n1 B.t0 299.455
R412 B.n1 B.t2 227.134
R413 B.n6 B.n5 182.814
R414 B.n2 B.n0 163.771
R415 B.n2 B.n1 139.294
R416 B.n4 B.n3 120.597
R417 B.n7 B.n4 72.544
R418 B.n4 B.n2 7.325
R419 B.n7 B.n6 4.65
R420 B.n7 B 0.046
R421 a_1666_101.t0 a_1666_101.n1 93.333
R422 a_1666_101.n4 a_1666_101.n2 79.092
R423 a_1666_101.t0 a_1666_101.n0 8.137
R424 a_1666_101.n4 a_1666_101.n3 4.614
R425 a_1666_101.t0 a_1666_101.n4 0.111
R426 SUM.n8 SUM.n7 327.32
R427 SUM.n5 SUM.n4 305.581
R428 SUM.n5 SUM.n0 260.107
R429 SUM.n8 SUM.n6 260.107
R430 SUM.n4 SUM.n3 30
R431 SUM.n2 SUM.n1 24.383
R432 SUM.n4 SUM.n2 23.684
R433 SUM.n0 SUM.t5 14.282
R434 SUM.n0 SUM.t3 14.282
R435 SUM.n6 SUM.t0 14.282
R436 SUM.n6 SUM.t1 14.282
R437 SUM SUM.n8 7.007
R438 SUM.n9 SUM.n5 4.65
R439 SUM.n9 SUM 0.046
R440 GND.n116 GND.n115 237.558
R441 GND.n149 GND.n148 237.558
R442 GND.n61 GND.n60 237.558
R443 GND.n182 GND.n181 237.558
R444 GND.n31 GND.n30 237.558
R445 GND.n28 GND.n27 210.82
R446 GND.n118 GND.n117 210.82
R447 GND.n151 GND.n150 210.82
R448 GND.n184 GND.n183 210.82
R449 GND.n58 GND.n57 210.82
R450 GND.n47 GND.n46 172.612
R451 GND.n79 GND.n78 166.605
R452 GND.n96 GND.n95 151.605
R453 GND.n12 GND.n11 92.5
R454 GND.n3 GND.t2 45.414
R455 GND.n19 GND.n18 40.414
R456 GND.n3 GND.n2 39.307
R457 GND.n162 GND.n161 37.582
R458 GND.n129 GND.n128 37.582
R459 GND.t4 GND.n159 32.601
R460 GND.t3 GND.n126 32.601
R461 GND.n95 GND.n94 28.421
R462 GND.n95 GND.n93 25.263
R463 GND.n93 GND.n92 24.383
R464 GND.n20 GND.n19 23.961
R465 GND.n4 GND.n3 23.77
R466 GND.n78 GND.n76 23.03
R467 GND.n159 GND.n158 21.734
R468 GND.n126 GND.n125 21.734
R469 GND.n5 GND.n4 20.705
R470 GND.n14 GND.n13 20.705
R471 GND.n21 GND.n20 20.705
R472 GND.n174 GND.n173 20.705
R473 GND.n168 GND.n167 20.705
R474 GND.n163 GND.n162 20.705
R475 GND.n141 GND.n140 20.705
R476 GND.n135 GND.n134 20.705
R477 GND.n130 GND.n129 20.705
R478 GND.n173 GND.n172 19.952
R479 GND.n140 GND.n139 19.952
R480 GND.n29 GND.n28 18.953
R481 GND.n119 GND.n118 18.953
R482 GND.n152 GND.n151 18.953
R483 GND.n185 GND.n184 18.953
R484 GND.n59 GND.n58 18.953
R485 GND.n161 GND.t4 15.644
R486 GND.n128 GND.t3 15.644
R487 GND.n32 GND.n29 14.864
R488 GND.n62 GND.n59 14.864
R489 GND.n186 GND.n185 14.864
R490 GND.n153 GND.n152 14.864
R491 GND.n120 GND.n119 14.864
R492 GND.n161 GND.n160 13.541
R493 GND.n128 GND.n127 13.541
R494 GND.n90 GND.n89 9.154
R495 GND.n98 GND.n97 9.154
R496 GND.n101 GND.n100 9.154
R497 GND.n104 GND.n103 9.154
R498 GND.n107 GND.n106 9.154
R499 GND.n110 GND.n109 9.154
R500 GND.n113 GND.n112 9.154
R501 GND.n120 GND.n116 9.154
R502 GND.n131 GND.n122 9.154
R503 GND.n137 GND.n136 9.154
R504 GND.n143 GND.n142 9.154
R505 GND.n146 GND.n145 9.154
R506 GND.n153 GND.n149 9.154
R507 GND.n164 GND.n155 9.154
R508 GND.n170 GND.n169 9.154
R509 GND.n176 GND.n175 9.154
R510 GND.n179 GND.n178 9.154
R511 GND.n186 GND.n182 9.154
R512 GND.n84 GND.n83 9.154
R513 GND.n81 GND.n80 9.154
R514 GND.n74 GND.n73 9.154
R515 GND.n71 GND.n70 9.154
R516 GND.n68 GND.n67 9.154
R517 GND.n65 GND.n64 9.154
R518 GND.n62 GND.n61 9.154
R519 GND.n55 GND.n54 9.154
R520 GND.n52 GND.n51 9.154
R521 GND.n49 GND.n48 9.154
R522 GND.n44 GND.n43 9.154
R523 GND.n41 GND.n40 9.154
R524 GND.n38 GND.n37 9.154
R525 GND.n35 GND.n34 9.154
R526 GND.n32 GND.n31 9.154
R527 GND.n25 GND.n24 9.154
R528 GND.n22 GND.n17 9.154
R529 GND.n15 GND.n9 9.154
R530 GND.n7 GND.n6 9.154
R531 GND.n78 GND.n77 8.128
R532 GND.n8 GND.n1 4.795
R533 GND.n88 GND.n87 4.65
R534 GND.n8 GND.n7 4.65
R535 GND.n16 GND.n15 4.65
R536 GND.n23 GND.n22 4.65
R537 GND.n26 GND.n25 4.65
R538 GND.n33 GND.n32 4.65
R539 GND.n36 GND.n35 4.65
R540 GND.n39 GND.n38 4.65
R541 GND.n42 GND.n41 4.65
R542 GND.n45 GND.n44 4.65
R543 GND.n50 GND.n49 4.65
R544 GND.n53 GND.n52 4.65
R545 GND.n56 GND.n55 4.65
R546 GND.n63 GND.n62 4.65
R547 GND.n66 GND.n65 4.65
R548 GND.n69 GND.n68 4.65
R549 GND.n72 GND.n71 4.65
R550 GND.n75 GND.n74 4.65
R551 GND.n82 GND.n81 4.65
R552 GND.n85 GND.n84 4.65
R553 GND.n187 GND.n186 4.65
R554 GND.n180 GND.n179 4.65
R555 GND.n177 GND.n176 4.65
R556 GND.n171 GND.n170 4.65
R557 GND.n165 GND.n164 4.65
R558 GND.n154 GND.n153 4.65
R559 GND.n147 GND.n146 4.65
R560 GND.n144 GND.n143 4.65
R561 GND.n138 GND.n137 4.65
R562 GND.n132 GND.n131 4.65
R563 GND.n121 GND.n120 4.65
R564 GND.n114 GND.n113 4.65
R565 GND.n111 GND.n110 4.65
R566 GND.n108 GND.n107 4.65
R567 GND.n105 GND.n104 4.65
R568 GND.n102 GND.n101 4.65
R569 GND.n99 GND.n98 4.65
R570 GND.n91 GND.n90 4.65
R571 GND.n157 GND.n156 4.504
R572 GND.n124 GND.n123 4.504
R573 GND.n22 GND.n21 4.129
R574 GND.n49 GND.n47 4.129
R575 GND.n81 GND.n79 4.129
R576 GND.n176 GND.n174 4.129
R577 GND.n143 GND.n141 4.129
R578 GND.n98 GND.n96 4.129
R579 GND.n7 GND.n5 3.716
R580 GND.n164 GND.n163 3.716
R581 GND.n131 GND.n130 3.716
R582 GND.t4 GND.n157 2.452
R583 GND.t3 GND.n124 2.452
R584 GND.n11 GND.n10 1.935
R585 GND.n1 GND.n0 0.474
R586 GND.n87 GND.n86 0.474
R587 GND.n13 GND.n12 0.376
R588 GND.n167 GND.n166 0.376
R589 GND.n134 GND.n133 0.376
R590 GND.n33 GND.n26 0.29
R591 GND.n63 GND.n56 0.29
R592 GND.n187 GND.n180 0.29
R593 GND.n154 GND.n147 0.29
R594 GND.n121 GND.n114 0.29
R595 GND.n88 GND 0.207
R596 GND.n15 GND.n14 0.206
R597 GND.n170 GND.n168 0.206
R598 GND.n137 GND.n135 0.206
R599 GND.n45 GND.n42 0.181
R600 GND.n75 GND.n72 0.181
R601 GND.n105 GND.n102 0.181
R602 GND.n16 GND.n8 0.157
R603 GND.n23 GND.n16 0.157
R604 GND.n177 GND.n171 0.157
R605 GND.n171 GND.n165 0.157
R606 GND.n144 GND.n138 0.157
R607 GND.n138 GND.n132 0.157
R608 GND.n26 GND.n23 0.145
R609 GND.n36 GND.n33 0.145
R610 GND.n39 GND.n36 0.145
R611 GND.n42 GND.n39 0.145
R612 GND.n50 GND.n45 0.145
R613 GND.n53 GND.n50 0.145
R614 GND.n56 GND.n53 0.145
R615 GND.n66 GND.n63 0.145
R616 GND.n69 GND.n66 0.145
R617 GND.n72 GND.n69 0.145
R618 GND.n82 GND.n75 0.145
R619 GND.n85 GND.n82 0.145
R620 GND.n180 GND.n177 0.145
R621 GND.n165 GND.n154 0.145
R622 GND.n147 GND.n144 0.145
R623 GND.n132 GND.n121 0.145
R624 GND.n114 GND.n111 0.145
R625 GND.n111 GND.n108 0.145
R626 GND.n108 GND.n105 0.145
R627 GND.n102 GND.n99 0.145
R628 GND.n99 GND.n91 0.145
R629 GND.n91 GND.n88 0.145
R630 GND GND.n187 0.078
R631 GND GND.n85 0.066
R632 a_1917_990.n0 a_1917_990.t5 477.179
R633 a_1917_990.n0 a_1917_990.t4 406.485
R634 a_1917_990.n4 a_1917_990.t3 312.917
R635 a_1917_990.n4 a_1917_990.n3 260.115
R636 a_1917_990.n6 a_1917_990.n5 215.563
R637 a_1917_990.n5 a_1917_990.n0 156.869
R638 a_1917_990.n5 a_1917_990.n4 83.576
R639 a_1917_990.n3 a_1917_990.n2 22.578
R640 a_1917_990.t2 a_1917_990.n6 14.282
R641 a_1917_990.n6 a_1917_990.t1 14.282
R642 a_1917_990.n3 a_1917_990.n1 8.58
R643 a_2332_101.n11 a_2332_101.n10 68.43
R644 a_2332_101.n3 a_2332_101.n2 62.817
R645 a_2332_101.n7 a_2332_101.n6 38.626
R646 a_2332_101.n6 a_2332_101.n5 35.955
R647 a_2332_101.n3 a_2332_101.n1 26.202
R648 a_2332_101.t0 a_2332_101.n3 19.737
R649 a_2332_101.t1 a_2332_101.n8 8.137
R650 a_2332_101.t0 a_2332_101.n4 7.273
R651 a_2332_101.t0 a_2332_101.n0 6.109
R652 a_2332_101.t1 a_2332_101.n7 4.864
R653 a_2332_101.t0 a_2332_101.n12 2.074
R654 a_2332_101.n12 a_2332_101.t1 0.937
R655 a_2332_101.t1 a_2332_101.n11 0.763
R656 a_2332_101.n11 a_2332_101.n9 0.185
R657 a_2351_1051.n0 a_2351_1051.t2 228.369
R658 a_2351_1051.n0 a_2351_1051.t0 219.778
R659 a_2351_1051.n1 a_2351_1051.n0 42.29
R660 a_2351_1051.n1 a_2351_1051.t3 14.282
R661 a_2351_1051.t1 a_2351_1051.n1 14.282
R662 a_1685_1051.t1 a_1685_1051.n1 228.371
R663 a_1685_1051.n1 a_1685_1051.t3 219.777
R664 a_1685_1051.n1 a_1685_1051.n0 42.29
R665 a_1685_1051.n0 a_1685_1051.t0 14.282
R666 a_1685_1051.n0 a_1685_1051.t2 14.282
R667 a_112_101.n3 a_112_101.n1 42.788
R668 a_112_101.t0 a_112_101.n0 8.137
R669 a_112_101.n3 a_112_101.n2 4.665
R670 a_112_101.t0 a_112_101.n3 0.06
C9 VDD GND 5.85fF
C10 a_112_101.n0 GND 0.05fF
C11 a_112_101.n1 GND 0.11fF
C12 a_112_101.n2 GND 0.04fF
C13 a_112_101.n3 GND 0.16fF
C14 a_1685_1051.n0 GND 0.22fF
C15 a_1685_1051.n1 GND 0.50fF
C16 a_2351_1051.n0 GND 0.50fF
C17 a_2351_1051.n1 GND 0.22fF
C18 a_2332_101.n0 GND 0.02fF
C19 a_2332_101.n1 GND 0.09fF
C20 a_2332_101.n2 GND 0.08fF
C21 a_2332_101.n3 GND 0.03fF
C22 a_2332_101.n4 GND 0.01fF
C23 a_2332_101.n5 GND 0.04fF
C24 a_2332_101.n6 GND 0.04fF
C25 a_2332_101.n7 GND 0.02fF
C26 a_2332_101.n8 GND 0.05fF
C27 a_2332_101.n9 GND 0.15fF
C28 a_2332_101.n10 GND 0.08fF
C29 a_2332_101.n11 GND 0.08fF
C30 a_2332_101.n12 GND 0.01fF
C31 a_1917_990.n0 GND 0.58fF
C32 a_1917_990.n1 GND 0.07fF
C33 a_1917_990.n2 GND 0.09fF
C34 a_1917_990.n3 GND 0.29fF
C35 a_1917_990.n4 GND 1.80fF
C36 a_1917_990.n5 GND 2.26fF
C37 a_1917_990.n6 GND 0.94fF
C38 SUM.n0 GND 0.91fF
C39 SUM.n1 GND 0.07fF
C40 SUM.n2 GND 0.09fF
C41 SUM.n3 GND 0.06fF
C42 SUM.n4 GND 0.37fF
C43 SUM.n5 GND 1.05fF
C44 SUM.n6 GND 0.91fF
C45 SUM.n7 GND 0.56fF
C46 SUM.n8 GND 1.24fF
C47 SUM.n9 GND 0.05fF
C48 a_1666_101.n0 GND 0.05fF
C49 a_1666_101.n1 GND 0.02fF
C50 a_1666_101.n2 GND 0.12fF
C51 a_1666_101.n3 GND 0.04fF
C52 a_1666_101.n4 GND 0.17fF
C53 a_1295_209.n0 GND 0.52fF
C54 a_1295_209.n1 GND 1.42fF
C55 a_1295_209.n2 GND 0.06fF
C56 a_1295_209.n3 GND 0.08fF
C57 a_1295_209.n4 GND 0.05fF
C58 a_1295_209.n5 GND 0.27fF
C59 a_1295_209.n6 GND 1.69fF
C60 a_1295_209.n7 GND 0.94fF
C61 VDD.n1 GND 0.03fF
C62 VDD.n2 GND 0.10fF
C63 VDD.n3 GND 0.03fF
C64 VDD.n4 GND 0.02fF
C65 VDD.n5 GND 0.06fF
C66 VDD.n6 GND 0.02fF
C67 VDD.n7 GND 0.02fF
C68 VDD.n8 GND 0.02fF
C69 VDD.n9 GND 0.02fF
C70 VDD.n10 GND 0.02fF
C71 VDD.n11 GND 0.02fF
C72 VDD.n12 GND 0.02fF
C73 VDD.n13 GND 0.02fF
C74 VDD.n14 GND 0.03fF
C75 VDD.n15 GND 0.01fF
C76 VDD.n20 GND 0.44fF
C77 VDD.n21 GND 0.26fF
C78 VDD.n22 GND 0.02fF
C79 VDD.n23 GND 0.03fF
C80 VDD.n24 GND 0.06fF
C81 VDD.n25 GND 0.19fF
C82 VDD.n26 GND 0.01fF
C83 VDD.n27 GND 0.01fF
C84 VDD.n28 GND 0.06fF
C85 VDD.n29 GND 0.16fF
C86 VDD.n30 GND 0.01fF
C87 VDD.n31 GND 0.02fF
C88 VDD.n32 GND 0.02fF
C89 VDD.n33 GND 0.19fF
C90 VDD.n34 GND 0.01fF
C91 VDD.n35 GND 0.06fF
C92 VDD.n36 GND 0.01fF
C93 VDD.n37 GND 0.02fF
C94 VDD.n38 GND 0.26fF
C95 VDD.n39 GND 0.01fF
C96 VDD.n40 GND 0.02fF
C97 VDD.n41 GND 0.03fF
C98 VDD.n42 GND 0.05fF
C99 VDD.n43 GND 0.02fF
C100 VDD.n44 GND 0.02fF
C101 VDD.n45 GND 0.02fF
C102 VDD.n46 GND 0.02fF
C103 VDD.n47 GND 0.02fF
C104 VDD.n48 GND 0.02fF
C105 VDD.n49 GND 0.02fF
C106 VDD.n50 GND 0.02fF
C107 VDD.n51 GND 0.02fF
C108 VDD.n52 GND 0.02fF
C109 VDD.n53 GND 0.02fF
C110 VDD.n54 GND 0.03fF
C111 VDD.n55 GND 0.02fF
C112 VDD.n56 GND 0.17fF
C113 VDD.n57 GND 0.02fF
C114 VDD.n58 GND 0.02fF
C115 VDD.n60 GND 0.02fF
C116 VDD.n64 GND 0.26fF
C117 VDD.n65 GND 0.26fF
C118 VDD.n66 GND 0.01fF
C119 VDD.n67 GND 0.02fF
C120 VDD.n68 GND 0.03fF
C121 VDD.n69 GND 0.23fF
C122 VDD.n70 GND 0.01fF
C123 VDD.n71 GND 0.02fF
C124 VDD.n72 GND 0.02fF
C125 VDD.n73 GND 0.16fF
C126 VDD.n74 GND 0.01fF
C127 VDD.n75 GND 0.02fF
C128 VDD.n76 GND 0.02fF
C129 VDD.n77 GND 0.01fF
C130 VDD.n78 GND 0.02fF
C131 VDD.n79 GND 0.02fF
C132 VDD.n80 GND 0.13fF
C133 VDD.n81 GND 0.01fF
C134 VDD.n82 GND 0.02fF
C135 VDD.n83 GND 0.02fF
C136 VDD.n84 GND 0.07fF
C137 VDD.n85 GND 0.05fF
C138 VDD.n86 GND 0.16fF
C139 VDD.n87 GND 0.01fF
C140 VDD.n88 GND 0.02fF
C141 VDD.n89 GND 0.02fF
C142 VDD.n90 GND 0.24fF
C143 VDD.n91 GND 0.01fF
C144 VDD.n92 GND 0.02fF
C145 VDD.n93 GND 0.02fF
C146 VDD.n94 GND 0.26fF
C147 VDD.n95 GND 0.01fF
C148 VDD.n96 GND 0.02fF
C149 VDD.n97 GND 0.03fF
C150 VDD.n98 GND 0.20fF
C151 VDD.n99 GND 0.02fF
C152 VDD.n100 GND 0.02fF
C153 VDD.n101 GND 0.02fF
C154 VDD.n102 GND 0.06fF
C155 VDD.n103 GND 0.02fF
C156 VDD.n104 GND 0.02fF
C157 VDD.n105 GND 0.02fF
C158 VDD.n106 GND 0.02fF
C159 VDD.n107 GND 0.02fF
C160 VDD.n108 GND 0.02fF
C161 VDD.n109 GND 0.02fF
C162 VDD.n110 GND 0.02fF
C163 VDD.n111 GND 0.02fF
C164 VDD.n112 GND 0.02fF
C165 VDD.n113 GND 0.03fF
C166 VDD.n114 GND 0.02fF
C167 VDD.n115 GND 0.02fF
C168 VDD.n119 GND 0.26fF
C169 VDD.n120 GND 0.26fF
C170 VDD.n121 GND 0.01fF
C171 VDD.n122 GND 0.02fF
C172 VDD.n123 GND 0.03fF
C173 VDD.n124 GND 0.23fF
C174 VDD.n125 GND 0.01fF
C175 VDD.n126 GND 0.02fF
C176 VDD.n127 GND 0.02fF
C177 VDD.n128 GND 0.16fF
C178 VDD.n129 GND 0.01fF
C179 VDD.n130 GND 0.02fF
C180 VDD.n131 GND 0.02fF
C181 VDD.n132 GND 0.01fF
C182 VDD.n133 GND 0.02fF
C183 VDD.n134 GND 0.02fF
C184 VDD.n135 GND 0.13fF
C185 VDD.n136 GND 0.01fF
C186 VDD.n137 GND 0.02fF
C187 VDD.n138 GND 0.02fF
C188 VDD.n139 GND 0.07fF
C189 VDD.n140 GND 0.05fF
C190 VDD.n141 GND 0.16fF
C191 VDD.n142 GND 0.01fF
C192 VDD.n143 GND 0.02fF
C193 VDD.n144 GND 0.02fF
C194 VDD.n145 GND 0.24fF
C195 VDD.n146 GND 0.01fF
C196 VDD.n147 GND 0.02fF
C197 VDD.n148 GND 0.02fF
C198 VDD.n149 GND 0.13fF
C199 VDD.n150 GND 0.02fF
C200 VDD.n151 GND 0.02fF
C201 VDD.n152 GND 0.06fF
C202 VDD.n153 GND 0.02fF
C203 VDD.n154 GND 0.02fF
C204 VDD.n155 GND 0.02fF
C205 VDD.n156 GND 0.02fF
C206 VDD.n157 GND 0.02fF
C207 VDD.n158 GND 0.02fF
C208 VDD.n159 GND 0.02fF
C209 VDD.n160 GND 0.02fF
C210 VDD.n161 GND 0.03fF
C211 VDD.n162 GND 0.03fF
C212 VDD.n163 GND 0.02fF
C213 VDD.n167 GND 0.44fF
C214 VDD.n168 GND 0.26fF
C215 VDD.n169 GND 0.02fF
C216 VDD.n170 GND 0.03fF
C217 VDD.n171 GND 0.03fF
C218 VDD.n172 GND 0.06fF
C219 VDD.n173 GND 0.24fF
C220 VDD.n174 GND 0.01fF
C221 VDD.n175 GND 0.01fF
C222 VDD.n176 GND 0.02fF
C223 VDD.n177 GND 0.16fF
C224 VDD.n178 GND 0.01fF
C225 VDD.n179 GND 0.02fF
C226 VDD.n180 GND 0.02fF
C227 VDD.n181 GND 0.13fF
C228 VDD.n182 GND 0.01fF
C229 VDD.n183 GND 0.02fF
C230 VDD.n184 GND 0.02fF
C231 VDD.n185 GND 0.08fF
C232 VDD.n186 GND 0.05fF
C233 VDD.n187 GND 0.01fF
C234 VDD.n188 GND 0.02fF
C235 VDD.n189 GND 0.02fF
C236 VDD.n190 GND 0.16fF
C237 VDD.n191 GND 0.01fF
C238 VDD.n192 GND 0.02fF
C239 VDD.n193 GND 0.02fF
C240 VDD.n194 GND 0.06fF
C241 VDD.n195 GND 0.23fF
C242 VDD.n196 GND 0.01fF
C243 VDD.n197 GND 0.01fF
C244 VDD.n198 GND 0.02fF
C245 VDD.n199 GND 0.26fF
C246 VDD.n200 GND 0.01fF
C247 VDD.n201 GND 0.02fF
C248 VDD.n202 GND 0.03fF
C249 VDD.n203 GND 0.05fF
C250 VDD.n204 GND 0.02fF
C251 VDD.n205 GND 0.02fF
C252 VDD.n206 GND 0.02fF
C253 VDD.n207 GND 0.02fF
C254 VDD.n208 GND 0.02fF
C255 VDD.n209 GND 0.02fF
C256 VDD.n210 GND 0.02fF
C257 VDD.n211 GND 0.02fF
C258 VDD.n212 GND 0.02fF
C259 VDD.n213 GND 0.02fF
C260 VDD.n214 GND 0.02fF
C261 VDD.n215 GND 0.03fF
C262 VDD.n216 GND 0.02fF
C263 VDD.n219 GND 0.02fF
C264 VDD.n221 GND 0.02fF
C265 VDD.n222 GND 0.17fF
C266 VDD.n223 GND 0.02fF
C267 VDD.n225 GND 0.26fF
C268 VDD.n226 GND 0.26fF
C269 VDD.n227 GND 0.01fF
C270 VDD.n228 GND 0.02fF
C271 VDD.n229 GND 0.03fF