magic
tech sky130A
magscale 1 2
timestamp 1647327697
<< nmos >>
tri 146 222 162 238 se
rect 162 222 192 276
tri 56 192 86 222 se
rect 86 192 192 222
rect 56 92 86 192
tri 86 176 102 192 nw
tri 146 176 162 192 ne
tri 86 92 102 108 sw
tri 146 92 162 108 se
rect 162 92 192 192
tri 56 62 86 92 ne
rect 86 62 162 92
tri 162 62 192 92 nw
<< ndiff >>
rect 0 238 162 276
rect 0 222 146 238
tri 146 222 162 238 nw
rect 0 189 56 222
tri 56 192 86 222 nw
rect 0 155 10 189
rect 44 155 56 189
rect 0 121 56 155
rect 0 87 10 121
rect 44 87 56 121
tri 86 176 102 192 se
rect 102 176 146 192
tri 146 176 162 192 sw
rect 86 144 162 176
rect 86 110 107 144
rect 141 110 162 144
rect 86 108 162 110
tri 86 92 102 108 ne
rect 102 92 146 108
tri 146 92 162 108 nw
rect 192 189 248 276
rect 192 155 204 189
rect 238 155 248 189
rect 192 121 248 155
rect 0 62 56 87
tri 56 62 86 92 sw
tri 162 62 192 92 se
rect 192 87 204 121
rect 238 87 248 121
rect 192 62 248 87
rect 0 50 248 62
rect 0 16 10 50
rect 44 16 107 50
rect 141 16 204 50
rect 238 16 248 50
rect 0 0 248 16
<< ndiffc >>
rect 10 155 44 189
rect 10 87 44 121
rect 107 110 141 144
rect 204 155 238 189
rect 204 87 238 121
rect 10 16 44 50
rect 107 16 141 50
rect 204 16 238 50
<< poly >>
rect 162 276 192 309
<< locali >>
rect 10 189 44 205
rect 204 189 238 205
rect 10 121 44 155
rect 107 144 141 160
rect 107 94 141 110
rect 204 121 238 155
rect 10 50 44 87
rect 204 50 238 87
rect 44 16 107 50
rect 141 16 204 50
rect 10 0 44 16
rect 204 0 238 16
<< end >>
