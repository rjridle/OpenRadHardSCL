* HSPICE file created from tmp.ext - technology: sky130A

.option scale=5000u

.subckt tmp CLK SN Q QN D VDD VSS
X0 VDD a_217_1051 a_1905_1051 VDD sky130_fd_pr__pfet_01v8 ad=236400 pd=9582 as=0 ps=0 w=400 l=30 M=2
X1 a_343_411 a_217_1051 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=400 l=30 M=2
X2 a_1265_990 CLK VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=400 l=30 M=2
X3 VDD a_343_411 QN VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=23200 ps=916 w=400 l=30 M=2
X4 VSS CLK a_2702_101 VSS sky130_fd_pr__nfet_01v8 ad=42528 pd=1872 as=0 ps=0 w=598 l=30
X5 a_1265_990 a_1905_1051 a_2702_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=598 l=30
X6 VDD a_1905_1051 a_1265_990 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=400 l=30 M=2
X7 a_343_411 a_1265_990 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=400 l=30 M=2
X8 VDD a_1265_990 a_1905_1051 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=400 l=30 M=2
X9 a_1905_1051 SN a_2000_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=598 l=30
X10 VDD a_1265_990 Q VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=34800 ps=1374 w=400 l=30 M=2
X11 Q QN a_3628_210 VSS sky130_fd_pr__nfet_01v8 ad=7088 pd=312 as=0 ps=0 w=598 l=30
X12 VDD D a_217_1051 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=400 l=30 M=2
X13 VDD SN a_1905_1051 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=400 l=30 M=2
X14 a_343_411 a_1265_990 a_1038_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=598 l=30
X15 VDD SN Q VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=400 l=30 M=2
X16 VDD QN Q VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=400 l=30 M=2
X17 a_3628_210 a_1265_990 a_3347_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=600 l=30
X18 VDD a_343_411 a_217_1051 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=400 l=30 M=2
X19 VDD CLK a_343_411 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=400 l=30 M=2
X20 QN Q VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=400 l=30 M=2
X21 VSS a_343_411 a_4330_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=598 l=30
X22 QN Q a_4330_101 VSS sky130_fd_pr__nfet_01v8 ad=7088 pd=312 as=0 ps=0 w=598 l=30
X23 a_1038_210 a_217_1051 a_757_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=600 l=30
X24 VSS CLK a_757_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=598 l=30
X25 VSS D a_112_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=598 l=30
X26 a_217_1051 a_343_411 a_112_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=598 l=30
X27 a_2000_210 a_1265_990 a_1719_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=600 l=30
X28 VSS SN a_3347_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=598 l=30
X29 VSS a_217_1051 a_1719_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=598 l=30
C0 a_343_411 VDD 3.15fF
C1 VDD CLK 2.46fF
C2 QN VDD 2.15fF
C3 a_1905_1051 VDD 2.83fF
C4 a_217_1051 VDD 2.51fF
C5 a_1265_990 VDD 2.71fF
C6 Q VDD 2.83fF
.ends

** hspice subcircuit dictionary
