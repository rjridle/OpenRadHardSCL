magic
tech sky130
magscale 1 2
timestamp 1651261323
<< nwell >>
rect 55 1505 89 1539
<< pwell >>
rect 55 13 89 47
<< metal1 >>
rect -31 1492 2251 1554
rect 131 871 165 905
rect 1611 723 1645 757
rect 2055 575 2089 609
rect -31 0 2251 62
use xnor2x1_pcell  xnor2x1_pcell_0 pcells
timestamp 1651260581
transform 1 0 0 0 1 0
box -84 0 2304 1575
use li1_M1_contact  li1_M1_contact_0 pcells
timestamp 1648061256
transform 1 0 2072 0 1 592
box -53 -33 29 33
<< labels >>
rlabel metal1 1611 723 1645 757 1 Y
port 1 nsew signal output
rlabel metal1 131 871 165 905 1 A
port 2 nsew signal input
rlabel metal1 2055 575 2089 609 1 B
port 3 nsew signal input
rlabel metal1 -31 1492 2251 1554 1 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 -31 0 2251 62 1 VGND
port 5 nsew ground bidirectional abutment
rlabel nwell 55 1505 89 1539 1 VPB
port 6 nsew power bidirectional
rlabel pwell 55 13 89 47 1 VNB
port 7 nsew ground bidirectional
<< end >>
