* SPICE3 file created from NAND2X1.ext - technology: sky130A

.subckt NAND2X1 Y A B VDD GND
X0 VDD.t3 A.t0 Y.t1 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X1 VDD.t7 B.t0 Y.t4  ��48 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X2 GND A.t1 a_112_101.t0 GND sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=0p ps=0u w=0u l=0u
X3 Y.t0 A.t2 VDD.t1 ���48 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X4 Y.t2 B.t1 VDD.t5  ��48 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X5 Y B.t2 a_112_101.t1 GND sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=0p ps=0u w=0u l=0u
C0 B Y 0.26fF
C1 B VDD 0.32fF
C2 B A 0.27fF
C3 Y VDD 1.82fF
C4 Y A 0.10fF
C5 A VDD 0.33fF
R0 A.n0 A.t0 480.392
R1 A.n0 A.t2 403.272
R2 A.n1 A.t1 385.063
R3 A.n1 A.n0 143.429
R4 A A.n1 4.65
R5 Y.n4 Y.n3 299.461
R6 Y.n4 Y.n2 187.858
R7 Y.n2 Y.n1 157.964
R8 Y.n2 Y.n0 91.706
R9 Y.n0 Y.t4 14.282
R10 Y.n0 Y.t2 14.282
R11 Y.n1 Y.t1 14.282
R12 Y.n1 Y.t0 14.282
R13 Y Y.n4 4.65
R14 VDD.n24 VDD.t7 143.754
R15 VDD.n62 VDD.t1 135.17
R16 VDD.n34 VDD.n33 129.472
R17 VDD.n47 VDD.n46 92.5
R18 VDD.n45 VDD.n44 92.5
R19 VDD.n43 VDD.n42 92.5
R20 VDD.n41 VDD.n40 92.5
R21 VDD.n49 VDD.n48 92.5
R22 VDD.n14 VDD.n1 92.5
R23 VDD.n5 VDD.n4 92.5
R24 VDD.n7 VDD.n6 92.5
R25 VDD.n9 VDD.n8 92.5
R26 VDD.n11 VDD.n10 92.5
R27 VDD.n13 VDD.n12 92.5
R28 VDD.n21 VDD.n20 92.059
R29 VDD.n58 VDD.n57 92.059
R30 VDD.n20 VDD.n16 67.194
R31 VDD.n20 VDD.n17 67.194
R32 VDD.n20 VDD.n18 67.194
R33 VDD.n20 VDD.n19 67.194
R34 VDD.n5 VDD.n3 44.141
R35 VDD.n3 VDD.n2 44.107
R36 VDD.n20 VDD.n15 41.052
R37 VDD.n56 VDD.n54 39.742
R38 VDD.n56 VDD.n55 39.742
R39 VDD.n53 VDD.n52 39.742
R40 VDD.n1 VDD.n0 30.923
R41 VDD.n57 VDD.n56 26.38
R42 VDD.n57 VDD.n53 26.38
R43 VDD.n57 VDD.n51 26.38
R44 VDD.n57 VDD.n50 26.38
R45 VDD.n60 VDD.n49 22.915
R46 VDD.n23 VDD.n14 22.915
R47 VDD.n29  ��48 20.457
R48 VDD.n67 ���48 17.9
R49 VDD.n49 VDD.n47 14.864
R50 VDD.n47 VDD.n45 14.864
R51 VDD.n45 VDD.n43 14.864
R52 VDD.n43 VDD.n41 14.864
R53 VDD.n41 VDD.n39 14.864
R54 VDD.n39 VDD.n38 14.864
R55 VDD.n14 VDD.n13 14.864
R56 VDD.n13 VDD.n11 14.864
R57 VDD.n11 VDD.n9 14.864
R58 VDD.n9 VDD.n7 14.864
R59 VDD.n7 VDD.n5 14.864
R60 VDD.n33 VDD.t5 14.282
R61 VDD.n33 VDD.t3 14.282
R62 VDD.n36 VDD.n34 9.083
R63 VDD.n23 VDD.n22 8.855
R64 VDD.n22 VDD.n21 8.855
R65 VDD.n27 VDD.n26 8.855
R66 VDD.n26 VDD.n25 8.855
R67 VDD.n31 VDD.n30 8.855
R68 VDD.n30 VDD.n29 8.855
R69 VDD.n36 VDD.n35 8.855
R70 VDD.n35  ��48 8.855
R71 VDD.n73 VDD.n72 8.855
R72 VDD.n72 VDD.n71 8.855
R73 VDD.n69 VDD.n68 8.855
R74 VDD.n68 VDD.n67 8.855
R75 VDD.n65 VDD.n64 8.855
R76 VDD.n64 VDD.n63 8.855
R77 VDD.n60 VDD.n59 8.855
R78 VDD.n59 VDD.n58 8.855
R79 VDD.n32 VDD.n31 4.65
R80 VDD.n37 VDD.n36 4.65
R81 VDD.n74 VDD.n73 4.65
R82 VDD.n70 VDD.n69 4.65
R83 VDD.n66 VDD.n65 4.65
R84 VDD.n61 VDD.n60 4.65
R85 VDD.n28 VDD.n23 2.933
R86 VDD.n65 VDD.n62 2.89
R87 VDD.n28 VDD.n27 2.844
R88 VDD.n71 VDD.t2 2.557
R89 VDD.n27 VDD.n24 2.477
R90 VDD.n32 VDD.n28 1.063
R91 VDD.n61 VDD 0.207
R92 VDD.n37 VDD.n32 0.145
R93 VDD.n74 VDD.n70 0.145
R94 VDD.n70 VDD.n66 0.145
R95 VDD.n66 VDD.n61 0.145
R96 VDD VDD.n37 0.09
R97 VDD VDD.n74 0.09
R98 B.n0 B.t0 472.359
R99 B.n0 B.t1 384.527
R100 B.n1 B.t2 314.896
R101 B.n1 B.n0 182.814
R102 B B.n1 4.65
R103 a_112_101.n10 a_112_101.n9 93.333
R104 a_112_101.n12 a_112_101.n11 68.43
R105 a_112_101.n3 a_112_101.n2 51.907
R106 a_112_101.n3 a_112_101.n1 51.594
R107 a_112_101.t0 a_112_101.n3 38.864
R108 a_112_101.n7 a_112_101.n6 38.626
R109 a_112_101.n6 a_112_101.n5 35.955
R110 a_112_101.t1 a_112_101.n8 8.137
R111 a_112_101.t0 a_112_101.n0 6.109
R112 a_112_101.t1 a_112_101.n7 4.864
R113 a_112_101.t0 a_112_101.n4 3.871
R114 a_112_101.t0 a_112_101.n13 2.535
R115 a_112_101.n13 a_112_101.t1 1.145
R116 a_112_101.t1 a_112_101.n12 0.763
R117 a_112_101.n12 a_112_101.n10 0.185
R118 GND.n17 GND.n16 172.612
R119 GND.n14 GND.n13 9.154
R120 GND.n19 GND.n18 9.154
R121 GND.n22 GND.n21 9.154
R122 GND.n8 GND.n7 9.154
R123 GND.n5 GND.n4 9.154
R124 GND.n2 GND.n1 9.154
R125 GND.n12 GND.n11 4.65
R126 GND.