magic
tech sky130A
magscale 1 2
timestamp 1648248471
<< nwell >>
rect 84 1555 878 1575
rect 84 1501 904 1555
rect 84 1421 878 1501
rect 84 1408 316 1421
rect 317 1408 878 1421
rect 84 1376 878 1408
rect 84 1358 526 1376
rect 527 1358 878 1376
rect 84 903 878 1358
rect 83 832 878 903
<< pdiffc >>
rect 147 1377 181 1411
rect 235 1377 269 1411
rect 323 1377 357 1411
rect 411 1377 445 1413
rect 499 1377 533 1411
rect 235 1105 269 1139
rect 411 1105 445 1139
<< psubdiff >>
rect 31 571 635 572
rect 31 510 940 571
rect 31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 343 47
rect 377 13 415 47
rect 449 13 513 47
rect 547 13 585 47
rect 619 13 657 47
rect 691 13 729 47
rect 763 13 801 47
rect 835 13 873 47
rect 907 13 931 47
<< nsubdiff >>
rect 31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 343 1539
rect 377 1505 415 1539
rect 449 1505 513 1539
rect 547 1505 585 1539
rect 619 1505 657 1539
rect 691 1505 729 1539
rect 763 1505 801 1539
rect 835 1505 873 1539
rect 907 1505 931 1539
rect 31 868 931 930
<< psubdiffcont >>
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 343 13 377 47
rect 415 13 449 47
rect 513 13 547 47
rect 585 13 619 47
rect 657 13 691 47
rect 729 13 763 47
rect 801 13 835 47
rect 873 13 907 47
<< nsubdiffcont >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 343 1505 377 1539
rect 415 1505 449 1539
rect 513 1505 547 1539
rect 585 1505 619 1539
rect 657 1505 691 1539
rect 729 1505 763 1539
rect 801 1505 835 1539
rect 873 1505 907 1539
<< poly >>
rect 771 990 814 1020
rect 164 411 206 441
rect 164 403 194 411
rect 358 410 388 434
rect 768 403 798 441
<< locali >>
rect 31 1539 931 1554
rect 31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 343 1539
rect 377 1505 415 1539
rect 449 1505 513 1539
rect 547 1505 585 1539
rect 619 1505 657 1539
rect 691 1505 729 1539
rect 763 1505 801 1539
rect 835 1505 873 1539
rect 907 1505 931 1539
rect 31 1492 931 1505
rect 147 1411 181 1492
rect 147 1343 181 1377
rect 235 1411 269 1445
rect 235 1343 269 1377
rect 323 1411 357 1492
rect 323 1343 357 1377
rect 411 1413 445 1429
rect 411 1343 445 1377
rect 499 1411 533 1492
rect 499 1359 533 1377
rect 607 1411 817 1445
rect 607 1359 641 1411
rect 783 1359 817 1411
rect 235 1139 269 1158
rect 411 1139 445 1173
rect 607 1105 641 1167
rect 235 1071 641 1105
rect 695 1105 729 1164
rect 695 1071 757 1105
rect 205 461 239 954
rect 353 469 387 988
rect 353 461 357 469
rect 409 339 616 373
rect 723 361 757 1071
rect 797 461 831 970
rect 409 261 443 339
rect 215 62 249 195
rect 713 62 747 186
rect 31 47 931 62
rect 31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 343 47
rect 377 13 415 47
rect 449 13 513 47
rect 547 13 585 47
rect 619 13 657 47
rect 691 13 729 47
rect 763 13 801 47
rect 835 13 873 47
rect 907 13 931 47
rect 31 0 931 13
<< viali >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 343 1505 377 1539
rect 415 1505 449 1539
rect 513 1505 547 1539
rect 585 1505 619 1539
rect 657 1505 691 1539
rect 729 1505 763 1539
rect 801 1505 835 1539
rect 873 1505 907 1539
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 343 13 377 47
rect 415 13 449 47
rect 513 13 547 47
rect 585 13 619 47
rect 657 13 691 47
rect 729 13 763 47
rect 801 13 835 47
rect 873 13 907 47
<< metal1 >>
rect 31 1539 931 1554
rect 31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 343 1539
rect 377 1505 415 1539
rect 449 1505 513 1539
rect 547 1505 585 1539
rect 619 1505 657 1539
rect 691 1505 729 1539
rect 763 1505 801 1539
rect 835 1505 873 1539
rect 907 1505 931 1539
rect 31 1492 931 1505
rect 769 871 1062 905
rect 31 47 931 62
rect 31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 343 47
rect 377 13 415 47
rect 449 13 513 47
rect 547 13 585 47
rect 619 13 657 47
rect 691 13 729 47
rect 763 13 801 47
rect 835 13 873 47
rect 907 13 931 47
rect 31 0 931 13
use poly_li1_contact  poly_li1_contact_1
timestamp 1648060378
transform 0 1 223 -1 0 445
box -32 -28 34 26
use diff_ring_side  diff_ring_side_1
timestamp 1648063806
transform 1 0 0 0 1 0
box -84 0 84 1575
use poly_li1_contact  poly_li1_contact_0
timestamp 1648060378
transform 0 1 223 -1 0 988
box -32 -28 34 26
use pmos2_1  pmos2_1_0
timestamp 1647326732
transform 1 0 49 0 1 1450
box 52 -460 352 37
use nmos_bottom  nmos_bottom_0
timestamp 1648062456
transform -1 0 356 0 1 101
box 0 0 248 302
use poly_li1_contact  poly_li1_contact_2
timestamp 1648060378
transform 0 -1 369 1 0 443
box -32 -28 34 26
use pmos2_1  pmos2_1_1
timestamp 1647326732
transform 1 0 225 0 1 1450
box 52 -460 352 37
use poly_li1_contact  poly_li1_contact_3
timestamp 1648060378
transform 0 1 387 -1 0 988
box -32 -28 34 26
use nmos_top_trim1  nmos_top_trim1_0
timestamp 1648061897
transform -1 0 550 0 1 101
box 0 0 248 309
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform 1 0 1110 0 1 888
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform -1 0 740 0 -1 888
box -53 -33 29 33
use poly_li1_contact  poly_li1_contact_5
timestamp 1648060378
transform 0 -1 813 1 0 443
box -32 -28 34 26
use poly_li1_contact  poly_li1_contact_4
timestamp 1648060378
transform 0 1 815 -1 0 988
box -32 -28 34 26
use nmos_bottom  nmos_bottom_1
timestamp 1648062456
transform 1 0 606 0 1 101
box 0 0 248 302
use pmos2_1  pmos2_1_2
timestamp 1647326732
transform 1 0 509 0 1 1450
box 52 -460 352 37
use invx1_pcell  invx1_pcell_0
timestamp 1648064504
transform 1 0 962 0 1 0
box -84 0 528 1575
<< end >>
