magic
tech sky130A
magscale 1 2
timestamp 1643179348
<< nwell >>
rect -159 761 399 1355
rect -76 760 356 761
rect -20 758 356 760
<< ndiff >>
rect 102 270 136 291
<< psubdiff >>
rect -61 491 299 553
rect -61 13 -37 47
rect -3 13 31 47
rect 65 13 100 47
rect 134 13 174 47
rect 208 13 242 47
rect 276 13 299 47
<< nsubdiff >>
rect -61 1283 -44 1317
rect -10 1283 24 1317
rect 58 1283 92 1317
rect 126 1283 160 1317
rect 195 1283 229 1317
rect 264 1283 299 1317
rect -61 795 299 857
<< psubdiffcont >>
rect -37 13 -3 47
rect 31 13 65 47
rect 100 13 134 47
rect 174 13 208 47
rect 242 13 276 47
<< nsubdiffcont >>
rect -44 1283 -10 1317
rect 24 1283 58 1317
rect 92 1283 126 1317
rect 160 1283 195 1317
rect 229 1283 264 1317
<< poly >>
rect 44 915 93 945
rect 56 401 86 467
<< locali >>
rect -61 1317 299 1332
rect -61 1283 -44 1317
rect -10 1283 24 1317
rect 58 1283 92 1317
rect 126 1283 160 1317
rect 195 1283 229 1317
rect 264 1283 299 1317
rect -61 1270 299 1283
rect 14 1269 48 1270
rect 190 1269 224 1270
rect 102 270 136 1007
rect 10 62 44 101
rect 194 62 228 101
rect -61 47 299 62
rect -61 13 -37 47
rect -3 13 31 47
rect 65 13 100 47
rect 134 13 174 47
rect 208 13 242 47
rect 276 13 299 47
rect -61 0 299 13
<< viali >>
rect -44 1283 -10 1317
rect 24 1283 58 1317
rect 92 1283 126 1317
rect 160 1283 195 1317
rect 229 1283 264 1317
rect -37 13 -3 47
rect 31 13 65 47
rect 100 13 134 47
rect 174 13 208 47
rect 242 13 276 47
<< metal1 >>
rect -61 1317 299 1332
rect -61 1283 -44 1317
rect -10 1283 24 1317
rect 58 1283 92 1317
rect 126 1283 160 1317
rect 195 1283 229 1317
rect 264 1283 299 1317
rect -61 1270 299 1283
rect 16 471 50 889
rect 16 456 42 471
rect -61 47 299 62
rect -61 13 -37 47
rect -3 13 31 47
rect 65 13 100 47
rect 134 13 174 47
rect 208 13 242 47
rect 276 13 299 47
rect -61 0 299 13
use M1_M2_contact  M1_M2_contact_0 pcells
timestamp 1643168619
transform 1 0 -64 0 1 2
box 64 391 130 473
use M1_M2_contact  M1_M2_contact_1
timestamp 1643168619
transform 1 0 -64 0 1 480
box 64 391 130 473
use nmos_top_left  nmos_top_left_0 pcells
timestamp 1643177486
transform 1 0 45 0 1 165
box -45 -64 193 238
use pmos  pmos_0 pcells
timestamp 1643179034
transform 1 0 4 0 1 1227
box -36 -312 264 42
use diff_ring_side  diff_ring_side_0 ./pcells
timestamp 1643172873
transform 1 0 405 0 1 0
box -159 0 9 1353
use diff_ring_side  diff_ring_side_1
timestamp 1643172873
transform 1 0 -17 0 1 0
box -159 0 9 1353
<< labels >>
rlabel metal1 161 1325 161 1325 1 VDD
port 1 n
rlabel metal1 153 31 153 31 1 VSS
port 4 n
<< end >>
