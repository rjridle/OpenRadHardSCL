magic
tech sky130A
magscale 1 2
timestamp 1649530812
<< nwell >>
rect -84 832 1490 1575
<< nmos >>
rect 147 318 177 379
tri 177 318 193 334 sw
rect 447 318 477 379
rect 147 288 253 318
tri 253 288 283 318 sw
rect 147 187 177 288
tri 177 272 193 288 nw
tri 237 272 253 288 ne
tri 177 187 193 203 sw
tri 237 187 253 203 se
rect 253 187 283 288
tri 342 288 372 318 se
rect 372 288 477 318
rect 342 194 372 288
tri 372 272 388 288 nw
tri 431 272 447 288 ne
tri 372 194 388 210 sw
tri 431 194 447 210 se
rect 447 194 477 288
tri 147 157 177 187 ne
rect 177 157 253 187
tri 253 157 283 187 nw
tri 342 164 372 194 ne
rect 372 164 447 194
tri 447 164 477 194 nw
rect 649 326 679 379
tri 679 326 695 342 sw
rect 649 296 755 326
tri 755 296 785 326 sw
rect 649 195 679 296
tri 679 280 695 296 nw
tri 739 280 755 296 ne
tri 679 195 695 211 sw
tri 739 195 755 211 se
rect 755 195 785 296
tri 649 165 679 195 ne
rect 679 165 755 195
tri 755 165 785 195 nw
rect 1117 324 1147 377
tri 1147 324 1163 340 sw
rect 1117 294 1223 324
tri 1223 294 1253 324 sw
rect 1117 193 1147 294
tri 1147 278 1163 294 nw
tri 1207 278 1223 294 ne
tri 1147 193 1163 209 sw
tri 1207 193 1223 209 se
rect 1223 193 1253 294
tri 1117 163 1147 193 ne
rect 1147 163 1223 193
tri 1223 163 1253 193 nw
<< pmos >>
rect 247 1050 277 1450
rect 335 1050 365 1450
rect 423 1050 453 1450
rect 511 1050 541 1450
rect 599 1050 629 1450
rect 687 1050 717 1450
rect 1125 1050 1155 1450
rect 1213 1050 1243 1450
<< ndiff >>
rect 91 363 147 379
rect 91 329 101 363
rect 135 329 147 363
rect 91 291 147 329
rect 177 363 447 379
rect 177 334 198 363
tri 177 318 193 334 ne
rect 193 329 198 334
rect 232 329 295 363
rect 329 329 392 363
rect 426 329 447 363
rect 193 318 447 329
rect 477 363 533 379
rect 477 329 489 363
rect 523 329 533 363
rect 91 257 101 291
rect 135 257 147 291
tri 253 288 283 318 ne
rect 283 291 342 318
rect 91 223 147 257
rect 91 189 101 223
rect 135 189 147 223
rect 91 157 147 189
tri 177 272 193 288 se
rect 193 272 237 288
tri 237 272 253 288 sw
rect 177 238 253 272
rect 177 204 198 238
rect 232 204 253 238
rect 177 203 253 204
tri 177 187 193 203 ne
rect 193 187 237 203
tri 237 187 253 203 nw
rect 283 257 295 291
rect 329 257 342 291
tri 342 288 372 318 nw
rect 283 223 342 257
rect 283 189 295 223
rect 329 189 342 223
tri 372 272 388 288 se
rect 388 272 431 288
tri 431 272 447 288 sw
rect 372 244 447 272
rect 372 210 393 244
rect 427 210 447 244
tri 372 194 388 210 ne
rect 388 194 431 210
tri 431 194 447 210 nw
tri 147 157 177 187 sw
tri 253 157 283 187 se
rect 283 164 342 189
tri 342 164 372 194 sw
tri 447 164 477 194 se
rect 477 164 533 329
rect 283 157 533 164
rect 91 153 533 157
rect 91 119 101 153
rect 135 119 295 153
rect 329 119 392 153
rect 426 119 489 153
rect 523 119 533 153
rect 91 103 533 119
rect 593 363 649 379
rect 593 329 603 363
rect 637 329 649 363
rect 593 291 649 329
rect 679 342 841 379
tri 679 326 695 342 ne
rect 695 326 841 342
tri 755 296 785 326 ne
rect 593 257 603 291
rect 637 257 649 291
rect 593 223 649 257
rect 593 189 603 223
rect 637 189 649 223
tri 679 280 695 296 se
rect 695 280 739 296
tri 739 280 755 296 sw
rect 679 247 755 280
rect 679 213 700 247
rect 734 213 755 247
rect 679 211 755 213
tri 679 195 695 211 ne
rect 695 195 739 211
tri 739 195 755 211 nw
rect 785 291 841 326
rect 785 257 797 291
rect 831 257 841 291
rect 785 223 841 257
rect 593 165 649 189
tri 649 165 679 195 sw
tri 755 165 785 195 se
rect 785 189 797 223
rect 831 189 841 223
rect 785 165 841 189
rect 593 153 841 165
rect 593 119 603 153
rect 637 119 700 153
rect 734 119 797 153
rect 831 119 841 153
rect 593 103 841 119
rect 1061 361 1117 377
rect 1061 327 1071 361
rect 1105 327 1117 361
rect 1061 289 1117 327
rect 1147 361 1307 377
rect 1147 340 1265 361
tri 1147 324 1163 340 ne
rect 1163 327 1265 340
rect 1299 327 1307 361
rect 1163 324 1307 327
tri 1223 294 1253 324 ne
rect 1061 255 1071 289
rect 1105 255 1117 289
rect 1061 221 1117 255
rect 1061 187 1071 221
rect 1105 187 1117 221
tri 1147 278 1163 294 se
rect 1163 278 1207 294
tri 1207 278 1223 294 sw
rect 1147 245 1223 278
rect 1147 211 1167 245
rect 1201 211 1223 245
rect 1147 209 1223 211
tri 1147 193 1163 209 ne
rect 1163 193 1207 209
tri 1207 193 1223 209 nw
rect 1253 289 1307 324
rect 1253 255 1265 289
rect 1299 255 1307 289
rect 1253 221 1307 255
rect 1061 163 1117 187
tri 1117 163 1147 193 sw
tri 1223 163 1253 193 se
rect 1253 187 1265 221
rect 1299 187 1307 221
rect 1253 163 1307 187
rect 1061 151 1307 163
rect 1061 117 1071 151
rect 1105 117 1167 151
rect 1201 117 1265 151
rect 1299 117 1307 151
rect 1061 101 1307 117
<< pdiff >>
rect 191 1412 247 1450
rect 191 1378 201 1412
rect 235 1378 247 1412
rect 191 1344 247 1378
rect 191 1310 201 1344
rect 235 1310 247 1344
rect 191 1276 247 1310
rect 191 1242 201 1276
rect 235 1242 247 1276
rect 191 1208 247 1242
rect 191 1174 201 1208
rect 235 1174 247 1208
rect 191 1139 247 1174
rect 191 1105 201 1139
rect 235 1105 247 1139
rect 191 1050 247 1105
rect 277 1412 335 1450
rect 277 1378 289 1412
rect 323 1378 335 1412
rect 277 1344 335 1378
rect 277 1310 289 1344
rect 323 1310 335 1344
rect 277 1276 335 1310
rect 277 1242 289 1276
rect 323 1242 335 1276
rect 277 1208 335 1242
rect 277 1174 289 1208
rect 323 1174 335 1208
rect 277 1139 335 1174
rect 277 1105 289 1139
rect 323 1105 335 1139
rect 277 1050 335 1105
rect 365 1412 423 1450
rect 365 1378 377 1412
rect 411 1378 423 1412
rect 365 1344 423 1378
rect 365 1310 377 1344
rect 411 1310 423 1344
rect 365 1276 423 1310
rect 365 1242 377 1276
rect 411 1242 423 1276
rect 365 1208 423 1242
rect 365 1174 377 1208
rect 411 1174 423 1208
rect 365 1050 423 1174
rect 453 1412 511 1450
rect 453 1378 465 1412
rect 499 1378 511 1412
rect 453 1344 511 1378
rect 453 1310 465 1344
rect 499 1310 511 1344
rect 453 1276 511 1310
rect 453 1242 465 1276
rect 499 1242 511 1276
rect 453 1208 511 1242
rect 453 1174 465 1208
rect 499 1174 511 1208
rect 453 1139 511 1174
rect 453 1105 465 1139
rect 499 1105 511 1139
rect 453 1050 511 1105
rect 541 1412 599 1450
rect 541 1378 553 1412
rect 587 1378 599 1412
rect 541 1344 599 1378
rect 541 1310 553 1344
rect 587 1310 599 1344
rect 541 1276 599 1310
rect 541 1242 553 1276
rect 587 1242 599 1276
rect 541 1208 599 1242
rect 541 1174 553 1208
rect 587 1174 599 1208
rect 541 1050 599 1174
rect 629 1412 687 1450
rect 629 1378 641 1412
rect 675 1378 687 1412
rect 629 1344 687 1378
rect 629 1310 641 1344
rect 675 1310 687 1344
rect 629 1276 687 1310
rect 629 1242 641 1276
rect 675 1242 687 1276
rect 629 1208 687 1242
rect 629 1174 641 1208
rect 675 1174 687 1208
rect 629 1139 687 1174
rect 629 1105 641 1139
rect 675 1105 687 1139
rect 629 1050 687 1105
rect 717 1412 771 1450
rect 717 1378 729 1412
rect 763 1378 771 1412
rect 717 1344 771 1378
rect 717 1310 729 1344
rect 763 1310 771 1344
rect 717 1276 771 1310
rect 717 1242 729 1276
rect 763 1242 771 1276
rect 717 1208 771 1242
rect 717 1174 729 1208
rect 763 1174 771 1208
rect 717 1050 771 1174
rect 1069 1412 1125 1450
rect 1069 1378 1079 1412
rect 1113 1378 1125 1412
rect 1069 1344 1125 1378
rect 1069 1310 1079 1344
rect 1113 1310 1125 1344
rect 1069 1276 1125 1310
rect 1069 1242 1079 1276
rect 1113 1242 1125 1276
rect 1069 1208 1125 1242
rect 1069 1174 1079 1208
rect 1113 1174 1125 1208
rect 1069 1139 1125 1174
rect 1069 1105 1079 1139
rect 1113 1105 1125 1139
rect 1069 1050 1125 1105
rect 1155 1412 1213 1450
rect 1155 1378 1167 1412
rect 1201 1378 1213 1412
rect 1155 1344 1213 1378
rect 1155 1310 1167 1344
rect 1201 1310 1213 1344
rect 1155 1276 1213 1310
rect 1155 1242 1167 1276
rect 1201 1242 1213 1276
rect 1155 1208 1213 1242
rect 1155 1174 1167 1208
rect 1201 1174 1213 1208
rect 1155 1139 1213 1174
rect 1155 1105 1167 1139
rect 1201 1105 1213 1139
rect 1155 1050 1213 1105
rect 1243 1412 1297 1450
rect 1243 1378 1255 1412
rect 1289 1378 1297 1412
rect 1243 1344 1297 1378
rect 1243 1310 1255 1344
rect 1289 1310 1297 1344
rect 1243 1276 1297 1310
rect 1243 1242 1255 1276
rect 1289 1242 1297 1276
rect 1243 1208 1297 1242
rect 1243 1174 1255 1208
rect 1289 1174 1297 1208
rect 1243 1139 1297 1174
rect 1243 1105 1255 1139
rect 1289 1105 1297 1139
rect 1243 1050 1297 1105
<< ndiffc >>
rect 101 329 135 363
rect 198 329 232 363
rect 295 329 329 363
rect 392 329 426 363
rect 489 329 523 363
rect 101 257 135 291
rect 101 189 135 223
rect 198 204 232 238
rect 295 257 329 291
rect 295 189 329 223
rect 393 210 427 244
rect 101 119 135 153
rect 295 119 329 153
rect 392 119 426 153
rect 489 119 523 153
rect 603 329 637 363
rect 603 257 637 291
rect 603 189 637 223
rect 700 213 734 247
rect 797 257 831 291
rect 797 189 831 223
rect 603 119 637 153
rect 700 119 734 153
rect 797 119 831 153
rect 1071 327 1105 361
rect 1265 327 1299 361
rect 1071 255 1105 289
rect 1071 187 1105 221
rect 1167 211 1201 245
rect 1265 255 1299 289
rect 1265 187 1299 221
rect 1071 117 1105 151
rect 1167 117 1201 151
rect 1265 117 1299 151
<< pdiffc >>
rect 201 1378 235 1412
rect 201 1310 235 1344
rect 201 1242 235 1276
rect 201 1174 235 1208
rect 201 1105 235 1139
rect 289 1378 323 1412
rect 289 1310 323 1344
rect 289 1242 323 1276
rect 289 1174 323 1208
rect 289 1105 323 1139
rect 377 1378 411 1412
rect 377 1310 411 1344
rect 377 1242 411 1276
rect 377 1174 411 1208
rect 465 1378 499 1412
rect 465 1310 499 1344
rect 465 1242 499 1276
rect 465 1174 499 1208
rect 465 1105 499 1139
rect 553 1378 587 1412
rect 553 1310 587 1344
rect 553 1242 587 1276
rect 553 1174 587 1208
rect 641 1378 675 1412
rect 641 1310 675 1344
rect 641 1242 675 1276
rect 641 1174 675 1208
rect 641 1105 675 1139
rect 729 1378 763 1412
rect 729 1310 763 1344
rect 729 1242 763 1276
rect 729 1174 763 1208
rect 1079 1378 1113 1412
rect 1079 1310 1113 1344
rect 1079 1242 1113 1276
rect 1079 1174 1113 1208
rect 1079 1105 1113 1139
rect 1167 1378 1201 1412
rect 1167 1310 1201 1344
rect 1167 1242 1201 1276
rect 1167 1174 1201 1208
rect 1167 1105 1201 1139
rect 1255 1378 1289 1412
rect 1255 1310 1289 1344
rect 1255 1242 1289 1276
rect 1255 1174 1289 1208
rect 1255 1105 1289 1139
<< psubdiff >>
rect -31 546 1437 572
rect -31 512 -17 546
rect 17 512 945 546
rect 979 512 1389 546
rect 1423 512 1437 546
rect -31 510 1437 512
rect -31 474 31 510
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect -31 368 -17 402
rect 17 368 31 402
rect 931 474 993 510
rect 931 440 945 474
rect 979 440 993 474
rect 931 402 993 440
rect 1375 474 1437 510
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect 931 368 945 402
rect 979 368 993 402
rect 1375 440 1389 474
rect 1423 440 1437 474
rect 1375 402 1437 440
rect 931 330 993 368
rect 931 296 945 330
rect 979 296 993 330
rect 931 258 993 296
rect 931 224 945 258
rect 979 224 993 258
rect 931 186 993 224
rect 931 152 945 186
rect 979 152 993 186
rect 931 114 993 152
rect -31 47 31 80
rect 931 80 945 114
rect 979 80 993 114
rect 1375 368 1389 402
rect 1423 368 1437 402
rect 1375 330 1437 368
rect 1375 296 1389 330
rect 1423 296 1437 330
rect 1375 258 1437 296
rect 1375 224 1389 258
rect 1423 224 1437 258
rect 1375 186 1437 224
rect 1375 152 1389 186
rect 1423 152 1437 186
rect 1375 114 1437 152
rect 931 47 993 80
rect 1375 80 1389 114
rect 1423 80 1437 114
rect 1375 47 1437 80
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 343 47
rect 377 13 415 47
rect 449 13 513 47
rect 547 13 585 47
rect 619 13 657 47
rect 691 13 729 47
rect 763 13 801 47
rect 835 13 873 47
rect 907 13 1017 47
rect 1051 13 1089 47
rect 1123 13 1167 47
rect 1201 13 1245 47
rect 1279 13 1317 47
rect 1351 13 1437 47
rect -31 11 31 13
rect 931 11 993 13
rect 1375 11 1437 13
<< nsubdiff >>
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 343 1539
rect 377 1505 415 1539
rect 449 1505 513 1539
rect 547 1505 585 1539
rect 619 1505 657 1539
rect 691 1505 729 1539
rect 763 1505 801 1539
rect 835 1505 873 1539
rect 907 1505 1017 1539
rect 1051 1505 1089 1539
rect 1123 1505 1167 1539
rect 1201 1505 1245 1539
rect 1279 1505 1317 1539
rect 1351 1505 1437 1539
rect -31 1470 31 1505
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect 931 1470 993 1505
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect -31 1038 31 1076
rect 931 1436 945 1470
rect 979 1436 993 1470
rect 1375 1470 1437 1505
rect 931 1398 993 1436
rect 931 1364 945 1398
rect 979 1364 993 1398
rect 931 1326 993 1364
rect 931 1292 945 1326
rect 979 1292 993 1326
rect 931 1254 993 1292
rect 931 1220 945 1254
rect 979 1220 993 1254
rect 931 1182 993 1220
rect 931 1148 945 1182
rect 979 1148 993 1182
rect 931 1110 993 1148
rect 931 1076 945 1110
rect 979 1076 993 1110
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect 931 1038 993 1076
rect 1375 1436 1389 1470
rect 1423 1436 1437 1470
rect 1375 1398 1437 1436
rect 1375 1364 1389 1398
rect 1423 1364 1437 1398
rect 1375 1326 1437 1364
rect 1375 1292 1389 1326
rect 1423 1292 1437 1326
rect 1375 1254 1437 1292
rect 1375 1220 1389 1254
rect 1423 1220 1437 1254
rect 1375 1182 1437 1220
rect 1375 1148 1389 1182
rect 1423 1148 1437 1182
rect 1375 1110 1437 1148
rect 1375 1076 1389 1110
rect 1423 1076 1437 1110
rect 931 1004 945 1038
rect 979 1004 993 1038
rect 931 966 993 1004
rect -31 930 31 932
rect 931 932 945 966
rect 979 932 993 966
rect 1375 1038 1437 1076
rect 1375 1004 1389 1038
rect 1423 1004 1437 1038
rect 1375 966 1437 1004
rect 931 930 993 932
rect 1375 932 1389 966
rect 1423 932 1437 966
rect 1375 930 1437 932
rect -31 868 1437 930
<< psubdiffcont >>
rect -17 512 17 546
rect 945 512 979 546
rect 1389 512 1423 546
rect -17 440 17 474
rect -17 368 17 402
rect 945 440 979 474
rect -17 296 17 330
rect -17 224 17 258
rect -17 152 17 186
rect -17 80 17 114
rect 945 368 979 402
rect 1389 440 1423 474
rect 945 296 979 330
rect 945 224 979 258
rect 945 152 979 186
rect 945 80 979 114
rect 1389 368 1423 402
rect 1389 296 1423 330
rect 1389 224 1423 258
rect 1389 152 1423 186
rect 1389 80 1423 114
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 343 13 377 47
rect 415 13 449 47
rect 513 13 547 47
rect 585 13 619 47
rect 657 13 691 47
rect 729 13 763 47
rect 801 13 835 47
rect 873 13 907 47
rect 1017 13 1051 47
rect 1089 13 1123 47
rect 1167 13 1201 47
rect 1245 13 1279 47
rect 1317 13 1351 47
<< nsubdiffcont >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 343 1505 377 1539
rect 415 1505 449 1539
rect 513 1505 547 1539
rect 585 1505 619 1539
rect 657 1505 691 1539
rect 729 1505 763 1539
rect 801 1505 835 1539
rect 873 1505 907 1539
rect 1017 1505 1051 1539
rect 1089 1505 1123 1539
rect 1167 1505 1201 1539
rect 1245 1505 1279 1539
rect 1317 1505 1351 1539
rect -17 1436 17 1470
rect -17 1364 17 1398
rect -17 1292 17 1326
rect -17 1220 17 1254
rect -17 1148 17 1182
rect -17 1076 17 1110
rect 945 1436 979 1470
rect 945 1364 979 1398
rect 945 1292 979 1326
rect 945 1220 979 1254
rect 945 1148 979 1182
rect 945 1076 979 1110
rect -17 1004 17 1038
rect -17 932 17 966
rect 1389 1436 1423 1470
rect 1389 1364 1423 1398
rect 1389 1292 1423 1326
rect 1389 1220 1423 1254
rect 1389 1148 1423 1182
rect 1389 1076 1423 1110
rect 945 1004 979 1038
rect 945 932 979 966
rect 1389 1004 1423 1038
rect 1389 932 1423 966
<< poly >>
rect 247 1450 277 1476
rect 335 1450 365 1476
rect 423 1450 453 1476
rect 511 1450 541 1476
rect 599 1450 629 1476
rect 687 1450 717 1476
rect 1125 1450 1155 1476
rect 1213 1450 1243 1476
rect 247 1019 277 1050
rect 335 1019 365 1050
rect 423 1019 453 1050
rect 511 1019 541 1050
rect 195 1003 365 1019
rect 195 969 205 1003
rect 239 989 365 1003
rect 417 1003 541 1019
rect 239 969 249 989
rect 195 953 249 969
rect 417 969 427 1003
rect 461 989 541 1003
rect 599 1019 629 1050
rect 687 1019 717 1050
rect 599 1003 717 1019
rect 599 989 649 1003
rect 461 969 471 989
rect 417 953 471 969
rect 639 969 649 989
rect 683 989 717 1003
rect 1125 1019 1155 1050
rect 1213 1019 1243 1050
rect 683 969 693 989
rect 639 953 693 969
rect 1083 1003 1243 1019
rect 1083 969 1093 1003
rect 1127 989 1243 1003
rect 1127 969 1137 989
rect 1083 953 1137 969
rect 195 461 249 477
rect 195 441 205 461
rect 147 427 205 441
rect 239 427 249 461
rect 147 411 249 427
rect 417 461 471 477
rect 417 427 427 461
rect 461 441 471 461
rect 639 461 693 477
rect 461 427 477 441
rect 417 411 477 427
rect 639 427 649 461
rect 683 427 693 461
rect 639 411 693 427
rect 147 379 177 411
rect 447 379 477 411
rect 649 379 679 411
rect 1083 461 1137 477
rect 1083 427 1093 461
rect 1127 441 1137 461
rect 1127 427 1147 441
rect 1083 411 1147 427
rect 1117 377 1147 411
<< polycont >>
rect 205 969 239 1003
rect 427 969 461 1003
rect 649 969 683 1003
rect 1093 969 1127 1003
rect 205 427 239 461
rect 427 427 461 461
rect 649 427 683 461
rect 1093 427 1127 461
<< locali >>
rect -31 1539 1437 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 343 1539
rect 377 1505 415 1539
rect 449 1505 513 1539
rect 547 1505 585 1539
rect 619 1505 657 1539
rect 691 1505 729 1539
rect 763 1505 801 1539
rect 835 1505 873 1539
rect 907 1505 1017 1539
rect 1051 1505 1089 1539
rect 1123 1505 1167 1539
rect 1201 1505 1245 1539
rect 1279 1505 1317 1539
rect 1351 1505 1437 1539
rect -31 1492 1437 1505
rect -31 1470 31 1492
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect 201 1412 235 1492
rect 201 1344 235 1378
rect 201 1276 235 1310
rect 201 1208 235 1242
rect 201 1139 235 1174
rect 201 1089 235 1105
rect 289 1412 323 1450
rect 289 1344 323 1378
rect 289 1276 323 1310
rect 289 1208 323 1242
rect 289 1139 323 1174
rect 377 1412 411 1492
rect 377 1344 411 1378
rect 377 1276 411 1310
rect 377 1208 411 1242
rect 377 1157 411 1174
rect 465 1412 499 1450
rect 465 1344 499 1378
rect 465 1276 499 1310
rect 465 1208 499 1242
rect 289 1094 323 1105
rect 465 1139 499 1174
rect 553 1412 587 1492
rect 553 1344 587 1378
rect 553 1276 587 1310
rect 553 1208 587 1242
rect 553 1157 587 1174
rect 641 1412 675 1450
rect 641 1344 675 1378
rect 641 1276 675 1310
rect 641 1208 675 1242
rect 465 1094 499 1105
rect 641 1139 675 1174
rect 729 1412 763 1492
rect 729 1344 763 1378
rect 729 1276 763 1310
rect 729 1208 763 1242
rect 729 1157 763 1174
rect 931 1470 993 1492
rect 931 1436 945 1470
rect 979 1436 993 1470
rect 931 1398 993 1436
rect 931 1364 945 1398
rect 979 1364 993 1398
rect 931 1326 993 1364
rect 931 1292 945 1326
rect 979 1292 993 1326
rect 931 1254 993 1292
rect 931 1220 945 1254
rect 979 1220 993 1254
rect 931 1182 993 1220
rect 641 1094 675 1105
rect 931 1148 945 1182
rect 979 1148 993 1182
rect 931 1110 993 1148
rect -31 1038 31 1076
rect 289 1060 831 1094
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect -31 868 31 932
rect 205 1003 239 1019
rect 205 831 239 969
rect -31 546 31 572
rect -31 512 -17 546
rect 17 512 31 546
rect -31 474 31 512
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect 205 461 239 797
rect 205 411 239 427
rect 427 1003 461 1019
rect 427 757 461 969
rect 427 461 461 723
rect 427 411 461 427
rect 649 1003 683 1019
rect 649 683 683 969
rect 649 461 683 649
rect 649 411 683 427
rect 797 683 831 1060
rect 931 1076 945 1110
rect 979 1076 993 1110
rect 1079 1412 1113 1492
rect 1079 1344 1113 1378
rect 1079 1276 1113 1310
rect 1079 1208 1113 1242
rect 1079 1139 1113 1174
rect 1079 1083 1113 1105
rect 1167 1412 1201 1450
rect 1167 1344 1201 1378
rect 1167 1276 1201 1310
rect 1167 1208 1201 1242
rect 1167 1139 1201 1174
rect 931 1038 993 1076
rect 931 1004 945 1038
rect 979 1004 993 1038
rect 931 966 993 1004
rect 931 932 945 966
rect 979 932 993 966
rect 931 868 993 932
rect 1093 1003 1127 1019
rect -31 368 -17 402
rect 17 368 31 402
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect 101 363 135 379
rect 295 363 329 379
rect 489 363 523 379
rect 135 329 198 363
rect 232 329 295 363
rect 329 329 392 363
rect 426 329 489 363
rect 101 291 135 329
rect 101 223 135 257
rect 295 291 329 329
rect 489 313 523 329
rect 603 363 637 379
rect 797 378 831 649
rect 1093 683 1127 969
rect 1167 979 1201 1105
rect 1255 1412 1289 1492
rect 1255 1344 1289 1378
rect 1255 1276 1289 1310
rect 1255 1208 1289 1242
rect 1255 1139 1289 1174
rect 1255 1083 1289 1105
rect 1375 1470 1437 1492
rect 1375 1436 1389 1470
rect 1423 1436 1437 1470
rect 1375 1398 1437 1436
rect 1375 1364 1389 1398
rect 1423 1364 1437 1398
rect 1375 1326 1437 1364
rect 1375 1292 1389 1326
rect 1423 1292 1437 1326
rect 1375 1254 1437 1292
rect 1375 1220 1389 1254
rect 1423 1220 1437 1254
rect 1375 1182 1437 1220
rect 1375 1148 1389 1182
rect 1423 1148 1437 1182
rect 1375 1110 1437 1148
rect 1375 1076 1389 1110
rect 1423 1076 1437 1110
rect 1375 1038 1437 1076
rect 1375 1004 1389 1038
rect 1423 1004 1437 1038
rect 1167 945 1275 979
rect 603 291 637 329
rect 101 153 135 189
rect 101 103 135 119
rect 198 238 232 254
rect -31 62 31 80
rect 198 62 232 204
rect 295 223 329 257
rect 393 244 427 260
rect 603 244 637 257
rect 427 223 637 244
rect 427 210 603 223
rect 393 194 427 210
rect 295 153 329 189
rect 700 344 831 378
rect 931 546 993 572
rect 931 512 945 546
rect 979 512 993 546
rect 931 474 993 512
rect 931 440 945 474
rect 979 440 993 474
rect 931 402 993 440
rect 1093 461 1127 649
rect 1241 683 1275 945
rect 1375 966 1437 1004
rect 1375 932 1389 966
rect 1423 932 1437 966
rect 1375 868 1437 932
rect 1241 461 1275 649
rect 1093 411 1127 427
rect 1167 427 1275 461
rect 1375 546 1437 572
rect 1375 512 1389 546
rect 1423 512 1437 546
rect 1375 474 1437 512
rect 1375 440 1389 474
rect 1423 440 1437 474
rect 931 368 945 402
rect 979 368 993 402
rect 700 247 734 344
rect 931 330 993 368
rect 700 197 734 213
rect 797 291 831 307
rect 797 223 831 257
rect 489 153 523 169
rect 329 119 392 153
rect 426 119 489 153
rect 295 103 329 119
rect 489 103 523 119
rect 603 153 637 189
rect 797 153 831 189
rect 637 119 700 153
rect 734 119 797 153
rect 603 103 637 119
rect 797 103 831 119
rect 931 296 945 330
rect 979 296 993 330
rect 931 258 993 296
rect 931 224 945 258
rect 979 224 993 258
rect 931 186 993 224
rect 931 152 945 186
rect 979 152 993 186
rect 931 114 993 152
rect 931 80 945 114
rect 979 80 993 114
rect 931 62 993 80
rect 1071 361 1105 377
rect 1071 289 1105 327
rect 1071 221 1105 255
rect 1167 245 1201 427
rect 1375 402 1437 440
rect 1167 195 1201 211
rect 1265 361 1299 377
rect 1265 289 1299 327
rect 1265 221 1299 255
rect 1071 151 1105 187
rect 1265 151 1299 187
rect 1105 117 1167 151
rect 1201 117 1265 151
rect 1071 62 1105 117
rect 1168 62 1202 117
rect 1265 62 1299 117
rect 1375 368 1389 402
rect 1423 368 1437 402
rect 1375 330 1437 368
rect 1375 296 1389 330
rect 1423 296 1437 330
rect 1375 258 1437 296
rect 1375 224 1389 258
rect 1423 224 1437 258
rect 1375 186 1437 224
rect 1375 152 1389 186
rect 1423 152 1437 186
rect 1375 114 1437 152
rect 1375 80 1389 114
rect 1423 80 1437 114
rect 1375 62 1437 80
rect -31 47 1437 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 343 47
rect 377 13 415 47
rect 449 13 513 47
rect 547 13 585 47
rect 619 13 657 47
rect 691 13 729 47
rect 763 13 801 47
rect 835 13 873 47
rect 907 13 1017 47
rect 1051 13 1089 47
rect 1123 13 1167 47
rect 1201 13 1245 47
rect 1279 13 1317 47
rect 1351 13 1437 47
rect -31 0 1437 13
<< viali >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 343 1505 377 1539
rect 415 1505 449 1539
rect 513 1505 547 1539
rect 585 1505 619 1539
rect 657 1505 691 1539
rect 729 1505 763 1539
rect 801 1505 835 1539
rect 873 1505 907 1539
rect 1017 1505 1051 1539
rect 1089 1505 1123 1539
rect 1167 1505 1201 1539
rect 1245 1505 1279 1539
rect 1317 1505 1351 1539
rect 205 797 239 831
rect 427 723 461 757
rect 649 649 683 683
rect 797 649 831 683
rect 1093 649 1127 683
rect 1241 649 1275 683
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 343 13 377 47
rect 415 13 449 47
rect 513 13 547 47
rect 585 13 619 47
rect 657 13 691 47
rect 729 13 763 47
rect 801 13 835 47
rect 873 13 907 47
rect 1017 13 1051 47
rect 1089 13 1123 47
rect 1167 13 1201 47
rect 1245 13 1279 47
rect 1317 13 1351 47
<< metal1 >>
rect -31 1539 1437 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 343 1539
rect 377 1505 415 1539
rect 449 1505 513 1539
rect 547 1505 585 1539
rect 619 1505 657 1539
rect 691 1505 729 1539
rect 763 1505 801 1539
rect 835 1505 873 1539
rect 907 1505 1017 1539
rect 1051 1505 1089 1539
rect 1123 1505 1167 1539
rect 1201 1505 1245 1539
rect 1279 1505 1317 1539
rect 1351 1505 1437 1539
rect -31 1492 1437 1505
rect 199 831 245 837
rect 169 797 205 831
rect 239 797 251 831
rect 199 791 245 797
rect 421 757 467 763
rect 391 723 427 757
rect 461 723 473 757
rect 421 717 467 723
rect 643 683 689 689
rect 791 683 837 689
rect 1087 683 1133 689
rect 1235 683 1281 689
rect 613 649 649 683
rect 683 649 695 683
rect 785 649 797 683
rect 831 649 1093 683
rect 1127 649 1139 683
rect 1229 649 1241 683
rect 1275 649 1311 683
rect 643 643 689 649
rect 791 643 837 649
rect 1087 643 1133 649
rect 1235 643 1281 649
rect -31 47 1437 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 343 47
rect 377 13 415 47
rect 449 13 513 47
rect 547 13 585 47
rect 619 13 657 47
rect 691 13 729 47
rect 763 13 801 47
rect 835 13 873 47
rect 907 13 1017 47
rect 1051 13 1089 47
rect 1123 13 1167 47
rect 1201 13 1245 47
rect 1279 13 1317 47
rect 1351 13 1437 47
rect -31 0 1437 13
<< labels >>
rlabel metal1 1258 666 1258 666 1 Y
port 1 n
rlabel metal1 222 814 222 814 1 A
port 2 n
rlabel metal1 444 740 444 740 1 B
port 3 n
rlabel metal1 666 666 666 666 1 C
port 4 n
rlabel metal1 72 1522 72 1522 1 VDD
port 5 n
rlabel metal1 72 30 72 30 1 VSS
port 6 n
<< end >>
