* SPICE3 file created from AND2X1.ext - technology: sky130A

.subckt AND2X1 Y A B VDD GND
X0 VDD.t9 A.t0 a_217_1050.t2 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X1 Y.t2 a_217_1050.t5 VDD.t5  �S�e sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X2 VDD.t1 B.t0 a_217_1050.t0 �S�e sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X3 GND A.t1 a_112_101.t0 GND sky130_fd_pr__nfet_01v8 ad=1.3199p pd=9.67u as=0p ps=0u w=0u l=0u
X4 a_217_1050.t3 A.t2 VDD.t7  �S�e sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X5 a_217_1050.t4 B.t1 VDD.t11 �S�e sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X6 VDD.t3 a_217_1050.t7 Y.t1  �S�e sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X7 Y a_217_1050.t6 GND.t0 GND sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=0p ps=0u w=0u l=0u
C0 Y VDD 1.07fF
C1 A VDD 0.33fF
C2 B A 0.27fF
C3 B VDD 0.32fF
R0 A.n0 A.t0 480.392
R1 A.n0 A.t2 403.272
R2 A.n1 A.t1 385.063
R3 A.n1 A.n0 143.429
R4 A A.n1 4.65
R5 a_217_1050.n3 a_217_1050.t7 512.525
R6 a_217_1050.n3 a_217_1050.t5 371.139
R7 a_217_1050.n7 a_217_1050.n5 284.244
R8 a_217_1050.n4 a_217_1050.t6 282.852
R9 a_217_1050.n4 a_217_1050.n3 247.347
R10 a_217_1050.n5 a_217_1050.n2 187.858
R11 a_217_1050.n2 a_217_1050.n1 157.964
R12 a_217_1050.n2 a_217_1050.n0 91.706
R13 a_217_1050.n7 a_217_1050.n6 15.218
R14 a_217_1050.n0 a_217_1050.t0 14.282
R15 a_217_1050.n0 a_217_1050.t4 14.282
R16 a_217_1050.n1 a_217_1050.t2 14.282
R17 a_217_1050.n1 a_217_1050.t3 14.282
R18 a_217_1050.n8 a_217_1050.n7 12.014
R19 a_217_1050.n5 a_217_1050.n4 10.343
R20 VDD.n66 VDD.n55 144.705
R21 VDD.n114 VDD.t1 143.754
R22 VDD.n92 VDD.t7 135.17
R23 VDD.n35 VDD.t5 135.17
R24 VDD.n24 VDD.t3 135.17
R25 VDD.n106 VDD.n105 129.472
R26 VDD.n51 VDD.n50 92.5
R27 VDD.n49 VDD.n48 92.5
R28 VDD.n47 VDD.n46 92.5
R29 VDD.n45 VDD.n44 92.5
R30 VDD.n53 VDD.n52 92.5
R31 VDD.n80 VDD.n79 92.5
R32 VDD.n78 VDD.n77 92.5
R33 VDD.n76 VDD.n75 92.5
R34 VDD.n74 VDD.n73 92.5
R35 VDD.n82 VDD.n81 92.5
R36 VDD.n14 VDD.n1 92.5
R37 VDD.n5 VDD.n4 92.5
R38 VDD.n7 VDD.n6 92.5
R39 VDD.n9 VDD.n8 92.5
R40 VDD.n11 VDD.n10 92.5
R41 VDD.n13 VDD.n12 92.5
R42 VDD.n21 VDD.n20 92.059
R43 VDD.n65 VDD.n64 92.059
R44 VDD.n88 VDD.n87 92.059
R45 VDD.n20 VDD.n16 67.194
R46 VDD.n20 VDD.n17 67.194
R47 VDD.n20 VDD.n18 67.194
R48 VDD.n20 VDD.n19 67.194
R49 VDD.n72 VDD.n71 44.141
R50 VDD.n5 VDD.n3 44.141
R51 VDD.n71 VDD.n69 44.107
R52 VDD.n3 VDD.n2 44.107
R53 VDD.n25  �S�e 43.472
R54 VDD.n33  �S�e 43.472
R55 VDD.n20 VDD.n15 41.052
R56 VDD.n84 VDD.n83 39.742
R57 VDD.n63 VDD.n60 39.742
R58 VDD.n63 VDD.n62 39.742
R59 VDD.n59 VDD.n58 39.742
R60 VDD.n71 VDD.n70 38
R61 VDD.n62 VDD.n61 36.774
R62 VDD.n1 VDD.n0 30.923
R63 VDD.n87 VDD.n85 26.38
R64 VDD.n87 VDD.n84 26.38
R65 VDD.n87 VDD.n86 26.38
R66 VDD.n64 VDD.n63 26.38
R67 VDD.n64 VDD.n59 26.38
R68 VDD.n64 VDD.n57 26.38
R69 VDD.n64 VDD.n56 26.38
R70 VDD.n90 VDD.n82 22.915
R71 VDD.n23 VDD.n14 22.915
R72 VDD.n110 �S�e 20.457
R73 VDD.n97  �S�e 17.9
R74 VDD.n82 VDD.n80 14.864
R75 VDD.n80 VDD.n78 14.864
R76 VDD.n78 VDD.n76 14.864
R77 VDD.n76 VDD.n74 14.864
R78 VDD.n74 VDD.n72 14.864
R79 VDD.n53 VDD.n51 14.864
R80 VDD.n51 VDD.n49 14.864
R81 VDD.n49 VDD.n47 14.864
R82 VDD.n47 VDD.n45 14.864
R83 VDD.n45 VDD.n43 14.864
R84 VDD.n43 VDD.n42 14.864
R85 VDD.n14 VDD.n13 14.864
R86 VDD.n13 VDD.n11 14.864
R87 VDD.n11 VDD.n9 14.864
R88 VDD.n9 VDD.n7 14.864
R89 VDD.n7 VDD.n5 14.864
R90 VDD.n67 VDD.n54 14.864
R91 VDD.n105 VDD.t11 14.282
R92 VDD.n105 VDD.t9 14.282
R93 VDD.n108 VDD.n106 9.083
R94 VDD.n23 VDD.n22 8.855
R95 VDD.n22 VDD.n21 8.855
R96 VDD.n27 VDD.n26 8.855
R97 VDD.n26 VDD.n25 8.855
R98 VDD.n31 VDD.n30 8.855
R99 VDD.n30 VDD.n29 8.855
R100 VDD.n36 VDD.n34 8.855
R101 VDD.n34 VDD.n33 8.855
R102 VDD.n40 VDD.n39 8.855
R103 VDD.n39 VDD.n38 8.855
R104 VDD.n67 VDD.n66 8.855
R105 VDD.n66 VDD.n65 8.855
R106 VDD.n117 VDD.n116 8.855
R107 VDD.n116 VDD.n115 8.855
R108 VDD.n112 VDD.n111 8.855
R109 VDD.n111 VDD.n110 8.855
R110 VDD.n108 VDD.n107 8.855
R111 VDD.n107 �S�e 8.855
R112 VDD.n103 VDD.n102 8.855
R113 VDD.n102 VDD.n101 8.855
R114 VDD.n99 VDD.n98 8.855
R115 VDD.n98 VDD.n97 8.855
R116 VDD.n95 VDD.n94 8.855
R117 VDD.n94 VDD.n93 8.855
R118 VDD.n90 VDD.n89 8.855
R119 VDD.n89 VDD.n88 8.855
R120 VDD.n54 VDD.n53 8.051
R121 VDD.n28 VDD.n23 4.795
R122 VDD.n28 VDD.n27 4.65
R123 VDD.n32 VDD.n31 4.65
R124 VDD.n37 VDD.n36 4.65
R125 VDD.n41 VDD.n40 4.65
R126 VDD.n68 VDD.n67 4.65
R127 VDD.n118 VDD.n117 4.65
R128 VDD.n113 VDD.n112 4.65
R129 VDD.n109 VDD.n108 4.65
R130 VDD.n104 VDD.n103 4.65
R131 VDD.n100 VDD.n99 4.65
R132 VDD.n96 VDD.n95 4.65
R133 VDD.n91 VDD.n90 4.65
R134 VDD.n95 VDD.n92 2.89
R135 VDD.n101 VDD.t8 2.557
R136 VDD.n117 VDD.n114 2.477
R137 VDD.n27 VDD.n24 2.064
R138 VDD.n36 VDD.n35 2.064
R139 VDD.n68 VDD.n41 0.29
R140 VDD.n91 VDD 0.207
R141 VDD.n109 VDD.n104 0.181
R142 VDD.n32 VDD.n28 0.157
R143 VDD.n37 VDD.n32 0.157
R144 VDD.n41 VDD.n37 0.145
R145 VDD.n118 VDD.n113 0.145
R146 VDD.n113 VDD.n109 0.145
R147 VDD.n104 VDD.n100 0.145
R148 VDD.n100 VDD.n96 0.145
R149 VDD.n96 VDD.n91 0.145
R150 VDD VDD.n68 0.078
R151 VDD VDD.n118 0.066
R152 Y.n5 Y.n4 272.451
R153 Y.n5 Y.n0 271.281
R154 Y.n4 Y.n3 30
R155 Y.n2 Y.n1 24.383
R156 Y.n4 Y.n2 23.684
R157 Y.n0 Y.t1 14.282
R158 Y.n0 Y.t2 14.282
R159 Y Y.n5 4.65
R160 GND.n32 GND.n31 237.558
R161 GND.n29 GND.n28 210.82
R162 GND.n45 GND.n44 151.605
R163 GND.n21 GND.n20 37.582
R164 GND.t0 GND.n18 32.601
R165 GND.n44 GND.n43 28.421
R166 GND.n44 GND.n42 25.263
R167 GND.n42 GND.n41 24.383
R168 GND.n18 GND.n17 21.734
R169 GND.n4 GND.n3 20.705
R170 GND.n10 GND.n9 20.705
R171 GND.n22 GND.n21 20.705
R172 GND.n3 GND.n2 19.952
R173 GND.n30 GND.n29 18.953
R174 GND.n20 GND.t0 15.644
R175 GND.n33 GND.n30 14.864
R176 GND.n20 GND.n19 13.541
R177 GND.n39 GND.n38 9.154
R178 GND.n47 GND.n46 9.154
R179 GND.n50 GND.n49 9.154
R180 GND.n53 GND.n52 9.154
R181 GND.n56 GND.n55 9.154
R182 GND.n59 GND.n58 9.154
R183 GND.n33 GND.n32 9.154
R184 GND.n26 GND.n25 9.154
R185 GND.n23 GND.n14 9.154
R186 GND.n12 GND.n11 9.154
R187 GND.n6 GND.n5 9.154
R188 GND.n7 GND.n1 4.795
R189 GND.n37 GND.n36 4.65
R190 GND.n7 GND.n6 4.65
R191 GND.n13 GND.n12 4.65
R192 GND.n24 GND.n23 4.65
R193 GND.n27 GND.n26 4.65
R194 GND.n34 GND.n33 4.65
R195 GND.n60 GND.n59 4.65
R196 GND.n57 GND.n56 4.65
R197 GND.n54 GND.n53 4.65
R198 GND.n51 GND.n50 4.65
R199 GND.n48 GND.n47 4.65
R200 GND.n40 GND.n39 4.65
R201 GND.n16 GND.n15 4.504
R202 GND.n6 GND.n4 4.129
R203 GND.n47 GND.n45 4.129
R204 GND.n23 GND.n22 3.716
R205 GND.t0 GND.n16 2.452
R206 GND.n1 GND.n0 0.474
R207 GND.n36 GND.n35 0.474
R208 GND.n9 GND.n8 0.376
R209 GND.n34 GND.n27 0.29
R210 GND.n37 GND 0.207
R211 GND.n12 GND.n10 0.206
R212 GND.n54 GND.n51 0.181
R213 GND.n13 GND.n7 0.157
R214 GND.n24 GND.n13 0.157
R215 GND.n27 GND.n24 0.145
R216 GND.n60 GND.n57 0.145
R217 GND.n57 GND.n54 0.145
R218 GND.n51 GND.n48 0.145
R219 GND.n48 GND.n40 0.145
R220 GND.n40 GND.n37 0.145
R221 GND GND.n34 0.078
R222 GND GND.n60 0.066
R223 B.n0 B.t0 472.359
R224 B.n0 B.t1 384.527
R225 B.n1 B.t2 314.896
R226 B.n1 B.n0 182.814
R227 B B.n1 4.65
R228 a_112_101.n3 a_112_101.n1 42.788
R229 a_112_101.t0 a_112_101.n0 8.137
R230 a_112_101.n3 a_112_101.n2 4.665
R231 a_112_101.t0 a_112_101.n3 0.06
C4 VDD GND 2.00fF
C5 a_112_101.n0 GND 0.05fF
C6 a_112_101.n1 GND 0.11fF
C7 a_112_101.n2 GND 0.04fF
C8 a_112_101.n3 GND 0.16fF
C9 Y.n0 GND 0.65fF
C10 Y.n1 GND 0.04fF
C11 Y.n2 GND 0.05fF
C12 Y.n3 GND 0.03fF
C13 Y.n4 GND 0.19fF
C14 Y.n5 GND 0.63fF
C15 VDD.n1 GND 0.02fF
C16 VDD.n2 GND 0.07fF
C17 VDD.n3 GND 0.02fF
C18 VDD.n4 GND 0.02fF
C19 VDD.n5 GND 0.04fF
C20 VDD.n6 GND 0.02fF
C21 VDD.n7 GND 0.02fF
C22 VDD.n8 GND 0.02fF
C23 VDD.n9 GND 0.02fF
C24 VDD.n10 GND 0.02fF
C25 VDD.n11 GND 0.02fF
C26 VDD.n12 GND 0.02fF
C27 VDD.n13 GND 0.02fF
C28 VDD.n14 GND 0.03fF
C29 VDD.n15 GND 0.01fF
C30 VDD.n20 GND 0.33fF
C31 VDD.n21 GND 0.20fF
C32 VDD.n22 GND 0.01fF
C33 VDD.n23 GND 0.02fF
C34 VDD.n24 GND 0.05fF
C35 VDD.n25 GND 0.15fF
C36 VDD.n26 GND 0.01fF
C37 VDD.n27 GND 0.01fF
C38 VDD.n28 GND 0.05fF
C39 VDD.n29 GND 0.12fF
C40 VDD.n30 GND 0.01fF
C41 VDD.n31 GND 0.02fF
C42 VDD.n32 GND 0.02fF
C43 VDD.n33 GND 0.15fF
C44 VDD.n34 GND 0.01f