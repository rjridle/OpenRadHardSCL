magic
tech sky130A
magscale 1 2
timestamp 1648504834
<< nwell >>
rect 55 1505 89 1539
<< psubdiffcont >>
rect 55 13 89 47
<< nsubdiffcont >>
rect 55 1505 89 1539
<< viali >>
rect 55 1505 89 1539
rect 55 13 89 47
<< metal1 >>
rect 1090 945 12712 979
rect 13264 945 14484 979
rect 14523 871 15567 905
rect 4087 797 4562 831
rect 8973 797 9440 831
rect 13857 797 14318 831
rect 16929 797 16963 831
rect 8334 723 15039 757
rect 3496 649 15837 683
rect 205 575 10003 609
rect 2055 427 13468 461
use li1_M1_contact  li1_M1_contact_3 pcells
timestamp 1648061256
transform -1 0 3478 0 -1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_7
timestamp 1648061256
transform -1 0 222 0 -1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_4
timestamp 1648061256
transform -1 0 4070 0 -1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_6
timestamp 1648061256
transform 1 0 4736 0 1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_5
timestamp 1648061256
transform 1 0 4588 0 1 814
box -53 -33 29 33
use dffsnqx1  dffsnqx1_1 pcells
timestamp 1648501217
transform 1 0 4884 0 1 0
box -84 0 4968 1575
use dffsnqx1  dffsnqx1_0
timestamp 1648501217
transform 1 0 0 0 1 0
box -84 0 4968 1575
use li1_M1_contact  li1_M1_contact_15
timestamp 1648061256
transform -1 0 5106 0 -1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_12
timestamp 1648061256
transform -1 0 8362 0 -1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_13
timestamp 1648061256
transform 1 0 9620 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_10
timestamp 1648061256
transform 1 0 9472 0 1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_9
timestamp 1648061256
transform -1 0 8954 0 -1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_8
timestamp 1648061256
transform 1 0 9990 0 1 592
box -53 -33 29 33
use dffsnqx1  dffsnqx1_2
timestamp 1648501217
transform 1 0 9768 0 1 0
box -84 0 4968 1575
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform -1 0 13246 0 -1 962
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_2
timestamp 1648061256
transform -1 0 14504 0 -1 888
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform 1 0 14504 0 1 962
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_11
timestamp 1648061256
transform -1 0 13838 0 -1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_19
timestamp 1648061256
transform 1 0 14356 0 1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_14
timestamp 1648061256
transform 1 0 15022 0 -1 740
box -53 -33 29 33
use voter3x1_pcell  voter3x1_pcell_0 pcells
timestamp 1648490579
transform 1 0 14652 0 1 0
box -84 0 2526 1575
use li1_M1_contact  li1_M1_contact_16
timestamp 1648061256
transform 1 0 15836 0 -1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_17
timestamp 1648061256
transform -1 0 16946 0 -1 814
box -53 -33 29 33
<< labels >>
rlabel metal1 16929 797 16963 831 1 Q
port 1 n
rlabel metal1 205 575 239 609 1 D
port 2 n
rlabel metal1 1093 945 1127 979 1 CLK
port 3 n
rlabel metal1 2055 427 2089 461 1 SN
port 4 n
rlabel metal1 72 1522 72 1522 1 VDD
port 5 n
rlabel metal1 72 30 72 30 1 VSS
port 6 n
<< end >>
