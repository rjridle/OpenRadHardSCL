magic
tech sky130A
magscale 1 2
timestamp 1648328097
<< nwell >>
rect -84 832 1712 1575
<< nmos >>
rect 164 316 194 377
tri 194 316 210 332 sw
rect 358 324 388 377
tri 388 324 404 340 sw
rect 164 286 270 316
tri 270 286 300 316 sw
rect 358 294 464 324
tri 464 294 494 324 sw
rect 164 185 194 286
tri 194 270 210 286 nw
tri 254 270 270 286 ne
tri 194 185 210 201 sw
tri 254 185 270 201 se
rect 270 185 300 286
rect 358 193 388 294
tri 388 278 404 294 nw
tri 448 278 464 294 ne
tri 388 193 404 209 sw
tri 448 193 464 209 se
rect 464 193 494 294
tri 164 155 194 185 ne
rect 194 155 270 185
tri 270 155 300 185 nw
tri 358 163 388 193 ne
rect 388 163 464 193
tri 464 163 494 193 nw
rect 662 324 692 377
tri 692 324 708 340 sw
rect 662 294 768 324
tri 768 294 798 324 sw
rect 662 193 692 294
tri 692 278 708 294 nw
tri 752 278 768 294 ne
tri 692 193 708 209 sw
tri 752 193 768 209 se
rect 768 193 798 294
rect 856 316 886 377
tri 886 316 902 332 sw
rect 856 286 962 316
tri 962 286 992 316 sw
tri 662 163 692 193 ne
rect 692 163 768 193
tri 768 163 798 193 nw
rect 856 185 886 286
tri 886 270 902 286 nw
tri 946 270 962 286 ne
tri 886 185 902 201 sw
tri 946 185 962 201 se
rect 962 185 992 286
tri 856 155 886 185 ne
rect 886 155 962 185
tri 962 155 992 185 nw
rect 1339 324 1369 377
tri 1369 324 1385 340 sw
rect 1339 294 1445 324
tri 1445 294 1475 324 sw
rect 1339 193 1369 294
tri 1369 278 1385 294 nw
tri 1429 278 1445 294 ne
tri 1369 193 1385 209 sw
tri 1429 193 1445 209 se
rect 1445 193 1475 294
tri 1339 163 1369 193 ne
rect 1369 163 1445 193
tri 1445 163 1475 193 nw
<< pmos >>
rect 193 1051 223 1451
rect 281 1051 311 1451
rect 369 1051 399 1451
rect 457 1051 487 1451
rect 545 1051 575 1451
rect 633 1051 663 1451
rect 829 1051 859 1451
rect 917 1051 947 1451
rect 1347 1050 1377 1450
rect 1435 1050 1465 1450
<< ndiff >>
rect 108 361 164 377
rect 108 327 118 361
rect 152 327 164 361
rect 108 289 164 327
rect 194 361 358 377
rect 194 332 215 361
tri 194 316 210 332 ne
rect 210 327 215 332
rect 249 327 312 361
rect 346 327 358 361
rect 210 316 358 327
rect 388 340 550 377
tri 388 324 404 340 ne
rect 404 324 550 340
rect 108 255 118 289
rect 152 255 164 289
tri 270 286 300 316 ne
rect 300 289 358 316
tri 464 294 494 324 ne
rect 108 221 164 255
rect 108 187 118 221
rect 152 187 164 221
rect 108 155 164 187
tri 194 270 210 286 se
rect 210 270 254 286
tri 254 270 270 286 sw
rect 194 236 270 270
rect 194 202 215 236
rect 249 202 270 236
rect 194 201 270 202
tri 194 185 210 201 ne
rect 210 185 254 201
tri 254 185 270 201 nw
rect 300 255 312 289
rect 346 255 358 289
rect 300 221 358 255
rect 300 187 312 221
rect 346 187 358 221
tri 388 278 404 294 se
rect 404 278 448 294
tri 448 278 464 294 sw
rect 388 245 464 278
rect 388 211 409 245
rect 443 211 464 245
rect 388 209 464 211
tri 388 193 404 209 ne
rect 404 193 448 209
tri 448 193 464 209 nw
rect 494 289 550 324
rect 494 255 506 289
rect 540 255 550 289
rect 494 221 550 255
tri 164 155 194 185 sw
tri 270 155 300 185 se
rect 300 163 358 187
tri 358 163 388 193 sw
tri 464 163 494 193 se
rect 494 187 506 221
rect 540 187 550 221
rect 494 163 550 187
rect 300 155 550 163
rect 108 151 550 155
rect 108 117 118 151
rect 152 117 312 151
rect 346 117 409 151
rect 443 117 506 151
rect 540 117 550 151
rect 108 101 550 117
rect 606 361 662 377
rect 606 327 616 361
rect 650 327 662 361
rect 606 289 662 327
rect 692 361 856 377
rect 692 340 810 361
tri 692 324 708 340 ne
rect 708 327 810 340
rect 844 327 856 361
rect 708 324 856 327
tri 768 294 798 324 ne
rect 606 255 616 289
rect 650 255 662 289
rect 606 221 662 255
rect 606 187 616 221
rect 650 187 662 221
tri 692 278 708 294 se
rect 708 278 752 294
tri 752 278 768 294 sw
rect 692 245 768 278
rect 692 211 713 245
rect 747 211 768 245
rect 692 209 768 211
tri 692 193 708 209 ne
rect 708 193 752 209
tri 752 193 768 209 nw
rect 798 289 856 324
rect 886 361 1048 377
rect 886 332 907 361
tri 886 316 902 332 ne
rect 902 327 907 332
rect 941 327 1004 361
rect 1038 327 1048 361
rect 902 316 1048 327
rect 798 255 810 289
rect 844 255 856 289
tri 962 286 992 316 ne
rect 992 289 1048 316
rect 798 221 856 255
rect 606 163 662 187
tri 662 163 692 193 sw
tri 768 163 798 193 se
rect 798 187 810 221
rect 844 187 856 221
rect 798 163 856 187
tri 886 270 902 286 se
rect 902 270 946 286
tri 946 270 962 286 sw
rect 886 236 962 270
rect 886 202 907 236
rect 941 202 962 236
rect 886 201 962 202
tri 886 185 902 201 ne
rect 902 185 946 201
tri 946 185 962 201 nw
rect 992 255 1004 289
rect 1038 255 1048 289
rect 992 221 1048 255
rect 992 187 1004 221
rect 1038 187 1048 221
rect 606 155 856 163
tri 856 155 886 185 sw
tri 962 155 992 185 se
rect 992 155 1048 187
rect 606 151 1048 155
rect 606 117 616 151
rect 650 117 713 151
rect 747 117 810 151
rect 844 117 1004 151
rect 1038 117 1048 151
rect 606 101 1048 117
rect 1283 361 1339 377
rect 1283 327 1293 361
rect 1327 327 1339 361
rect 1283 289 1339 327
rect 1369 361 1529 377
rect 1369 340 1487 361
tri 1369 324 1385 340 ne
rect 1385 327 1487 340
rect 1521 327 1529 361
rect 1385 324 1529 327
tri 1445 294 1475 324 ne
rect 1283 255 1293 289
rect 1327 255 1339 289
rect 1283 221 1339 255
rect 1283 187 1293 221
rect 1327 187 1339 221
tri 1369 278 1385 294 se
rect 1385 278 1429 294
tri 1429 278 1445 294 sw
rect 1369 245 1445 278
rect 1369 211 1389 245
rect 1423 211 1445 245
rect 1369 209 1445 211
tri 1369 193 1385 209 ne
rect 1385 193 1429 209
tri 1429 193 1445 209 nw
rect 1475 289 1529 324
rect 1475 255 1487 289
rect 1521 255 1529 289
rect 1475 221 1529 255
rect 1283 163 1339 187
tri 1339 163 1369 193 sw
tri 1445 163 1475 193 se
rect 1475 187 1487 221
rect 1521 187 1529 221
rect 1475 163 1529 187
rect 1283 151 1529 163
rect 1283 117 1293 151
rect 1327 117 1389 151
rect 1423 117 1487 151
rect 1521 117 1529 151
rect 1283 101 1529 117
<< pdiff >>
rect 137 1411 193 1451
rect 137 1377 147 1411
rect 181 1377 193 1411
rect 137 1343 193 1377
rect 137 1309 147 1343
rect 181 1309 193 1343
rect 137 1275 193 1309
rect 137 1241 147 1275
rect 181 1241 193 1275
rect 137 1207 193 1241
rect 137 1173 147 1207
rect 181 1173 193 1207
rect 137 1051 193 1173
rect 223 1411 281 1451
rect 223 1377 235 1411
rect 269 1377 281 1411
rect 223 1343 281 1377
rect 223 1309 235 1343
rect 269 1309 281 1343
rect 223 1275 281 1309
rect 223 1241 235 1275
rect 269 1241 281 1275
rect 223 1207 281 1241
rect 223 1173 235 1207
rect 269 1173 281 1207
rect 223 1139 281 1173
rect 223 1105 235 1139
rect 269 1105 281 1139
rect 223 1051 281 1105
rect 311 1411 369 1451
rect 311 1377 323 1411
rect 357 1377 369 1411
rect 311 1343 369 1377
rect 311 1309 323 1343
rect 357 1309 369 1343
rect 311 1275 369 1309
rect 311 1241 323 1275
rect 357 1241 369 1275
rect 311 1207 369 1241
rect 311 1173 323 1207
rect 357 1173 369 1207
rect 311 1051 369 1173
rect 399 1413 457 1451
rect 399 1377 411 1413
rect 445 1377 457 1413
rect 399 1343 457 1377
rect 399 1309 411 1343
rect 445 1309 457 1343
rect 399 1275 457 1309
rect 399 1241 411 1275
rect 445 1241 457 1275
rect 399 1207 457 1241
rect 399 1173 411 1207
rect 445 1173 457 1207
rect 399 1139 457 1173
rect 399 1105 411 1139
rect 445 1105 457 1139
rect 399 1051 457 1105
rect 487 1411 545 1451
rect 487 1377 499 1411
rect 533 1377 545 1411
rect 487 1343 545 1377
rect 487 1309 499 1343
rect 533 1309 545 1343
rect 487 1275 545 1309
rect 487 1241 499 1275
rect 533 1241 545 1275
rect 487 1207 545 1241
rect 487 1173 499 1207
rect 533 1173 545 1207
rect 487 1051 545 1173
rect 575 1343 633 1451
rect 575 1309 587 1343
rect 621 1309 633 1343
rect 575 1275 633 1309
rect 575 1241 587 1275
rect 621 1241 633 1275
rect 575 1207 633 1241
rect 575 1173 587 1207
rect 621 1173 633 1207
rect 575 1051 633 1173
rect 663 1411 717 1451
rect 663 1377 675 1411
rect 709 1377 717 1411
rect 663 1343 717 1377
rect 663 1309 675 1343
rect 709 1309 717 1343
rect 663 1275 717 1309
rect 663 1241 675 1275
rect 709 1241 717 1275
rect 663 1207 717 1241
rect 663 1173 675 1207
rect 709 1173 717 1207
rect 663 1051 717 1173
rect 773 1411 829 1451
rect 773 1377 783 1411
rect 817 1377 829 1411
rect 773 1343 829 1377
rect 773 1309 783 1343
rect 817 1309 829 1343
rect 773 1275 829 1309
rect 773 1241 783 1275
rect 817 1241 829 1275
rect 773 1207 829 1241
rect 773 1173 783 1207
rect 817 1173 829 1207
rect 773 1051 829 1173
rect 859 1343 917 1451
rect 859 1309 871 1343
rect 905 1309 917 1343
rect 859 1275 917 1309
rect 859 1241 871 1275
rect 905 1241 917 1275
rect 859 1207 917 1241
rect 859 1173 871 1207
rect 905 1173 917 1207
rect 859 1051 917 1173
rect 947 1411 1001 1451
rect 947 1377 959 1411
rect 993 1377 1001 1411
rect 947 1343 1001 1377
rect 947 1309 959 1343
rect 993 1309 1001 1343
rect 947 1275 1001 1309
rect 947 1241 959 1275
rect 993 1241 1001 1275
rect 947 1207 1001 1241
rect 947 1173 959 1207
rect 993 1173 1001 1207
rect 947 1051 1001 1173
rect 1291 1412 1347 1450
rect 1291 1378 1301 1412
rect 1335 1378 1347 1412
rect 1291 1344 1347 1378
rect 1291 1310 1301 1344
rect 1335 1310 1347 1344
rect 1291 1276 1347 1310
rect 1291 1242 1301 1276
rect 1335 1242 1347 1276
rect 1291 1208 1347 1242
rect 1291 1174 1301 1208
rect 1335 1174 1347 1208
rect 1291 1139 1347 1174
rect 1291 1105 1301 1139
rect 1335 1105 1347 1139
rect 1291 1050 1347 1105
rect 1377 1412 1435 1450
rect 1377 1378 1389 1412
rect 1423 1378 1435 1412
rect 1377 1344 1435 1378
rect 1377 1310 1389 1344
rect 1423 1310 1435 1344
rect 1377 1276 1435 1310
rect 1377 1242 1389 1276
rect 1423 1242 1435 1276
rect 1377 1208 1435 1242
rect 1377 1174 1389 1208
rect 1423 1174 1435 1208
rect 1377 1139 1435 1174
rect 1377 1105 1389 1139
rect 1423 1105 1435 1139
rect 1377 1050 1435 1105
rect 1465 1412 1519 1450
rect 1465 1378 1477 1412
rect 1511 1378 1519 1412
rect 1465 1344 1519 1378
rect 1465 1310 1477 1344
rect 1511 1310 1519 1344
rect 1465 1276 1519 1310
rect 1465 1242 1477 1276
rect 1511 1242 1519 1276
rect 1465 1208 1519 1242
rect 1465 1174 1477 1208
rect 1511 1174 1519 1208
rect 1465 1139 1519 1174
rect 1465 1105 1477 1139
rect 1511 1105 1519 1139
rect 1465 1050 1519 1105
<< ndiffc >>
rect 118 327 152 361
rect 215 327 249 361
rect 312 327 346 361
rect 118 255 152 289
rect 118 187 152 221
rect 215 202 249 236
rect 312 255 346 289
rect 312 187 346 221
rect 409 211 443 245
rect 506 255 540 289
rect 506 187 540 221
rect 118 117 152 151
rect 312 117 346 151
rect 409 117 443 151
rect 506 117 540 151
rect 616 327 650 361
rect 810 327 844 361
rect 616 255 650 289
rect 616 187 650 221
rect 713 211 747 245
rect 907 327 941 361
rect 1004 327 1038 361
rect 810 255 844 289
rect 810 187 844 221
rect 907 202 941 236
rect 1004 255 1038 289
rect 1004 187 1038 221
rect 616 117 650 151
rect 713 117 747 151
rect 810 117 844 151
rect 1004 117 1038 151
rect 1293 327 1327 361
rect 1487 327 1521 361
rect 1293 255 1327 289
rect 1293 187 1327 221
rect 1389 211 1423 245
rect 1487 255 1521 289
rect 1487 187 1521 221
rect 1293 117 1327 151
rect 1389 117 1423 151
rect 1487 117 1521 151
<< pdiffc >>
rect 147 1377 181 1411
rect 147 1309 181 1343
rect 147 1241 181 1275
rect 147 1173 181 1207
rect 235 1377 269 1411
rect 235 1309 269 1343
rect 235 1241 269 1275
rect 235 1173 269 1207
rect 235 1105 269 1139
rect 323 1377 357 1411
rect 323 1309 357 1343
rect 323 1241 357 1275
rect 323 1173 357 1207
rect 411 1377 445 1413
rect 411 1309 445 1343
rect 411 1241 445 1275
rect 411 1173 445 1207
rect 411 1105 445 1139
rect 499 1377 533 1411
rect 499 1309 533 1343
rect 499 1241 533 1275
rect 499 1173 533 1207
rect 587 1309 621 1343
rect 587 1241 621 1275
rect 587 1173 621 1207
rect 675 1377 709 1411
rect 675 1309 709 1343
rect 675 1241 709 1275
rect 675 1173 709 1207
rect 783 1377 817 1411
rect 783 1309 817 1343
rect 783 1241 817 1275
rect 783 1173 817 1207
rect 871 1309 905 1343
rect 871 1241 905 1275
rect 871 1173 905 1207
rect 959 1377 993 1411
rect 959 1309 993 1343
rect 959 1241 993 1275
rect 959 1173 993 1207
rect 1301 1378 1335 1412
rect 1301 1310 1335 1344
rect 1301 1242 1335 1276
rect 1301 1174 1335 1208
rect 1301 1105 1335 1139
rect 1389 1378 1423 1412
rect 1389 1310 1423 1344
rect 1389 1242 1423 1276
rect 1389 1174 1423 1208
rect 1389 1105 1423 1139
rect 1477 1378 1511 1412
rect 1477 1310 1511 1344
rect 1477 1242 1511 1276
rect 1477 1174 1511 1208
rect 1477 1105 1511 1139
<< psubdiff >>
rect -31 546 1659 572
rect -31 512 -17 546
rect 17 512 1167 546
rect 1201 512 1611 546
rect 1645 512 1659 546
rect -31 510 1659 512
rect -31 474 31 510
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect -31 368 -17 402
rect 17 368 31 402
rect 1153 474 1215 510
rect 1153 440 1167 474
rect 1201 440 1215 474
rect 1153 402 1215 440
rect 1597 474 1659 510
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect 1153 368 1167 402
rect 1201 368 1215 402
rect 1597 440 1611 474
rect 1645 440 1659 474
rect 1597 402 1659 440
rect 1153 330 1215 368
rect 1153 296 1167 330
rect 1201 296 1215 330
rect 1153 258 1215 296
rect 1153 224 1167 258
rect 1201 224 1215 258
rect 1153 186 1215 224
rect 1153 152 1167 186
rect 1201 152 1215 186
rect 1153 114 1215 152
rect -31 47 31 80
rect 1153 80 1167 114
rect 1201 80 1215 114
rect 1597 368 1611 402
rect 1645 368 1659 402
rect 1597 330 1659 368
rect 1597 296 1611 330
rect 1645 296 1659 330
rect 1597 258 1659 296
rect 1597 224 1611 258
rect 1645 224 1659 258
rect 1597 186 1659 224
rect 1597 152 1611 186
rect 1645 152 1659 186
rect 1597 114 1659 152
rect 1153 47 1215 80
rect 1597 80 1611 114
rect 1645 80 1659 114
rect 1597 47 1659 80
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 343 47
rect 377 13 415 47
rect 449 13 487 47
rect 521 13 585 47
rect 619 13 663 47
rect 697 13 735 47
rect 769 13 807 47
rect 841 13 879 47
rect 913 13 951 47
rect 985 13 1023 47
rect 1057 13 1095 47
rect 1129 13 1239 47
rect 1273 13 1311 47
rect 1345 13 1389 47
rect 1423 13 1467 47
rect 1501 13 1539 47
rect 1573 13 1659 47
rect -31 11 31 13
rect 1153 11 1215 13
rect 1597 11 1659 13
<< nsubdiff >>
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 343 1539
rect 377 1505 415 1539
rect 449 1505 487 1539
rect 521 1505 585 1539
rect 619 1505 663 1539
rect 697 1505 735 1539
rect 769 1505 807 1539
rect 841 1505 879 1539
rect 913 1505 951 1539
rect 985 1505 1023 1539
rect 1057 1505 1095 1539
rect 1129 1505 1239 1539
rect 1273 1505 1311 1539
rect 1345 1505 1389 1539
rect 1423 1505 1467 1539
rect 1501 1505 1539 1539
rect 1573 1505 1659 1539
rect -31 1470 31 1505
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect 1153 1470 1215 1505
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect -31 1038 31 1076
rect 1153 1436 1167 1470
rect 1201 1436 1215 1470
rect 1597 1470 1659 1505
rect 1153 1398 1215 1436
rect 1153 1364 1167 1398
rect 1201 1364 1215 1398
rect 1153 1326 1215 1364
rect 1153 1292 1167 1326
rect 1201 1292 1215 1326
rect 1153 1254 1215 1292
rect 1153 1220 1167 1254
rect 1201 1220 1215 1254
rect 1153 1182 1215 1220
rect 1153 1148 1167 1182
rect 1201 1148 1215 1182
rect 1153 1110 1215 1148
rect 1153 1076 1167 1110
rect 1201 1076 1215 1110
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect 1153 1038 1215 1076
rect 1597 1436 1611 1470
rect 1645 1436 1659 1470
rect 1597 1398 1659 1436
rect 1597 1364 1611 1398
rect 1645 1364 1659 1398
rect 1597 1326 1659 1364
rect 1597 1292 1611 1326
rect 1645 1292 1659 1326
rect 1597 1254 1659 1292
rect 1597 1220 1611 1254
rect 1645 1220 1659 1254
rect 1597 1182 1659 1220
rect 1597 1148 1611 1182
rect 1645 1148 1659 1182
rect 1597 1110 1659 1148
rect 1597 1076 1611 1110
rect 1645 1076 1659 1110
rect 1153 1004 1167 1038
rect 1201 1004 1215 1038
rect 1153 966 1215 1004
rect -31 930 31 932
rect 1153 932 1167 966
rect 1201 932 1215 966
rect 1597 1038 1659 1076
rect 1597 1004 1611 1038
rect 1645 1004 1659 1038
rect 1597 966 1659 1004
rect 1153 930 1215 932
rect 1597 932 1611 966
rect 1645 932 1659 966
rect 1597 930 1659 932
rect -31 868 1659 930
<< psubdiffcont >>
rect -17 512 17 546
rect 1167 512 1201 546
rect 1611 512 1645 546
rect -17 440 17 474
rect -17 368 17 402
rect 1167 440 1201 474
rect -17 296 17 330
rect -17 224 17 258
rect -17 152 17 186
rect -17 80 17 114
rect 1167 368 1201 402
rect 1611 440 1645 474
rect 1167 296 1201 330
rect 1167 224 1201 258
rect 1167 152 1201 186
rect 1167 80 1201 114
rect 1611 368 1645 402
rect 1611 296 1645 330
rect 1611 224 1645 258
rect 1611 152 1645 186
rect 1611 80 1645 114
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 343 13 377 47
rect 415 13 449 47
rect 487 13 521 47
rect 585 13 619 47
rect 663 13 697 47
rect 735 13 769 47
rect 807 13 841 47
rect 879 13 913 47
rect 951 13 985 47
rect 1023 13 1057 47
rect 1095 13 1129 47
rect 1239 13 1273 47
rect 1311 13 1345 47
rect 1389 13 1423 47
rect 1467 13 1501 47
rect 1539 13 1573 47
<< nsubdiffcont >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 343 1505 377 1539
rect 415 1505 449 1539
rect 487 1505 521 1539
rect 585 1505 619 1539
rect 663 1505 697 1539
rect 735 1505 769 1539
rect 807 1505 841 1539
rect 879 1505 913 1539
rect 951 1505 985 1539
rect 1023 1505 1057 1539
rect 1095 1505 1129 1539
rect 1239 1505 1273 1539
rect 1311 1505 1345 1539
rect 1389 1505 1423 1539
rect 1467 1505 1501 1539
rect 1539 1505 1573 1539
rect -17 1436 17 1470
rect -17 1364 17 1398
rect -17 1292 17 1326
rect -17 1220 17 1254
rect -17 1148 17 1182
rect -17 1076 17 1110
rect 1167 1436 1201 1470
rect 1167 1364 1201 1398
rect 1167 1292 1201 1326
rect 1167 1220 1201 1254
rect 1167 1148 1201 1182
rect 1167 1076 1201 1110
rect -17 1004 17 1038
rect -17 932 17 966
rect 1611 1436 1645 1470
rect 1611 1364 1645 1398
rect 1611 1292 1645 1326
rect 1611 1220 1645 1254
rect 1611 1148 1645 1182
rect 1611 1076 1645 1110
rect 1167 1004 1201 1038
rect 1167 932 1201 966
rect 1611 1004 1645 1038
rect 1611 932 1645 966
<< poly >>
rect 193 1451 223 1477
rect 281 1451 311 1477
rect 369 1451 399 1477
rect 457 1451 487 1477
rect 545 1451 575 1477
rect 633 1451 663 1477
rect 829 1451 859 1477
rect 917 1451 947 1477
rect 1347 1450 1377 1476
rect 1435 1450 1465 1476
rect 193 1020 223 1051
rect 281 1020 311 1051
rect 369 1020 399 1051
rect 457 1020 487 1051
rect 193 1004 311 1020
rect 193 990 205 1004
rect 195 970 205 990
rect 239 990 311 1004
rect 359 1004 487 1020
rect 239 970 249 990
rect 195 954 249 970
rect 359 970 369 1004
rect 403 990 487 1004
rect 545 1020 575 1051
rect 633 1020 663 1051
rect 829 1020 859 1051
rect 917 1020 947 1051
rect 545 1004 693 1020
rect 545 990 649 1004
rect 403 970 413 990
rect 359 954 413 970
rect 639 970 649 990
rect 683 970 693 1004
rect 829 1004 947 1020
rect 829 990 871 1004
rect 639 954 693 970
rect 861 970 871 990
rect 905 990 947 1004
rect 1347 1019 1377 1050
rect 1435 1019 1465 1050
rect 905 970 915 990
rect 861 954 915 970
rect 1305 1003 1465 1019
rect 1305 969 1315 1003
rect 1349 989 1465 1003
rect 1349 969 1359 989
rect 1305 953 1359 969
rect 195 461 249 477
rect 195 441 205 461
rect 164 427 205 441
rect 239 427 249 461
rect 164 411 249 427
rect 343 461 397 477
rect 343 427 353 461
rect 387 427 397 461
rect 343 411 397 427
rect 639 461 693 477
rect 639 427 649 461
rect 683 427 693 461
rect 861 461 915 477
rect 861 444 871 461
rect 639 411 693 427
rect 856 427 871 444
rect 905 427 915 461
rect 856 411 915 427
rect 164 377 194 411
rect 358 377 388 411
rect 662 377 692 411
rect 856 377 886 411
rect 1305 461 1359 477
rect 1305 427 1315 461
rect 1349 441 1359 461
rect 1349 427 1369 441
rect 1305 411 1369 427
rect 1339 377 1369 411
<< polycont >>
rect 205 970 239 1004
rect 369 970 403 1004
rect 649 970 683 1004
rect 871 970 905 1004
rect 1315 969 1349 1003
rect 205 427 239 461
rect 353 427 387 461
rect 649 427 683 461
rect 871 427 905 461
rect 1315 427 1349 461
<< locali >>
rect -31 1539 1659 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 343 1539
rect 377 1505 415 1539
rect 449 1505 487 1539
rect 521 1505 585 1539
rect 619 1505 663 1539
rect 697 1505 735 1539
rect 769 1505 807 1539
rect 841 1505 879 1539
rect 913 1505 951 1539
rect 985 1505 1023 1539
rect 1057 1505 1095 1539
rect 1129 1505 1239 1539
rect 1273 1505 1311 1539
rect 1345 1505 1389 1539
rect 1423 1505 1467 1539
rect 1501 1505 1539 1539
rect 1573 1505 1659 1539
rect -31 1492 1659 1505
rect -31 1470 31 1492
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect 147 1411 181 1492
rect 147 1343 181 1377
rect 147 1275 181 1309
rect 147 1207 181 1241
rect 147 1157 181 1173
rect 235 1411 269 1445
rect 235 1343 269 1377
rect 235 1275 269 1309
rect 235 1207 269 1241
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect -31 1038 31 1076
rect 235 1139 269 1173
rect 323 1411 357 1492
rect 323 1343 357 1377
rect 323 1275 357 1309
rect 323 1207 357 1241
rect 323 1157 357 1173
rect 411 1413 445 1429
rect 411 1343 445 1377
rect 411 1275 445 1309
rect 411 1207 445 1241
rect 235 1071 269 1105
rect 411 1139 445 1173
rect 499 1411 533 1492
rect 499 1343 533 1377
rect 675 1411 709 1492
rect 1153 1470 1215 1492
rect 499 1275 533 1309
rect 499 1207 533 1241
rect 499 1157 533 1173
rect 587 1343 621 1359
rect 587 1275 621 1309
rect 587 1207 621 1241
rect 587 1105 621 1173
rect 675 1343 709 1377
rect 675 1275 709 1309
rect 675 1207 709 1241
rect 675 1157 709 1173
rect 783 1411 993 1445
rect 783 1343 817 1377
rect 783 1275 817 1309
rect 783 1207 817 1241
rect 783 1105 817 1173
rect 871 1343 905 1359
rect 871 1275 905 1309
rect 871 1207 905 1241
rect 871 1157 905 1173
rect 959 1343 993 1377
rect 959 1275 993 1309
rect 959 1207 993 1241
rect 959 1157 993 1173
rect 1153 1436 1167 1470
rect 1201 1436 1215 1470
rect 1153 1398 1215 1436
rect 1153 1364 1167 1398
rect 1201 1364 1215 1398
rect 1153 1326 1215 1364
rect 1153 1292 1167 1326
rect 1201 1292 1215 1326
rect 1153 1254 1215 1292
rect 1153 1220 1167 1254
rect 1201 1220 1215 1254
rect 1153 1182 1215 1220
rect 411 1071 817 1105
rect 1153 1148 1167 1182
rect 1201 1148 1215 1182
rect 1153 1110 1215 1148
rect 1153 1076 1167 1110
rect 1201 1076 1215 1110
rect 1301 1412 1335 1492
rect 1301 1344 1335 1378
rect 1301 1276 1335 1310
rect 1301 1208 1335 1242
rect 1301 1139 1335 1174
rect 1301 1083 1335 1105
rect 1389 1412 1423 1450
rect 1389 1344 1423 1378
rect 1389 1276 1423 1310
rect 1389 1208 1423 1242
rect 1389 1139 1423 1174
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect 1153 1038 1215 1076
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect -31 868 31 932
rect 205 1004 239 1020
rect 369 1004 403 1020
rect 205 609 239 970
rect -31 546 31 572
rect -31 512 -17 546
rect 17 512 31 546
rect -31 474 31 512
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect 205 461 239 575
rect 205 411 239 427
rect 353 970 369 988
rect 353 954 403 970
rect 649 1004 683 1020
rect 353 683 387 954
rect 353 461 387 649
rect 353 411 387 427
rect 649 757 683 970
rect 649 461 683 723
rect 871 1004 905 1020
rect 871 831 905 970
rect 1153 1004 1167 1038
rect 1201 1004 1215 1038
rect 1153 966 1215 1004
rect 1153 932 1167 966
rect 1201 932 1215 966
rect 1153 868 1215 932
rect 1315 1003 1349 1019
rect 649 411 683 427
rect 723 535 757 551
rect -31 368 -17 402
rect 17 368 31 402
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect 118 361 152 377
rect 312 361 346 377
rect 616 373 650 377
rect 152 327 215 361
rect 249 327 312 361
rect 118 289 152 327
rect 118 221 152 255
rect 312 289 346 327
rect 118 151 152 187
rect 118 101 152 117
rect 215 236 249 252
rect -31 62 31 80
rect 215 62 249 202
rect 312 221 346 255
rect 409 361 650 373
rect 409 339 616 361
rect 409 245 443 339
rect 409 195 443 211
rect 506 289 540 305
rect 506 221 540 255
rect 312 151 346 187
rect 506 151 540 187
rect 346 117 409 151
rect 443 117 506 151
rect 312 101 346 117
rect 506 101 540 117
rect 616 289 650 327
rect 723 262 757 501
rect 871 461 905 797
rect 871 411 905 427
rect 1153 546 1215 572
rect 1153 512 1167 546
rect 1201 512 1215 546
rect 1153 474 1215 512
rect 1153 440 1167 474
rect 1201 440 1215 474
rect 1153 402 1215 440
rect 1315 535 1349 969
rect 1389 979 1423 1105
rect 1477 1412 1511 1492
rect 1477 1344 1511 1378
rect 1477 1276 1511 1310
rect 1477 1208 1511 1242
rect 1477 1139 1511 1174
rect 1477 1083 1511 1105
rect 1597 1470 1659 1492
rect 1597 1436 1611 1470
rect 1645 1436 1659 1470
rect 1597 1398 1659 1436
rect 1597 1364 1611 1398
rect 1645 1364 1659 1398
rect 1597 1326 1659 1364
rect 1597 1292 1611 1326
rect 1645 1292 1659 1326
rect 1597 1254 1659 1292
rect 1597 1220 1611 1254
rect 1645 1220 1659 1254
rect 1597 1182 1659 1220
rect 1597 1148 1611 1182
rect 1645 1148 1659 1182
rect 1597 1110 1659 1148
rect 1597 1076 1611 1110
rect 1645 1076 1659 1110
rect 1597 1038 1659 1076
rect 1597 1004 1611 1038
rect 1645 1004 1659 1038
rect 1389 945 1497 979
rect 1315 461 1349 501
rect 1463 831 1497 945
rect 1597 966 1659 1004
rect 1597 932 1611 966
rect 1645 932 1659 966
rect 1597 868 1659 932
rect 1463 461 1497 797
rect 1315 411 1349 427
rect 1389 427 1497 461
rect 1597 546 1659 572
rect 1597 512 1611 546
rect 1645 512 1659 546
rect 1597 474 1659 512
rect 1597 440 1611 474
rect 1645 440 1659 474
rect 616 221 650 255
rect 713 245 757 262
rect 747 213 757 245
rect 810 361 844 377
rect 1004 361 1038 377
rect 844 327 907 361
rect 941 327 1004 361
rect 810 289 844 327
rect 810 221 844 255
rect 1004 289 1038 327
rect 713 195 747 211
rect 616 151 650 187
rect 810 151 844 187
rect 650 117 713 151
rect 747 117 810 151
rect 616 101 650 117
rect 810 101 844 117
rect 907 236 941 252
rect 907 62 941 202
rect 1004 221 1038 255
rect 1004 151 1038 187
rect 1004 101 1038 117
rect 1153 368 1167 402
rect 1201 368 1215 402
rect 1153 330 1215 368
rect 1153 296 1167 330
rect 1201 296 1215 330
rect 1153 258 1215 296
rect 1153 224 1167 258
rect 1201 224 1215 258
rect 1153 186 1215 224
rect 1153 152 1167 186
rect 1201 152 1215 186
rect 1153 114 1215 152
rect 1153 80 1167 114
rect 1201 80 1215 114
rect 1153 62 1215 80
rect 1293 361 1327 377
rect 1293 289 1327 327
rect 1293 221 1327 255
rect 1389 245 1423 427
rect 1597 402 1659 440
rect 1389 195 1423 211
rect 1487 361 1521 377
rect 1487 289 1521 327
rect 1487 221 1521 255
rect 1293 151 1327 187
rect 1487 151 1521 187
rect 1327 117 1389 151
rect 1423 117 1487 151
rect 1293 62 1327 117
rect 1390 62 1424 117
rect 1487 62 1521 117
rect 1597 368 1611 402
rect 1645 368 1659 402
rect 1597 330 1659 368
rect 1597 296 1611 330
rect 1645 296 1659 330
rect 1597 258 1659 296
rect 1597 224 1611 258
rect 1645 224 1659 258
rect 1597 186 1659 224
rect 1597 152 1611 186
rect 1645 152 1659 186
rect 1597 114 1659 152
rect 1597 80 1611 114
rect 1645 80 1659 114
rect 1597 62 1659 80
rect -31 47 1659 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 343 47
rect 377 13 415 47
rect 449 13 487 47
rect 521 13 585 47
rect 619 13 663 47
rect 697 13 735 47
rect 769 13 807 47
rect 841 13 879 47
rect 913 13 951 47
rect 985 13 1023 47
rect 1057 13 1095 47
rect 1129 13 1239 47
rect 1273 13 1311 47
rect 1345 13 1389 47
rect 1423 13 1467 47
rect 1501 13 1539 47
rect 1573 13 1659 47
rect -31 0 1659 13
<< viali >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 343 1505 377 1539
rect 415 1505 449 1539
rect 487 1505 521 1539
rect 585 1505 619 1539
rect 663 1505 697 1539
rect 735 1505 769 1539
rect 807 1505 841 1539
rect 879 1505 913 1539
rect 951 1505 985 1539
rect 1023 1505 1057 1539
rect 1095 1505 1129 1539
rect 1239 1505 1273 1539
rect 1311 1505 1345 1539
rect 1389 1505 1423 1539
rect 1467 1505 1501 1539
rect 1539 1505 1573 1539
rect 205 575 239 609
rect 353 649 387 683
rect 649 723 683 757
rect 871 797 905 831
rect 723 501 757 535
rect 1315 501 1349 535
rect 1463 797 1497 831
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 343 13 377 47
rect 415 13 449 47
rect 487 13 521 47
rect 585 13 619 47
rect 663 13 697 47
rect 735 13 769 47
rect 807 13 841 47
rect 879 13 913 47
rect 951 13 985 47
rect 1023 13 1057 47
rect 1095 13 1129 47
rect 1239 13 1273 47
rect 1311 13 1345 47
rect 1389 13 1423 47
rect 1467 13 1501 47
rect 1539 13 1573 47
<< metal1 >>
rect -31 1539 1659 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 343 1539
rect 377 1505 415 1539
rect 449 1505 487 1539
rect 521 1505 585 1539
rect 619 1505 663 1539
rect 697 1505 735 1539
rect 769 1505 807 1539
rect 841 1505 879 1539
rect 913 1505 951 1539
rect 985 1505 1023 1539
rect 1057 1505 1095 1539
rect 1129 1505 1239 1539
rect 1273 1505 1311 1539
rect 1345 1505 1389 1539
rect 1423 1505 1467 1539
rect 1501 1505 1539 1539
rect 1573 1505 1659 1539
rect -31 1492 1659 1505
rect 865 831 911 837
rect 1457 831 1503 837
rect 835 797 871 831
rect 905 797 917 831
rect 1451 797 1463 831
rect 1497 797 1533 831
rect 865 791 911 797
rect 1457 791 1503 797
rect 643 757 689 763
rect 613 723 649 757
rect 683 723 695 757
rect 643 717 689 723
rect 347 683 393 689
rect 317 649 353 683
rect 387 649 399 683
rect 347 643 393 649
rect 199 609 245 615
rect 169 575 205 609
rect 239 575 251 609
rect 199 569 245 575
rect 717 535 763 541
rect 1309 535 1355 541
rect 711 501 723 535
rect 757 501 1315 535
rect 1349 501 1361 535
rect 717 495 763 501
rect 1309 495 1355 501
rect -31 47 1659 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 343 47
rect 377 13 415 47
rect 449 13 487 47
rect 521 13 585 47
rect 619 13 663 47
rect 697 13 735 47
rect 769 13 807 47
rect 841 13 879 47
rect 913 13 951 47
rect 985 13 1023 47
rect 1057 13 1095 47
rect 1129 13 1239 47
rect 1273 13 1311 47
rect 1345 13 1389 47
rect 1423 13 1467 47
rect 1501 13 1539 47
rect 1573 13 1659 47
rect -31 0 1659 13
<< labels >>
rlabel metal1 1463 797 1497 831 1 Y
port 1 n
rlabel metal1 871 797 905 831 1 A
port 2 n
rlabel metal1 353 649 387 683 1 B
port 3 n
rlabel metal1 205 575 239 609 1 C
port 4 n
rlabel metal1 649 723 683 757 1 D
port 5 n
rlabel metal1 55 1505 89 1539 1 VDD
port 6 n
rlabel metal1 55 13 89 47 1 VSS
port 7 n
rlabel space 205 461 239 970 1 aoa4x1_pcell_0/C
rlabel space 353 461 387 988 1 aoa4x1_pcell_0/B
rlabel space 871 461 905 970 1 aoa4x1_pcell_0/A
rlabel space 649 461 683 970 1 aoa4x1_pcell_0/D
rlabel space 1463 427 1497 979 1 aoa4x1_pcell_0/Y
<< end >>
