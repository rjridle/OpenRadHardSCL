magic
tech sky130A
magscale 1 2
timestamp 1648751685
<< nwell >>
rect 55 1505 89 1539
<< psubdiffcont >>
rect 55 13 89 47
<< nsubdiffcont >>
rect 55 1505 89 1539
<< viali >>
rect 55 1505 89 1539
rect 55 13 89 47
<< metal1 >>
rect 427 945 461 979
rect 3349 978 11270 979
rect 479 947 11270 978
rect 3349 945 11270 947
rect 12079 945 12450 979
rect 13006 945 13775 979
rect 3495 797 3827 831
rect 6691 797 7477 831
rect 7741 797 8114 831
rect 11931 797 13041 831
rect 3348 649 14068 683
rect 7639 501 13263 535
rect 1279 427 9942 461
use li1_M1_contact  li1_M1_contact_9 pcells
timestamp 1648061256
transform -1 0 3478 0 -1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_10
timestamp 1648061256
transform 1 0 3848 0 1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform -1 0 3330 0 -1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform -1 0 4144 0 -1 666
box -53 -33 29 33
use dffx1_pcell  dffx1_pcell_0 pcells
timestamp 1648742316
transform 1 0 0 0 1 0
box -84 0 4376 1575
use dffx1_pcell  dffx1_pcell_1
timestamp 1648742316
transform 1 0 4292 0 1 0
box -84 0 4376 1575
use li1_M1_contact  li1_M1_contact_11
timestamp 1648061256
transform -1 0 7770 0 -1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_12
timestamp 1648061256
transform 1 0 8140 0 1 814
box -53 -33 29 33
use dffx1_pcell  dffx1_pcell_2
timestamp 1648742316
transform 1 0 8584 0 1 0
box -84 0 4376 1575
use li1_M1_contact  li1_M1_contact_3
timestamp 1648061256
transform 1 0 8436 0 1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_4
timestamp 1648061256
transform -1 0 7622 0 -1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_8
timestamp 1648061256
transform 1 0 13246 0 -1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_7
timestamp 1648061256
transform 1 0 13024 0 -1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_5
timestamp 1648061256
transform -1 0 12062 0 -1 962
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_6
timestamp 1648061256
transform 1 0 12432 0 1 962
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_15
timestamp 1648061256
transform -1 0 12728 0 1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_13
timestamp 1648061256
transform -1 0 11914 0 -1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_2
timestamp 1648061256
transform 1 0 14060 0 -1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_16
timestamp 1648061256
transform -1 0 15170 0 -1 814
box -53 -33 29 33
use voter3x1_pcell  voter3x1_pcell_0 pcells
timestamp 1648740352
transform 1 0 12876 0 1 0
box -84 0 2526 1575
<< labels >>
rlabel metal1 1315 427 1349 461 1 D
port 2 n
rlabel metal1 427 945 461 979 1 CLK
port 3 n
rlabel metal1 72 1522 72 1522 1 VDD
port 4 n
rlabel metal1 72 30 72 30 1 VSS
port 5 n
rlabel metal1 15153 797 15187 831 1 Q
port 1 n
<< end >>
