magic
tech sky130A
magscale 1 2
timestamp 1651071491
<< metal1 >>
rect -31 1492 1363 1554
rect 1167 797 1201 831
rect 1019 723 1053 757
rect 353 649 387 683
rect 205 575 239 609
rect -31 0 1363 62
use aoi3x1_pcell  aoi3x1_pcell_0 pcells
timestamp 1648661061
transform 1 0 0 0 1 0
box -84 0 1416 1575
use li1_M1_contact  li1_M1_contact_1 pcells
timestamp 1648061256
transform 1 0 222 0 1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform 1 0 370 0 1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_2
timestamp 1648061256
transform 1 0 1036 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_3
timestamp 1648061256
transform -1 0 1184 0 -1 814
box -53 -33 29 33
<< labels >>
rlabel metal1 1167 797 1201 831 1 YN
port 1 n
rlabel metal1 205 575 239 609 1 A
port 2 n
rlabel metal1 353 649 387 683 1 B
port 3 n
rlabel metal1 1019 723 1053 757 1 C
port 4 n
rlabel metal1 -31 1492 1363 1554 1 VDD
port 5 n
rlabel metal1 -31 0 1363 62 1 GND
port 6 n
<< end >>
