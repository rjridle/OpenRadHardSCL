* SPICE3 file created from DFFSNX1.ext - technology: sky130A

.subckt DFFSNX1 CLK SN Q QN D VDD VSS
X0 VDD D a_217_1050# VDD sky130_fd_pr__pfet_01v8 ad=1.182p pd=9.582u as=0p ps=0u w=2u l=0.15u M=2
X1 VDD SN a_1905_1050# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X2 VDD SN Q VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.74p ps=1.374u w=2u l=0.15u M=2
X3 a_1265_989# a_1905_1050# a_2702_101# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X4 a_1905_1050# a_217_1050# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X5 VDD QN Q VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X6 VDD a_343_411# a_217_1050# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X7 VDD CLK a_343_411# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X8 a_1905_1050# SN a_2000_210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X9 VDD a_217_1050# a_343_411# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X10 QN Q VDD VDD sky130_fd_pr__pfet_01v8 ad=1.16p pd=9.16u as=0p ps=0u w=2u l=0.15u M=2
X11 VDD CLK a_1265_989# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X12 Q QN a_3628_210# VSS sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=0p ps=0u w=3u l=0.15u
X13 VSS a_343_411# a_4330_101# VSS sky130_fd_pr__nfet_01v8 ad=1.0746p pd=9.42u as=0p ps=0u w=3u l=0.15u
X14 a_343_411# a_1265_989# a_1038_210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X15 Q a_1265_989# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X16 VSS CLK a_757_103# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X17 VDD a_1265_989# a_343_411# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X18 VSS D a_112_101# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X19 a_3628_210# a_1265_989# a_3347_103# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X20 VSS SN a_3347_103# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X21 a_1905_1050# a_1265_989# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X22 VSS a_217_1050# a_1719_103# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X23 QN Q a_4330_101# VSS sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=0p ps=0u w=3u l=0.15u
X24 a_1038_210# a_217_1050# a_757_103# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X25 VDD a_343_411# QN VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X26 VSS CLK a_2702_101# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X27 a_217_1050# a_343_411# a_112_101# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X28 VDD a_1905_1050# a_1265_989# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X29 a_2000_210# a_1265_989# a_1719_103# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
C0 VDD CLK 2.46fF
C1 QN VDD 2.14fF
C2 a_1905_1050# VDD 2.82fF
C3 a_217_1050# VDD 2.50fF
C4 a_1265_989# VDD 2.71fF
C5 Q VDD 2.82fF
C6 a_343_411# VDD 3.14fF
C7 VDD VSS 7.98fF
.ends
