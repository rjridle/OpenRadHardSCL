magic
tech sky130
magscale 1 2
timestamp 1651261209
<< nwell >>
rect 55 1505 89 1539
<< pwell >>
rect 55 13 89 47
<< psubdiffcont >>
rect 55 13 89 47
<< nsubdiffcont >>
rect 55 1505 89 1539
<< viali >>
rect 55 1505 89 1539
rect 55 13 89 47
<< metal1 >>
rect -31 1539 17125 1554
rect -31 1505 55 1539
rect 89 1505 17125 1539
rect -31 1492 17125 1505
rect 1090 945 12712 979
rect 13561 945 13878 979
rect 3813 871 4132 905
rect 8629 871 8975 905
rect 13413 871 15028 905
rect 16929 797 16963 831
rect 8522 723 14821 757
rect 3606 649 15819 683
rect 2047 501 14146 535
rect 205 427 239 461
rect 240 427 10019 461
rect -31 47 17125 62
rect -31 13 55 47
rect 89 13 17125 47
rect -31 0 17125 13
use dffsnx1_pcell  dffsnx1_pcell_0 pcells
timestamp 1651259636
transform 1 0 0 0 1 0
box -84 0 4968 1575
use dffsnx1_pcell  dffsnx1_pcell_1
timestamp 1651259636
transform 1 0 4884 0 1 0
box -84 0 4968 1575
use li1_M1_contact  li1_M1_contact_12 pcells
timestamp 1648061256
transform -1 0 4736 0 -1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_18
timestamp 1648061256
transform 1 0 4144 0 1 888
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_13
timestamp 1648061256
transform -1 0 3774 0 -1 888
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_20
timestamp 1648061256
transform -1 0 3626 0 -1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_5
timestamp 1648061256
transform 1 0 4588 0 1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_7
timestamp 1648061256
transform -1 0 222 0 -1 444
box -53 -33 29 33
use dffsnx1_pcell  dffsnx1_pcell_2
timestamp 1651259636
transform 1 0 9768 0 1 0
box -84 0 4968 1575
use li1_M1_contact  li1_M1_contact_9
timestamp 1648061256
transform 1 0 9620 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_4
timestamp 1648061256
transform 1 0 9028 0 1 888
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_3
timestamp 1648061256
transform -1 0 8658 0 -1 888
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_6
timestamp 1648061256
transform -1 0 8510 0 -1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_15
timestamp 1648061256
transform -1 0 5106 0 -1 444
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_8
timestamp 1648061256
transform 1 0 9990 0 1 444
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_10
timestamp 1648061256
transform 1 0 9472 0 1 814
box -53 -33 29 33
use voter3x1_pcell  voter3x1_pcell_0 pcells
timestamp 1651259615
transform 1 0 14652 0 1 0
box -84 0 2526 1575
use li1_M1_contact  li1_M1_contact_14
timestamp 1648061256
transform 1 0 14800 0 -1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_2
timestamp 1648061256
transform -1 0 13542 0 -1 962
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform 1 0 13912 0 1 962
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_11
timestamp 1648061256
transform 1 0 14504 0 1 888
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform -1 0 13394 0 -1 888
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_19
timestamp 1648061256
transform 1 0 14356 0 1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_16
timestamp 1648061256
transform 1 0 15836 0 -1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_17
timestamp 1648061256
transform -1 0 16946 0 -1 814
box -53 -33 29 33
<< labels >>
rlabel metal1 16929 797 16963 831 1 Q
port 1 nsew signal output
rlabel metal1 205 427 239 461 1 D
port 2 nsew signal input
rlabel metal1 1093 945 1127 979 1 CLK
port 3 nsew signal input
rlabel metal1 2055 501 2089 535 1 SN
port 4 nsew signal input
rlabel metal1 -31 1492 17125 1554 1 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 -31 0 17125 62 1 VGND
port 6 nsew ground bidirectional abutment
rlabel nwell 55 1505 89 1539 1 VPB
port 7 nsew power bidirectional
rlabel pwell 55 13 89 47 1 VNB
port 8 nsew ground bidirectional
<< end >>
