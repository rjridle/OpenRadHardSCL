magic
tech sky130A
magscale 1 2
timestamp 1649361818
<< nwell >>
rect -84 832 5856 1575
<< nmos >>
rect 147 318 177 379
tri 177 318 193 334 sw
rect 447 318 477 379
rect 147 288 253 318
tri 253 288 283 318 sw
rect 147 187 177 288
tri 177 272 193 288 nw
tri 237 272 253 288 ne
tri 177 187 193 203 sw
tri 237 187 253 203 se
rect 253 187 283 288
tri 342 288 372 318 se
rect 372 288 477 318
rect 342 194 372 288
tri 372 272 388 288 nw
tri 431 272 447 288 ne
tri 372 194 388 210 sw
tri 431 194 447 210 se
rect 447 194 477 288
tri 147 157 177 187 ne
rect 177 157 253 187
tri 253 157 283 187 nw
tri 342 164 372 194 ne
rect 372 164 447 194
tri 447 164 477 194 nw
rect 649 326 679 379
tri 679 326 695 342 sw
rect 649 296 755 326
tri 755 296 785 326 sw
rect 649 195 679 296
tri 679 280 695 296 nw
tri 739 280 755 296 ne
tri 679 195 695 211 sw
tri 739 195 755 211 se
rect 755 195 785 296
tri 649 165 679 195 ne
rect 679 165 755 195
tri 755 165 785 195 nw
rect 1109 318 1139 379
tri 1139 318 1155 334 sw
rect 1409 318 1439 379
rect 1109 288 1215 318
tri 1215 288 1245 318 sw
rect 1109 187 1139 288
tri 1139 272 1155 288 nw
tri 1199 272 1215 288 ne
tri 1139 187 1155 203 sw
tri 1199 187 1215 203 se
rect 1215 187 1245 288
tri 1304 288 1334 318 se
rect 1334 288 1439 318
rect 1304 194 1334 288
tri 1334 272 1350 288 nw
tri 1393 272 1409 288 ne
tri 1334 194 1350 210 sw
tri 1393 194 1409 210 se
rect 1409 194 1439 288
tri 1109 157 1139 187 ne
rect 1139 157 1215 187
tri 1215 157 1245 187 nw
tri 1304 164 1334 194 ne
rect 1334 164 1409 194
tri 1409 164 1439 194 nw
rect 1611 326 1641 379
tri 1641 326 1657 342 sw
rect 1611 296 1717 326
tri 1717 296 1747 326 sw
rect 1611 195 1641 296
tri 1641 280 1657 296 nw
tri 1701 280 1717 296 ne
tri 1641 195 1657 211 sw
tri 1701 195 1717 211 se
rect 1717 195 1747 296
tri 1611 165 1641 195 ne
rect 1641 165 1717 195
tri 1717 165 1747 195 nw
rect 2071 318 2101 379
tri 2101 318 2117 334 sw
rect 2371 318 2401 379
rect 2071 288 2177 318
tri 2177 288 2207 318 sw
rect 2071 187 2101 288
tri 2101 272 2117 288 nw
tri 2161 272 2177 288 ne
tri 2101 187 2117 203 sw
tri 2161 187 2177 203 se
rect 2177 187 2207 288
tri 2266 288 2296 318 se
rect 2296 288 2401 318
rect 2266 194 2296 288
tri 2296 272 2312 288 nw
tri 2355 272 2371 288 ne
tri 2296 194 2312 210 sw
tri 2355 194 2371 210 se
rect 2371 194 2401 288
tri 2071 157 2101 187 ne
rect 2101 157 2177 187
tri 2177 157 2207 187 nw
tri 2266 164 2296 194 ne
rect 2296 164 2371 194
tri 2371 164 2401 194 nw
rect 2573 326 2603 379
tri 2603 326 2619 342 sw
rect 2573 296 2679 326
tri 2679 296 2709 326 sw
rect 2573 195 2603 296
tri 2603 280 2619 296 nw
tri 2663 280 2679 296 ne
tri 2603 195 2619 211 sw
tri 2663 195 2679 211 se
rect 2679 195 2709 296
tri 2573 165 2603 195 ne
rect 2603 165 2679 195
tri 2679 165 2709 195 nw
rect 3033 318 3063 379
tri 3063 318 3079 334 sw
rect 3333 318 3363 379
rect 3033 288 3139 318
tri 3139 288 3169 318 sw
rect 3033 187 3063 288
tri 3063 272 3079 288 nw
tri 3123 272 3139 288 ne
tri 3063 187 3079 203 sw
tri 3123 187 3139 203 se
rect 3139 187 3169 288
tri 3228 288 3258 318 se
rect 3258 288 3363 318
rect 3228 194 3258 288
tri 3258 272 3274 288 nw
tri 3317 272 3333 288 ne
tri 3258 194 3274 210 sw
tri 3317 194 3333 210 se
rect 3333 194 3363 288
tri 3033 157 3063 187 ne
rect 3063 157 3139 187
tri 3139 157 3169 187 nw
tri 3228 164 3258 194 ne
rect 3258 164 3333 194
tri 3333 164 3363 194 nw
rect 3535 326 3565 379
tri 3565 326 3581 342 sw
rect 3535 296 3641 326
tri 3641 296 3671 326 sw
rect 3535 195 3565 296
tri 3565 280 3581 296 nw
tri 3625 280 3641 296 ne
tri 3565 195 3581 211 sw
tri 3625 195 3641 211 se
rect 3641 195 3671 296
tri 3535 165 3565 195 ne
rect 3565 165 3641 195
tri 3641 165 3671 195 nw
rect 3995 318 4025 379
tri 4025 318 4041 334 sw
rect 4295 318 4325 379
rect 3995 288 4101 318
tri 4101 288 4131 318 sw
rect 3995 187 4025 288
tri 4025 272 4041 288 nw
tri 4085 272 4101 288 ne
tri 4025 187 4041 203 sw
tri 4085 187 4101 203 se
rect 4101 187 4131 288
tri 4190 288 4220 318 se
rect 4220 288 4325 318
rect 4190 194 4220 288
tri 4220 272 4236 288 nw
tri 4279 272 4295 288 ne
tri 4220 194 4236 210 sw
tri 4279 194 4295 210 se
rect 4295 194 4325 288
tri 3995 157 4025 187 ne
rect 4025 157 4101 187
tri 4101 157 4131 187 nw
tri 4190 164 4220 194 ne
rect 4220 164 4295 194
tri 4295 164 4325 194 nw
rect 4497 326 4527 379
tri 4527 326 4543 342 sw
rect 4497 296 4603 326
tri 4603 296 4633 326 sw
rect 4497 195 4527 296
tri 4527 280 4543 296 nw
tri 4587 280 4603 296 ne
tri 4527 195 4543 211 sw
tri 4587 195 4603 211 se
rect 4603 195 4633 296
tri 4497 165 4527 195 ne
rect 4527 165 4603 195
tri 4603 165 4633 195 nw
rect 4957 318 4987 379
tri 4987 318 5003 334 sw
rect 5257 318 5287 379
rect 4957 288 5063 318
tri 5063 288 5093 318 sw
rect 4957 187 4987 288
tri 4987 272 5003 288 nw
tri 5047 272 5063 288 ne
tri 4987 187 5003 203 sw
tri 5047 187 5063 203 se
rect 5063 187 5093 288
tri 5152 288 5182 318 se
rect 5182 288 5287 318
rect 5152 194 5182 288
tri 5182 272 5198 288 nw
tri 5241 272 5257 288 ne
tri 5182 194 5198 210 sw
tri 5241 194 5257 210 se
rect 5257 194 5287 288
tri 4957 157 4987 187 ne
rect 4987 157 5063 187
tri 5063 157 5093 187 nw
tri 5152 164 5182 194 ne
rect 5182 164 5257 194
tri 5257 164 5287 194 nw
rect 5459 326 5489 379
tri 5489 326 5505 342 sw
rect 5459 296 5565 326
tri 5565 296 5595 326 sw
rect 5459 195 5489 296
tri 5489 280 5505 296 nw
tri 5549 280 5565 296 ne
tri 5489 195 5505 211 sw
tri 5549 195 5565 211 se
rect 5565 195 5595 296
tri 5459 165 5489 195 ne
rect 5489 165 5565 195
tri 5565 165 5595 195 nw
<< pmos >>
rect 247 1050 277 1450
rect 335 1050 365 1450
rect 423 1050 453 1450
rect 511 1050 541 1450
rect 599 1050 629 1450
rect 687 1050 717 1450
rect 1209 1050 1239 1450
rect 1297 1050 1327 1450
rect 1385 1050 1415 1450
rect 1473 1050 1503 1450
rect 1561 1050 1591 1450
rect 1649 1050 1679 1450
rect 2171 1050 2201 1450
rect 2259 1050 2289 1450
rect 2347 1050 2377 1450
rect 2435 1050 2465 1450
rect 2523 1050 2553 1450
rect 2611 1050 2641 1450
rect 3133 1050 3163 1450
rect 3221 1050 3251 1450
rect 3309 1050 3339 1450
rect 3397 1050 3427 1450
rect 3485 1050 3515 1450
rect 3573 1050 3603 1450
rect 4095 1050 4125 1450
rect 4183 1050 4213 1450
rect 4271 1050 4301 1450
rect 4359 1050 4389 1450
rect 4447 1050 4477 1450
rect 4535 1050 4565 1450
rect 5057 1050 5087 1450
rect 5145 1050 5175 1450
rect 5233 1050 5263 1450
rect 5321 1050 5351 1450
rect 5409 1050 5439 1450
rect 5497 1050 5527 1450
<< ndiff >>
rect 91 363 147 379
rect 91 329 101 363
rect 135 329 147 363
rect 91 291 147 329
rect 177 363 447 379
rect 177 334 198 363
tri 177 318 193 334 ne
rect 193 329 198 334
rect 232 329 295 363
rect 329 329 392 363
rect 426 329 447 363
rect 193 318 447 329
rect 477 363 533 379
rect 477 329 489 363
rect 523 329 533 363
rect 91 257 101 291
rect 135 257 147 291
tri 253 288 283 318 ne
rect 283 291 342 318
rect 91 223 147 257
rect 91 189 101 223
rect 135 189 147 223
rect 91 157 147 189
tri 177 272 193 288 se
rect 193 272 237 288
tri 237 272 253 288 sw
rect 177 238 253 272
rect 177 204 198 238
rect 232 204 253 238
rect 177 203 253 204
tri 177 187 193 203 ne
rect 193 187 237 203
tri 237 187 253 203 nw
rect 283 257 295 291
rect 329 257 342 291
tri 342 288 372 318 nw
rect 283 223 342 257
rect 283 189 295 223
rect 329 189 342 223
tri 372 272 388 288 se
rect 388 272 431 288
tri 431 272 447 288 sw
rect 372 244 447 272
rect 372 210 393 244
rect 427 210 447 244
tri 372 194 388 210 ne
rect 388 194 431 210
tri 431 194 447 210 nw
tri 147 157 177 187 sw
tri 253 157 283 187 se
rect 283 164 342 189
tri 342 164 372 194 sw
tri 447 164 477 194 se
rect 477 164 533 329
rect 283 157 533 164
rect 91 153 533 157
rect 91 119 101 153
rect 135 119 295 153
rect 329 119 392 153
rect 426 119 489 153
rect 523 119 533 153
rect 91 103 533 119
rect 593 363 649 379
rect 593 329 603 363
rect 637 329 649 363
rect 593 291 649 329
rect 679 342 841 379
tri 679 326 695 342 ne
rect 695 326 841 342
tri 755 296 785 326 ne
rect 593 257 603 291
rect 637 257 649 291
rect 593 223 649 257
rect 593 189 603 223
rect 637 189 649 223
tri 679 280 695 296 se
rect 695 280 739 296
tri 739 280 755 296 sw
rect 679 247 755 280
rect 679 213 700 247
rect 734 213 755 247
rect 679 211 755 213
tri 679 195 695 211 ne
rect 695 195 739 211
tri 739 195 755 211 nw
rect 785 291 841 326
rect 785 257 797 291
rect 831 257 841 291
rect 785 223 841 257
rect 593 165 649 189
tri 649 165 679 195 sw
tri 755 165 785 195 se
rect 785 189 797 223
rect 831 189 841 223
rect 785 165 841 189
rect 593 153 841 165
rect 593 119 603 153
rect 637 119 700 153
rect 734 119 797 153
rect 831 119 841 153
rect 593 103 841 119
rect 1053 363 1109 379
rect 1053 329 1063 363
rect 1097 329 1109 363
rect 1053 291 1109 329
rect 1139 363 1409 379
rect 1139 334 1160 363
tri 1139 318 1155 334 ne
rect 1155 329 1160 334
rect 1194 329 1257 363
rect 1291 329 1354 363
rect 1388 329 1409 363
rect 1155 318 1409 329
rect 1439 363 1495 379
rect 1439 329 1451 363
rect 1485 329 1495 363
rect 1053 257 1063 291
rect 1097 257 1109 291
tri 1215 288 1245 318 ne
rect 1245 291 1304 318
rect 1053 223 1109 257
rect 1053 189 1063 223
rect 1097 189 1109 223
rect 1053 157 1109 189
tri 1139 272 1155 288 se
rect 1155 272 1199 288
tri 1199 272 1215 288 sw
rect 1139 238 1215 272
rect 1139 204 1160 238
rect 1194 204 1215 238
rect 1139 203 1215 204
tri 1139 187 1155 203 ne
rect 1155 187 1199 203
tri 1199 187 1215 203 nw
rect 1245 257 1257 291
rect 1291 257 1304 291
tri 1304 288 1334 318 nw
rect 1245 223 1304 257
rect 1245 189 1257 223
rect 1291 189 1304 223
tri 1334 272 1350 288 se
rect 1350 272 1393 288
tri 1393 272 1409 288 sw
rect 1334 244 1409 272
rect 1334 210 1355 244
rect 1389 210 1409 244
tri 1334 194 1350 210 ne
rect 1350 194 1393 210
tri 1393 194 1409 210 nw
tri 1109 157 1139 187 sw
tri 1215 157 1245 187 se
rect 1245 164 1304 189
tri 1304 164 1334 194 sw
tri 1409 164 1439 194 se
rect 1439 164 1495 329
rect 1245 157 1495 164
rect 1053 153 1495 157
rect 1053 119 1063 153
rect 1097 119 1257 153
rect 1291 119 1354 153
rect 1388 119 1451 153
rect 1485 119 1495 153
rect 1053 103 1495 119
rect 1555 363 1611 379
rect 1555 329 1565 363
rect 1599 329 1611 363
rect 1555 291 1611 329
rect 1641 342 1803 379
tri 1641 326 1657 342 ne
rect 1657 326 1803 342
tri 1717 296 1747 326 ne
rect 1555 257 1565 291
rect 1599 257 1611 291
rect 1555 223 1611 257
rect 1555 189 1565 223
rect 1599 189 1611 223
tri 1641 280 1657 296 se
rect 1657 280 1701 296
tri 1701 280 1717 296 sw
rect 1641 247 1717 280
rect 1641 213 1662 247
rect 1696 213 1717 247
rect 1641 211 1717 213
tri 1641 195 1657 211 ne
rect 1657 195 1701 211
tri 1701 195 1717 211 nw
rect 1747 291 1803 326
rect 1747 257 1759 291
rect 1793 257 1803 291
rect 1747 223 1803 257
rect 1555 165 1611 189
tri 1611 165 1641 195 sw
tri 1717 165 1747 195 se
rect 1747 189 1759 223
rect 1793 189 1803 223
rect 1747 165 1803 189
rect 1555 153 1803 165
rect 1555 119 1565 153
rect 1599 119 1662 153
rect 1696 119 1759 153
rect 1793 119 1803 153
rect 1555 103 1803 119
rect 2015 363 2071 379
rect 2015 329 2025 363
rect 2059 329 2071 363
rect 2015 291 2071 329
rect 2101 363 2371 379
rect 2101 334 2122 363
tri 2101 318 2117 334 ne
rect 2117 329 2122 334
rect 2156 329 2219 363
rect 2253 329 2316 363
rect 2350 329 2371 363
rect 2117 318 2371 329
rect 2401 363 2457 379
rect 2401 329 2413 363
rect 2447 329 2457 363
rect 2015 257 2025 291
rect 2059 257 2071 291
tri 2177 288 2207 318 ne
rect 2207 291 2266 318
rect 2015 223 2071 257
rect 2015 189 2025 223
rect 2059 189 2071 223
rect 2015 157 2071 189
tri 2101 272 2117 288 se
rect 2117 272 2161 288
tri 2161 272 2177 288 sw
rect 2101 238 2177 272
rect 2101 204 2122 238
rect 2156 204 2177 238
rect 2101 203 2177 204
tri 2101 187 2117 203 ne
rect 2117 187 2161 203
tri 2161 187 2177 203 nw
rect 2207 257 2219 291
rect 2253 257 2266 291
tri 2266 288 2296 318 nw
rect 2207 223 2266 257
rect 2207 189 2219 223
rect 2253 189 2266 223
tri 2296 272 2312 288 se
rect 2312 272 2355 288
tri 2355 272 2371 288 sw
rect 2296 244 2371 272
rect 2296 210 2317 244
rect 2351 210 2371 244
tri 2296 194 2312 210 ne
rect 2312 194 2355 210
tri 2355 194 2371 210 nw
tri 2071 157 2101 187 sw
tri 2177 157 2207 187 se
rect 2207 164 2266 189
tri 2266 164 2296 194 sw
tri 2371 164 2401 194 se
rect 2401 164 2457 329
rect 2207 157 2457 164
rect 2015 153 2457 157
rect 2015 119 2025 153
rect 2059 119 2219 153
rect 2253 119 2316 153
rect 2350 119 2413 153
rect 2447 119 2457 153
rect 2015 103 2457 119
rect 2517 363 2573 379
rect 2517 329 2527 363
rect 2561 329 2573 363
rect 2517 291 2573 329
rect 2603 342 2765 379
tri 2603 326 2619 342 ne
rect 2619 326 2765 342
tri 2679 296 2709 326 ne
rect 2517 257 2527 291
rect 2561 257 2573 291
rect 2517 223 2573 257
rect 2517 189 2527 223
rect 2561 189 2573 223
tri 2603 280 2619 296 se
rect 2619 280 2663 296
tri 2663 280 2679 296 sw
rect 2603 247 2679 280
rect 2603 213 2624 247
rect 2658 213 2679 247
rect 2603 211 2679 213
tri 2603 195 2619 211 ne
rect 2619 195 2663 211
tri 2663 195 2679 211 nw
rect 2709 291 2765 326
rect 2709 257 2721 291
rect 2755 257 2765 291
rect 2709 223 2765 257
rect 2517 165 2573 189
tri 2573 165 2603 195 sw
tri 2679 165 2709 195 se
rect 2709 189 2721 223
rect 2755 189 2765 223
rect 2709 165 2765 189
rect 2517 153 2765 165
rect 2517 119 2527 153
rect 2561 119 2624 153
rect 2658 119 2721 153
rect 2755 119 2765 153
rect 2517 103 2765 119
rect 2977 363 3033 379
rect 2977 329 2987 363
rect 3021 329 3033 363
rect 2977 291 3033 329
rect 3063 363 3333 379
rect 3063 334 3084 363
tri 3063 318 3079 334 ne
rect 3079 329 3084 334
rect 3118 329 3181 363
rect 3215 329 3278 363
rect 3312 329 3333 363
rect 3079 318 3333 329
rect 3363 363 3419 379
rect 3363 329 3375 363
rect 3409 329 3419 363
rect 2977 257 2987 291
rect 3021 257 3033 291
tri 3139 288 3169 318 ne
rect 3169 291 3228 318
rect 2977 223 3033 257
rect 2977 189 2987 223
rect 3021 189 3033 223
rect 2977 157 3033 189
tri 3063 272 3079 288 se
rect 3079 272 3123 288
tri 3123 272 3139 288 sw
rect 3063 238 3139 272
rect 3063 204 3084 238
rect 3118 204 3139 238
rect 3063 203 3139 204
tri 3063 187 3079 203 ne
rect 3079 187 3123 203
tri 3123 187 3139 203 nw
rect 3169 257 3181 291
rect 3215 257 3228 291
tri 3228 288 3258 318 nw
rect 3169 223 3228 257
rect 3169 189 3181 223
rect 3215 189 3228 223
tri 3258 272 3274 288 se
rect 3274 272 3317 288
tri 3317 272 3333 288 sw
rect 3258 244 3333 272
rect 3258 210 3279 244
rect 3313 210 3333 244
tri 3258 194 3274 210 ne
rect 3274 194 3317 210
tri 3317 194 3333 210 nw
tri 3033 157 3063 187 sw
tri 3139 157 3169 187 se
rect 3169 164 3228 189
tri 3228 164 3258 194 sw
tri 3333 164 3363 194 se
rect 3363 164 3419 329
rect 3169 157 3419 164
rect 2977 153 3419 157
rect 2977 119 2987 153
rect 3021 119 3181 153
rect 3215 119 3278 153
rect 3312 119 3375 153
rect 3409 119 3419 153
rect 2977 103 3419 119
rect 3479 363 3535 379
rect 3479 329 3489 363
rect 3523 329 3535 363
rect 3479 291 3535 329
rect 3565 342 3727 379
tri 3565 326 3581 342 ne
rect 3581 326 3727 342
tri 3641 296 3671 326 ne
rect 3479 257 3489 291
rect 3523 257 3535 291
rect 3479 223 3535 257
rect 3479 189 3489 223
rect 3523 189 3535 223
tri 3565 280 3581 296 se
rect 3581 280 3625 296
tri 3625 280 3641 296 sw
rect 3565 247 3641 280
rect 3565 213 3586 247
rect 3620 213 3641 247
rect 3565 211 3641 213
tri 3565 195 3581 211 ne
rect 3581 195 3625 211
tri 3625 195 3641 211 nw
rect 3671 291 3727 326
rect 3671 257 3683 291
rect 3717 257 3727 291
rect 3671 223 3727 257
rect 3479 165 3535 189
tri 3535 165 3565 195 sw
tri 3641 165 3671 195 se
rect 3671 189 3683 223
rect 3717 189 3727 223
rect 3671 165 3727 189
rect 3479 153 3727 165
rect 3479 119 3489 153
rect 3523 119 3586 153
rect 3620 119 3683 153
rect 3717 119 3727 153
rect 3479 103 3727 119
rect 3939 363 3995 379
rect 3939 329 3949 363
rect 3983 329 3995 363
rect 3939 291 3995 329
rect 4025 363 4295 379
rect 4025 334 4046 363
tri 4025 318 4041 334 ne
rect 4041 329 4046 334
rect 4080 329 4143 363
rect 4177 329 4240 363
rect 4274 329 4295 363
rect 4041 318 4295 329
rect 4325 363 4381 379
rect 4325 329 4337 363
rect 4371 329 4381 363
rect 3939 257 3949 291
rect 3983 257 3995 291
tri 4101 288 4131 318 ne
rect 4131 291 4190 318
rect 3939 223 3995 257
rect 3939 189 3949 223
rect 3983 189 3995 223
rect 3939 157 3995 189
tri 4025 272 4041 288 se
rect 4041 272 4085 288
tri 4085 272 4101 288 sw
rect 4025 238 4101 272
rect 4025 204 4046 238
rect 4080 204 4101 238
rect 4025 203 4101 204
tri 4025 187 4041 203 ne
rect 4041 187 4085 203
tri 4085 187 4101 203 nw
rect 4131 257 4143 291
rect 4177 257 4190 291
tri 4190 288 4220 318 nw
rect 4131 223 4190 257
rect 4131 189 4143 223
rect 4177 189 4190 223
tri 4220 272 4236 288 se
rect 4236 272 4279 288
tri 4279 272 4295 288 sw
rect 4220 244 4295 272
rect 4220 210 4241 244
rect 4275 210 4295 244
tri 4220 194 4236 210 ne
rect 4236 194 4279 210
tri 4279 194 4295 210 nw
tri 3995 157 4025 187 sw
tri 4101 157 4131 187 se
rect 4131 164 4190 189
tri 4190 164 4220 194 sw
tri 4295 164 4325 194 se
rect 4325 164 4381 329
rect 4131 157 4381 164
rect 3939 153 4381 157
rect 3939 119 3949 153
rect 3983 119 4143 153
rect 4177 119 4240 153
rect 4274 119 4337 153
rect 4371 119 4381 153
rect 3939 103 4381 119
rect 4441 363 4497 379
rect 4441 329 4451 363
rect 4485 329 4497 363
rect 4441 291 4497 329
rect 4527 342 4689 379
tri 4527 326 4543 342 ne
rect 4543 326 4689 342
tri 4603 296 4633 326 ne
rect 4441 257 4451 291
rect 4485 257 4497 291
rect 4441 223 4497 257
rect 4441 189 4451 223
rect 4485 189 4497 223
tri 4527 280 4543 296 se
rect 4543 280 4587 296
tri 4587 280 4603 296 sw
rect 4527 247 4603 280
rect 4527 213 4548 247
rect 4582 213 4603 247
rect 4527 211 4603 213
tri 4527 195 4543 211 ne
rect 4543 195 4587 211
tri 4587 195 4603 211 nw
rect 4633 291 4689 326
rect 4633 257 4645 291
rect 4679 257 4689 291
rect 4633 223 4689 257
rect 4441 165 4497 189
tri 4497 165 4527 195 sw
tri 4603 165 4633 195 se
rect 4633 189 4645 223
rect 4679 189 4689 223
rect 4633 165 4689 189
rect 4441 153 4689 165
rect 4441 119 4451 153
rect 4485 119 4548 153
rect 4582 119 4645 153
rect 4679 119 4689 153
rect 4441 103 4689 119
rect 4901 363 4957 379
rect 4901 329 4911 363
rect 4945 329 4957 363
rect 4901 291 4957 329
rect 4987 363 5257 379
rect 4987 334 5008 363
tri 4987 318 5003 334 ne
rect 5003 329 5008 334
rect 5042 329 5105 363
rect 5139 329 5202 363
rect 5236 329 5257 363
rect 5003 318 5257 329
rect 5287 363 5343 379
rect 5287 329 5299 363
rect 5333 329 5343 363
rect 4901 257 4911 291
rect 4945 257 4957 291
tri 5063 288 5093 318 ne
rect 5093 291 5152 318
rect 4901 223 4957 257
rect 4901 189 4911 223
rect 4945 189 4957 223
rect 4901 157 4957 189
tri 4987 272 5003 288 se
rect 5003 272 5047 288
tri 5047 272 5063 288 sw
rect 4987 238 5063 272
rect 4987 204 5008 238
rect 5042 204 5063 238
rect 4987 203 5063 204
tri 4987 187 5003 203 ne
rect 5003 187 5047 203
tri 5047 187 5063 203 nw
rect 5093 257 5105 291
rect 5139 257 5152 291
tri 5152 288 5182 318 nw
rect 5093 223 5152 257
rect 5093 189 5105 223
rect 5139 189 5152 223
tri 5182 272 5198 288 se
rect 5198 272 5241 288
tri 5241 272 5257 288 sw
rect 5182 244 5257 272
rect 5182 210 5203 244
rect 5237 210 5257 244
tri 5182 194 5198 210 ne
rect 5198 194 5241 210
tri 5241 194 5257 210 nw
tri 4957 157 4987 187 sw
tri 5063 157 5093 187 se
rect 5093 164 5152 189
tri 5152 164 5182 194 sw
tri 5257 164 5287 194 se
rect 5287 164 5343 329
rect 5093 157 5343 164
rect 4901 153 5343 157
rect 4901 119 4911 153
rect 4945 119 5105 153
rect 5139 119 5202 153
rect 5236 119 5299 153
rect 5333 119 5343 153
rect 4901 103 5343 119
rect 5403 363 5459 379
rect 5403 329 5413 363
rect 5447 329 5459 363
rect 5403 291 5459 329
rect 5489 342 5651 379
tri 5489 326 5505 342 ne
rect 5505 326 5651 342
tri 5565 296 5595 326 ne
rect 5403 257 5413 291
rect 5447 257 5459 291
rect 5403 223 5459 257
rect 5403 189 5413 223
rect 5447 189 5459 223
tri 5489 280 5505 296 se
rect 5505 280 5549 296
tri 5549 280 5565 296 sw
rect 5489 247 5565 280
rect 5489 213 5510 247
rect 5544 213 5565 247
rect 5489 211 5565 213
tri 5489 195 5505 211 ne
rect 5505 195 5549 211
tri 5549 195 5565 211 nw
rect 5595 291 5651 326
rect 5595 257 5607 291
rect 5641 257 5651 291
rect 5595 223 5651 257
rect 5403 165 5459 189
tri 5459 165 5489 195 sw
tri 5565 165 5595 195 se
rect 5595 189 5607 223
rect 5641 189 5651 223
rect 5595 165 5651 189
rect 5403 153 5651 165
rect 5403 119 5413 153
rect 5447 119 5510 153
rect 5544 119 5607 153
rect 5641 119 5651 153
rect 5403 103 5651 119
<< pdiff >>
rect 191 1412 247 1450
rect 191 1378 201 1412
rect 235 1378 247 1412
rect 191 1344 247 1378
rect 191 1310 201 1344
rect 235 1310 247 1344
rect 191 1276 247 1310
rect 191 1242 201 1276
rect 235 1242 247 1276
rect 191 1208 247 1242
rect 191 1174 201 1208
rect 235 1174 247 1208
rect 191 1139 247 1174
rect 191 1105 201 1139
rect 235 1105 247 1139
rect 191 1050 247 1105
rect 277 1412 335 1450
rect 277 1378 289 1412
rect 323 1378 335 1412
rect 277 1344 335 1378
rect 277 1310 289 1344
rect 323 1310 335 1344
rect 277 1276 335 1310
rect 277 1242 289 1276
rect 323 1242 335 1276
rect 277 1208 335 1242
rect 277 1174 289 1208
rect 323 1174 335 1208
rect 277 1139 335 1174
rect 277 1105 289 1139
rect 323 1105 335 1139
rect 277 1050 335 1105
rect 365 1412 423 1450
rect 365 1378 377 1412
rect 411 1378 423 1412
rect 365 1344 423 1378
rect 365 1310 377 1344
rect 411 1310 423 1344
rect 365 1276 423 1310
rect 365 1242 377 1276
rect 411 1242 423 1276
rect 365 1208 423 1242
rect 365 1174 377 1208
rect 411 1174 423 1208
rect 365 1050 423 1174
rect 453 1412 511 1450
rect 453 1378 465 1412
rect 499 1378 511 1412
rect 453 1344 511 1378
rect 453 1310 465 1344
rect 499 1310 511 1344
rect 453 1276 511 1310
rect 453 1242 465 1276
rect 499 1242 511 1276
rect 453 1208 511 1242
rect 453 1174 465 1208
rect 499 1174 511 1208
rect 453 1139 511 1174
rect 453 1105 465 1139
rect 499 1105 511 1139
rect 453 1050 511 1105
rect 541 1412 599 1450
rect 541 1378 553 1412
rect 587 1378 599 1412
rect 541 1344 599 1378
rect 541 1310 553 1344
rect 587 1310 599 1344
rect 541 1276 599 1310
rect 541 1242 553 1276
rect 587 1242 599 1276
rect 541 1208 599 1242
rect 541 1174 553 1208
rect 587 1174 599 1208
rect 541 1050 599 1174
rect 629 1412 687 1450
rect 629 1378 641 1412
rect 675 1378 687 1412
rect 629 1344 687 1378
rect 629 1310 641 1344
rect 675 1310 687 1344
rect 629 1276 687 1310
rect 629 1242 641 1276
rect 675 1242 687 1276
rect 629 1208 687 1242
rect 629 1174 641 1208
rect 675 1174 687 1208
rect 629 1139 687 1174
rect 629 1105 641 1139
rect 675 1105 687 1139
rect 629 1050 687 1105
rect 717 1412 771 1450
rect 717 1378 729 1412
rect 763 1378 771 1412
rect 717 1344 771 1378
rect 717 1310 729 1344
rect 763 1310 771 1344
rect 717 1276 771 1310
rect 717 1242 729 1276
rect 763 1242 771 1276
rect 717 1208 771 1242
rect 717 1174 729 1208
rect 763 1174 771 1208
rect 717 1050 771 1174
rect 1153 1412 1209 1450
rect 1153 1378 1163 1412
rect 1197 1378 1209 1412
rect 1153 1344 1209 1378
rect 1153 1310 1163 1344
rect 1197 1310 1209 1344
rect 1153 1276 1209 1310
rect 1153 1242 1163 1276
rect 1197 1242 1209 1276
rect 1153 1208 1209 1242
rect 1153 1174 1163 1208
rect 1197 1174 1209 1208
rect 1153 1139 1209 1174
rect 1153 1105 1163 1139
rect 1197 1105 1209 1139
rect 1153 1050 1209 1105
rect 1239 1412 1297 1450
rect 1239 1378 1251 1412
rect 1285 1378 1297 1412
rect 1239 1344 1297 1378
rect 1239 1310 1251 1344
rect 1285 1310 1297 1344
rect 1239 1276 1297 1310
rect 1239 1242 1251 1276
rect 1285 1242 1297 1276
rect 1239 1208 1297 1242
rect 1239 1174 1251 1208
rect 1285 1174 1297 1208
rect 1239 1139 1297 1174
rect 1239 1105 1251 1139
rect 1285 1105 1297 1139
rect 1239 1050 1297 1105
rect 1327 1412 1385 1450
rect 1327 1378 1339 1412
rect 1373 1378 1385 1412
rect 1327 1344 1385 1378
rect 1327 1310 1339 1344
rect 1373 1310 1385 1344
rect 1327 1276 1385 1310
rect 1327 1242 1339 1276
rect 1373 1242 1385 1276
rect 1327 1208 1385 1242
rect 1327 1174 1339 1208
rect 1373 1174 1385 1208
rect 1327 1050 1385 1174
rect 1415 1412 1473 1450
rect 1415 1378 1427 1412
rect 1461 1378 1473 1412
rect 1415 1344 1473 1378
rect 1415 1310 1427 1344
rect 1461 1310 1473 1344
rect 1415 1276 1473 1310
rect 1415 1242 1427 1276
rect 1461 1242 1473 1276
rect 1415 1208 1473 1242
rect 1415 1174 1427 1208
rect 1461 1174 1473 1208
rect 1415 1139 1473 1174
rect 1415 1105 1427 1139
rect 1461 1105 1473 1139
rect 1415 1050 1473 1105
rect 1503 1412 1561 1450
rect 1503 1378 1515 1412
rect 1549 1378 1561 1412
rect 1503 1344 1561 1378
rect 1503 1310 1515 1344
rect 1549 1310 1561 1344
rect 1503 1276 1561 1310
rect 1503 1242 1515 1276
rect 1549 1242 1561 1276
rect 1503 1208 1561 1242
rect 1503 1174 1515 1208
rect 1549 1174 1561 1208
rect 1503 1050 1561 1174
rect 1591 1412 1649 1450
rect 1591 1378 1603 1412
rect 1637 1378 1649 1412
rect 1591 1344 1649 1378
rect 1591 1310 1603 1344
rect 1637 1310 1649 1344
rect 1591 1276 1649 1310
rect 1591 1242 1603 1276
rect 1637 1242 1649 1276
rect 1591 1208 1649 1242
rect 1591 1174 1603 1208
rect 1637 1174 1649 1208
rect 1591 1139 1649 1174
rect 1591 1105 1603 1139
rect 1637 1105 1649 1139
rect 1591 1050 1649 1105
rect 1679 1412 1733 1450
rect 1679 1378 1691 1412
rect 1725 1378 1733 1412
rect 1679 1344 1733 1378
rect 1679 1310 1691 1344
rect 1725 1310 1733 1344
rect 1679 1276 1733 1310
rect 1679 1242 1691 1276
rect 1725 1242 1733 1276
rect 1679 1208 1733 1242
rect 1679 1174 1691 1208
rect 1725 1174 1733 1208
rect 1679 1050 1733 1174
rect 2115 1412 2171 1450
rect 2115 1378 2125 1412
rect 2159 1378 2171 1412
rect 2115 1344 2171 1378
rect 2115 1310 2125 1344
rect 2159 1310 2171 1344
rect 2115 1276 2171 1310
rect 2115 1242 2125 1276
rect 2159 1242 2171 1276
rect 2115 1208 2171 1242
rect 2115 1174 2125 1208
rect 2159 1174 2171 1208
rect 2115 1139 2171 1174
rect 2115 1105 2125 1139
rect 2159 1105 2171 1139
rect 2115 1050 2171 1105
rect 2201 1412 2259 1450
rect 2201 1378 2213 1412
rect 2247 1378 2259 1412
rect 2201 1344 2259 1378
rect 2201 1310 2213 1344
rect 2247 1310 2259 1344
rect 2201 1276 2259 1310
rect 2201 1242 2213 1276
rect 2247 1242 2259 1276
rect 2201 1208 2259 1242
rect 2201 1174 2213 1208
rect 2247 1174 2259 1208
rect 2201 1139 2259 1174
rect 2201 1105 2213 1139
rect 2247 1105 2259 1139
rect 2201 1050 2259 1105
rect 2289 1412 2347 1450
rect 2289 1378 2301 1412
rect 2335 1378 2347 1412
rect 2289 1344 2347 1378
rect 2289 1310 2301 1344
rect 2335 1310 2347 1344
rect 2289 1276 2347 1310
rect 2289 1242 2301 1276
rect 2335 1242 2347 1276
rect 2289 1208 2347 1242
rect 2289 1174 2301 1208
rect 2335 1174 2347 1208
rect 2289 1050 2347 1174
rect 2377 1412 2435 1450
rect 2377 1378 2389 1412
rect 2423 1378 2435 1412
rect 2377 1344 2435 1378
rect 2377 1310 2389 1344
rect 2423 1310 2435 1344
rect 2377 1276 2435 1310
rect 2377 1242 2389 1276
rect 2423 1242 2435 1276
rect 2377 1208 2435 1242
rect 2377 1174 2389 1208
rect 2423 1174 2435 1208
rect 2377 1139 2435 1174
rect 2377 1105 2389 1139
rect 2423 1105 2435 1139
rect 2377 1050 2435 1105
rect 2465 1412 2523 1450
rect 2465 1378 2477 1412
rect 2511 1378 2523 1412
rect 2465 1344 2523 1378
rect 2465 1310 2477 1344
rect 2511 1310 2523 1344
rect 2465 1276 2523 1310
rect 2465 1242 2477 1276
rect 2511 1242 2523 1276
rect 2465 1208 2523 1242
rect 2465 1174 2477 1208
rect 2511 1174 2523 1208
rect 2465 1050 2523 1174
rect 2553 1412 2611 1450
rect 2553 1378 2565 1412
rect 2599 1378 2611 1412
rect 2553 1344 2611 1378
rect 2553 1310 2565 1344
rect 2599 1310 2611 1344
rect 2553 1276 2611 1310
rect 2553 1242 2565 1276
rect 2599 1242 2611 1276
rect 2553 1208 2611 1242
rect 2553 1174 2565 1208
rect 2599 1174 2611 1208
rect 2553 1139 2611 1174
rect 2553 1105 2565 1139
rect 2599 1105 2611 1139
rect 2553 1050 2611 1105
rect 2641 1412 2695 1450
rect 2641 1378 2653 1412
rect 2687 1378 2695 1412
rect 2641 1344 2695 1378
rect 2641 1310 2653 1344
rect 2687 1310 2695 1344
rect 2641 1276 2695 1310
rect 2641 1242 2653 1276
rect 2687 1242 2695 1276
rect 2641 1208 2695 1242
rect 2641 1174 2653 1208
rect 2687 1174 2695 1208
rect 2641 1050 2695 1174
rect 3077 1412 3133 1450
rect 3077 1378 3087 1412
rect 3121 1378 3133 1412
rect 3077 1344 3133 1378
rect 3077 1310 3087 1344
rect 3121 1310 3133 1344
rect 3077 1276 3133 1310
rect 3077 1242 3087 1276
rect 3121 1242 3133 1276
rect 3077 1208 3133 1242
rect 3077 1174 3087 1208
rect 3121 1174 3133 1208
rect 3077 1139 3133 1174
rect 3077 1105 3087 1139
rect 3121 1105 3133 1139
rect 3077 1050 3133 1105
rect 3163 1412 3221 1450
rect 3163 1378 3175 1412
rect 3209 1378 3221 1412
rect 3163 1344 3221 1378
rect 3163 1310 3175 1344
rect 3209 1310 3221 1344
rect 3163 1276 3221 1310
rect 3163 1242 3175 1276
rect 3209 1242 3221 1276
rect 3163 1208 3221 1242
rect 3163 1174 3175 1208
rect 3209 1174 3221 1208
rect 3163 1139 3221 1174
rect 3163 1105 3175 1139
rect 3209 1105 3221 1139
rect 3163 1050 3221 1105
rect 3251 1412 3309 1450
rect 3251 1378 3263 1412
rect 3297 1378 3309 1412
rect 3251 1344 3309 1378
rect 3251 1310 3263 1344
rect 3297 1310 3309 1344
rect 3251 1276 3309 1310
rect 3251 1242 3263 1276
rect 3297 1242 3309 1276
rect 3251 1208 3309 1242
rect 3251 1174 3263 1208
rect 3297 1174 3309 1208
rect 3251 1050 3309 1174
rect 3339 1412 3397 1450
rect 3339 1378 3351 1412
rect 3385 1378 3397 1412
rect 3339 1344 3397 1378
rect 3339 1310 3351 1344
rect 3385 1310 3397 1344
rect 3339 1276 3397 1310
rect 3339 1242 3351 1276
rect 3385 1242 3397 1276
rect 3339 1208 3397 1242
rect 3339 1174 3351 1208
rect 3385 1174 3397 1208
rect 3339 1139 3397 1174
rect 3339 1105 3351 1139
rect 3385 1105 3397 1139
rect 3339 1050 3397 1105
rect 3427 1412 3485 1450
rect 3427 1378 3439 1412
rect 3473 1378 3485 1412
rect 3427 1344 3485 1378
rect 3427 1310 3439 1344
rect 3473 1310 3485 1344
rect 3427 1276 3485 1310
rect 3427 1242 3439 1276
rect 3473 1242 3485 1276
rect 3427 1208 3485 1242
rect 3427 1174 3439 1208
rect 3473 1174 3485 1208
rect 3427 1050 3485 1174
rect 3515 1412 3573 1450
rect 3515 1378 3527 1412
rect 3561 1378 3573 1412
rect 3515 1344 3573 1378
rect 3515 1310 3527 1344
rect 3561 1310 3573 1344
rect 3515 1276 3573 1310
rect 3515 1242 3527 1276
rect 3561 1242 3573 1276
rect 3515 1208 3573 1242
rect 3515 1174 3527 1208
rect 3561 1174 3573 1208
rect 3515 1139 3573 1174
rect 3515 1105 3527 1139
rect 3561 1105 3573 1139
rect 3515 1050 3573 1105
rect 3603 1412 3657 1450
rect 3603 1378 3615 1412
rect 3649 1378 3657 1412
rect 3603 1344 3657 1378
rect 3603 1310 3615 1344
rect 3649 1310 3657 1344
rect 3603 1276 3657 1310
rect 3603 1242 3615 1276
rect 3649 1242 3657 1276
rect 3603 1208 3657 1242
rect 3603 1174 3615 1208
rect 3649 1174 3657 1208
rect 3603 1050 3657 1174
rect 4039 1412 4095 1450
rect 4039 1378 4049 1412
rect 4083 1378 4095 1412
rect 4039 1344 4095 1378
rect 4039 1310 4049 1344
rect 4083 1310 4095 1344
rect 4039 1276 4095 1310
rect 4039 1242 4049 1276
rect 4083 1242 4095 1276
rect 4039 1208 4095 1242
rect 4039 1174 4049 1208
rect 4083 1174 4095 1208
rect 4039 1139 4095 1174
rect 4039 1105 4049 1139
rect 4083 1105 4095 1139
rect 4039 1050 4095 1105
rect 4125 1412 4183 1450
rect 4125 1378 4137 1412
rect 4171 1378 4183 1412
rect 4125 1344 4183 1378
rect 4125 1310 4137 1344
rect 4171 1310 4183 1344
rect 4125 1276 4183 1310
rect 4125 1242 4137 1276
rect 4171 1242 4183 1276
rect 4125 1208 4183 1242
rect 4125 1174 4137 1208
rect 4171 1174 4183 1208
rect 4125 1139 4183 1174
rect 4125 1105 4137 1139
rect 4171 1105 4183 1139
rect 4125 1050 4183 1105
rect 4213 1412 4271 1450
rect 4213 1378 4225 1412
rect 4259 1378 4271 1412
rect 4213 1344 4271 1378
rect 4213 1310 4225 1344
rect 4259 1310 4271 1344
rect 4213 1276 4271 1310
rect 4213 1242 4225 1276
rect 4259 1242 4271 1276
rect 4213 1208 4271 1242
rect 4213 1174 4225 1208
rect 4259 1174 4271 1208
rect 4213 1050 4271 1174
rect 4301 1412 4359 1450
rect 4301 1378 4313 1412
rect 4347 1378 4359 1412
rect 4301 1344 4359 1378
rect 4301 1310 4313 1344
rect 4347 1310 4359 1344
rect 4301 1276 4359 1310
rect 4301 1242 4313 1276
rect 4347 1242 4359 1276
rect 4301 1208 4359 1242
rect 4301 1174 4313 1208
rect 4347 1174 4359 1208
rect 4301 1139 4359 1174
rect 4301 1105 4313 1139
rect 4347 1105 4359 1139
rect 4301 1050 4359 1105
rect 4389 1412 4447 1450
rect 4389 1378 4401 1412
rect 4435 1378 4447 1412
rect 4389 1344 4447 1378
rect 4389 1310 4401 1344
rect 4435 1310 4447 1344
rect 4389 1276 4447 1310
rect 4389 1242 4401 1276
rect 4435 1242 4447 1276
rect 4389 1208 4447 1242
rect 4389 1174 4401 1208
rect 4435 1174 4447 1208
rect 4389 1050 4447 1174
rect 4477 1412 4535 1450
rect 4477 1378 4489 1412
rect 4523 1378 4535 1412
rect 4477 1344 4535 1378
rect 4477 1310 4489 1344
rect 4523 1310 4535 1344
rect 4477 1276 4535 1310
rect 4477 1242 4489 1276
rect 4523 1242 4535 1276
rect 4477 1208 4535 1242
rect 4477 1174 4489 1208
rect 4523 1174 4535 1208
rect 4477 1139 4535 1174
rect 4477 1105 4489 1139
rect 4523 1105 4535 1139
rect 4477 1050 4535 1105
rect 4565 1412 4619 1450
rect 4565 1378 4577 1412
rect 4611 1378 4619 1412
rect 4565 1344 4619 1378
rect 4565 1310 4577 1344
rect 4611 1310 4619 1344
rect 4565 1276 4619 1310
rect 4565 1242 4577 1276
rect 4611 1242 4619 1276
rect 4565 1208 4619 1242
rect 4565 1174 4577 1208
rect 4611 1174 4619 1208
rect 4565 1050 4619 1174
rect 5001 1412 5057 1450
rect 5001 1378 5011 1412
rect 5045 1378 5057 1412
rect 5001 1344 5057 1378
rect 5001 1310 5011 1344
rect 5045 1310 5057 1344
rect 5001 1276 5057 1310
rect 5001 1242 5011 1276
rect 5045 1242 5057 1276
rect 5001 1208 5057 1242
rect 5001 1174 5011 1208
rect 5045 1174 5057 1208
rect 5001 1139 5057 1174
rect 5001 1105 5011 1139
rect 5045 1105 5057 1139
rect 5001 1050 5057 1105
rect 5087 1412 5145 1450
rect 5087 1378 5099 1412
rect 5133 1378 5145 1412
rect 5087 1344 5145 1378
rect 5087 1310 5099 1344
rect 5133 1310 5145 1344
rect 5087 1276 5145 1310
rect 5087 1242 5099 1276
rect 5133 1242 5145 1276
rect 5087 1208 5145 1242
rect 5087 1174 5099 1208
rect 5133 1174 5145 1208
rect 5087 1139 5145 1174
rect 5087 1105 5099 1139
rect 5133 1105 5145 1139
rect 5087 1050 5145 1105
rect 5175 1412 5233 1450
rect 5175 1378 5187 1412
rect 5221 1378 5233 1412
rect 5175 1344 5233 1378
rect 5175 1310 5187 1344
rect 5221 1310 5233 1344
rect 5175 1276 5233 1310
rect 5175 1242 5187 1276
rect 5221 1242 5233 1276
rect 5175 1208 5233 1242
rect 5175 1174 5187 1208
rect 5221 1174 5233 1208
rect 5175 1050 5233 1174
rect 5263 1412 5321 1450
rect 5263 1378 5275 1412
rect 5309 1378 5321 1412
rect 5263 1344 5321 1378
rect 5263 1310 5275 1344
rect 5309 1310 5321 1344
rect 5263 1276 5321 1310
rect 5263 1242 5275 1276
rect 5309 1242 5321 1276
rect 5263 1208 5321 1242
rect 5263 1174 5275 1208
rect 5309 1174 5321 1208
rect 5263 1139 5321 1174
rect 5263 1105 5275 1139
rect 5309 1105 5321 1139
rect 5263 1050 5321 1105
rect 5351 1412 5409 1450
rect 5351 1378 5363 1412
rect 5397 1378 5409 1412
rect 5351 1344 5409 1378
rect 5351 1310 5363 1344
rect 5397 1310 5409 1344
rect 5351 1276 5409 1310
rect 5351 1242 5363 1276
rect 5397 1242 5409 1276
rect 5351 1208 5409 1242
rect 5351 1174 5363 1208
rect 5397 1174 5409 1208
rect 5351 1050 5409 1174
rect 5439 1412 5497 1450
rect 5439 1378 5451 1412
rect 5485 1378 5497 1412
rect 5439 1344 5497 1378
rect 5439 1310 5451 1344
rect 5485 1310 5497 1344
rect 5439 1276 5497 1310
rect 5439 1242 5451 1276
rect 5485 1242 5497 1276
rect 5439 1208 5497 1242
rect 5439 1174 5451 1208
rect 5485 1174 5497 1208
rect 5439 1139 5497 1174
rect 5439 1105 5451 1139
rect 5485 1105 5497 1139
rect 5439 1050 5497 1105
rect 5527 1412 5581 1450
rect 5527 1378 5539 1412
rect 5573 1378 5581 1412
rect 5527 1344 5581 1378
rect 5527 1310 5539 1344
rect 5573 1310 5581 1344
rect 5527 1276 5581 1310
rect 5527 1242 5539 1276
rect 5573 1242 5581 1276
rect 5527 1208 5581 1242
rect 5527 1174 5539 1208
rect 5573 1174 5581 1208
rect 5527 1050 5581 1174
<< ndiffc >>
rect 101 329 135 363
rect 198 329 232 363
rect 295 329 329 363
rect 392 329 426 363
rect 489 329 523 363
rect 101 257 135 291
rect 101 189 135 223
rect 198 204 232 238
rect 295 257 329 291
rect 295 189 329 223
rect 393 210 427 244
rect 101 119 135 153
rect 295 119 329 153
rect 392 119 426 153
rect 489 119 523 153
rect 603 329 637 363
rect 603 257 637 291
rect 603 189 637 223
rect 700 213 734 247
rect 797 257 831 291
rect 797 189 831 223
rect 603 119 637 153
rect 700 119 734 153
rect 797 119 831 153
rect 1063 329 1097 363
rect 1160 329 1194 363
rect 1257 329 1291 363
rect 1354 329 1388 363
rect 1451 329 1485 363
rect 1063 257 1097 291
rect 1063 189 1097 223
rect 1160 204 1194 238
rect 1257 257 1291 291
rect 1257 189 1291 223
rect 1355 210 1389 244
rect 1063 119 1097 153
rect 1257 119 1291 153
rect 1354 119 1388 153
rect 1451 119 1485 153
rect 1565 329 1599 363
rect 1565 257 1599 291
rect 1565 189 1599 223
rect 1662 213 1696 247
rect 1759 257 1793 291
rect 1759 189 1793 223
rect 1565 119 1599 153
rect 1662 119 1696 153
rect 1759 119 1793 153
rect 2025 329 2059 363
rect 2122 329 2156 363
rect 2219 329 2253 363
rect 2316 329 2350 363
rect 2413 329 2447 363
rect 2025 257 2059 291
rect 2025 189 2059 223
rect 2122 204 2156 238
rect 2219 257 2253 291
rect 2219 189 2253 223
rect 2317 210 2351 244
rect 2025 119 2059 153
rect 2219 119 2253 153
rect 2316 119 2350 153
rect 2413 119 2447 153
rect 2527 329 2561 363
rect 2527 257 2561 291
rect 2527 189 2561 223
rect 2624 213 2658 247
rect 2721 257 2755 291
rect 2721 189 2755 223
rect 2527 119 2561 153
rect 2624 119 2658 153
rect 2721 119 2755 153
rect 2987 329 3021 363
rect 3084 329 3118 363
rect 3181 329 3215 363
rect 3278 329 3312 363
rect 3375 329 3409 363
rect 2987 257 3021 291
rect 2987 189 3021 223
rect 3084 204 3118 238
rect 3181 257 3215 291
rect 3181 189 3215 223
rect 3279 210 3313 244
rect 2987 119 3021 153
rect 3181 119 3215 153
rect 3278 119 3312 153
rect 3375 119 3409 153
rect 3489 329 3523 363
rect 3489 257 3523 291
rect 3489 189 3523 223
rect 3586 213 3620 247
rect 3683 257 3717 291
rect 3683 189 3717 223
rect 3489 119 3523 153
rect 3586 119 3620 153
rect 3683 119 3717 153
rect 3949 329 3983 363
rect 4046 329 4080 363
rect 4143 329 4177 363
rect 4240 329 4274 363
rect 4337 329 4371 363
rect 3949 257 3983 291
rect 3949 189 3983 223
rect 4046 204 4080 238
rect 4143 257 4177 291
rect 4143 189 4177 223
rect 4241 210 4275 244
rect 3949 119 3983 153
rect 4143 119 4177 153
rect 4240 119 4274 153
rect 4337 119 4371 153
rect 4451 329 4485 363
rect 4451 257 4485 291
rect 4451 189 4485 223
rect 4548 213 4582 247
rect 4645 257 4679 291
rect 4645 189 4679 223
rect 4451 119 4485 153
rect 4548 119 4582 153
rect 4645 119 4679 153
rect 4911 329 4945 363
rect 5008 329 5042 363
rect 5105 329 5139 363
rect 5202 329 5236 363
rect 5299 329 5333 363
rect 4911 257 4945 291
rect 4911 189 4945 223
rect 5008 204 5042 238
rect 5105 257 5139 291
rect 5105 189 5139 223
rect 5203 210 5237 244
rect 4911 119 4945 153
rect 5105 119 5139 153
rect 5202 119 5236 153
rect 5299 119 5333 153
rect 5413 329 5447 363
rect 5413 257 5447 291
rect 5413 189 5447 223
rect 5510 213 5544 247
rect 5607 257 5641 291
rect 5607 189 5641 223
rect 5413 119 5447 153
rect 5510 119 5544 153
rect 5607 119 5641 153
<< pdiffc >>
rect 201 1378 235 1412
rect 201 1310 235 1344
rect 201 1242 235 1276
rect 201 1174 235 1208
rect 201 1105 235 1139
rect 289 1378 323 1412
rect 289 1310 323 1344
rect 289 1242 323 1276
rect 289 1174 323 1208
rect 289 1105 323 1139
rect 377 1378 411 1412
rect 377 1310 411 1344
rect 377 1242 411 1276
rect 377 1174 411 1208
rect 465 1378 499 1412
rect 465 1310 499 1344
rect 465 1242 499 1276
rect 465 1174 499 1208
rect 465 1105 499 1139
rect 553 1378 587 1412
rect 553 1310 587 1344
rect 553 1242 587 1276
rect 553 1174 587 1208
rect 641 1378 675 1412
rect 641 1310 675 1344
rect 641 1242 675 1276
rect 641 1174 675 1208
rect 641 1105 675 1139
rect 729 1378 763 1412
rect 729 1310 763 1344
rect 729 1242 763 1276
rect 729 1174 763 1208
rect 1163 1378 1197 1412
rect 1163 1310 1197 1344
rect 1163 1242 1197 1276
rect 1163 1174 1197 1208
rect 1163 1105 1197 1139
rect 1251 1378 1285 1412
rect 1251 1310 1285 1344
rect 1251 1242 1285 1276
rect 1251 1174 1285 1208
rect 1251 1105 1285 1139
rect 1339 1378 1373 1412
rect 1339 1310 1373 1344
rect 1339 1242 1373 1276
rect 1339 1174 1373 1208
rect 1427 1378 1461 1412
rect 1427 1310 1461 1344
rect 1427 1242 1461 1276
rect 1427 1174 1461 1208
rect 1427 1105 1461 1139
rect 1515 1378 1549 1412
rect 1515 1310 1549 1344
rect 1515 1242 1549 1276
rect 1515 1174 1549 1208
rect 1603 1378 1637 1412
rect 1603 1310 1637 1344
rect 1603 1242 1637 1276
rect 1603 1174 1637 1208
rect 1603 1105 1637 1139
rect 1691 1378 1725 1412
rect 1691 1310 1725 1344
rect 1691 1242 1725 1276
rect 1691 1174 1725 1208
rect 2125 1378 2159 1412
rect 2125 1310 2159 1344
rect 2125 1242 2159 1276
rect 2125 1174 2159 1208
rect 2125 1105 2159 1139
rect 2213 1378 2247 1412
rect 2213 1310 2247 1344
rect 2213 1242 2247 1276
rect 2213 1174 2247 1208
rect 2213 1105 2247 1139
rect 2301 1378 2335 1412
rect 2301 1310 2335 1344
rect 2301 1242 2335 1276
rect 2301 1174 2335 1208
rect 2389 1378 2423 1412
rect 2389 1310 2423 1344
rect 2389 1242 2423 1276
rect 2389 1174 2423 1208
rect 2389 1105 2423 1139
rect 2477 1378 2511 1412
rect 2477 1310 2511 1344
rect 2477 1242 2511 1276
rect 2477 1174 2511 1208
rect 2565 1378 2599 1412
rect 2565 1310 2599 1344
rect 2565 1242 2599 1276
rect 2565 1174 2599 1208
rect 2565 1105 2599 1139
rect 2653 1378 2687 1412
rect 2653 1310 2687 1344
rect 2653 1242 2687 1276
rect 2653 1174 2687 1208
rect 3087 1378 3121 1412
rect 3087 1310 3121 1344
rect 3087 1242 3121 1276
rect 3087 1174 3121 1208
rect 3087 1105 3121 1139
rect 3175 1378 3209 1412
rect 3175 1310 3209 1344
rect 3175 1242 3209 1276
rect 3175 1174 3209 1208
rect 3175 1105 3209 1139
rect 3263 1378 3297 1412
rect 3263 1310 3297 1344
rect 3263 1242 3297 1276
rect 3263 1174 3297 1208
rect 3351 1378 3385 1412
rect 3351 1310 3385 1344
rect 3351 1242 3385 1276
rect 3351 1174 3385 1208
rect 3351 1105 3385 1139
rect 3439 1378 3473 1412
rect 3439 1310 3473 1344
rect 3439 1242 3473 1276
rect 3439 1174 3473 1208
rect 3527 1378 3561 1412
rect 3527 1310 3561 1344
rect 3527 1242 3561 1276
rect 3527 1174 3561 1208
rect 3527 1105 3561 1139
rect 3615 1378 3649 1412
rect 3615 1310 3649 1344
rect 3615 1242 3649 1276
rect 3615 1174 3649 1208
rect 4049 1378 4083 1412
rect 4049 1310 4083 1344
rect 4049 1242 4083 1276
rect 4049 1174 4083 1208
rect 4049 1105 4083 1139
rect 4137 1378 4171 1412
rect 4137 1310 4171 1344
rect 4137 1242 4171 1276
rect 4137 1174 4171 1208
rect 4137 1105 4171 1139
rect 4225 1378 4259 1412
rect 4225 1310 4259 1344
rect 4225 1242 4259 1276
rect 4225 1174 4259 1208
rect 4313 1378 4347 1412
rect 4313 1310 4347 1344
rect 4313 1242 4347 1276
rect 4313 1174 4347 1208
rect 4313 1105 4347 1139
rect 4401 1378 4435 1412
rect 4401 1310 4435 1344
rect 4401 1242 4435 1276
rect 4401 1174 4435 1208
rect 4489 1378 4523 1412
rect 4489 1310 4523 1344
rect 4489 1242 4523 1276
rect 4489 1174 4523 1208
rect 4489 1105 4523 1139
rect 4577 1378 4611 1412
rect 4577 1310 4611 1344
rect 4577 1242 4611 1276
rect 4577 1174 4611 1208
rect 5011 1378 5045 1412
rect 5011 1310 5045 1344
rect 5011 1242 5045 1276
rect 5011 1174 5045 1208
rect 5011 1105 5045 1139
rect 5099 1378 5133 1412
rect 5099 1310 5133 1344
rect 5099 1242 5133 1276
rect 5099 1174 5133 1208
rect 5099 1105 5133 1139
rect 5187 1378 5221 1412
rect 5187 1310 5221 1344
rect 5187 1242 5221 1276
rect 5187 1174 5221 1208
rect 5275 1378 5309 1412
rect 5275 1310 5309 1344
rect 5275 1242 5309 1276
rect 5275 1174 5309 1208
rect 5275 1105 5309 1139
rect 5363 1378 5397 1412
rect 5363 1310 5397 1344
rect 5363 1242 5397 1276
rect 5363 1174 5397 1208
rect 5451 1378 5485 1412
rect 5451 1310 5485 1344
rect 5451 1242 5485 1276
rect 5451 1174 5485 1208
rect 5451 1105 5485 1139
rect 5539 1378 5573 1412
rect 5539 1310 5573 1344
rect 5539 1242 5573 1276
rect 5539 1174 5573 1208
<< psubdiff >>
rect -31 546 5803 572
rect -31 512 -17 546
rect 17 512 945 546
rect 979 512 1907 546
rect 1941 512 2869 546
rect 2903 512 3831 546
rect 3865 512 4793 546
rect 4827 512 5755 546
rect 5789 512 5803 546
rect -31 510 5803 512
rect -31 474 31 510
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect -31 368 -17 402
rect 17 368 31 402
rect 931 474 993 510
rect 931 440 945 474
rect 979 440 993 474
rect 931 402 993 440
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect 931 368 945 402
rect 979 368 993 402
rect 1893 474 1955 510
rect 1893 440 1907 474
rect 1941 440 1955 474
rect 1893 402 1955 440
rect 931 330 993 368
rect 931 296 945 330
rect 979 296 993 330
rect 931 258 993 296
rect 931 224 945 258
rect 979 224 993 258
rect 931 186 993 224
rect 931 152 945 186
rect 979 152 993 186
rect 931 114 993 152
rect -31 47 31 80
rect 931 80 945 114
rect 979 80 993 114
rect 1893 368 1907 402
rect 1941 368 1955 402
rect 2855 474 2917 510
rect 2855 440 2869 474
rect 2903 440 2917 474
rect 2855 402 2917 440
rect 1893 330 1955 368
rect 1893 296 1907 330
rect 1941 296 1955 330
rect 1893 258 1955 296
rect 1893 224 1907 258
rect 1941 224 1955 258
rect 1893 186 1955 224
rect 1893 152 1907 186
rect 1941 152 1955 186
rect 1893 114 1955 152
rect 931 47 993 80
rect 1893 80 1907 114
rect 1941 80 1955 114
rect 2855 368 2869 402
rect 2903 368 2917 402
rect 3817 474 3879 510
rect 3817 440 3831 474
rect 3865 440 3879 474
rect 3817 402 3879 440
rect 2855 330 2917 368
rect 2855 296 2869 330
rect 2903 296 2917 330
rect 2855 258 2917 296
rect 2855 224 2869 258
rect 2903 224 2917 258
rect 2855 186 2917 224
rect 2855 152 2869 186
rect 2903 152 2917 186
rect 2855 114 2917 152
rect 1893 47 1955 80
rect 2855 80 2869 114
rect 2903 80 2917 114
rect 3817 368 3831 402
rect 3865 368 3879 402
rect 4779 474 4841 510
rect 4779 440 4793 474
rect 4827 440 4841 474
rect 4779 402 4841 440
rect 3817 330 3879 368
rect 3817 296 3831 330
rect 3865 296 3879 330
rect 3817 258 3879 296
rect 3817 224 3831 258
rect 3865 224 3879 258
rect 3817 186 3879 224
rect 3817 152 3831 186
rect 3865 152 3879 186
rect 3817 114 3879 152
rect 2855 47 2917 80
rect 3817 80 3831 114
rect 3865 80 3879 114
rect 4779 368 4793 402
rect 4827 368 4841 402
rect 5741 474 5803 510
rect 5741 440 5755 474
rect 5789 440 5803 474
rect 5741 402 5803 440
rect 4779 330 4841 368
rect 4779 296 4793 330
rect 4827 296 4841 330
rect 4779 258 4841 296
rect 4779 224 4793 258
rect 4827 224 4841 258
rect 4779 186 4841 224
rect 4779 152 4793 186
rect 4827 152 4841 186
rect 4779 114 4841 152
rect 3817 47 3879 80
rect 4779 80 4793 114
rect 4827 80 4841 114
rect 5741 368 5755 402
rect 5789 368 5803 402
rect 5741 330 5803 368
rect 5741 296 5755 330
rect 5789 296 5803 330
rect 5741 258 5803 296
rect 5741 224 5755 258
rect 5789 224 5803 258
rect 5741 186 5803 224
rect 5741 152 5755 186
rect 5789 152 5803 186
rect 5741 114 5803 152
rect 4779 47 4841 80
rect 5741 80 5755 114
rect 5789 80 5803 114
rect 5741 47 5803 80
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 343 47
rect 377 13 415 47
rect 449 13 513 47
rect 547 13 585 47
rect 619 13 657 47
rect 691 13 729 47
rect 763 13 801 47
rect 835 13 873 47
rect 907 13 1017 47
rect 1051 13 1089 47
rect 1123 13 1161 47
rect 1195 13 1233 47
rect 1267 13 1305 47
rect 1339 13 1377 47
rect 1411 13 1475 47
rect 1509 13 1547 47
rect 1581 13 1619 47
rect 1653 13 1691 47
rect 1725 13 1763 47
rect 1797 13 1835 47
rect 1869 13 1979 47
rect 2013 13 2051 47
rect 2085 13 2123 47
rect 2157 13 2195 47
rect 2229 13 2267 47
rect 2301 13 2339 47
rect 2373 13 2437 47
rect 2471 13 2509 47
rect 2543 13 2581 47
rect 2615 13 2653 47
rect 2687 13 2725 47
rect 2759 13 2797 47
rect 2831 13 2941 47
rect 2975 13 3013 47
rect 3047 13 3085 47
rect 3119 13 3157 47
rect 3191 13 3229 47
rect 3263 13 3301 47
rect 3335 13 3399 47
rect 3433 13 3471 47
rect 3505 13 3543 47
rect 3577 13 3615 47
rect 3649 13 3687 47
rect 3721 13 3759 47
rect 3793 13 3903 47
rect 3937 13 3975 47
rect 4009 13 4047 47
rect 4081 13 4119 47
rect 4153 13 4191 47
rect 4225 13 4263 47
rect 4297 13 4361 47
rect 4395 13 4433 47
rect 4467 13 4505 47
rect 4539 13 4577 47
rect 4611 13 4649 47
rect 4683 13 4721 47
rect 4755 13 4865 47
rect 4899 13 4937 47
rect 4971 13 5009 47
rect 5043 13 5081 47
rect 5115 13 5153 47
rect 5187 13 5225 47
rect 5259 13 5323 47
rect 5357 13 5395 47
rect 5429 13 5467 47
rect 5501 13 5539 47
rect 5573 13 5611 47
rect 5645 13 5683 47
rect 5717 13 5803 47
rect -31 11 31 13
rect 931 11 993 13
rect 1893 11 1955 13
rect 2855 11 2917 13
rect 3817 11 3879 13
rect 4779 11 4841 13
rect 5741 11 5803 13
<< nsubdiff >>
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 343 1539
rect 377 1505 415 1539
rect 449 1505 513 1539
rect 547 1505 585 1539
rect 619 1505 657 1539
rect 691 1505 729 1539
rect 763 1505 801 1539
rect 835 1505 873 1539
rect 907 1505 1017 1539
rect 1051 1505 1089 1539
rect 1123 1505 1161 1539
rect 1195 1505 1233 1539
rect 1267 1505 1305 1539
rect 1339 1505 1377 1539
rect 1411 1505 1475 1539
rect 1509 1505 1547 1539
rect 1581 1505 1619 1539
rect 1653 1505 1691 1539
rect 1725 1505 1763 1539
rect 1797 1505 1835 1539
rect 1869 1505 1979 1539
rect 2013 1505 2051 1539
rect 2085 1505 2123 1539
rect 2157 1505 2195 1539
rect 2229 1505 2267 1539
rect 2301 1505 2339 1539
rect 2373 1505 2437 1539
rect 2471 1505 2509 1539
rect 2543 1505 2581 1539
rect 2615 1505 2653 1539
rect 2687 1505 2725 1539
rect 2759 1505 2797 1539
rect 2831 1505 2941 1539
rect 2975 1505 3013 1539
rect 3047 1505 3085 1539
rect 3119 1505 3157 1539
rect 3191 1505 3229 1539
rect 3263 1505 3301 1539
rect 3335 1505 3399 1539
rect 3433 1505 3471 1539
rect 3505 1505 3543 1539
rect 3577 1505 3615 1539
rect 3649 1505 3687 1539
rect 3721 1505 3759 1539
rect 3793 1505 3903 1539
rect 3937 1505 3975 1539
rect 4009 1505 4047 1539
rect 4081 1505 4119 1539
rect 4153 1505 4191 1539
rect 4225 1505 4263 1539
rect 4297 1505 4361 1539
rect 4395 1505 4433 1539
rect 4467 1505 4505 1539
rect 4539 1505 4577 1539
rect 4611 1505 4649 1539
rect 4683 1505 4721 1539
rect 4755 1505 4865 1539
rect 4899 1505 4937 1539
rect 4971 1505 5009 1539
rect 5043 1505 5081 1539
rect 5115 1505 5153 1539
rect 5187 1505 5225 1539
rect 5259 1505 5323 1539
rect 5357 1505 5395 1539
rect 5429 1505 5467 1539
rect 5501 1505 5539 1539
rect 5573 1505 5611 1539
rect 5645 1505 5683 1539
rect 5717 1505 5803 1539
rect -31 1470 31 1505
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect 931 1470 993 1505
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect -31 1038 31 1076
rect 931 1436 945 1470
rect 979 1436 993 1470
rect 1893 1470 1955 1505
rect 931 1398 993 1436
rect 931 1364 945 1398
rect 979 1364 993 1398
rect 931 1326 993 1364
rect 931 1292 945 1326
rect 979 1292 993 1326
rect 931 1254 993 1292
rect 931 1220 945 1254
rect 979 1220 993 1254
rect 931 1182 993 1220
rect 931 1148 945 1182
rect 979 1148 993 1182
rect 931 1110 993 1148
rect 931 1076 945 1110
rect 979 1076 993 1110
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect 931 1038 993 1076
rect 1893 1436 1907 1470
rect 1941 1436 1955 1470
rect 2855 1470 2917 1505
rect 1893 1398 1955 1436
rect 1893 1364 1907 1398
rect 1941 1364 1955 1398
rect 1893 1326 1955 1364
rect 1893 1292 1907 1326
rect 1941 1292 1955 1326
rect 1893 1254 1955 1292
rect 1893 1220 1907 1254
rect 1941 1220 1955 1254
rect 1893 1182 1955 1220
rect 1893 1148 1907 1182
rect 1941 1148 1955 1182
rect 1893 1110 1955 1148
rect 1893 1076 1907 1110
rect 1941 1076 1955 1110
rect 931 1004 945 1038
rect 979 1004 993 1038
rect 931 966 993 1004
rect -31 930 31 932
rect 931 932 945 966
rect 979 932 993 966
rect 1893 1038 1955 1076
rect 2855 1436 2869 1470
rect 2903 1436 2917 1470
rect 3817 1470 3879 1505
rect 2855 1398 2917 1436
rect 2855 1364 2869 1398
rect 2903 1364 2917 1398
rect 2855 1326 2917 1364
rect 2855 1292 2869 1326
rect 2903 1292 2917 1326
rect 2855 1254 2917 1292
rect 2855 1220 2869 1254
rect 2903 1220 2917 1254
rect 2855 1182 2917 1220
rect 2855 1148 2869 1182
rect 2903 1148 2917 1182
rect 2855 1110 2917 1148
rect 2855 1076 2869 1110
rect 2903 1076 2917 1110
rect 1893 1004 1907 1038
rect 1941 1004 1955 1038
rect 1893 966 1955 1004
rect 931 930 993 932
rect 1893 932 1907 966
rect 1941 932 1955 966
rect 2855 1038 2917 1076
rect 3817 1436 3831 1470
rect 3865 1436 3879 1470
rect 4779 1470 4841 1505
rect 3817 1398 3879 1436
rect 3817 1364 3831 1398
rect 3865 1364 3879 1398
rect 3817 1326 3879 1364
rect 3817 1292 3831 1326
rect 3865 1292 3879 1326
rect 3817 1254 3879 1292
rect 3817 1220 3831 1254
rect 3865 1220 3879 1254
rect 3817 1182 3879 1220
rect 3817 1148 3831 1182
rect 3865 1148 3879 1182
rect 3817 1110 3879 1148
rect 3817 1076 3831 1110
rect 3865 1076 3879 1110
rect 2855 1004 2869 1038
rect 2903 1004 2917 1038
rect 2855 966 2917 1004
rect 1893 930 1955 932
rect 2855 932 2869 966
rect 2903 932 2917 966
rect 3817 1038 3879 1076
rect 4779 1436 4793 1470
rect 4827 1436 4841 1470
rect 5741 1470 5803 1505
rect 4779 1398 4841 1436
rect 4779 1364 4793 1398
rect 4827 1364 4841 1398
rect 4779 1326 4841 1364
rect 4779 1292 4793 1326
rect 4827 1292 4841 1326
rect 4779 1254 4841 1292
rect 4779 1220 4793 1254
rect 4827 1220 4841 1254
rect 4779 1182 4841 1220
rect 4779 1148 4793 1182
rect 4827 1148 4841 1182
rect 4779 1110 4841 1148
rect 4779 1076 4793 1110
rect 4827 1076 4841 1110
rect 3817 1004 3831 1038
rect 3865 1004 3879 1038
rect 3817 966 3879 1004
rect 2855 930 2917 932
rect 3817 932 3831 966
rect 3865 932 3879 966
rect 4779 1038 4841 1076
rect 5741 1436 5755 1470
rect 5789 1436 5803 1470
rect 5741 1398 5803 1436
rect 5741 1364 5755 1398
rect 5789 1364 5803 1398
rect 5741 1326 5803 1364
rect 5741 1292 5755 1326
rect 5789 1292 5803 1326
rect 5741 1254 5803 1292
rect 5741 1220 5755 1254
rect 5789 1220 5803 1254
rect 5741 1182 5803 1220
rect 5741 1148 5755 1182
rect 5789 1148 5803 1182
rect 5741 1110 5803 1148
rect 5741 1076 5755 1110
rect 5789 1076 5803 1110
rect 4779 1004 4793 1038
rect 4827 1004 4841 1038
rect 4779 966 4841 1004
rect 3817 930 3879 932
rect 4779 932 4793 966
rect 4827 932 4841 966
rect 5741 1038 5803 1076
rect 5741 1004 5755 1038
rect 5789 1004 5803 1038
rect 5741 966 5803 1004
rect 4779 930 4841 932
rect 5741 932 5755 966
rect 5789 932 5803 966
rect 5741 930 5803 932
rect -31 868 5803 930
<< psubdiffcont >>
rect -17 512 17 546
rect 945 512 979 546
rect 1907 512 1941 546
rect 2869 512 2903 546
rect 3831 512 3865 546
rect 4793 512 4827 546
rect 5755 512 5789 546
rect -17 440 17 474
rect -17 368 17 402
rect 945 440 979 474
rect -17 296 17 330
rect -17 224 17 258
rect -17 152 17 186
rect -17 80 17 114
rect 945 368 979 402
rect 1907 440 1941 474
rect 945 296 979 330
rect 945 224 979 258
rect 945 152 979 186
rect 945 80 979 114
rect 1907 368 1941 402
rect 2869 440 2903 474
rect 1907 296 1941 330
rect 1907 224 1941 258
rect 1907 152 1941 186
rect 1907 80 1941 114
rect 2869 368 2903 402
rect 3831 440 3865 474
rect 2869 296 2903 330
rect 2869 224 2903 258
rect 2869 152 2903 186
rect 2869 80 2903 114
rect 3831 368 3865 402
rect 4793 440 4827 474
rect 3831 296 3865 330
rect 3831 224 3865 258
rect 3831 152 3865 186
rect 3831 80 3865 114
rect 4793 368 4827 402
rect 5755 440 5789 474
rect 4793 296 4827 330
rect 4793 224 4827 258
rect 4793 152 4827 186
rect 4793 80 4827 114
rect 5755 368 5789 402
rect 5755 296 5789 330
rect 5755 224 5789 258
rect 5755 152 5789 186
rect 5755 80 5789 114
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 343 13 377 47
rect 415 13 449 47
rect 513 13 547 47
rect 585 13 619 47
rect 657 13 691 47
rect 729 13 763 47
rect 801 13 835 47
rect 873 13 907 47
rect 1017 13 1051 47
rect 1089 13 1123 47
rect 1161 13 1195 47
rect 1233 13 1267 47
rect 1305 13 1339 47
rect 1377 13 1411 47
rect 1475 13 1509 47
rect 1547 13 1581 47
rect 1619 13 1653 47
rect 1691 13 1725 47
rect 1763 13 1797 47
rect 1835 13 1869 47
rect 1979 13 2013 47
rect 2051 13 2085 47
rect 2123 13 2157 47
rect 2195 13 2229 47
rect 2267 13 2301 47
rect 2339 13 2373 47
rect 2437 13 2471 47
rect 2509 13 2543 47
rect 2581 13 2615 47
rect 2653 13 2687 47
rect 2725 13 2759 47
rect 2797 13 2831 47
rect 2941 13 2975 47
rect 3013 13 3047 47
rect 3085 13 3119 47
rect 3157 13 3191 47
rect 3229 13 3263 47
rect 3301 13 3335 47
rect 3399 13 3433 47
rect 3471 13 3505 47
rect 3543 13 3577 47
rect 3615 13 3649 47
rect 3687 13 3721 47
rect 3759 13 3793 47
rect 3903 13 3937 47
rect 3975 13 4009 47
rect 4047 13 4081 47
rect 4119 13 4153 47
rect 4191 13 4225 47
rect 4263 13 4297 47
rect 4361 13 4395 47
rect 4433 13 4467 47
rect 4505 13 4539 47
rect 4577 13 4611 47
rect 4649 13 4683 47
rect 4721 13 4755 47
rect 4865 13 4899 47
rect 4937 13 4971 47
rect 5009 13 5043 47
rect 5081 13 5115 47
rect 5153 13 5187 47
rect 5225 13 5259 47
rect 5323 13 5357 47
rect 5395 13 5429 47
rect 5467 13 5501 47
rect 5539 13 5573 47
rect 5611 13 5645 47
rect 5683 13 5717 47
<< nsubdiffcont >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 343 1505 377 1539
rect 415 1505 449 1539
rect 513 1505 547 1539
rect 585 1505 619 1539
rect 657 1505 691 1539
rect 729 1505 763 1539
rect 801 1505 835 1539
rect 873 1505 907 1539
rect 1017 1505 1051 1539
rect 1089 1505 1123 1539
rect 1161 1505 1195 1539
rect 1233 1505 1267 1539
rect 1305 1505 1339 1539
rect 1377 1505 1411 1539
rect 1475 1505 1509 1539
rect 1547 1505 1581 1539
rect 1619 1505 1653 1539
rect 1691 1505 1725 1539
rect 1763 1505 1797 1539
rect 1835 1505 1869 1539
rect 1979 1505 2013 1539
rect 2051 1505 2085 1539
rect 2123 1505 2157 1539
rect 2195 1505 2229 1539
rect 2267 1505 2301 1539
rect 2339 1505 2373 1539
rect 2437 1505 2471 1539
rect 2509 1505 2543 1539
rect 2581 1505 2615 1539
rect 2653 1505 2687 1539
rect 2725 1505 2759 1539
rect 2797 1505 2831 1539
rect 2941 1505 2975 1539
rect 3013 1505 3047 1539
rect 3085 1505 3119 1539
rect 3157 1505 3191 1539
rect 3229 1505 3263 1539
rect 3301 1505 3335 1539
rect 3399 1505 3433 1539
rect 3471 1505 3505 1539
rect 3543 1505 3577 1539
rect 3615 1505 3649 1539
rect 3687 1505 3721 1539
rect 3759 1505 3793 1539
rect 3903 1505 3937 1539
rect 3975 1505 4009 1539
rect 4047 1505 4081 1539
rect 4119 1505 4153 1539
rect 4191 1505 4225 1539
rect 4263 1505 4297 1539
rect 4361 1505 4395 1539
rect 4433 1505 4467 1539
rect 4505 1505 4539 1539
rect 4577 1505 4611 1539
rect 4649 1505 4683 1539
rect 4721 1505 4755 1539
rect 4865 1505 4899 1539
rect 4937 1505 4971 1539
rect 5009 1505 5043 1539
rect 5081 1505 5115 1539
rect 5153 1505 5187 1539
rect 5225 1505 5259 1539
rect 5323 1505 5357 1539
rect 5395 1505 5429 1539
rect 5467 1505 5501 1539
rect 5539 1505 5573 1539
rect 5611 1505 5645 1539
rect 5683 1505 5717 1539
rect -17 1436 17 1470
rect -17 1364 17 1398
rect -17 1292 17 1326
rect -17 1220 17 1254
rect -17 1148 17 1182
rect -17 1076 17 1110
rect 945 1436 979 1470
rect 945 1364 979 1398
rect 945 1292 979 1326
rect 945 1220 979 1254
rect 945 1148 979 1182
rect 945 1076 979 1110
rect -17 1004 17 1038
rect -17 932 17 966
rect 1907 1436 1941 1470
rect 1907 1364 1941 1398
rect 1907 1292 1941 1326
rect 1907 1220 1941 1254
rect 1907 1148 1941 1182
rect 1907 1076 1941 1110
rect 945 1004 979 1038
rect 945 932 979 966
rect 2869 1436 2903 1470
rect 2869 1364 2903 1398
rect 2869 1292 2903 1326
rect 2869 1220 2903 1254
rect 2869 1148 2903 1182
rect 2869 1076 2903 1110
rect 1907 1004 1941 1038
rect 1907 932 1941 966
rect 3831 1436 3865 1470
rect 3831 1364 3865 1398
rect 3831 1292 3865 1326
rect 3831 1220 3865 1254
rect 3831 1148 3865 1182
rect 3831 1076 3865 1110
rect 2869 1004 2903 1038
rect 2869 932 2903 966
rect 4793 1436 4827 1470
rect 4793 1364 4827 1398
rect 4793 1292 4827 1326
rect 4793 1220 4827 1254
rect 4793 1148 4827 1182
rect 4793 1076 4827 1110
rect 3831 1004 3865 1038
rect 3831 932 3865 966
rect 5755 1436 5789 1470
rect 5755 1364 5789 1398
rect 5755 1292 5789 1326
rect 5755 1220 5789 1254
rect 5755 1148 5789 1182
rect 5755 1076 5789 1110
rect 4793 1004 4827 1038
rect 4793 932 4827 966
rect 5755 1004 5789 1038
rect 5755 932 5789 966
<< poly >>
rect 247 1450 277 1476
rect 335 1450 365 1476
rect 423 1450 453 1476
rect 511 1450 541 1476
rect 599 1450 629 1476
rect 687 1450 717 1476
rect 1209 1450 1239 1476
rect 1297 1450 1327 1476
rect 1385 1450 1415 1476
rect 1473 1450 1503 1476
rect 1561 1450 1591 1476
rect 1649 1450 1679 1476
rect 247 1019 277 1050
rect 335 1019 365 1050
rect 423 1019 453 1050
rect 511 1019 541 1050
rect 195 1003 365 1019
rect 195 969 205 1003
rect 239 989 365 1003
rect 417 1003 541 1019
rect 239 969 249 989
rect 195 953 249 969
rect 417 969 427 1003
rect 461 989 541 1003
rect 599 1019 629 1050
rect 687 1019 717 1050
rect 599 1003 717 1019
rect 599 989 649 1003
rect 461 969 471 989
rect 417 953 471 969
rect 639 969 649 989
rect 683 989 717 1003
rect 2171 1450 2201 1476
rect 2259 1450 2289 1476
rect 2347 1450 2377 1476
rect 2435 1450 2465 1476
rect 2523 1450 2553 1476
rect 2611 1450 2641 1476
rect 1209 1019 1239 1050
rect 1297 1019 1327 1050
rect 1385 1019 1415 1050
rect 1473 1019 1503 1050
rect 683 969 693 989
rect 639 953 693 969
rect 1157 1003 1327 1019
rect 1157 969 1167 1003
rect 1201 989 1327 1003
rect 1379 1003 1503 1019
rect 1201 969 1211 989
rect 1157 953 1211 969
rect 1379 969 1389 1003
rect 1423 989 1503 1003
rect 1561 1019 1591 1050
rect 1649 1019 1679 1050
rect 1561 1003 1679 1019
rect 1561 989 1611 1003
rect 1423 969 1433 989
rect 1379 953 1433 969
rect 1601 969 1611 989
rect 1645 989 1679 1003
rect 3133 1450 3163 1476
rect 3221 1450 3251 1476
rect 3309 1450 3339 1476
rect 3397 1450 3427 1476
rect 3485 1450 3515 1476
rect 3573 1450 3603 1476
rect 2171 1019 2201 1050
rect 2259 1019 2289 1050
rect 2347 1019 2377 1050
rect 2435 1019 2465 1050
rect 1645 969 1655 989
rect 1601 953 1655 969
rect 2119 1003 2289 1019
rect 2119 969 2129 1003
rect 2163 989 2289 1003
rect 2341 1003 2465 1019
rect 2163 969 2173 989
rect 2119 953 2173 969
rect 2341 969 2351 1003
rect 2385 989 2465 1003
rect 2523 1019 2553 1050
rect 2611 1019 2641 1050
rect 2523 1003 2641 1019
rect 2523 989 2573 1003
rect 2385 969 2395 989
rect 2341 953 2395 969
rect 2563 969 2573 989
rect 2607 989 2641 1003
rect 4095 1450 4125 1476
rect 4183 1450 4213 1476
rect 4271 1450 4301 1476
rect 4359 1450 4389 1476
rect 4447 1450 4477 1476
rect 4535 1450 4565 1476
rect 3133 1019 3163 1050
rect 3221 1019 3251 1050
rect 3309 1019 3339 1050
rect 3397 1019 3427 1050
rect 2607 969 2617 989
rect 2563 953 2617 969
rect 3081 1003 3251 1019
rect 3081 969 3091 1003
rect 3125 989 3251 1003
rect 3303 1003 3427 1019
rect 3125 969 3135 989
rect 3081 953 3135 969
rect 3303 969 3313 1003
rect 3347 989 3427 1003
rect 3485 1019 3515 1050
rect 3573 1019 3603 1050
rect 3485 1003 3603 1019
rect 3485 989 3535 1003
rect 3347 969 3357 989
rect 3303 953 3357 969
rect 3525 969 3535 989
rect 3569 989 3603 1003
rect 5057 1450 5087 1476
rect 5145 1450 5175 1476
rect 5233 1450 5263 1476
rect 5321 1450 5351 1476
rect 5409 1450 5439 1476
rect 5497 1450 5527 1476
rect 4095 1019 4125 1050
rect 4183 1019 4213 1050
rect 4271 1019 4301 1050
rect 4359 1019 4389 1050
rect 3569 969 3579 989
rect 3525 953 3579 969
rect 4043 1003 4213 1019
rect 4043 969 4053 1003
rect 4087 989 4213 1003
rect 4265 1003 4389 1019
rect 4087 969 4097 989
rect 4043 953 4097 969
rect 4265 969 4275 1003
rect 4309 989 4389 1003
rect 4447 1019 4477 1050
rect 4535 1019 4565 1050
rect 4447 1003 4565 1019
rect 4447 989 4497 1003
rect 4309 969 4319 989
rect 4265 953 4319 969
rect 4487 969 4497 989
rect 4531 989 4565 1003
rect 5057 1019 5087 1050
rect 5145 1019 5175 1050
rect 5233 1019 5263 1050
rect 5321 1019 5351 1050
rect 4531 969 4541 989
rect 4487 953 4541 969
rect 5005 1003 5175 1019
rect 5005 969 5015 1003
rect 5049 989 5175 1003
rect 5227 1003 5351 1019
rect 5049 969 5059 989
rect 5005 953 5059 969
rect 5227 969 5237 1003
rect 5271 989 5351 1003
rect 5409 1019 5439 1050
rect 5497 1019 5527 1050
rect 5409 1003 5527 1019
rect 5409 989 5459 1003
rect 5271 969 5281 989
rect 5227 953 5281 969
rect 5449 969 5459 989
rect 5493 989 5527 1003
rect 5493 969 5503 989
rect 5449 953 5503 969
rect 195 461 249 477
rect 195 441 205 461
rect 147 427 205 441
rect 239 427 249 461
rect 147 411 249 427
rect 417 461 471 477
rect 417 427 427 461
rect 461 441 471 461
rect 639 461 693 477
rect 461 427 477 441
rect 417 411 477 427
rect 639 427 649 461
rect 683 427 693 461
rect 639 411 693 427
rect 1157 461 1211 477
rect 1157 441 1167 461
rect 147 379 177 411
rect 447 379 477 411
rect 649 379 679 411
rect 1109 427 1167 441
rect 1201 427 1211 461
rect 1109 411 1211 427
rect 1379 461 1433 477
rect 1379 427 1389 461
rect 1423 441 1433 461
rect 1601 461 1655 477
rect 1423 427 1439 441
rect 1379 411 1439 427
rect 1601 427 1611 461
rect 1645 427 1655 461
rect 1601 411 1655 427
rect 2119 461 2173 477
rect 2119 441 2129 461
rect 1109 379 1139 411
rect 1409 379 1439 411
rect 1611 379 1641 411
rect 2071 427 2129 441
rect 2163 427 2173 461
rect 2071 411 2173 427
rect 2341 461 2395 477
rect 2341 427 2351 461
rect 2385 441 2395 461
rect 2563 461 2617 477
rect 2385 427 2401 441
rect 2341 411 2401 427
rect 2563 427 2573 461
rect 2607 427 2617 461
rect 2563 411 2617 427
rect 3081 461 3135 477
rect 3081 441 3091 461
rect 2071 379 2101 411
rect 2371 379 2401 411
rect 2573 379 2603 411
rect 3033 427 3091 441
rect 3125 427 3135 461
rect 3033 411 3135 427
rect 3303 461 3357 477
rect 3303 427 3313 461
rect 3347 441 3357 461
rect 3525 461 3579 477
rect 3347 427 3363 441
rect 3303 411 3363 427
rect 3525 427 3535 461
rect 3569 427 3579 461
rect 3525 411 3579 427
rect 4043 461 4097 477
rect 4043 441 4053 461
rect 3033 379 3063 411
rect 3333 379 3363 411
rect 3535 379 3565 411
rect 3995 427 4053 441
rect 4087 427 4097 461
rect 3995 411 4097 427
rect 4265 461 4319 477
rect 4265 427 4275 461
rect 4309 441 4319 461
rect 4487 461 4541 477
rect 4309 427 4325 441
rect 4265 411 4325 427
rect 4487 427 4497 461
rect 4531 427 4541 461
rect 4487 411 4541 427
rect 5005 461 5059 477
rect 5005 441 5015 461
rect 3995 379 4025 411
rect 4295 379 4325 411
rect 4497 379 4527 411
rect 4957 427 5015 441
rect 5049 427 5059 461
rect 4957 411 5059 427
rect 5227 461 5281 477
rect 5227 427 5237 461
rect 5271 441 5281 461
rect 5449 461 5503 477
rect 5271 427 5287 441
rect 5227 411 5287 427
rect 5449 427 5459 461
rect 5493 427 5503 461
rect 5449 411 5503 427
rect 4957 379 4987 411
rect 5257 379 5287 411
rect 5459 379 5489 411
<< polycont >>
rect 205 969 239 1003
rect 427 969 461 1003
rect 649 969 683 1003
rect 1167 969 1201 1003
rect 1389 969 1423 1003
rect 1611 969 1645 1003
rect 2129 969 2163 1003
rect 2351 969 2385 1003
rect 2573 969 2607 1003
rect 3091 969 3125 1003
rect 3313 969 3347 1003
rect 3535 969 3569 1003
rect 4053 969 4087 1003
rect 4275 969 4309 1003
rect 4497 969 4531 1003
rect 5015 969 5049 1003
rect 5237 969 5271 1003
rect 5459 969 5493 1003
rect 205 427 239 461
rect 427 427 461 461
rect 649 427 683 461
rect 1167 427 1201 461
rect 1389 427 1423 461
rect 1611 427 1645 461
rect 2129 427 2163 461
rect 2351 427 2385 461
rect 2573 427 2607 461
rect 3091 427 3125 461
rect 3313 427 3347 461
rect 3535 427 3569 461
rect 4053 427 4087 461
rect 4275 427 4309 461
rect 4497 427 4531 461
rect 5015 427 5049 461
rect 5237 427 5271 461
rect 5459 427 5493 461
<< locali >>
rect -31 1539 5803 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 343 1539
rect 377 1505 415 1539
rect 449 1505 513 1539
rect 547 1505 585 1539
rect 619 1505 657 1539
rect 691 1505 729 1539
rect 763 1505 801 1539
rect 835 1505 873 1539
rect 907 1505 1017 1539
rect 1051 1505 1089 1539
rect 1123 1505 1161 1539
rect 1195 1505 1233 1539
rect 1267 1505 1305 1539
rect 1339 1505 1377 1539
rect 1411 1505 1475 1539
rect 1509 1505 1547 1539
rect 1581 1505 1619 1539
rect 1653 1505 1691 1539
rect 1725 1505 1763 1539
rect 1797 1505 1835 1539
rect 1869 1505 1979 1539
rect 2013 1505 2051 1539
rect 2085 1505 2123 1539
rect 2157 1505 2195 1539
rect 2229 1505 2267 1539
rect 2301 1505 2339 1539
rect 2373 1505 2437 1539
rect 2471 1505 2509 1539
rect 2543 1505 2581 1539
rect 2615 1505 2653 1539
rect 2687 1505 2725 1539
rect 2759 1505 2797 1539
rect 2831 1505 2941 1539
rect 2975 1505 3013 1539
rect 3047 1505 3085 1539
rect 3119 1505 3157 1539
rect 3191 1505 3229 1539
rect 3263 1505 3301 1539
rect 3335 1505 3399 1539
rect 3433 1505 3471 1539
rect 3505 1505 3543 1539
rect 3577 1505 3615 1539
rect 3649 1505 3687 1539
rect 3721 1505 3759 1539
rect 3793 1505 3903 1539
rect 3937 1505 3975 1539
rect 4009 1505 4047 1539
rect 4081 1505 4119 1539
rect 4153 1505 4191 1539
rect 4225 1505 4263 1539
rect 4297 1505 4361 1539
rect 4395 1505 4433 1539
rect 4467 1505 4505 1539
rect 4539 1505 4577 1539
rect 4611 1505 4649 1539
rect 4683 1505 4721 1539
rect 4755 1505 4865 1539
rect 4899 1505 4937 1539
rect 4971 1505 5009 1539
rect 5043 1505 5081 1539
rect 5115 1505 5153 1539
rect 5187 1505 5225 1539
rect 5259 1505 5323 1539
rect 5357 1505 5395 1539
rect 5429 1505 5467 1539
rect 5501 1505 5539 1539
rect 5573 1505 5611 1539
rect 5645 1505 5683 1539
rect 5717 1505 5803 1539
rect -31 1492 5803 1505
rect -31 1470 31 1492
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect 201 1412 235 1492
rect 201 1344 235 1378
rect 201 1276 235 1310
rect 201 1208 235 1242
rect 201 1139 235 1174
rect 201 1089 235 1105
rect 289 1412 323 1450
rect 289 1344 323 1378
rect 289 1276 323 1310
rect 289 1208 323 1242
rect 289 1139 323 1174
rect 377 1412 411 1492
rect 377 1344 411 1378
rect 377 1276 411 1310
rect 377 1208 411 1242
rect 377 1157 411 1174
rect 465 1412 499 1450
rect 465 1344 499 1378
rect 465 1276 499 1310
rect 465 1208 499 1242
rect 289 1094 323 1105
rect 465 1139 499 1174
rect 553 1412 587 1492
rect 553 1344 587 1378
rect 553 1276 587 1310
rect 553 1208 587 1242
rect 553 1157 587 1174
rect 641 1412 675 1450
rect 641 1344 675 1378
rect 641 1276 675 1310
rect 641 1208 675 1242
rect 465 1094 499 1105
rect 641 1139 675 1174
rect 729 1412 763 1492
rect 729 1344 763 1378
rect 729 1276 763 1310
rect 729 1208 763 1242
rect 729 1157 763 1174
rect 931 1470 993 1492
rect 931 1436 945 1470
rect 979 1436 993 1470
rect 931 1398 993 1436
rect 931 1364 945 1398
rect 979 1364 993 1398
rect 931 1326 993 1364
rect 931 1292 945 1326
rect 979 1292 993 1326
rect 931 1254 993 1292
rect 931 1220 945 1254
rect 979 1220 993 1254
rect 931 1182 993 1220
rect 641 1094 675 1105
rect 931 1148 945 1182
rect 979 1148 993 1182
rect 931 1110 993 1148
rect -31 1038 31 1076
rect 289 1060 831 1094
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect -31 868 31 932
rect 205 1003 239 1019
rect 205 609 239 969
rect -31 546 31 572
rect -31 512 -17 546
rect 17 512 31 546
rect -31 474 31 512
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect 205 461 239 575
rect 205 411 239 427
rect 427 1003 461 1019
rect 427 905 461 969
rect 427 461 461 871
rect 427 411 461 427
rect 649 1003 683 1019
rect 649 757 683 969
rect 649 461 683 723
rect 649 411 683 427
rect 797 610 831 1060
rect 931 1076 945 1110
rect 979 1076 993 1110
rect 1163 1412 1197 1492
rect 1163 1344 1197 1378
rect 1163 1276 1197 1310
rect 1163 1208 1197 1242
rect 1163 1139 1197 1174
rect 1163 1089 1197 1105
rect 1251 1412 1285 1450
rect 1251 1344 1285 1378
rect 1251 1276 1285 1310
rect 1251 1208 1285 1242
rect 1251 1139 1285 1174
rect 1339 1412 1373 1492
rect 1339 1344 1373 1378
rect 1339 1276 1373 1310
rect 1339 1208 1373 1242
rect 1339 1157 1373 1174
rect 1427 1412 1461 1450
rect 1427 1344 1461 1378
rect 1427 1276 1461 1310
rect 1427 1208 1461 1242
rect 1251 1094 1285 1105
rect 1427 1139 1461 1174
rect 1515 1412 1549 1492
rect 1515 1344 1549 1378
rect 1515 1276 1549 1310
rect 1515 1208 1549 1242
rect 1515 1157 1549 1174
rect 1603 1412 1637 1450
rect 1603 1344 1637 1378
rect 1603 1276 1637 1310
rect 1603 1208 1637 1242
rect 1427 1094 1461 1105
rect 1603 1139 1637 1174
rect 1691 1412 1725 1492
rect 1691 1344 1725 1378
rect 1691 1276 1725 1310
rect 1691 1208 1725 1242
rect 1691 1157 1725 1174
rect 1893 1470 1955 1492
rect 1893 1436 1907 1470
rect 1941 1436 1955 1470
rect 1893 1398 1955 1436
rect 1893 1364 1907 1398
rect 1941 1364 1955 1398
rect 1893 1326 1955 1364
rect 1893 1292 1907 1326
rect 1941 1292 1955 1326
rect 1893 1254 1955 1292
rect 1893 1220 1907 1254
rect 1941 1220 1955 1254
rect 1893 1182 1955 1220
rect 1603 1094 1637 1105
rect 1893 1148 1907 1182
rect 1941 1148 1955 1182
rect 1893 1110 1955 1148
rect 931 1038 993 1076
rect 1251 1060 1793 1094
rect 931 1004 945 1038
rect 979 1004 993 1038
rect 931 966 993 1004
rect 931 932 945 966
rect 979 932 993 966
rect 931 868 993 932
rect 1167 1003 1201 1019
rect -31 368 -17 402
rect 17 368 31 402
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect 101 363 135 379
rect 295 363 329 379
rect 489 363 523 379
rect 135 329 198 363
rect 232 329 295 363
rect 329 329 392 363
rect 426 329 489 363
rect 101 291 135 329
rect 101 223 135 257
rect 295 291 329 329
rect 489 313 523 329
rect 603 363 637 379
rect 797 378 831 576
rect 1167 610 1201 969
rect 603 291 637 329
rect 101 153 135 189
rect 101 103 135 119
rect 198 238 232 254
rect -31 62 31 80
rect 198 62 232 204
rect 295 223 329 257
rect 393 244 427 260
rect 603 244 637 257
rect 427 223 637 244
rect 427 210 603 223
rect 393 194 427 210
rect 295 153 329 189
rect 700 344 831 378
rect 931 546 993 572
rect 931 512 945 546
rect 979 512 993 546
rect 931 474 993 512
rect 931 440 945 474
rect 979 440 993 474
rect 931 402 993 440
rect 1167 461 1201 576
rect 1167 411 1201 427
rect 1389 1003 1423 1019
rect 1389 683 1423 969
rect 1611 1003 1645 1019
rect 1611 847 1645 969
rect 1610 831 1645 847
rect 1644 797 1645 831
rect 1610 781 1645 797
rect 1389 461 1423 649
rect 1389 411 1423 427
rect 1611 461 1645 781
rect 1611 411 1645 427
rect 1759 757 1793 1060
rect 1893 1076 1907 1110
rect 1941 1076 1955 1110
rect 2125 1412 2159 1492
rect 2125 1344 2159 1378
rect 2125 1276 2159 1310
rect 2125 1208 2159 1242
rect 2125 1139 2159 1174
rect 2125 1089 2159 1105
rect 2213 1412 2247 1450
rect 2213 1344 2247 1378
rect 2213 1276 2247 1310
rect 2213 1208 2247 1242
rect 2213 1139 2247 1174
rect 2301 1412 2335 1492
rect 2301 1344 2335 1378
rect 2301 1276 2335 1310
rect 2301 1208 2335 1242
rect 2301 1157 2335 1174
rect 2389 1412 2423 1450
rect 2389 1344 2423 1378
rect 2389 1276 2423 1310
rect 2389 1208 2423 1242
rect 2213 1094 2247 1105
rect 2389 1139 2423 1174
rect 2477 1412 2511 1492
rect 2477 1344 2511 1378
rect 2477 1276 2511 1310
rect 2477 1208 2511 1242
rect 2477 1157 2511 1174
rect 2565 1412 2599 1450
rect 2565 1344 2599 1378
rect 2565 1276 2599 1310
rect 2565 1208 2599 1242
rect 2389 1094 2423 1105
rect 2565 1139 2599 1174
rect 2653 1412 2687 1492
rect 2653 1344 2687 1378
rect 2653 1276 2687 1310
rect 2653 1208 2687 1242
rect 2653 1157 2687 1174
rect 2855 1470 2917 1492
rect 2855 1436 2869 1470
rect 2903 1436 2917 1470
rect 2855 1398 2917 1436
rect 2855 1364 2869 1398
rect 2903 1364 2917 1398
rect 2855 1326 2917 1364
rect 2855 1292 2869 1326
rect 2903 1292 2917 1326
rect 2855 1254 2917 1292
rect 2855 1220 2869 1254
rect 2903 1220 2917 1254
rect 2855 1182 2917 1220
rect 2565 1094 2599 1105
rect 2855 1148 2869 1182
rect 2903 1148 2917 1182
rect 2855 1110 2917 1148
rect 1893 1038 1955 1076
rect 2213 1060 2755 1094
rect 1893 1004 1907 1038
rect 1941 1004 1955 1038
rect 1893 966 1955 1004
rect 1893 932 1907 966
rect 1941 932 1955 966
rect 1893 868 1955 932
rect 2129 1003 2163 1019
rect 931 368 945 402
rect 979 368 993 402
rect 700 247 734 344
rect 931 330 993 368
rect 700 197 734 213
rect 797 291 831 307
rect 797 223 831 257
rect 489 153 523 169
rect 329 119 392 153
rect 426 119 489 153
rect 295 103 329 119
rect 489 103 523 119
rect 603 153 637 189
rect 797 153 831 189
rect 637 119 700 153
rect 734 119 797 153
rect 603 103 637 119
rect 797 103 831 119
rect 931 296 945 330
rect 979 296 993 330
rect 931 258 993 296
rect 931 224 945 258
rect 979 224 993 258
rect 931 186 993 224
rect 931 152 945 186
rect 979 152 993 186
rect 931 114 993 152
rect 931 80 945 114
rect 979 80 993 114
rect 1063 363 1097 379
rect 1257 363 1291 379
rect 1451 363 1485 379
rect 1097 329 1160 363
rect 1194 329 1257 363
rect 1291 329 1354 363
rect 1388 329 1451 363
rect 1063 291 1097 329
rect 1063 223 1097 257
rect 1257 291 1291 329
rect 1451 313 1485 329
rect 1565 363 1599 379
rect 1759 378 1793 723
rect 2129 610 2163 969
rect 1565 291 1599 329
rect 1063 153 1097 189
rect 1063 103 1097 119
rect 1160 238 1194 254
rect 931 62 993 80
rect 1160 62 1194 204
rect 1257 223 1291 257
rect 1355 244 1389 260
rect 1565 244 1599 257
rect 1389 223 1599 244
rect 1389 210 1565 223
rect 1355 194 1389 210
rect 1257 153 1291 189
rect 1662 344 1793 378
rect 1893 546 1955 572
rect 1893 512 1907 546
rect 1941 512 1955 546
rect 1893 474 1955 512
rect 1893 440 1907 474
rect 1941 440 1955 474
rect 1893 402 1955 440
rect 2129 461 2163 576
rect 2129 411 2163 427
rect 2351 1003 2385 1019
rect 2351 536 2385 969
rect 2351 461 2385 502
rect 2351 411 2385 427
rect 2573 1003 2607 1019
rect 2573 831 2607 969
rect 2573 461 2607 797
rect 2573 411 2607 427
rect 2721 609 2755 1060
rect 2855 1076 2869 1110
rect 2903 1076 2917 1110
rect 3087 1412 3121 1492
rect 3087 1344 3121 1378
rect 3087 1276 3121 1310
rect 3087 1208 3121 1242
rect 3087 1139 3121 1174
rect 3087 1089 3121 1105
rect 3175 1412 3209 1450
rect 3175 1344 3209 1378
rect 3175 1276 3209 1310
rect 3175 1208 3209 1242
rect 3175 1139 3209 1174
rect 3263 1412 3297 1492
rect 3263 1344 3297 1378
rect 3263 1276 3297 1310
rect 3263 1208 3297 1242
rect 3263 1157 3297 1174
rect 3351 1412 3385 1450
rect 3351 1344 3385 1378
rect 3351 1276 3385 1310
rect 3351 1208 3385 1242
rect 3175 1094 3209 1105
rect 3351 1139 3385 1174
rect 3439 1412 3473 1492
rect 3439 1344 3473 1378
rect 3439 1276 3473 1310
rect 3439 1208 3473 1242
rect 3439 1157 3473 1174
rect 3527 1412 3561 1450
rect 3527 1344 3561 1378
rect 3527 1276 3561 1310
rect 3527 1208 3561 1242
rect 3351 1094 3385 1105
rect 3527 1139 3561 1174
rect 3615 1412 3649 1492
rect 3615 1344 3649 1378
rect 3615 1276 3649 1310
rect 3615 1208 3649 1242
rect 3615 1157 3649 1174
rect 3817 1470 3879 1492
rect 3817 1436 3831 1470
rect 3865 1436 3879 1470
rect 3817 1398 3879 1436
rect 3817 1364 3831 1398
rect 3865 1364 3879 1398
rect 3817 1326 3879 1364
rect 3817 1292 3831 1326
rect 3865 1292 3879 1326
rect 3817 1254 3879 1292
rect 3817 1220 3831 1254
rect 3865 1220 3879 1254
rect 3817 1182 3879 1220
rect 3527 1094 3561 1105
rect 3817 1148 3831 1182
rect 3865 1148 3879 1182
rect 3817 1110 3879 1148
rect 2855 1038 2917 1076
rect 3175 1060 3717 1094
rect 2855 1004 2869 1038
rect 2903 1004 2917 1038
rect 2855 966 2917 1004
rect 2855 932 2869 966
rect 2903 932 2917 966
rect 2855 868 2917 932
rect 3091 1003 3125 1019
rect 1893 368 1907 402
rect 1941 368 1955 402
rect 1662 247 1696 344
rect 1893 330 1955 368
rect 1662 197 1696 213
rect 1759 291 1793 307
rect 1759 223 1793 257
rect 1451 153 1485 169
rect 1291 119 1354 153
rect 1388 119 1451 153
rect 1257 103 1291 119
rect 1451 103 1485 119
rect 1565 153 1599 189
rect 1759 153 1793 189
rect 1599 119 1662 153
rect 1696 119 1759 153
rect 1565 103 1599 119
rect 1759 103 1793 119
rect 1893 296 1907 330
rect 1941 296 1955 330
rect 1893 258 1955 296
rect 1893 224 1907 258
rect 1941 224 1955 258
rect 1893 186 1955 224
rect 1893 152 1907 186
rect 1941 152 1955 186
rect 1893 114 1955 152
rect 1893 80 1907 114
rect 1941 80 1955 114
rect 2025 363 2059 379
rect 2219 363 2253 379
rect 2413 363 2447 379
rect 2059 329 2122 363
rect 2156 329 2219 363
rect 2253 329 2316 363
rect 2350 329 2413 363
rect 2025 291 2059 329
rect 2025 223 2059 257
rect 2219 291 2253 329
rect 2413 313 2447 329
rect 2527 363 2561 379
rect 2721 378 2755 575
rect 3091 609 3125 969
rect 2527 291 2561 329
rect 2025 153 2059 189
rect 2025 103 2059 119
rect 2122 238 2156 254
rect 1893 62 1955 80
rect 2122 62 2156 204
rect 2219 223 2253 257
rect 2317 244 2351 260
rect 2527 244 2561 257
rect 2351 223 2561 244
rect 2351 210 2527 223
rect 2317 194 2351 210
rect 2219 153 2253 189
rect 2624 344 2755 378
rect 2855 546 2917 572
rect 2855 512 2869 546
rect 2903 512 2917 546
rect 2855 474 2917 512
rect 2855 440 2869 474
rect 2903 440 2917 474
rect 2855 402 2917 440
rect 3091 461 3125 575
rect 3091 411 3125 427
rect 3313 1003 3347 1019
rect 3313 683 3347 969
rect 3313 461 3347 649
rect 3313 411 3347 427
rect 3535 1003 3569 1019
rect 3535 905 3569 969
rect 3535 461 3569 871
rect 3535 411 3569 427
rect 3683 831 3717 1060
rect 3817 1076 3831 1110
rect 3865 1076 3879 1110
rect 4049 1412 4083 1492
rect 4049 1344 4083 1378
rect 4049 1276 4083 1310
rect 4049 1208 4083 1242
rect 4049 1139 4083 1174
rect 4049 1089 4083 1105
rect 4137 1412 4171 1450
rect 4137 1344 4171 1378
rect 4137 1276 4171 1310
rect 4137 1208 4171 1242
rect 4137 1139 4171 1174
rect 4225 1412 4259 1492
rect 4225 1344 4259 1378
rect 4225 1276 4259 1310
rect 4225 1208 4259 1242
rect 4225 1157 4259 1174
rect 4313 1412 4347 1450
rect 4313 1344 4347 1378
rect 4313 1276 4347 1310
rect 4313 1208 4347 1242
rect 4137 1094 4171 1105
rect 4313 1139 4347 1174
rect 4401 1412 4435 1492
rect 4401 1344 4435 1378
rect 4401 1276 4435 1310
rect 4401 1208 4435 1242
rect 4401 1157 4435 1174
rect 4489 1412 4523 1450
rect 4489 1344 4523 1378
rect 4489 1276 4523 1310
rect 4489 1208 4523 1242
rect 4313 1094 4347 1105
rect 4489 1139 4523 1174
rect 4577 1412 4611 1492
rect 4577 1344 4611 1378
rect 4577 1276 4611 1310
rect 4577 1208 4611 1242
rect 4577 1157 4611 1174
rect 4779 1470 4841 1492
rect 4779 1436 4793 1470
rect 4827 1436 4841 1470
rect 4779 1398 4841 1436
rect 4779 1364 4793 1398
rect 4827 1364 4841 1398
rect 4779 1326 4841 1364
rect 4779 1292 4793 1326
rect 4827 1292 4841 1326
rect 4779 1254 4841 1292
rect 4779 1220 4793 1254
rect 4827 1220 4841 1254
rect 4779 1182 4841 1220
rect 4489 1094 4523 1105
rect 4779 1148 4793 1182
rect 4827 1148 4841 1182
rect 4779 1110 4841 1148
rect 3817 1038 3879 1076
rect 4137 1060 4679 1094
rect 3817 1004 3831 1038
rect 3865 1004 3879 1038
rect 3817 966 3879 1004
rect 3817 932 3831 966
rect 3865 932 3879 966
rect 3817 868 3879 932
rect 4053 1003 4087 1019
rect 2855 368 2869 402
rect 2903 368 2917 402
rect 2624 247 2658 344
rect 2855 330 2917 368
rect 2624 197 2658 213
rect 2721 291 2755 307
rect 2721 223 2755 257
rect 2413 153 2447 169
rect 2253 119 2316 153
rect 2350 119 2413 153
rect 2219 103 2253 119
rect 2413 103 2447 119
rect 2527 153 2561 189
rect 2721 153 2755 189
rect 2561 119 2624 153
rect 2658 119 2721 153
rect 2527 103 2561 119
rect 2721 103 2755 119
rect 2855 296 2869 330
rect 2903 296 2917 330
rect 2855 258 2917 296
rect 2855 224 2869 258
rect 2903 224 2917 258
rect 2855 186 2917 224
rect 2855 152 2869 186
rect 2903 152 2917 186
rect 2855 114 2917 152
rect 2855 80 2869 114
rect 2903 80 2917 114
rect 2987 363 3021 379
rect 3181 363 3215 379
rect 3375 363 3409 379
rect 3021 329 3084 363
rect 3118 329 3181 363
rect 3215 329 3278 363
rect 3312 329 3375 363
rect 2987 291 3021 329
rect 2987 223 3021 257
rect 3181 291 3215 329
rect 3375 313 3409 329
rect 3489 363 3523 379
rect 3683 378 3717 797
rect 4053 757 4087 969
rect 3489 291 3523 329
rect 2987 153 3021 189
rect 2987 103 3021 119
rect 3084 238 3118 254
rect 2855 62 2917 80
rect 3084 62 3118 204
rect 3181 223 3215 257
rect 3279 244 3313 260
rect 3489 244 3523 257
rect 3313 223 3523 244
rect 3313 210 3489 223
rect 3279 194 3313 210
rect 3181 153 3215 189
rect 3586 344 3717 378
rect 3817 546 3879 572
rect 3817 512 3831 546
rect 3865 512 3879 546
rect 3817 474 3879 512
rect 3817 440 3831 474
rect 3865 440 3879 474
rect 3817 402 3879 440
rect 4053 461 4087 723
rect 4053 411 4087 427
rect 4275 1003 4309 1019
rect 4275 905 4309 969
rect 4275 461 4309 871
rect 4275 411 4309 427
rect 4497 1003 4531 1019
rect 4497 757 4531 969
rect 4497 461 4531 723
rect 4497 411 4531 427
rect 4645 683 4679 1060
rect 4779 1076 4793 1110
rect 4827 1076 4841 1110
rect 5011 1412 5045 1492
rect 5011 1344 5045 1378
rect 5011 1276 5045 1310
rect 5011 1208 5045 1242
rect 5011 1139 5045 1174
rect 5011 1089 5045 1105
rect 5099 1412 5133 1450
rect 5099 1344 5133 1378
rect 5099 1276 5133 1310
rect 5099 1208 5133 1242
rect 5099 1139 5133 1174
rect 5187 1412 5221 1492
rect 5187 1344 5221 1378
rect 5187 1276 5221 1310
rect 5187 1208 5221 1242
rect 5187 1157 5221 1174
rect 5275 1412 5309 1450
rect 5275 1344 5309 1378
rect 5275 1276 5309 1310
rect 5275 1208 5309 1242
rect 5099 1094 5133 1105
rect 5275 1139 5309 1174
rect 5363 1412 5397 1492
rect 5363 1344 5397 1378
rect 5363 1276 5397 1310
rect 5363 1208 5397 1242
rect 5363 1157 5397 1174
rect 5451 1412 5485 1450
rect 5451 1344 5485 1378
rect 5451 1276 5485 1310
rect 5451 1208 5485 1242
rect 5275 1094 5309 1105
rect 5451 1139 5485 1174
rect 5539 1412 5573 1492
rect 5539 1344 5573 1378
rect 5539 1276 5573 1310
rect 5539 1208 5573 1242
rect 5539 1157 5573 1174
rect 5741 1470 5803 1492
rect 5741 1436 5755 1470
rect 5789 1436 5803 1470
rect 5741 1398 5803 1436
rect 5741 1364 5755 1398
rect 5789 1364 5803 1398
rect 5741 1326 5803 1364
rect 5741 1292 5755 1326
rect 5789 1292 5803 1326
rect 5741 1254 5803 1292
rect 5741 1220 5755 1254
rect 5789 1220 5803 1254
rect 5741 1182 5803 1220
rect 5451 1094 5485 1105
rect 5741 1148 5755 1182
rect 5789 1148 5803 1182
rect 5741 1110 5803 1148
rect 4779 1038 4841 1076
rect 5099 1060 5641 1094
rect 4779 1004 4793 1038
rect 4827 1004 4841 1038
rect 4779 966 4841 1004
rect 4779 932 4793 966
rect 4827 932 4841 966
rect 4779 868 4841 932
rect 5015 1003 5049 1019
rect 3817 368 3831 402
rect 3865 368 3879 402
rect 3586 247 3620 344
rect 3817 330 3879 368
rect 3586 197 3620 213
rect 3683 291 3717 307
rect 3683 223 3717 257
rect 3375 153 3409 169
rect 3215 119 3278 153
rect 3312 119 3375 153
rect 3181 103 3215 119
rect 3375 103 3409 119
rect 3489 153 3523 189
rect 3683 153 3717 189
rect 3523 119 3586 153
rect 3620 119 3683 153
rect 3489 103 3523 119
rect 3683 103 3717 119
rect 3817 296 3831 330
rect 3865 296 3879 330
rect 3817 258 3879 296
rect 3817 224 3831 258
rect 3865 224 3879 258
rect 3817 186 3879 224
rect 3817 152 3831 186
rect 3865 152 3879 186
rect 3817 114 3879 152
rect 3817 80 3831 114
rect 3865 80 3879 114
rect 3949 363 3983 379
rect 4143 363 4177 379
rect 4337 363 4371 379
rect 3983 329 4046 363
rect 4080 329 4143 363
rect 4177 329 4240 363
rect 4274 329 4337 363
rect 3949 291 3983 329
rect 3949 223 3983 257
rect 4143 291 4177 329
rect 4337 313 4371 329
rect 4451 363 4485 379
rect 4645 378 4679 649
rect 5015 683 5049 969
rect 4451 291 4485 329
rect 3949 153 3983 189
rect 3949 103 3983 119
rect 4046 238 4080 254
rect 3817 62 3879 80
rect 4046 62 4080 204
rect 4143 223 4177 257
rect 4241 244 4275 260
rect 4451 244 4485 257
rect 4275 223 4485 244
rect 4275 210 4451 223
rect 4241 194 4275 210
rect 4143 153 4177 189
rect 4548 344 4679 378
rect 4779 546 4841 572
rect 4779 512 4793 546
rect 4827 512 4841 546
rect 4779 474 4841 512
rect 4779 440 4793 474
rect 4827 440 4841 474
rect 4779 402 4841 440
rect 5015 461 5049 649
rect 5015 411 5049 427
rect 5237 1003 5271 1019
rect 5237 535 5271 969
rect 5237 461 5271 501
rect 5237 411 5271 427
rect 5459 1003 5493 1019
rect 5459 831 5493 969
rect 5459 461 5493 797
rect 5459 411 5493 427
rect 5607 757 5641 1060
rect 5741 1076 5755 1110
rect 5789 1076 5803 1110
rect 5741 1038 5803 1076
rect 5741 1004 5755 1038
rect 5789 1004 5803 1038
rect 5741 966 5803 1004
rect 5741 932 5755 966
rect 5789 932 5803 966
rect 5741 868 5803 932
rect 4779 368 4793 402
rect 4827 368 4841 402
rect 4548 247 4582 344
rect 4779 330 4841 368
rect 4548 197 4582 213
rect 4645 291 4679 307
rect 4645 223 4679 257
rect 4337 153 4371 169
rect 4177 119 4240 153
rect 4274 119 4337 153
rect 4143 103 4177 119
rect 4337 103 4371 119
rect 4451 153 4485 189
rect 4645 153 4679 189
rect 4485 119 4548 153
rect 4582 119 4645 153
rect 4451 103 4485 119
rect 4645 103 4679 119
rect 4779 296 4793 330
rect 4827 296 4841 330
rect 4779 258 4841 296
rect 4779 224 4793 258
rect 4827 224 4841 258
rect 4779 186 4841 224
rect 4779 152 4793 186
rect 4827 152 4841 186
rect 4779 114 4841 152
rect 4779 80 4793 114
rect 4827 80 4841 114
rect 4911 363 4945 379
rect 5105 363 5139 379
rect 5299 363 5333 379
rect 4945 329 5008 363
rect 5042 329 5105 363
rect 5139 329 5202 363
rect 5236 329 5299 363
rect 4911 291 4945 329
rect 4911 223 4945 257
rect 5105 291 5139 329
rect 5299 313 5333 329
rect 5413 363 5447 379
rect 5607 378 5641 723
rect 5413 291 5447 329
rect 4911 153 4945 189
rect 4911 103 4945 119
rect 5008 238 5042 254
rect 4779 62 4841 80
rect 5008 62 5042 204
rect 5105 223 5139 257
rect 5203 244 5237 260
rect 5413 244 5447 257
rect 5237 223 5447 244
rect 5237 210 5413 223
rect 5203 194 5237 210
rect 5105 153 5139 189
rect 5510 344 5641 378
rect 5741 546 5803 572
rect 5741 512 5755 546
rect 5789 512 5803 546
rect 5741 474 5803 512
rect 5741 440 5755 474
rect 5789 440 5803 474
rect 5741 402 5803 440
rect 5741 368 5755 402
rect 5789 368 5803 402
rect 5510 247 5544 344
rect 5741 330 5803 368
rect 5510 197 5544 213
rect 5607 291 5641 307
rect 5607 223 5641 257
rect 5299 153 5333 169
rect 5139 119 5202 153
rect 5236 119 5299 153
rect 5105 103 5139 119
rect 5299 103 5333 119
rect 5413 153 5447 189
rect 5607 153 5641 189
rect 5447 119 5510 153
rect 5544 119 5607 153
rect 5413 103 5447 119
rect 5607 103 5641 119
rect 5741 296 5755 330
rect 5789 296 5803 330
rect 5741 258 5803 296
rect 5741 224 5755 258
rect 5789 224 5803 258
rect 5741 186 5803 224
rect 5741 152 5755 186
rect 5789 152 5803 186
rect 5741 114 5803 152
rect 5741 80 5755 114
rect 5789 80 5803 114
rect 5741 62 5803 80
rect -31 47 5803 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 343 47
rect 377 13 415 47
rect 449 13 513 47
rect 547 13 585 47
rect 619 13 657 47
rect 691 13 729 47
rect 763 13 801 47
rect 835 13 873 47
rect 907 13 1017 47
rect 1051 13 1089 47
rect 1123 13 1161 47
rect 1195 13 1233 47
rect 1267 13 1305 47
rect 1339 13 1377 47
rect 1411 13 1475 47
rect 1509 13 1547 47
rect 1581 13 1619 47
rect 1653 13 1691 47
rect 1725 13 1763 47
rect 1797 13 1835 47
rect 1869 13 1979 47
rect 2013 13 2051 47
rect 2085 13 2123 47
rect 2157 13 2195 47
rect 2229 13 2267 47
rect 2301 13 2339 47
rect 2373 13 2437 47
rect 2471 13 2509 47
rect 2543 13 2581 47
rect 2615 13 2653 47
rect 2687 13 2725 47
rect 2759 13 2797 47
rect 2831 13 2941 47
rect 2975 13 3013 47
rect 3047 13 3085 47
rect 3119 13 3157 47
rect 3191 13 3229 47
rect 3263 13 3301 47
rect 3335 13 3399 47
rect 3433 13 3471 47
rect 3505 13 3543 47
rect 3577 13 3615 47
rect 3649 13 3687 47
rect 3721 13 3759 47
rect 3793 13 3903 47
rect 3937 13 3975 47
rect 4009 13 4047 47
rect 4081 13 4119 47
rect 4153 13 4191 47
rect 4225 13 4263 47
rect 4297 13 4361 47
rect 4395 13 4433 47
rect 4467 13 4505 47
rect 4539 13 4577 47
rect 4611 13 4649 47
rect 4683 13 4721 47
rect 4755 13 4865 47
rect 4899 13 4937 47
rect 4971 13 5009 47
rect 5043 13 5081 47
rect 5115 13 5153 47
rect 5187 13 5225 47
rect 5259 13 5323 47
rect 5357 13 5395 47
rect 5429 13 5467 47
rect 5501 13 5539 47
rect 5573 13 5611 47
rect 5645 13 5683 47
rect 5717 13 5803 47
rect -31 0 5803 13
<< viali >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 343 1505 377 1539
rect 415 1505 449 1539
rect 513 1505 547 1539
rect 585 1505 619 1539
rect 657 1505 691 1539
rect 729 1505 763 1539
rect 801 1505 835 1539
rect 873 1505 907 1539
rect 1017 1505 1051 1539
rect 1089 1505 1123 1539
rect 1161 1505 1195 1539
rect 1233 1505 1267 1539
rect 1305 1505 1339 1539
rect 1377 1505 1411 1539
rect 1475 1505 1509 1539
rect 1547 1505 1581 1539
rect 1619 1505 1653 1539
rect 1691 1505 1725 1539
rect 1763 1505 1797 1539
rect 1835 1505 1869 1539
rect 1979 1505 2013 1539
rect 2051 1505 2085 1539
rect 2123 1505 2157 1539
rect 2195 1505 2229 1539
rect 2267 1505 2301 1539
rect 2339 1505 2373 1539
rect 2437 1505 2471 1539
rect 2509 1505 2543 1539
rect 2581 1505 2615 1539
rect 2653 1505 2687 1539
rect 2725 1505 2759 1539
rect 2797 1505 2831 1539
rect 2941 1505 2975 1539
rect 3013 1505 3047 1539
rect 3085 1505 3119 1539
rect 3157 1505 3191 1539
rect 3229 1505 3263 1539
rect 3301 1505 3335 1539
rect 3399 1505 3433 1539
rect 3471 1505 3505 1539
rect 3543 1505 3577 1539
rect 3615 1505 3649 1539
rect 3687 1505 3721 1539
rect 3759 1505 3793 1539
rect 3903 1505 3937 1539
rect 3975 1505 4009 1539
rect 4047 1505 4081 1539
rect 4119 1505 4153 1539
rect 4191 1505 4225 1539
rect 4263 1505 4297 1539
rect 4361 1505 4395 1539
rect 4433 1505 4467 1539
rect 4505 1505 4539 1539
rect 4577 1505 4611 1539
rect 4649 1505 4683 1539
rect 4721 1505 4755 1539
rect 4865 1505 4899 1539
rect 4937 1505 4971 1539
rect 5009 1505 5043 1539
rect 5081 1505 5115 1539
rect 5153 1505 5187 1539
rect 5225 1505 5259 1539
rect 5323 1505 5357 1539
rect 5395 1505 5429 1539
rect 5467 1505 5501 1539
rect 5539 1505 5573 1539
rect 5611 1505 5645 1539
rect 5683 1505 5717 1539
rect 205 575 239 609
rect 427 871 461 905
rect 649 723 683 757
rect 797 576 831 610
rect 1167 576 1201 610
rect 1610 797 1644 831
rect 1389 649 1423 683
rect 1759 723 1793 757
rect 2129 576 2163 610
rect 2351 502 2385 536
rect 2573 797 2607 831
rect 2721 575 2755 609
rect 3091 575 3125 609
rect 3313 649 3347 683
rect 3535 871 3569 905
rect 3683 797 3717 831
rect 4053 723 4087 757
rect 4275 871 4309 905
rect 4497 723 4531 757
rect 4645 649 4679 683
rect 5015 649 5049 683
rect 5237 501 5271 535
rect 5459 797 5493 831
rect 5607 723 5641 757
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 343 13 377 47
rect 415 13 449 47
rect 513 13 547 47
rect 585 13 619 47
rect 657 13 691 47
rect 729 13 763 47
rect 801 13 835 47
rect 873 13 907 47
rect 1017 13 1051 47
rect 1089 13 1123 47
rect 1161 13 1195 47
rect 1233 13 1267 47
rect 1305 13 1339 47
rect 1377 13 1411 47
rect 1475 13 1509 47
rect 1547 13 1581 47
rect 1619 13 1653 47
rect 1691 13 1725 47
rect 1763 13 1797 47
rect 1835 13 1869 47
rect 1979 13 2013 47
rect 2051 13 2085 47
rect 2123 13 2157 47
rect 2195 13 2229 47
rect 2267 13 2301 47
rect 2339 13 2373 47
rect 2437 13 2471 47
rect 2509 13 2543 47
rect 2581 13 2615 47
rect 2653 13 2687 47
rect 2725 13 2759 47
rect 2797 13 2831 47
rect 2941 13 2975 47
rect 3013 13 3047 47
rect 3085 13 3119 47
rect 3157 13 3191 47
rect 3229 13 3263 47
rect 3301 13 3335 47
rect 3399 13 3433 47
rect 3471 13 3505 47
rect 3543 13 3577 47
rect 3615 13 3649 47
rect 3687 13 3721 47
rect 3759 13 3793 47
rect 3903 13 3937 47
rect 3975 13 4009 47
rect 4047 13 4081 47
rect 4119 13 4153 47
rect 4191 13 4225 47
rect 4263 13 4297 47
rect 4361 13 4395 47
rect 4433 13 4467 47
rect 4505 13 4539 47
rect 4577 13 4611 47
rect 4649 13 4683 47
rect 4721 13 4755 47
rect 4865 13 4899 47
rect 4937 13 4971 47
rect 5009 13 5043 47
rect 5081 13 5115 47
rect 5153 13 5187 47
rect 5225 13 5259 47
rect 5323 13 5357 47
rect 5395 13 5429 47
rect 5467 13 5501 47
rect 5539 13 5573 47
rect 5611 13 5645 47
rect 5683 13 5717 47
<< metal1 >>
rect -31 1539 5803 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 343 1539
rect 377 1505 415 1539
rect 449 1505 513 1539
rect 547 1505 585 1539
rect 619 1505 657 1539
rect 691 1505 729 1539
rect 763 1505 801 1539
rect 835 1505 873 1539
rect 907 1505 1017 1539
rect 1051 1505 1089 1539
rect 1123 1505 1161 1539
rect 1195 1505 1233 1539
rect 1267 1505 1305 1539
rect 1339 1505 1377 1539
rect 1411 1505 1475 1539
rect 1509 1505 1547 1539
rect 1581 1505 1619 1539
rect 1653 1505 1691 1539
rect 1725 1505 1763 1539
rect 1797 1505 1835 1539
rect 1869 1505 1979 1539
rect 2013 1505 2051 1539
rect 2085 1505 2123 1539
rect 2157 1505 2195 1539
rect 2229 1505 2267 1539
rect 2301 1505 2339 1539
rect 2373 1505 2437 1539
rect 2471 1505 2509 1539
rect 2543 1505 2581 1539
rect 2615 1505 2653 1539
rect 2687 1505 2725 1539
rect 2759 1505 2797 1539
rect 2831 1505 2941 1539
rect 2975 1505 3013 1539
rect 3047 1505 3085 1539
rect 3119 1505 3157 1539
rect 3191 1505 3229 1539
rect 3263 1505 3301 1539
rect 3335 1505 3399 1539
rect 3433 1505 3471 1539
rect 3505 1505 3543 1539
rect 3577 1505 3615 1539
rect 3649 1505 3687 1539
rect 3721 1505 3759 1539
rect 3793 1505 3903 1539
rect 3937 1505 3975 1539
rect 4009 1505 4047 1539
rect 4081 1505 4119 1539
rect 4153 1505 4191 1539
rect 4225 1505 4263 1539
rect 4297 1505 4361 1539
rect 4395 1505 4433 1539
rect 4467 1505 4505 1539
rect 4539 1505 4577 1539
rect 4611 1505 4649 1539
rect 4683 1505 4721 1539
rect 4755 1505 4865 1539
rect 4899 1505 4937 1539
rect 4971 1505 5009 1539
rect 5043 1505 5081 1539
rect 5115 1505 5153 1539
rect 5187 1505 5225 1539
rect 5259 1505 5323 1539
rect 5357 1505 5395 1539
rect 5429 1505 5467 1539
rect 5501 1505 5539 1539
rect 5573 1505 5611 1539
rect 5645 1505 5683 1539
rect 5717 1505 5803 1539
rect -31 1492 5803 1505
rect 421 905 467 911
rect 3529 905 3575 911
rect 4269 905 4315 911
rect 415 871 427 905
rect 461 871 3535 905
rect 3569 871 4275 905
rect 4309 871 4321 905
rect 421 865 467 871
rect 3529 865 3575 871
rect 4269 865 4315 871
rect 1604 831 1650 837
rect 2567 831 2613 837
rect 3677 831 3723 837
rect 5453 831 5499 837
rect 1598 797 1610 831
rect 1644 797 2573 831
rect 2607 797 3683 831
rect 3717 797 5459 831
rect 5493 797 5505 831
rect 1604 791 1650 797
rect 2567 791 2613 797
rect 3677 791 3723 797
rect 5453 791 5499 797
rect 643 757 689 763
rect 1753 757 1799 763
rect 4047 757 4093 763
rect 4491 757 4537 763
rect 5601 757 5647 763
rect 637 723 649 757
rect 683 723 1759 757
rect 1793 723 4053 757
rect 4087 723 4099 757
rect 4485 723 4497 757
rect 4531 723 5607 757
rect 5641 723 5653 757
rect 643 717 689 723
rect 1753 717 1799 723
rect 4047 717 4093 723
rect 4491 717 4537 723
rect 5601 717 5647 723
rect 1383 683 1429 689
rect 3307 683 3353 689
rect 4639 683 4685 689
rect 5009 683 5055 689
rect 1377 649 1389 683
rect 1423 649 3313 683
rect 3347 649 3359 683
rect 4633 649 4645 683
rect 4679 649 5015 683
rect 5049 649 5061 683
rect 1383 643 1429 649
rect 3307 643 3353 649
rect 4639 643 4685 649
rect 5009 643 5055 649
rect 199 609 245 615
rect 791 610 837 616
rect 1161 610 1207 616
rect 2123 610 2169 616
rect 169 575 205 609
rect 239 575 251 609
rect 785 576 797 610
rect 831 576 1167 610
rect 1201 576 2129 610
rect 2163 576 2175 610
rect 2715 609 2761 615
rect 3085 609 3131 615
rect 199 569 245 575
rect 791 570 837 576
rect 1161 570 1207 576
rect 2123 570 2169 576
rect 2709 575 2721 609
rect 2755 575 3091 609
rect 3125 575 3137 609
rect 2715 569 2761 575
rect 3085 569 3131 575
rect 2345 536 2391 542
rect 2339 502 2351 536
rect 2385 535 2421 536
rect 5231 535 5277 541
rect 2385 502 5237 535
rect 2345 501 5237 502
rect 5271 501 5283 535
rect 2345 496 2391 501
rect 5231 495 5277 501
rect -31 47 5803 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 343 47
rect 377 13 415 47
rect 449 13 513 47
rect 547 13 585 47
rect 619 13 657 47
rect 691 13 729 47
rect 763 13 801 47
rect 835 13 873 47
rect 907 13 1017 47
rect 1051 13 1089 47
rect 1123 13 1161 47
rect 1195 13 1233 47
rect 1267 13 1305 47
rect 1339 13 1377 47
rect 1411 13 1475 47
rect 1509 13 1547 47
rect 1581 13 1619 47
rect 1653 13 1691 47
rect 1725 13 1763 47
rect 1797 13 1835 47
rect 1869 13 1979 47
rect 2013 13 2051 47
rect 2085 13 2123 47
rect 2157 13 2195 47
rect 2229 13 2267 47
rect 2301 13 2339 47
rect 2373 13 2437 47
rect 2471 13 2509 47
rect 2543 13 2581 47
rect 2615 13 2653 47
rect 2687 13 2725 47
rect 2759 13 2797 47
rect 2831 13 2941 47
rect 2975 13 3013 47
rect 3047 13 3085 47
rect 3119 13 3157 47
rect 3191 13 3229 47
rect 3263 13 3301 47
rect 3335 13 3399 47
rect 3433 13 3471 47
rect 3505 13 3543 47
rect 3577 13 3615 47
rect 3649 13 3687 47
rect 3721 13 3759 47
rect 3793 13 3903 47
rect 3937 13 3975 47
rect 4009 13 4047 47
rect 4081 13 4119 47
rect 4153 13 4191 47
rect 4225 13 4263 47
rect 4297 13 4361 47
rect 4395 13 4433 47
rect 4467 13 4505 47
rect 4539 13 4577 47
rect 4611 13 4649 47
rect 4683 13 4721 47
rect 4755 13 4865 47
rect 4899 13 4937 47
rect 4971 13 5009 47
rect 5043 13 5081 47
rect 5115 13 5153 47
rect 5187 13 5225 47
rect 5259 13 5323 47
rect 5357 13 5395 47
rect 5429 13 5467 47
rect 5501 13 5539 47
rect 5573 13 5611 47
rect 5645 13 5683 47
rect 5717 13 5803 47
rect -31 0 5803 13
<< labels >>
rlabel metal1 5607 723 5641 757 1 Q
port 1 n
rlabel metal1 4645 649 4679 683 1 QN
port 2 n
rlabel metal1 205 575 239 609 1 D
port 3 n
rlabel metal1 1389 649 1423 683 1 CLK
port 4 n
rlabel metal1 2351 502 2385 536 1 SN
port 5 n
rlabel metal1 427 871 461 905 1 RN
port 6 n
rlabel metal1 55 1505 89 1539 1 VDD
port 7 n
rlabel metal1 55 13 89 47 1 VSS
port 8 n
<< end >>
