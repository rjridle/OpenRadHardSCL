magic
tech sky130A
magscale 1 2
timestamp 1648742928
<< metal1 >>
rect 55 1505 89 1539
rect 427 945 461 979
rect 3349 797 4115 831
rect 4127 797 4161 831
rect 3497 723 3807 757
rect 3831 723 3865 757
rect 1315 649 1349 683
rect 55 13 89 47
use li1_M1_contact  li1_M1_contact_4 pcells
timestamp 1648061256
transform 1 0 1332 0 1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_8
timestamp 1648061256
transform -1 0 3330 0 -1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform 1 0 3848 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform -1 0 3478 0 -1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_15
timestamp 1648061256
transform 1 0 4144 0 1 814
box -53 -33 29 33
use dffx1_pcell  dffx1_pcell_0 pcells
timestamp 1648742316
transform 1 0 0 0 1 0
box -84 0 4376 1575
<< labels >>
rlabel metal1 4127 797 4161 831 1 Q
port 1 n
rlabel metal1 3831 723 3865 757 1 QN
port 2 n
rlabel metal1 1315 649 1349 683 1 D
port 3 n
rlabel metal1 427 945 461 979 1 CLK
port 4 n
rlabel metal1 55 1505 89 1539 1 VDD
port 5 n
rlabel metal1 55 13 89 47 1 VSS
port 6 n
<< end >>
