magic
tech sky130A
magscale 1 2
timestamp 1648506367
<< nwell >>
rect -84 832 18066 1575
<< nmos >>
rect 147 318 177 379
tri 177 318 193 334 sw
rect 447 318 477 379
rect 147 288 253 318
tri 253 288 283 318 sw
rect 147 187 177 288
tri 177 272 193 288 nw
tri 237 272 253 288 ne
tri 177 187 193 203 sw
tri 237 187 253 203 se
rect 253 187 283 288
tri 342 288 372 318 se
rect 372 288 477 318
rect 342 194 372 288
tri 372 272 388 288 nw
tri 431 272 447 288 ne
tri 372 194 388 210 sw
tri 431 194 447 210 se
rect 447 194 477 288
tri 147 157 177 187 ne
rect 177 157 253 187
tri 253 157 283 187 nw
tri 342 164 372 194 ne
rect 372 164 447 194
tri 447 164 477 194 nw
rect 649 326 679 379
tri 679 326 695 342 sw
rect 649 296 755 326
tri 755 296 785 326 sw
rect 649 195 679 296
tri 679 280 695 296 nw
tri 739 280 755 296 ne
tri 679 195 695 211 sw
tri 739 195 755 211 se
rect 755 195 785 296
tri 649 165 679 195 ne
rect 679 165 755 195
tri 755 165 785 195 nw
rect 1109 318 1139 379
tri 1139 318 1155 334 sw
rect 1409 318 1439 379
rect 1109 288 1215 318
tri 1215 288 1245 318 sw
rect 1109 187 1139 288
tri 1139 272 1155 288 nw
tri 1199 272 1215 288 ne
tri 1139 187 1155 203 sw
tri 1199 187 1215 203 se
rect 1215 187 1245 288
tri 1304 288 1334 318 se
rect 1334 288 1439 318
rect 1304 194 1334 288
tri 1334 272 1350 288 nw
tri 1393 272 1409 288 ne
tri 1334 194 1350 210 sw
tri 1393 194 1409 210 se
rect 1409 194 1439 288
tri 1109 157 1139 187 ne
rect 1139 157 1215 187
tri 1215 157 1245 187 nw
tri 1304 164 1334 194 ne
rect 1334 164 1409 194
tri 1409 164 1439 194 nw
rect 1611 326 1641 379
tri 1641 326 1657 342 sw
rect 1611 296 1717 326
tri 1717 296 1747 326 sw
rect 1611 195 1641 296
tri 1641 280 1657 296 nw
tri 1701 280 1717 296 ne
tri 1641 195 1657 211 sw
tri 1701 195 1717 211 se
rect 1717 195 1747 296
tri 1611 165 1641 195 ne
rect 1641 165 1717 195
tri 1717 165 1747 195 nw
rect 2092 316 2122 377
tri 2122 316 2138 332 sw
rect 2286 324 2316 377
tri 2316 324 2332 340 sw
rect 2092 286 2198 316
tri 2198 286 2228 316 sw
rect 2286 294 2392 324
tri 2392 294 2422 324 sw
rect 2092 185 2122 286
tri 2122 270 2138 286 nw
tri 2182 270 2198 286 ne
tri 2122 185 2138 201 sw
tri 2182 185 2198 201 se
rect 2198 185 2228 286
rect 2286 193 2316 294
tri 2316 278 2332 294 nw
tri 2376 278 2392 294 ne
tri 2316 193 2332 209 sw
tri 2376 193 2392 209 se
rect 2392 193 2422 294
tri 2092 155 2122 185 ne
rect 2122 155 2198 185
tri 2198 155 2228 185 nw
tri 2286 163 2316 193 ne
rect 2316 163 2392 193
tri 2392 163 2422 193 nw
rect 2737 318 2767 379
tri 2767 318 2783 334 sw
rect 3037 318 3067 379
rect 2737 288 2843 318
tri 2843 288 2873 318 sw
rect 2737 187 2767 288
tri 2767 272 2783 288 nw
tri 2827 272 2843 288 ne
tri 2767 187 2783 203 sw
tri 2827 187 2843 203 se
rect 2843 187 2873 288
tri 2932 288 2962 318 se
rect 2962 288 3067 318
rect 2932 194 2962 288
tri 2962 272 2978 288 nw
tri 3021 272 3037 288 ne
tri 2962 194 2978 210 sw
tri 3021 194 3037 210 se
rect 3037 194 3067 288
tri 2737 157 2767 187 ne
rect 2767 157 2843 187
tri 2843 157 2873 187 nw
tri 2932 164 2962 194 ne
rect 2962 164 3037 194
tri 3037 164 3067 194 nw
rect 3239 326 3269 379
tri 3269 326 3285 342 sw
rect 3239 296 3345 326
tri 3345 296 3375 326 sw
rect 3239 195 3269 296
tri 3269 280 3285 296 nw
tri 3329 280 3345 296 ne
tri 3269 195 3285 211 sw
tri 3329 195 3345 211 se
rect 3345 195 3375 296
tri 3239 165 3269 195 ne
rect 3269 165 3345 195
tri 3345 165 3375 195 nw
rect 3699 318 3729 379
tri 3729 318 3745 334 sw
rect 3999 318 4029 379
rect 3699 288 3805 318
tri 3805 288 3835 318 sw
rect 3699 187 3729 288
tri 3729 272 3745 288 nw
tri 3789 272 3805 288 ne
tri 3729 187 3745 203 sw
tri 3789 187 3805 203 se
rect 3805 187 3835 288
tri 3894 288 3924 318 se
rect 3924 288 4029 318
rect 3894 194 3924 288
tri 3924 272 3940 288 nw
tri 3983 272 3999 288 ne
tri 3924 194 3940 210 sw
tri 3983 194 3999 210 se
rect 3999 194 4029 288
tri 3699 157 3729 187 ne
rect 3729 157 3805 187
tri 3805 157 3835 187 nw
tri 3894 164 3924 194 ne
rect 3924 164 3999 194
tri 3999 164 4029 194 nw
rect 4201 326 4231 379
tri 4231 326 4247 342 sw
rect 4201 296 4307 326
tri 4307 296 4337 326 sw
rect 4201 195 4231 296
tri 4231 280 4247 296 nw
tri 4291 280 4307 296 ne
tri 4231 195 4247 211 sw
tri 4291 195 4307 211 se
rect 4307 195 4337 296
tri 4201 165 4231 195 ne
rect 4231 165 4307 195
tri 4307 165 4337 195 nw
rect 4682 316 4712 377
tri 4712 316 4728 332 sw
rect 4876 324 4906 377
tri 4906 324 4922 340 sw
rect 4682 286 4788 316
tri 4788 286 4818 316 sw
rect 4876 294 4982 324
tri 4982 294 5012 324 sw
rect 4682 185 4712 286
tri 4712 270 4728 286 nw
tri 4772 270 4788 286 ne
tri 4712 185 4728 201 sw
tri 4772 185 4788 201 se
rect 4788 185 4818 286
rect 4876 193 4906 294
tri 4906 278 4922 294 nw
tri 4966 278 4982 294 ne
tri 4906 193 4922 209 sw
tri 4966 193 4982 209 se
rect 4982 193 5012 294
tri 4682 155 4712 185 ne
rect 4712 155 4788 185
tri 4788 155 4818 185 nw
tri 4876 163 4906 193 ne
rect 4906 163 4982 193
tri 4982 163 5012 193 nw
rect 5327 318 5357 379
tri 5357 318 5373 334 sw
rect 5627 318 5657 379
rect 5327 288 5433 318
tri 5433 288 5463 318 sw
rect 5327 187 5357 288
tri 5357 272 5373 288 nw
tri 5417 272 5433 288 ne
tri 5357 187 5373 203 sw
tri 5417 187 5433 203 se
rect 5433 187 5463 288
tri 5522 288 5552 318 se
rect 5552 288 5657 318
rect 5522 194 5552 288
tri 5552 272 5568 288 nw
tri 5611 272 5627 288 ne
tri 5552 194 5568 210 sw
tri 5611 194 5627 210 se
rect 5627 194 5657 288
tri 5327 157 5357 187 ne
rect 5357 157 5433 187
tri 5433 157 5463 187 nw
tri 5522 164 5552 194 ne
rect 5552 164 5627 194
tri 5627 164 5657 194 nw
rect 5829 326 5859 379
tri 5859 326 5875 342 sw
rect 5829 296 5935 326
tri 5935 296 5965 326 sw
rect 5829 195 5859 296
tri 5859 280 5875 296 nw
tri 5919 280 5935 296 ne
tri 5859 195 5875 211 sw
tri 5919 195 5935 211 se
rect 5935 195 5965 296
tri 5829 165 5859 195 ne
rect 5859 165 5935 195
tri 5935 165 5965 195 nw
rect 6289 318 6319 379
tri 6319 318 6335 334 sw
rect 6589 318 6619 379
rect 6289 288 6395 318
tri 6395 288 6425 318 sw
rect 6289 187 6319 288
tri 6319 272 6335 288 nw
tri 6379 272 6395 288 ne
tri 6319 187 6335 203 sw
tri 6379 187 6395 203 se
rect 6395 187 6425 288
tri 6484 288 6514 318 se
rect 6514 288 6619 318
rect 6484 194 6514 288
tri 6514 272 6530 288 nw
tri 6573 272 6589 288 ne
tri 6514 194 6530 210 sw
tri 6573 194 6589 210 se
rect 6589 194 6619 288
tri 6289 157 6319 187 ne
rect 6319 157 6395 187
tri 6395 157 6425 187 nw
tri 6484 164 6514 194 ne
rect 6514 164 6589 194
tri 6589 164 6619 194 nw
rect 6791 326 6821 379
tri 6821 326 6837 342 sw
rect 6791 296 6897 326
tri 6897 296 6927 326 sw
rect 6791 195 6821 296
tri 6821 280 6837 296 nw
tri 6881 280 6897 296 ne
tri 6821 195 6837 211 sw
tri 6881 195 6897 211 se
rect 6897 195 6927 296
tri 6791 165 6821 195 ne
rect 6821 165 6897 195
tri 6897 165 6927 195 nw
rect 7272 316 7302 377
tri 7302 316 7318 332 sw
rect 7466 324 7496 377
tri 7496 324 7512 340 sw
rect 7272 286 7378 316
tri 7378 286 7408 316 sw
rect 7466 294 7572 324
tri 7572 294 7602 324 sw
rect 7272 185 7302 286
tri 7302 270 7318 286 nw
tri 7362 270 7378 286 ne
tri 7302 185 7318 201 sw
tri 7362 185 7378 201 se
rect 7378 185 7408 286
rect 7466 193 7496 294
tri 7496 278 7512 294 nw
tri 7556 278 7572 294 ne
tri 7496 193 7512 209 sw
tri 7556 193 7572 209 se
rect 7572 193 7602 294
tri 7272 155 7302 185 ne
rect 7302 155 7378 185
tri 7378 155 7408 185 nw
tri 7466 163 7496 193 ne
rect 7496 163 7572 193
tri 7572 163 7602 193 nw
rect 7917 318 7947 379
tri 7947 318 7963 334 sw
rect 8217 318 8247 379
rect 7917 288 8023 318
tri 8023 288 8053 318 sw
rect 7917 187 7947 288
tri 7947 272 7963 288 nw
tri 8007 272 8023 288 ne
tri 7947 187 7963 203 sw
tri 8007 187 8023 203 se
rect 8023 187 8053 288
tri 8112 288 8142 318 se
rect 8142 288 8247 318
rect 8112 194 8142 288
tri 8142 272 8158 288 nw
tri 8201 272 8217 288 ne
tri 8142 194 8158 210 sw
tri 8201 194 8217 210 se
rect 8217 194 8247 288
tri 7917 157 7947 187 ne
rect 7947 157 8023 187
tri 8023 157 8053 187 nw
tri 8112 164 8142 194 ne
rect 8142 164 8217 194
tri 8217 164 8247 194 nw
rect 8419 326 8449 379
tri 8449 326 8465 342 sw
rect 8419 296 8525 326
tri 8525 296 8555 326 sw
rect 8419 195 8449 296
tri 8449 280 8465 296 nw
tri 8509 280 8525 296 ne
tri 8449 195 8465 211 sw
tri 8509 195 8525 211 se
rect 8525 195 8555 296
tri 8419 165 8449 195 ne
rect 8449 165 8525 195
tri 8525 165 8555 195 nw
rect 8879 318 8909 379
tri 8909 318 8925 334 sw
rect 9179 318 9209 379
rect 8879 288 8985 318
tri 8985 288 9015 318 sw
rect 8879 187 8909 288
tri 8909 272 8925 288 nw
tri 8969 272 8985 288 ne
tri 8909 187 8925 203 sw
tri 8969 187 8985 203 se
rect 8985 187 9015 288
tri 9074 288 9104 318 se
rect 9104 288 9209 318
rect 9074 194 9104 288
tri 9104 272 9120 288 nw
tri 9163 272 9179 288 ne
tri 9104 194 9120 210 sw
tri 9163 194 9179 210 se
rect 9179 194 9209 288
tri 8879 157 8909 187 ne
rect 8909 157 8985 187
tri 8985 157 9015 187 nw
tri 9074 164 9104 194 ne
rect 9104 164 9179 194
tri 9179 164 9209 194 nw
rect 9381 326 9411 379
tri 9411 326 9427 342 sw
rect 9381 296 9487 326
tri 9487 296 9517 326 sw
rect 9381 195 9411 296
tri 9411 280 9427 296 nw
tri 9471 280 9487 296 ne
tri 9411 195 9427 211 sw
tri 9471 195 9487 211 se
rect 9487 195 9517 296
tri 9381 165 9411 195 ne
rect 9411 165 9487 195
tri 9487 165 9517 195 nw
rect 9862 316 9892 377
tri 9892 316 9908 332 sw
rect 10056 324 10086 377
tri 10086 324 10102 340 sw
rect 9862 286 9968 316
tri 9968 286 9998 316 sw
rect 10056 294 10162 324
tri 10162 294 10192 324 sw
rect 9862 185 9892 286
tri 9892 270 9908 286 nw
tri 9952 270 9968 286 ne
tri 9892 185 9908 201 sw
tri 9952 185 9968 201 se
rect 9968 185 9998 286
rect 10056 193 10086 294
tri 10086 278 10102 294 nw
tri 10146 278 10162 294 ne
tri 10086 193 10102 209 sw
tri 10146 193 10162 209 se
rect 10162 193 10192 294
tri 9862 155 9892 185 ne
rect 9892 155 9968 185
tri 9968 155 9998 185 nw
tri 10056 163 10086 193 ne
rect 10086 163 10162 193
tri 10162 163 10192 193 nw
rect 10507 318 10537 379
tri 10537 318 10553 334 sw
rect 10807 318 10837 379
rect 10507 288 10613 318
tri 10613 288 10643 318 sw
rect 10507 187 10537 288
tri 10537 272 10553 288 nw
tri 10597 272 10613 288 ne
tri 10537 187 10553 203 sw
tri 10597 187 10613 203 se
rect 10613 187 10643 288
tri 10702 288 10732 318 se
rect 10732 288 10837 318
rect 10702 194 10732 288
tri 10732 272 10748 288 nw
tri 10791 272 10807 288 ne
tri 10732 194 10748 210 sw
tri 10791 194 10807 210 se
rect 10807 194 10837 288
tri 10507 157 10537 187 ne
rect 10537 157 10613 187
tri 10613 157 10643 187 nw
tri 10702 164 10732 194 ne
rect 10732 164 10807 194
tri 10807 164 10837 194 nw
rect 11009 326 11039 379
tri 11039 326 11055 342 sw
rect 11009 296 11115 326
tri 11115 296 11145 326 sw
rect 11009 195 11039 296
tri 11039 280 11055 296 nw
tri 11099 280 11115 296 ne
tri 11039 195 11055 211 sw
tri 11099 195 11115 211 se
rect 11115 195 11145 296
tri 11009 165 11039 195 ne
rect 11039 165 11115 195
tri 11115 165 11145 195 nw
rect 11469 318 11499 379
tri 11499 318 11515 334 sw
rect 11769 318 11799 379
rect 11469 288 11575 318
tri 11575 288 11605 318 sw
rect 11469 187 11499 288
tri 11499 272 11515 288 nw
tri 11559 272 11575 288 ne
tri 11499 187 11515 203 sw
tri 11559 187 11575 203 se
rect 11575 187 11605 288
tri 11664 288 11694 318 se
rect 11694 288 11799 318
rect 11664 194 11694 288
tri 11694 272 11710 288 nw
tri 11753 272 11769 288 ne
tri 11694 194 11710 210 sw
tri 11753 194 11769 210 se
rect 11769 194 11799 288
tri 11469 157 11499 187 ne
rect 11499 157 11575 187
tri 11575 157 11605 187 nw
tri 11664 164 11694 194 ne
rect 11694 164 11769 194
tri 11769 164 11799 194 nw
rect 11971 326 12001 379
tri 12001 326 12017 342 sw
rect 11971 296 12077 326
tri 12077 296 12107 326 sw
rect 11971 195 12001 296
tri 12001 280 12017 296 nw
tri 12061 280 12077 296 ne
tri 12001 195 12017 211 sw
tri 12061 195 12077 211 se
rect 12077 195 12107 296
tri 11971 165 12001 195 ne
rect 12001 165 12077 195
tri 12077 165 12107 195 nw
rect 12452 316 12482 377
tri 12482 316 12498 332 sw
rect 12646 324 12676 377
tri 12676 324 12692 340 sw
rect 12452 286 12558 316
tri 12558 286 12588 316 sw
rect 12646 294 12752 324
tri 12752 294 12782 324 sw
rect 12452 185 12482 286
tri 12482 270 12498 286 nw
tri 12542 270 12558 286 ne
tri 12482 185 12498 201 sw
tri 12542 185 12558 201 se
rect 12558 185 12588 286
rect 12646 193 12676 294
tri 12676 278 12692 294 nw
tri 12736 278 12752 294 ne
tri 12676 193 12692 209 sw
tri 12736 193 12752 209 se
rect 12752 193 12782 294
tri 12452 155 12482 185 ne
rect 12482 155 12558 185
tri 12558 155 12588 185 nw
tri 12646 163 12676 193 ne
rect 12676 163 12752 193
tri 12752 163 12782 193 nw
rect 13097 318 13127 379
tri 13127 318 13143 334 sw
rect 13397 318 13427 379
rect 13097 288 13203 318
tri 13203 288 13233 318 sw
rect 13097 187 13127 288
tri 13127 272 13143 288 nw
tri 13187 272 13203 288 ne
tri 13127 187 13143 203 sw
tri 13187 187 13203 203 se
rect 13203 187 13233 288
tri 13292 288 13322 318 se
rect 13322 288 13427 318
rect 13292 194 13322 288
tri 13322 272 13338 288 nw
tri 13381 272 13397 288 ne
tri 13322 194 13338 210 sw
tri 13381 194 13397 210 se
rect 13397 194 13427 288
tri 13097 157 13127 187 ne
rect 13127 157 13203 187
tri 13203 157 13233 187 nw
tri 13292 164 13322 194 ne
rect 13322 164 13397 194
tri 13397 164 13427 194 nw
rect 13599 326 13629 379
tri 13629 326 13645 342 sw
rect 13599 296 13705 326
tri 13705 296 13735 326 sw
rect 13599 195 13629 296
tri 13629 280 13645 296 nw
tri 13689 280 13705 296 ne
tri 13629 195 13645 211 sw
tri 13689 195 13705 211 se
rect 13705 195 13735 296
tri 13599 165 13629 195 ne
rect 13629 165 13705 195
tri 13705 165 13735 195 nw
rect 14059 318 14089 379
tri 14089 318 14105 334 sw
rect 14359 318 14389 379
rect 14059 288 14165 318
tri 14165 288 14195 318 sw
rect 14059 187 14089 288
tri 14089 272 14105 288 nw
tri 14149 272 14165 288 ne
tri 14089 187 14105 203 sw
tri 14149 187 14165 203 se
rect 14165 187 14195 288
tri 14254 288 14284 318 se
rect 14284 288 14389 318
rect 14254 194 14284 288
tri 14284 272 14300 288 nw
tri 14343 272 14359 288 ne
tri 14284 194 14300 210 sw
tri 14343 194 14359 210 se
rect 14359 194 14389 288
tri 14059 157 14089 187 ne
rect 14089 157 14165 187
tri 14165 157 14195 187 nw
tri 14254 164 14284 194 ne
rect 14284 164 14359 194
tri 14359 164 14389 194 nw
rect 14561 326 14591 379
tri 14591 326 14607 342 sw
rect 14561 296 14667 326
tri 14667 296 14697 326 sw
rect 14561 195 14591 296
tri 14591 280 14607 296 nw
tri 14651 280 14667 296 ne
tri 14591 195 14607 211 sw
tri 14651 195 14667 211 se
rect 14667 195 14697 296
tri 14561 165 14591 195 ne
rect 14591 165 14667 195
tri 14667 165 14697 195 nw
rect 15042 316 15072 377
tri 15072 316 15088 332 sw
rect 15236 324 15266 377
tri 15266 324 15282 340 sw
rect 15042 286 15148 316
tri 15148 286 15178 316 sw
rect 15236 294 15342 324
tri 15342 294 15372 324 sw
rect 15042 185 15072 286
tri 15072 270 15088 286 nw
tri 15132 270 15148 286 ne
tri 15072 185 15088 201 sw
tri 15132 185 15148 201 se
rect 15148 185 15178 286
rect 15236 193 15266 294
tri 15266 278 15282 294 nw
tri 15326 278 15342 294 ne
tri 15266 193 15282 209 sw
tri 15326 193 15342 209 se
rect 15342 193 15372 294
tri 15042 155 15072 185 ne
rect 15072 155 15148 185
tri 15148 155 15178 185 nw
tri 15236 163 15266 193 ne
rect 15266 163 15342 193
tri 15342 163 15372 193 nw
rect 15708 316 15738 377
tri 15738 316 15754 332 sw
rect 15902 324 15932 377
tri 15932 324 15948 340 sw
rect 15708 286 15814 316
tri 15814 286 15844 316 sw
rect 15902 294 16008 324
tri 16008 294 16038 324 sw
rect 15708 185 15738 286
tri 15738 270 15754 286 nw
tri 15798 270 15814 286 ne
tri 15738 185 15754 201 sw
tri 15798 185 15814 201 se
rect 15814 185 15844 286
rect 15902 193 15932 294
tri 15932 278 15948 294 nw
tri 15992 278 16008 294 ne
tri 15932 193 15948 209 sw
tri 15992 193 16008 209 se
rect 16008 193 16038 294
tri 15708 155 15738 185 ne
rect 15738 155 15814 185
tri 15814 155 15844 185 nw
tri 15902 163 15932 193 ne
rect 15932 163 16008 193
tri 16008 163 16038 193 nw
rect 16374 316 16404 377
tri 16404 316 16420 332 sw
tri 16658 324 16674 340 se
rect 16674 324 16704 377
rect 16374 286 16480 316
tri 16480 286 16510 316 sw
tri 16568 294 16598 324 se
rect 16598 294 16704 324
rect 16374 185 16404 286
tri 16404 270 16420 286 nw
tri 16464 270 16480 286 ne
tri 16404 185 16420 201 sw
tri 16464 185 16480 201 se
rect 16480 185 16510 286
rect 16568 193 16598 294
tri 16598 278 16614 294 nw
tri 16658 278 16674 294 ne
tri 16598 193 16614 209 sw
tri 16658 193 16674 209 se
rect 16674 193 16704 294
tri 16374 155 16404 185 ne
rect 16404 155 16480 185
tri 16480 155 16510 185 nw
tri 16568 163 16598 193 ne
rect 16598 163 16674 193
tri 16674 163 16704 193 nw
rect 17040 316 17070 377
tri 17070 316 17086 332 sw
rect 17234 324 17264 377
tri 17264 324 17280 340 sw
rect 17040 286 17146 316
tri 17146 286 17176 316 sw
rect 17234 294 17340 324
tri 17340 294 17370 324 sw
rect 17040 185 17070 286
tri 17070 270 17086 286 nw
tri 17130 270 17146 286 ne
tri 17070 185 17086 201 sw
tri 17130 185 17146 201 se
rect 17146 185 17176 286
rect 17234 279 17265 294
tri 17265 279 17280 294 nw
tri 17324 279 17339 294 ne
rect 17339 279 17370 294
rect 17234 193 17264 279
tri 17264 193 17280 209 sw
tri 17324 193 17340 209 se
rect 17340 193 17370 279
tri 17040 155 17070 185 ne
rect 17070 155 17146 185
tri 17146 155 17176 185 nw
tri 17234 163 17264 193 ne
rect 17264 163 17340 193
tri 17340 163 17370 193 nw
rect 17693 324 17723 377
tri 17723 324 17739 340 sw
rect 17693 294 17799 324
tri 17799 294 17829 324 sw
rect 17693 193 17723 294
tri 17723 278 17739 294 nw
tri 17783 278 17799 294 ne
tri 17723 193 17739 209 sw
tri 17783 193 17799 209 se
rect 17799 193 17829 294
tri 17693 163 17723 193 ne
rect 17723 163 17799 193
tri 17799 163 17829 193 nw
<< pmos >>
rect 247 1050 277 1450
rect 335 1050 365 1450
rect 423 1050 453 1450
rect 511 1050 541 1450
rect 599 1050 629 1450
rect 687 1050 717 1450
rect 1209 1050 1239 1450
rect 1297 1050 1327 1450
rect 1385 1050 1415 1450
rect 1473 1050 1503 1450
rect 1561 1050 1591 1450
rect 1649 1050 1679 1450
rect 2111 1050 2141 1450
rect 2199 1050 2229 1450
rect 2287 1050 2317 1450
rect 2375 1050 2405 1450
rect 2837 1050 2867 1450
rect 2925 1050 2955 1450
rect 3013 1050 3043 1450
rect 3101 1050 3131 1450
rect 3189 1050 3219 1450
rect 3277 1050 3307 1450
rect 3799 1050 3829 1450
rect 3887 1050 3917 1450
rect 3975 1050 4005 1450
rect 4063 1050 4093 1450
rect 4151 1050 4181 1450
rect 4239 1050 4269 1450
rect 4701 1050 4731 1450
rect 4789 1050 4819 1450
rect 4877 1050 4907 1450
rect 4965 1050 4995 1450
rect 5427 1050 5457 1450
rect 5515 1050 5545 1450
rect 5603 1050 5633 1450
rect 5691 1050 5721 1450
rect 5779 1050 5809 1450
rect 5867 1050 5897 1450
rect 6389 1050 6419 1450
rect 6477 1050 6507 1450
rect 6565 1050 6595 1450
rect 6653 1050 6683 1450
rect 6741 1050 6771 1450
rect 6829 1050 6859 1450
rect 7291 1050 7321 1450
rect 7379 1050 7409 1450
rect 7467 1050 7497 1450
rect 7555 1050 7585 1450
rect 8017 1050 8047 1450
rect 8105 1050 8135 1450
rect 8193 1050 8223 1450
rect 8281 1050 8311 1450
rect 8369 1050 8399 1450
rect 8457 1050 8487 1450
rect 8979 1050 9009 1450
rect 9067 1050 9097 1450
rect 9155 1050 9185 1450
rect 9243 1050 9273 1450
rect 9331 1050 9361 1450
rect 9419 1050 9449 1450
rect 9881 1050 9911 1450
rect 9969 1050 9999 1450
rect 10057 1050 10087 1450
rect 10145 1050 10175 1450
rect 10607 1050 10637 1450
rect 10695 1050 10725 1450
rect 10783 1050 10813 1450
rect 10871 1050 10901 1450
rect 10959 1050 10989 1450
rect 11047 1050 11077 1450
rect 11569 1050 11599 1450
rect 11657 1050 11687 1450
rect 11745 1050 11775 1450
rect 11833 1050 11863 1450
rect 11921 1050 11951 1450
rect 12009 1050 12039 1450
rect 12471 1050 12501 1450
rect 12559 1050 12589 1450
rect 12647 1050 12677 1450
rect 12735 1050 12765 1450
rect 13197 1050 13227 1450
rect 13285 1050 13315 1450
rect 13373 1050 13403 1450
rect 13461 1050 13491 1450
rect 13549 1050 13579 1450
rect 13637 1050 13667 1450
rect 14159 1050 14189 1450
rect 14247 1050 14277 1450
rect 14335 1050 14365 1450
rect 14423 1050 14453 1450
rect 14511 1050 14541 1450
rect 14599 1050 14629 1450
rect 15061 1050 15091 1450
rect 15149 1050 15179 1450
rect 15237 1050 15267 1450
rect 15325 1050 15355 1450
rect 15727 1051 15757 1451
rect 15815 1051 15845 1451
rect 15903 1051 15933 1451
rect 15991 1051 16021 1451
rect 16391 1051 16421 1451
rect 16479 1051 16509 1451
rect 16567 1051 16597 1451
rect 16655 1051 16685 1451
rect 17059 1051 17089 1451
rect 17147 1051 17177 1451
rect 17235 1051 17265 1451
rect 17323 1051 17353 1451
rect 17701 1050 17731 1450
rect 17789 1050 17819 1450
<< ndiff >>
rect 91 363 147 379
rect 91 329 101 363
rect 135 329 147 363
rect 91 291 147 329
rect 177 363 447 379
rect 177 334 198 363
tri 177 318 193 334 ne
rect 193 329 198 334
rect 232 329 295 363
rect 329 329 392 363
rect 426 329 447 363
rect 193 318 447 329
rect 477 363 533 379
rect 477 329 489 363
rect 523 329 533 363
rect 91 257 101 291
rect 135 257 147 291
tri 253 288 283 318 ne
rect 283 291 342 318
rect 91 223 147 257
rect 91 189 101 223
rect 135 189 147 223
rect 91 157 147 189
tri 177 272 193 288 se
rect 193 272 237 288
tri 237 272 253 288 sw
rect 177 238 253 272
rect 177 204 198 238
rect 232 204 253 238
rect 177 203 253 204
tri 177 187 193 203 ne
rect 193 187 237 203
tri 237 187 253 203 nw
rect 283 257 295 291
rect 329 257 342 291
tri 342 288 372 318 nw
rect 283 223 342 257
rect 283 189 295 223
rect 329 189 342 223
tri 372 272 388 288 se
rect 388 272 431 288
tri 431 272 447 288 sw
rect 372 244 447 272
rect 372 210 393 244
rect 427 210 447 244
tri 372 194 388 210 ne
rect 388 194 431 210
tri 431 194 447 210 nw
tri 147 157 177 187 sw
tri 253 157 283 187 se
rect 283 164 342 189
tri 342 164 372 194 sw
tri 447 164 477 194 se
rect 477 164 533 329
rect 283 157 533 164
rect 91 153 533 157
rect 91 119 101 153
rect 135 119 295 153
rect 329 119 392 153
rect 426 119 489 153
rect 523 119 533 153
rect 91 103 533 119
rect 593 363 649 379
rect 593 329 603 363
rect 637 329 649 363
rect 593 291 649 329
rect 679 342 841 379
tri 679 326 695 342 ne
rect 695 326 841 342
tri 755 296 785 326 ne
rect 593 257 603 291
rect 637 257 649 291
rect 593 223 649 257
rect 593 189 603 223
rect 637 189 649 223
tri 679 280 695 296 se
rect 695 280 739 296
tri 739 280 755 296 sw
rect 679 247 755 280
rect 679 213 700 247
rect 734 213 755 247
rect 679 211 755 213
tri 679 195 695 211 ne
rect 695 195 739 211
tri 739 195 755 211 nw
rect 785 291 841 326
rect 785 257 797 291
rect 831 257 841 291
rect 785 223 841 257
rect 593 165 649 189
tri 649 165 679 195 sw
tri 755 165 785 195 se
rect 785 189 797 223
rect 831 189 841 223
rect 785 165 841 189
rect 593 153 841 165
rect 593 119 603 153
rect 637 119 700 153
rect 734 119 797 153
rect 831 119 841 153
rect 593 103 841 119
rect 1053 363 1109 379
rect 1053 329 1063 363
rect 1097 329 1109 363
rect 1053 291 1109 329
rect 1139 363 1409 379
rect 1139 334 1160 363
tri 1139 318 1155 334 ne
rect 1155 329 1160 334
rect 1194 329 1257 363
rect 1291 329 1354 363
rect 1388 329 1409 363
rect 1155 318 1409 329
rect 1439 363 1495 379
rect 1439 329 1451 363
rect 1485 329 1495 363
rect 1053 257 1063 291
rect 1097 257 1109 291
tri 1215 288 1245 318 ne
rect 1245 291 1304 318
rect 1053 223 1109 257
rect 1053 189 1063 223
rect 1097 189 1109 223
rect 1053 157 1109 189
tri 1139 272 1155 288 se
rect 1155 272 1199 288
tri 1199 272 1215 288 sw
rect 1139 238 1215 272
rect 1139 204 1160 238
rect 1194 204 1215 238
rect 1139 203 1215 204
tri 1139 187 1155 203 ne
rect 1155 187 1199 203
tri 1199 187 1215 203 nw
rect 1245 257 1257 291
rect 1291 257 1304 291
tri 1304 288 1334 318 nw
rect 1245 223 1304 257
rect 1245 189 1257 223
rect 1291 189 1304 223
tri 1334 272 1350 288 se
rect 1350 272 1393 288
tri 1393 272 1409 288 sw
rect 1334 244 1409 272
rect 1334 210 1355 244
rect 1389 210 1409 244
tri 1334 194 1350 210 ne
rect 1350 194 1393 210
tri 1393 194 1409 210 nw
tri 1109 157 1139 187 sw
tri 1215 157 1245 187 se
rect 1245 164 1304 189
tri 1304 164 1334 194 sw
tri 1409 164 1439 194 se
rect 1439 164 1495 329
rect 1245 157 1495 164
rect 1053 153 1495 157
rect 1053 119 1063 153
rect 1097 119 1257 153
rect 1291 119 1354 153
rect 1388 119 1451 153
rect 1485 119 1495 153
rect 1053 103 1495 119
rect 1555 363 1611 379
rect 1555 329 1565 363
rect 1599 329 1611 363
rect 1555 291 1611 329
rect 1641 342 1803 379
tri 1641 326 1657 342 ne
rect 1657 326 1803 342
tri 1717 296 1747 326 ne
rect 1555 257 1565 291
rect 1599 257 1611 291
rect 1555 223 1611 257
rect 1555 189 1565 223
rect 1599 189 1611 223
tri 1641 280 1657 296 se
rect 1657 280 1701 296
tri 1701 280 1717 296 sw
rect 1641 247 1717 280
rect 1641 213 1662 247
rect 1696 213 1717 247
rect 1641 211 1717 213
tri 1641 195 1657 211 ne
rect 1657 195 1701 211
tri 1701 195 1717 211 nw
rect 1747 291 1803 326
rect 1747 257 1759 291
rect 1793 257 1803 291
rect 1747 223 1803 257
rect 1555 165 1611 189
tri 1611 165 1641 195 sw
tri 1717 165 1747 195 se
rect 1747 189 1759 223
rect 1793 189 1803 223
rect 1747 165 1803 189
rect 1555 153 1803 165
rect 1555 119 1565 153
rect 1599 119 1662 153
rect 1696 119 1759 153
rect 1793 119 1803 153
rect 1555 103 1803 119
rect 2036 361 2092 377
rect 2036 327 2046 361
rect 2080 327 2092 361
rect 2036 289 2092 327
rect 2122 361 2286 377
rect 2122 332 2143 361
tri 2122 316 2138 332 ne
rect 2138 327 2143 332
rect 2177 327 2240 361
rect 2274 327 2286 361
rect 2138 316 2286 327
rect 2316 340 2478 377
tri 2316 324 2332 340 ne
rect 2332 324 2478 340
rect 2036 255 2046 289
rect 2080 255 2092 289
tri 2198 286 2228 316 ne
rect 2228 289 2286 316
tri 2392 294 2422 324 ne
rect 2036 221 2092 255
rect 2036 187 2046 221
rect 2080 187 2092 221
rect 2036 155 2092 187
tri 2122 270 2138 286 se
rect 2138 270 2182 286
tri 2182 270 2198 286 sw
rect 2122 236 2198 270
rect 2122 202 2143 236
rect 2177 202 2198 236
rect 2122 201 2198 202
tri 2122 185 2138 201 ne
rect 2138 185 2182 201
tri 2182 185 2198 201 nw
rect 2228 255 2240 289
rect 2274 255 2286 289
rect 2228 221 2286 255
rect 2228 187 2240 221
rect 2274 187 2286 221
tri 2316 278 2332 294 se
rect 2332 278 2376 294
tri 2376 278 2392 294 sw
rect 2316 245 2392 278
rect 2316 211 2337 245
rect 2371 211 2392 245
rect 2316 209 2392 211
tri 2316 193 2332 209 ne
rect 2332 193 2376 209
tri 2376 193 2392 209 nw
rect 2422 289 2478 324
rect 2422 255 2434 289
rect 2468 255 2478 289
rect 2422 221 2478 255
tri 2092 155 2122 185 sw
tri 2198 155 2228 185 se
rect 2228 163 2286 187
tri 2286 163 2316 193 sw
tri 2392 163 2422 193 se
rect 2422 187 2434 221
rect 2468 187 2478 221
rect 2422 163 2478 187
rect 2228 155 2478 163
rect 2036 151 2478 155
rect 2036 117 2046 151
rect 2080 117 2240 151
rect 2274 117 2337 151
rect 2371 117 2434 151
rect 2468 117 2478 151
rect 2036 101 2478 117
rect 2681 363 2737 379
rect 2681 329 2691 363
rect 2725 329 2737 363
rect 2681 291 2737 329
rect 2767 363 3037 379
rect 2767 334 2788 363
tri 2767 318 2783 334 ne
rect 2783 329 2788 334
rect 2822 329 2885 363
rect 2919 329 2982 363
rect 3016 329 3037 363
rect 2783 318 3037 329
rect 3067 363 3123 379
rect 3067 329 3079 363
rect 3113 329 3123 363
rect 2681 257 2691 291
rect 2725 257 2737 291
tri 2843 288 2873 318 ne
rect 2873 291 2932 318
rect 2681 223 2737 257
rect 2681 189 2691 223
rect 2725 189 2737 223
rect 2681 157 2737 189
tri 2767 272 2783 288 se
rect 2783 272 2827 288
tri 2827 272 2843 288 sw
rect 2767 238 2843 272
rect 2767 204 2788 238
rect 2822 204 2843 238
rect 2767 203 2843 204
tri 2767 187 2783 203 ne
rect 2783 187 2827 203
tri 2827 187 2843 203 nw
rect 2873 257 2885 291
rect 2919 257 2932 291
tri 2932 288 2962 318 nw
rect 2873 223 2932 257
rect 2873 189 2885 223
rect 2919 189 2932 223
tri 2962 272 2978 288 se
rect 2978 272 3021 288
tri 3021 272 3037 288 sw
rect 2962 244 3037 272
rect 2962 210 2983 244
rect 3017 210 3037 244
tri 2962 194 2978 210 ne
rect 2978 194 3021 210
tri 3021 194 3037 210 nw
tri 2737 157 2767 187 sw
tri 2843 157 2873 187 se
rect 2873 164 2932 189
tri 2932 164 2962 194 sw
tri 3037 164 3067 194 se
rect 3067 164 3123 329
rect 2873 157 3123 164
rect 2681 153 3123 157
rect 2681 119 2691 153
rect 2725 119 2885 153
rect 2919 119 2982 153
rect 3016 119 3079 153
rect 3113 119 3123 153
rect 2681 103 3123 119
rect 3183 363 3239 379
rect 3183 329 3193 363
rect 3227 329 3239 363
rect 3183 291 3239 329
rect 3269 342 3431 379
tri 3269 326 3285 342 ne
rect 3285 326 3431 342
tri 3345 296 3375 326 ne
rect 3183 257 3193 291
rect 3227 257 3239 291
rect 3183 223 3239 257
rect 3183 189 3193 223
rect 3227 189 3239 223
tri 3269 280 3285 296 se
rect 3285 280 3329 296
tri 3329 280 3345 296 sw
rect 3269 247 3345 280
rect 3269 213 3290 247
rect 3324 213 3345 247
rect 3269 211 3345 213
tri 3269 195 3285 211 ne
rect 3285 195 3329 211
tri 3329 195 3345 211 nw
rect 3375 291 3431 326
rect 3375 257 3387 291
rect 3421 257 3431 291
rect 3375 223 3431 257
rect 3183 165 3239 189
tri 3239 165 3269 195 sw
tri 3345 165 3375 195 se
rect 3375 189 3387 223
rect 3421 189 3431 223
rect 3375 165 3431 189
rect 3183 153 3431 165
rect 3183 119 3193 153
rect 3227 119 3290 153
rect 3324 119 3387 153
rect 3421 119 3431 153
rect 3183 103 3431 119
rect 3643 363 3699 379
rect 3643 329 3653 363
rect 3687 329 3699 363
rect 3643 291 3699 329
rect 3729 363 3999 379
rect 3729 334 3750 363
tri 3729 318 3745 334 ne
rect 3745 329 3750 334
rect 3784 329 3847 363
rect 3881 329 3944 363
rect 3978 329 3999 363
rect 3745 318 3999 329
rect 4029 363 4085 379
rect 4029 329 4041 363
rect 4075 329 4085 363
rect 3643 257 3653 291
rect 3687 257 3699 291
tri 3805 288 3835 318 ne
rect 3835 291 3894 318
rect 3643 223 3699 257
rect 3643 189 3653 223
rect 3687 189 3699 223
rect 3643 157 3699 189
tri 3729 272 3745 288 se
rect 3745 272 3789 288
tri 3789 272 3805 288 sw
rect 3729 238 3805 272
rect 3729 204 3750 238
rect 3784 204 3805 238
rect 3729 203 3805 204
tri 3729 187 3745 203 ne
rect 3745 187 3789 203
tri 3789 187 3805 203 nw
rect 3835 257 3847 291
rect 3881 257 3894 291
tri 3894 288 3924 318 nw
rect 3835 223 3894 257
rect 3835 189 3847 223
rect 3881 189 3894 223
tri 3924 272 3940 288 se
rect 3940 272 3983 288
tri 3983 272 3999 288 sw
rect 3924 244 3999 272
rect 3924 210 3945 244
rect 3979 210 3999 244
tri 3924 194 3940 210 ne
rect 3940 194 3983 210
tri 3983 194 3999 210 nw
tri 3699 157 3729 187 sw
tri 3805 157 3835 187 se
rect 3835 164 3894 189
tri 3894 164 3924 194 sw
tri 3999 164 4029 194 se
rect 4029 164 4085 329
rect 3835 157 4085 164
rect 3643 153 4085 157
rect 3643 119 3653 153
rect 3687 119 3847 153
rect 3881 119 3944 153
rect 3978 119 4041 153
rect 4075 119 4085 153
rect 3643 103 4085 119
rect 4145 363 4201 379
rect 4145 329 4155 363
rect 4189 329 4201 363
rect 4145 291 4201 329
rect 4231 342 4393 379
tri 4231 326 4247 342 ne
rect 4247 326 4393 342
tri 4307 296 4337 326 ne
rect 4145 257 4155 291
rect 4189 257 4201 291
rect 4145 223 4201 257
rect 4145 189 4155 223
rect 4189 189 4201 223
tri 4231 280 4247 296 se
rect 4247 280 4291 296
tri 4291 280 4307 296 sw
rect 4231 247 4307 280
rect 4231 213 4252 247
rect 4286 213 4307 247
rect 4231 211 4307 213
tri 4231 195 4247 211 ne
rect 4247 195 4291 211
tri 4291 195 4307 211 nw
rect 4337 291 4393 326
rect 4337 257 4349 291
rect 4383 257 4393 291
rect 4337 223 4393 257
rect 4145 165 4201 189
tri 4201 165 4231 195 sw
tri 4307 165 4337 195 se
rect 4337 189 4349 223
rect 4383 189 4393 223
rect 4337 165 4393 189
rect 4145 153 4393 165
rect 4145 119 4155 153
rect 4189 119 4252 153
rect 4286 119 4349 153
rect 4383 119 4393 153
rect 4145 103 4393 119
rect 4626 361 4682 377
rect 4626 327 4636 361
rect 4670 327 4682 361
rect 4626 289 4682 327
rect 4712 361 4876 377
rect 4712 332 4733 361
tri 4712 316 4728 332 ne
rect 4728 327 4733 332
rect 4767 327 4830 361
rect 4864 327 4876 361
rect 4728 316 4876 327
rect 4906 340 5068 377
tri 4906 324 4922 340 ne
rect 4922 324 5068 340
rect 4626 255 4636 289
rect 4670 255 4682 289
tri 4788 286 4818 316 ne
rect 4818 289 4876 316
tri 4982 294 5012 324 ne
rect 4626 221 4682 255
rect 4626 187 4636 221
rect 4670 187 4682 221
rect 4626 155 4682 187
tri 4712 270 4728 286 se
rect 4728 270 4772 286
tri 4772 270 4788 286 sw
rect 4712 236 4788 270
rect 4712 202 4733 236
rect 4767 202 4788 236
rect 4712 201 4788 202
tri 4712 185 4728 201 ne
rect 4728 185 4772 201
tri 4772 185 4788 201 nw
rect 4818 255 4830 289
rect 4864 255 4876 289
rect 4818 221 4876 255
rect 4818 187 4830 221
rect 4864 187 4876 221
tri 4906 278 4922 294 se
rect 4922 278 4966 294
tri 4966 278 4982 294 sw
rect 4906 245 4982 278
rect 4906 211 4927 245
rect 4961 211 4982 245
rect 4906 209 4982 211
tri 4906 193 4922 209 ne
rect 4922 193 4966 209
tri 4966 193 4982 209 nw
rect 5012 289 5068 324
rect 5012 255 5024 289
rect 5058 255 5068 289
rect 5012 221 5068 255
tri 4682 155 4712 185 sw
tri 4788 155 4818 185 se
rect 4818 163 4876 187
tri 4876 163 4906 193 sw
tri 4982 163 5012 193 se
rect 5012 187 5024 221
rect 5058 187 5068 221
rect 5012 163 5068 187
rect 4818 155 5068 163
rect 4626 151 5068 155
rect 4626 117 4636 151
rect 4670 117 4830 151
rect 4864 117 4927 151
rect 4961 117 5024 151
rect 5058 117 5068 151
rect 4626 101 5068 117
rect 5271 363 5327 379
rect 5271 329 5281 363
rect 5315 329 5327 363
rect 5271 291 5327 329
rect 5357 363 5627 379
rect 5357 334 5378 363
tri 5357 318 5373 334 ne
rect 5373 329 5378 334
rect 5412 329 5475 363
rect 5509 329 5572 363
rect 5606 329 5627 363
rect 5373 318 5627 329
rect 5657 363 5713 379
rect 5657 329 5669 363
rect 5703 329 5713 363
rect 5271 257 5281 291
rect 5315 257 5327 291
tri 5433 288 5463 318 ne
rect 5463 291 5522 318
rect 5271 223 5327 257
rect 5271 189 5281 223
rect 5315 189 5327 223
rect 5271 157 5327 189
tri 5357 272 5373 288 se
rect 5373 272 5417 288
tri 5417 272 5433 288 sw
rect 5357 238 5433 272
rect 5357 204 5378 238
rect 5412 204 5433 238
rect 5357 203 5433 204
tri 5357 187 5373 203 ne
rect 5373 187 5417 203
tri 5417 187 5433 203 nw
rect 5463 257 5475 291
rect 5509 257 5522 291
tri 5522 288 5552 318 nw
rect 5463 223 5522 257
rect 5463 189 5475 223
rect 5509 189 5522 223
tri 5552 272 5568 288 se
rect 5568 272 5611 288
tri 5611 272 5627 288 sw
rect 5552 244 5627 272
rect 5552 210 5573 244
rect 5607 210 5627 244
tri 5552 194 5568 210 ne
rect 5568 194 5611 210
tri 5611 194 5627 210 nw
tri 5327 157 5357 187 sw
tri 5433 157 5463 187 se
rect 5463 164 5522 189
tri 5522 164 5552 194 sw
tri 5627 164 5657 194 se
rect 5657 164 5713 329
rect 5463 157 5713 164
rect 5271 153 5713 157
rect 5271 119 5281 153
rect 5315 119 5475 153
rect 5509 119 5572 153
rect 5606 119 5669 153
rect 5703 119 5713 153
rect 5271 103 5713 119
rect 5773 363 5829 379
rect 5773 329 5783 363
rect 5817 329 5829 363
rect 5773 291 5829 329
rect 5859 342 6021 379
tri 5859 326 5875 342 ne
rect 5875 326 6021 342
tri 5935 296 5965 326 ne
rect 5773 257 5783 291
rect 5817 257 5829 291
rect 5773 223 5829 257
rect 5773 189 5783 223
rect 5817 189 5829 223
tri 5859 280 5875 296 se
rect 5875 280 5919 296
tri 5919 280 5935 296 sw
rect 5859 247 5935 280
rect 5859 213 5880 247
rect 5914 213 5935 247
rect 5859 211 5935 213
tri 5859 195 5875 211 ne
rect 5875 195 5919 211
tri 5919 195 5935 211 nw
rect 5965 291 6021 326
rect 5965 257 5977 291
rect 6011 257 6021 291
rect 5965 223 6021 257
rect 5773 165 5829 189
tri 5829 165 5859 195 sw
tri 5935 165 5965 195 se
rect 5965 189 5977 223
rect 6011 189 6021 223
rect 5965 165 6021 189
rect 5773 153 6021 165
rect 5773 119 5783 153
rect 5817 119 5880 153
rect 5914 119 5977 153
rect 6011 119 6021 153
rect 5773 103 6021 119
rect 6233 363 6289 379
rect 6233 329 6243 363
rect 6277 329 6289 363
rect 6233 291 6289 329
rect 6319 363 6589 379
rect 6319 334 6340 363
tri 6319 318 6335 334 ne
rect 6335 329 6340 334
rect 6374 329 6437 363
rect 6471 329 6534 363
rect 6568 329 6589 363
rect 6335 318 6589 329
rect 6619 363 6675 379
rect 6619 329 6631 363
rect 6665 329 6675 363
rect 6233 257 6243 291
rect 6277 257 6289 291
tri 6395 288 6425 318 ne
rect 6425 291 6484 318
rect 6233 223 6289 257
rect 6233 189 6243 223
rect 6277 189 6289 223
rect 6233 157 6289 189
tri 6319 272 6335 288 se
rect 6335 272 6379 288
tri 6379 272 6395 288 sw
rect 6319 238 6395 272
rect 6319 204 6340 238
rect 6374 204 6395 238
rect 6319 203 6395 204
tri 6319 187 6335 203 ne
rect 6335 187 6379 203
tri 6379 187 6395 203 nw
rect 6425 257 6437 291
rect 6471 257 6484 291
tri 6484 288 6514 318 nw
rect 6425 223 6484 257
rect 6425 189 6437 223
rect 6471 189 6484 223
tri 6514 272 6530 288 se
rect 6530 272 6573 288
tri 6573 272 6589 288 sw
rect 6514 244 6589 272
rect 6514 210 6535 244
rect 6569 210 6589 244
tri 6514 194 6530 210 ne
rect 6530 194 6573 210
tri 6573 194 6589 210 nw
tri 6289 157 6319 187 sw
tri 6395 157 6425 187 se
rect 6425 164 6484 189
tri 6484 164 6514 194 sw
tri 6589 164 6619 194 se
rect 6619 164 6675 329
rect 6425 157 6675 164
rect 6233 153 6675 157
rect 6233 119 6243 153
rect 6277 119 6437 153
rect 6471 119 6534 153
rect 6568 119 6631 153
rect 6665 119 6675 153
rect 6233 103 6675 119
rect 6735 363 6791 379
rect 6735 329 6745 363
rect 6779 329 6791 363
rect 6735 291 6791 329
rect 6821 342 6983 379
tri 6821 326 6837 342 ne
rect 6837 326 6983 342
tri 6897 296 6927 326 ne
rect 6735 257 6745 291
rect 6779 257 6791 291
rect 6735 223 6791 257
rect 6735 189 6745 223
rect 6779 189 6791 223
tri 6821 280 6837 296 se
rect 6837 280 6881 296
tri 6881 280 6897 296 sw
rect 6821 247 6897 280
rect 6821 213 6842 247
rect 6876 213 6897 247
rect 6821 211 6897 213
tri 6821 195 6837 211 ne
rect 6837 195 6881 211
tri 6881 195 6897 211 nw
rect 6927 291 6983 326
rect 6927 257 6939 291
rect 6973 257 6983 291
rect 6927 223 6983 257
rect 6735 165 6791 189
tri 6791 165 6821 195 sw
tri 6897 165 6927 195 se
rect 6927 189 6939 223
rect 6973 189 6983 223
rect 6927 165 6983 189
rect 6735 153 6983 165
rect 6735 119 6745 153
rect 6779 119 6842 153
rect 6876 119 6939 153
rect 6973 119 6983 153
rect 6735 103 6983 119
rect 7216 361 7272 377
rect 7216 327 7226 361
rect 7260 327 7272 361
rect 7216 289 7272 327
rect 7302 361 7466 377
rect 7302 332 7323 361
tri 7302 316 7318 332 ne
rect 7318 327 7323 332
rect 7357 327 7420 361
rect 7454 327 7466 361
rect 7318 316 7466 327
rect 7496 340 7658 377
tri 7496 324 7512 340 ne
rect 7512 324 7658 340
rect 7216 255 7226 289
rect 7260 255 7272 289
tri 7378 286 7408 316 ne
rect 7408 289 7466 316
tri 7572 294 7602 324 ne
rect 7216 221 7272 255
rect 7216 187 7226 221
rect 7260 187 7272 221
rect 7216 155 7272 187
tri 7302 270 7318 286 se
rect 7318 270 7362 286
tri 7362 270 7378 286 sw
rect 7302 236 7378 270
rect 7302 202 7323 236
rect 7357 202 7378 236
rect 7302 201 7378 202
tri 7302 185 7318 201 ne
rect 7318 185 7362 201
tri 7362 185 7378 201 nw
rect 7408 255 7420 289
rect 7454 255 7466 289
rect 7408 221 7466 255
rect 7408 187 7420 221
rect 7454 187 7466 221
tri 7496 278 7512 294 se
rect 7512 278 7556 294
tri 7556 278 7572 294 sw
rect 7496 245 7572 278
rect 7496 211 7517 245
rect 7551 211 7572 245
rect 7496 209 7572 211
tri 7496 193 7512 209 ne
rect 7512 193 7556 209
tri 7556 193 7572 209 nw
rect 7602 289 7658 324
rect 7602 255 7614 289
rect 7648 255 7658 289
rect 7602 221 7658 255
tri 7272 155 7302 185 sw
tri 7378 155 7408 185 se
rect 7408 163 7466 187
tri 7466 163 7496 193 sw
tri 7572 163 7602 193 se
rect 7602 187 7614 221
rect 7648 187 7658 221
rect 7602 163 7658 187
rect 7408 155 7658 163
rect 7216 151 7658 155
rect 7216 117 7226 151
rect 7260 117 7420 151
rect 7454 117 7517 151
rect 7551 117 7614 151
rect 7648 117 7658 151
rect 7216 101 7658 117
rect 7861 363 7917 379
rect 7861 329 7871 363
rect 7905 329 7917 363
rect 7861 291 7917 329
rect 7947 363 8217 379
rect 7947 334 7968 363
tri 7947 318 7963 334 ne
rect 7963 329 7968 334
rect 8002 329 8065 363
rect 8099 329 8162 363
rect 8196 329 8217 363
rect 7963 318 8217 329
rect 8247 363 8303 379
rect 8247 329 8259 363
rect 8293 329 8303 363
rect 7861 257 7871 291
rect 7905 257 7917 291
tri 8023 288 8053 318 ne
rect 8053 291 8112 318
rect 7861 223 7917 257
rect 7861 189 7871 223
rect 7905 189 7917 223
rect 7861 157 7917 189
tri 7947 272 7963 288 se
rect 7963 272 8007 288
tri 8007 272 8023 288 sw
rect 7947 238 8023 272
rect 7947 204 7968 238
rect 8002 204 8023 238
rect 7947 203 8023 204
tri 7947 187 7963 203 ne
rect 7963 187 8007 203
tri 8007 187 8023 203 nw
rect 8053 257 8065 291
rect 8099 257 8112 291
tri 8112 288 8142 318 nw
rect 8053 223 8112 257
rect 8053 189 8065 223
rect 8099 189 8112 223
tri 8142 272 8158 288 se
rect 8158 272 8201 288
tri 8201 272 8217 288 sw
rect 8142 244 8217 272
rect 8142 210 8163 244
rect 8197 210 8217 244
tri 8142 194 8158 210 ne
rect 8158 194 8201 210
tri 8201 194 8217 210 nw
tri 7917 157 7947 187 sw
tri 8023 157 8053 187 se
rect 8053 164 8112 189
tri 8112 164 8142 194 sw
tri 8217 164 8247 194 se
rect 8247 164 8303 329
rect 8053 157 8303 164
rect 7861 153 8303 157
rect 7861 119 7871 153
rect 7905 119 8065 153
rect 8099 119 8162 153
rect 8196 119 8259 153
rect 8293 119 8303 153
rect 7861 103 8303 119
rect 8363 363 8419 379
rect 8363 329 8373 363
rect 8407 329 8419 363
rect 8363 291 8419 329
rect 8449 342 8611 379
tri 8449 326 8465 342 ne
rect 8465 326 8611 342
tri 8525 296 8555 326 ne
rect 8363 257 8373 291
rect 8407 257 8419 291
rect 8363 223 8419 257
rect 8363 189 8373 223
rect 8407 189 8419 223
tri 8449 280 8465 296 se
rect 8465 280 8509 296
tri 8509 280 8525 296 sw
rect 8449 247 8525 280
rect 8449 213 8470 247
rect 8504 213 8525 247
rect 8449 211 8525 213
tri 8449 195 8465 211 ne
rect 8465 195 8509 211
tri 8509 195 8525 211 nw
rect 8555 291 8611 326
rect 8555 257 8567 291
rect 8601 257 8611 291
rect 8555 223 8611 257
rect 8363 165 8419 189
tri 8419 165 8449 195 sw
tri 8525 165 8555 195 se
rect 8555 189 8567 223
rect 8601 189 8611 223
rect 8555 165 8611 189
rect 8363 153 8611 165
rect 8363 119 8373 153
rect 8407 119 8470 153
rect 8504 119 8567 153
rect 8601 119 8611 153
rect 8363 103 8611 119
rect 8823 363 8879 379
rect 8823 329 8833 363
rect 8867 329 8879 363
rect 8823 291 8879 329
rect 8909 363 9179 379
rect 8909 334 8930 363
tri 8909 318 8925 334 ne
rect 8925 329 8930 334
rect 8964 329 9027 363
rect 9061 329 9124 363
rect 9158 329 9179 363
rect 8925 318 9179 329
rect 9209 363 9265 379
rect 9209 329 9221 363
rect 9255 329 9265 363
rect 8823 257 8833 291
rect 8867 257 8879 291
tri 8985 288 9015 318 ne
rect 9015 291 9074 318
rect 8823 223 8879 257
rect 8823 189 8833 223
rect 8867 189 8879 223
rect 8823 157 8879 189
tri 8909 272 8925 288 se
rect 8925 272 8969 288
tri 8969 272 8985 288 sw
rect 8909 238 8985 272
rect 8909 204 8930 238
rect 8964 204 8985 238
rect 8909 203 8985 204
tri 8909 187 8925 203 ne
rect 8925 187 8969 203
tri 8969 187 8985 203 nw
rect 9015 257 9027 291
rect 9061 257 9074 291
tri 9074 288 9104 318 nw
rect 9015 223 9074 257
rect 9015 189 9027 223
rect 9061 189 9074 223
tri 9104 272 9120 288 se
rect 9120 272 9163 288
tri 9163 272 9179 288 sw
rect 9104 244 9179 272
rect 9104 210 9125 244
rect 9159 210 9179 244
tri 9104 194 9120 210 ne
rect 9120 194 9163 210
tri 9163 194 9179 210 nw
tri 8879 157 8909 187 sw
tri 8985 157 9015 187 se
rect 9015 164 9074 189
tri 9074 164 9104 194 sw
tri 9179 164 9209 194 se
rect 9209 164 9265 329
rect 9015 157 9265 164
rect 8823 153 9265 157
rect 8823 119 8833 153
rect 8867 119 9027 153
rect 9061 119 9124 153
rect 9158 119 9221 153
rect 9255 119 9265 153
rect 8823 103 9265 119
rect 9325 363 9381 379
rect 9325 329 9335 363
rect 9369 329 9381 363
rect 9325 291 9381 329
rect 9411 342 9573 379
tri 9411 326 9427 342 ne
rect 9427 326 9573 342
tri 9487 296 9517 326 ne
rect 9325 257 9335 291
rect 9369 257 9381 291
rect 9325 223 9381 257
rect 9325 189 9335 223
rect 9369 189 9381 223
tri 9411 280 9427 296 se
rect 9427 280 9471 296
tri 9471 280 9487 296 sw
rect 9411 247 9487 280
rect 9411 213 9432 247
rect 9466 213 9487 247
rect 9411 211 9487 213
tri 9411 195 9427 211 ne
rect 9427 195 9471 211
tri 9471 195 9487 211 nw
rect 9517 291 9573 326
rect 9517 257 9529 291
rect 9563 257 9573 291
rect 9517 223 9573 257
rect 9325 165 9381 189
tri 9381 165 9411 195 sw
tri 9487 165 9517 195 se
rect 9517 189 9529 223
rect 9563 189 9573 223
rect 9517 165 9573 189
rect 9325 153 9573 165
rect 9325 119 9335 153
rect 9369 119 9432 153
rect 9466 119 9529 153
rect 9563 119 9573 153
rect 9325 103 9573 119
rect 9806 361 9862 377
rect 9806 327 9816 361
rect 9850 327 9862 361
rect 9806 289 9862 327
rect 9892 361 10056 377
rect 9892 332 9913 361
tri 9892 316 9908 332 ne
rect 9908 327 9913 332
rect 9947 327 10010 361
rect 10044 327 10056 361
rect 9908 316 10056 327
rect 10086 340 10248 377
tri 10086 324 10102 340 ne
rect 10102 324 10248 340
rect 9806 255 9816 289
rect 9850 255 9862 289
tri 9968 286 9998 316 ne
rect 9998 289 10056 316
tri 10162 294 10192 324 ne
rect 9806 221 9862 255
rect 9806 187 9816 221
rect 9850 187 9862 221
rect 9806 155 9862 187
tri 9892 270 9908 286 se
rect 9908 270 9952 286
tri 9952 270 9968 286 sw
rect 9892 236 9968 270
rect 9892 202 9913 236
rect 9947 202 9968 236
rect 9892 201 9968 202
tri 9892 185 9908 201 ne
rect 9908 185 9952 201
tri 9952 185 9968 201 nw
rect 9998 255 10010 289
rect 10044 255 10056 289
rect 9998 221 10056 255
rect 9998 187 10010 221
rect 10044 187 10056 221
tri 10086 278 10102 294 se
rect 10102 278 10146 294
tri 10146 278 10162 294 sw
rect 10086 245 10162 278
rect 10086 211 10107 245
rect 10141 211 10162 245
rect 10086 209 10162 211
tri 10086 193 10102 209 ne
rect 10102 193 10146 209
tri 10146 193 10162 209 nw
rect 10192 289 10248 324
rect 10192 255 10204 289
rect 10238 255 10248 289
rect 10192 221 10248 255
tri 9862 155 9892 185 sw
tri 9968 155 9998 185 se
rect 9998 163 10056 187
tri 10056 163 10086 193 sw
tri 10162 163 10192 193 se
rect 10192 187 10204 221
rect 10238 187 10248 221
rect 10192 163 10248 187
rect 9998 155 10248 163
rect 9806 151 10248 155
rect 9806 117 9816 151
rect 9850 117 10010 151
rect 10044 117 10107 151
rect 10141 117 10204 151
rect 10238 117 10248 151
rect 9806 101 10248 117
rect 10451 363 10507 379
rect 10451 329 10461 363
rect 10495 329 10507 363
rect 10451 291 10507 329
rect 10537 363 10807 379
rect 10537 334 10558 363
tri 10537 318 10553 334 ne
rect 10553 329 10558 334
rect 10592 329 10655 363
rect 10689 329 10752 363
rect 10786 329 10807 363
rect 10553 318 10807 329
rect 10837 363 10893 379
rect 10837 329 10849 363
rect 10883 329 10893 363
rect 10451 257 10461 291
rect 10495 257 10507 291
tri 10613 288 10643 318 ne
rect 10643 291 10702 318
rect 10451 223 10507 257
rect 10451 189 10461 223
rect 10495 189 10507 223
rect 10451 157 10507 189
tri 10537 272 10553 288 se
rect 10553 272 10597 288
tri 10597 272 10613 288 sw
rect 10537 238 10613 272
rect 10537 204 10558 238
rect 10592 204 10613 238
rect 10537 203 10613 204
tri 10537 187 10553 203 ne
rect 10553 187 10597 203
tri 10597 187 10613 203 nw
rect 10643 257 10655 291
rect 10689 257 10702 291
tri 10702 288 10732 318 nw
rect 10643 223 10702 257
rect 10643 189 10655 223
rect 10689 189 10702 223
tri 10732 272 10748 288 se
rect 10748 272 10791 288
tri 10791 272 10807 288 sw
rect 10732 244 10807 272
rect 10732 210 10753 244
rect 10787 210 10807 244
tri 10732 194 10748 210 ne
rect 10748 194 10791 210
tri 10791 194 10807 210 nw
tri 10507 157 10537 187 sw
tri 10613 157 10643 187 se
rect 10643 164 10702 189
tri 10702 164 10732 194 sw
tri 10807 164 10837 194 se
rect 10837 164 10893 329
rect 10643 157 10893 164
rect 10451 153 10893 157
rect 10451 119 10461 153
rect 10495 119 10655 153
rect 10689 119 10752 153
rect 10786 119 10849 153
rect 10883 119 10893 153
rect 10451 103 10893 119
rect 10953 363 11009 379
rect 10953 329 10963 363
rect 10997 329 11009 363
rect 10953 291 11009 329
rect 11039 342 11201 379
tri 11039 326 11055 342 ne
rect 11055 326 11201 342
tri 11115 296 11145 326 ne
rect 10953 257 10963 291
rect 10997 257 11009 291
rect 10953 223 11009 257
rect 10953 189 10963 223
rect 10997 189 11009 223
tri 11039 280 11055 296 se
rect 11055 280 11099 296
tri 11099 280 11115 296 sw
rect 11039 247 11115 280
rect 11039 213 11060 247
rect 11094 213 11115 247
rect 11039 211 11115 213
tri 11039 195 11055 211 ne
rect 11055 195 11099 211
tri 11099 195 11115 211 nw
rect 11145 291 11201 326
rect 11145 257 11157 291
rect 11191 257 11201 291
rect 11145 223 11201 257
rect 10953 165 11009 189
tri 11009 165 11039 195 sw
tri 11115 165 11145 195 se
rect 11145 189 11157 223
rect 11191 189 11201 223
rect 11145 165 11201 189
rect 10953 153 11201 165
rect 10953 119 10963 153
rect 10997 119 11060 153
rect 11094 119 11157 153
rect 11191 119 11201 153
rect 10953 103 11201 119
rect 11413 363 11469 379
rect 11413 329 11423 363
rect 11457 329 11469 363
rect 11413 291 11469 329
rect 11499 363 11769 379
rect 11499 334 11520 363
tri 11499 318 11515 334 ne
rect 11515 329 11520 334
rect 11554 329 11617 363
rect 11651 329 11714 363
rect 11748 329 11769 363
rect 11515 318 11769 329
rect 11799 363 11855 379
rect 11799 329 11811 363
rect 11845 329 11855 363
rect 11413 257 11423 291
rect 11457 257 11469 291
tri 11575 288 11605 318 ne
rect 11605 291 11664 318
rect 11413 223 11469 257
rect 11413 189 11423 223
rect 11457 189 11469 223
rect 11413 157 11469 189
tri 11499 272 11515 288 se
rect 11515 272 11559 288
tri 11559 272 11575 288 sw
rect 11499 238 11575 272
rect 11499 204 11520 238
rect 11554 204 11575 238
rect 11499 203 11575 204
tri 11499 187 11515 203 ne
rect 11515 187 11559 203
tri 11559 187 11575 203 nw
rect 11605 257 11617 291
rect 11651 257 11664 291
tri 11664 288 11694 318 nw
rect 11605 223 11664 257
rect 11605 189 11617 223
rect 11651 189 11664 223
tri 11694 272 11710 288 se
rect 11710 272 11753 288
tri 11753 272 11769 288 sw
rect 11694 244 11769 272
rect 11694 210 11715 244
rect 11749 210 11769 244
tri 11694 194 11710 210 ne
rect 11710 194 11753 210
tri 11753 194 11769 210 nw
tri 11469 157 11499 187 sw
tri 11575 157 11605 187 se
rect 11605 164 11664 189
tri 11664 164 11694 194 sw
tri 11769 164 11799 194 se
rect 11799 164 11855 329
rect 11605 157 11855 164
rect 11413 153 11855 157
rect 11413 119 11423 153
rect 11457 119 11617 153
rect 11651 119 11714 153
rect 11748 119 11811 153
rect 11845 119 11855 153
rect 11413 103 11855 119
rect 11915 363 11971 379
rect 11915 329 11925 363
rect 11959 329 11971 363
rect 11915 291 11971 329
rect 12001 342 12163 379
tri 12001 326 12017 342 ne
rect 12017 326 12163 342
tri 12077 296 12107 326 ne
rect 11915 257 11925 291
rect 11959 257 11971 291
rect 11915 223 11971 257
rect 11915 189 11925 223
rect 11959 189 11971 223
tri 12001 280 12017 296 se
rect 12017 280 12061 296
tri 12061 280 12077 296 sw
rect 12001 247 12077 280
rect 12001 213 12022 247
rect 12056 213 12077 247
rect 12001 211 12077 213
tri 12001 195 12017 211 ne
rect 12017 195 12061 211
tri 12061 195 12077 211 nw
rect 12107 291 12163 326
rect 12107 257 12119 291
rect 12153 257 12163 291
rect 12107 223 12163 257
rect 11915 165 11971 189
tri 11971 165 12001 195 sw
tri 12077 165 12107 195 se
rect 12107 189 12119 223
rect 12153 189 12163 223
rect 12107 165 12163 189
rect 11915 153 12163 165
rect 11915 119 11925 153
rect 11959 119 12022 153
rect 12056 119 12119 153
rect 12153 119 12163 153
rect 11915 103 12163 119
rect 12396 361 12452 377
rect 12396 327 12406 361
rect 12440 327 12452 361
rect 12396 289 12452 327
rect 12482 361 12646 377
rect 12482 332 12503 361
tri 12482 316 12498 332 ne
rect 12498 327 12503 332
rect 12537 327 12600 361
rect 12634 327 12646 361
rect 12498 316 12646 327
rect 12676 340 12838 377
tri 12676 324 12692 340 ne
rect 12692 324 12838 340
rect 12396 255 12406 289
rect 12440 255 12452 289
tri 12558 286 12588 316 ne
rect 12588 289 12646 316
tri 12752 294 12782 324 ne
rect 12396 221 12452 255
rect 12396 187 12406 221
rect 12440 187 12452 221
rect 12396 155 12452 187
tri 12482 270 12498 286 se
rect 12498 270 12542 286
tri 12542 270 12558 286 sw
rect 12482 236 12558 270
rect 12482 202 12503 236
rect 12537 202 12558 236
rect 12482 201 12558 202
tri 12482 185 12498 201 ne
rect 12498 185 12542 201
tri 12542 185 12558 201 nw
rect 12588 255 12600 289
rect 12634 255 12646 289
rect 12588 221 12646 255
rect 12588 187 12600 221
rect 12634 187 12646 221
tri 12676 278 12692 294 se
rect 12692 278 12736 294
tri 12736 278 12752 294 sw
rect 12676 245 12752 278
rect 12676 211 12697 245
rect 12731 211 12752 245
rect 12676 209 12752 211
tri 12676 193 12692 209 ne
rect 12692 193 12736 209
tri 12736 193 12752 209 nw
rect 12782 289 12838 324
rect 12782 255 12794 289
rect 12828 255 12838 289
rect 12782 221 12838 255
tri 12452 155 12482 185 sw
tri 12558 155 12588 185 se
rect 12588 163 12646 187
tri 12646 163 12676 193 sw
tri 12752 163 12782 193 se
rect 12782 187 12794 221
rect 12828 187 12838 221
rect 12782 163 12838 187
rect 12588 155 12838 163
rect 12396 151 12838 155
rect 12396 117 12406 151
rect 12440 117 12600 151
rect 12634 117 12697 151
rect 12731 117 12794 151
rect 12828 117 12838 151
rect 12396 101 12838 117
rect 13041 363 13097 379
rect 13041 329 13051 363
rect 13085 329 13097 363
rect 13041 291 13097 329
rect 13127 363 13397 379
rect 13127 334 13148 363
tri 13127 318 13143 334 ne
rect 13143 329 13148 334
rect 13182 329 13245 363
rect 13279 329 13342 363
rect 13376 329 13397 363
rect 13143 318 13397 329
rect 13427 363 13483 379
rect 13427 329 13439 363
rect 13473 329 13483 363
rect 13041 257 13051 291
rect 13085 257 13097 291
tri 13203 288 13233 318 ne
rect 13233 291 13292 318
rect 13041 223 13097 257
rect 13041 189 13051 223
rect 13085 189 13097 223
rect 13041 157 13097 189
tri 13127 272 13143 288 se
rect 13143 272 13187 288
tri 13187 272 13203 288 sw
rect 13127 238 13203 272
rect 13127 204 13148 238
rect 13182 204 13203 238
rect 13127 203 13203 204
tri 13127 187 13143 203 ne
rect 13143 187 13187 203
tri 13187 187 13203 203 nw
rect 13233 257 13245 291
rect 13279 257 13292 291
tri 13292 288 13322 318 nw
rect 13233 223 13292 257
rect 13233 189 13245 223
rect 13279 189 13292 223
tri 13322 272 13338 288 se
rect 13338 272 13381 288
tri 13381 272 13397 288 sw
rect 13322 244 13397 272
rect 13322 210 13343 244
rect 13377 210 13397 244
tri 13322 194 13338 210 ne
rect 13338 194 13381 210
tri 13381 194 13397 210 nw
tri 13097 157 13127 187 sw
tri 13203 157 13233 187 se
rect 13233 164 13292 189
tri 13292 164 13322 194 sw
tri 13397 164 13427 194 se
rect 13427 164 13483 329
rect 13233 157 13483 164
rect 13041 153 13483 157
rect 13041 119 13051 153
rect 13085 119 13245 153
rect 13279 119 13342 153
rect 13376 119 13439 153
rect 13473 119 13483 153
rect 13041 103 13483 119
rect 13543 363 13599 379
rect 13543 329 13553 363
rect 13587 329 13599 363
rect 13543 291 13599 329
rect 13629 342 13791 379
tri 13629 326 13645 342 ne
rect 13645 326 13791 342
tri 13705 296 13735 326 ne
rect 13543 257 13553 291
rect 13587 257 13599 291
rect 13543 223 13599 257
rect 13543 189 13553 223
rect 13587 189 13599 223
tri 13629 280 13645 296 se
rect 13645 280 13689 296
tri 13689 280 13705 296 sw
rect 13629 247 13705 280
rect 13629 213 13650 247
rect 13684 213 13705 247
rect 13629 211 13705 213
tri 13629 195 13645 211 ne
rect 13645 195 13689 211
tri 13689 195 13705 211 nw
rect 13735 291 13791 326
rect 13735 257 13747 291
rect 13781 257 13791 291
rect 13735 223 13791 257
rect 13543 165 13599 189
tri 13599 165 13629 195 sw
tri 13705 165 13735 195 se
rect 13735 189 13747 223
rect 13781 189 13791 223
rect 13735 165 13791 189
rect 13543 153 13791 165
rect 13543 119 13553 153
rect 13587 119 13650 153
rect 13684 119 13747 153
rect 13781 119 13791 153
rect 13543 103 13791 119
rect 14003 363 14059 379
rect 14003 329 14013 363
rect 14047 329 14059 363
rect 14003 291 14059 329
rect 14089 363 14359 379
rect 14089 334 14110 363
tri 14089 318 14105 334 ne
rect 14105 329 14110 334
rect 14144 329 14207 363
rect 14241 329 14304 363
rect 14338 329 14359 363
rect 14105 318 14359 329
rect 14389 363 14445 379
rect 14389 329 14401 363
rect 14435 329 14445 363
rect 14003 257 14013 291
rect 14047 257 14059 291
tri 14165 288 14195 318 ne
rect 14195 291 14254 318
rect 14003 223 14059 257
rect 14003 189 14013 223
rect 14047 189 14059 223
rect 14003 157 14059 189
tri 14089 272 14105 288 se
rect 14105 272 14149 288
tri 14149 272 14165 288 sw
rect 14089 238 14165 272
rect 14089 204 14110 238
rect 14144 204 14165 238
rect 14089 203 14165 204
tri 14089 187 14105 203 ne
rect 14105 187 14149 203
tri 14149 187 14165 203 nw
rect 14195 257 14207 291
rect 14241 257 14254 291
tri 14254 288 14284 318 nw
rect 14195 223 14254 257
rect 14195 189 14207 223
rect 14241 189 14254 223
tri 14284 272 14300 288 se
rect 14300 272 14343 288
tri 14343 272 14359 288 sw
rect 14284 244 14359 272
rect 14284 210 14305 244
rect 14339 210 14359 244
tri 14284 194 14300 210 ne
rect 14300 194 14343 210
tri 14343 194 14359 210 nw
tri 14059 157 14089 187 sw
tri 14165 157 14195 187 se
rect 14195 164 14254 189
tri 14254 164 14284 194 sw
tri 14359 164 14389 194 se
rect 14389 164 14445 329
rect 14195 157 14445 164
rect 14003 153 14445 157
rect 14003 119 14013 153
rect 14047 119 14207 153
rect 14241 119 14304 153
rect 14338 119 14401 153
rect 14435 119 14445 153
rect 14003 103 14445 119
rect 14505 363 14561 379
rect 14505 329 14515 363
rect 14549 329 14561 363
rect 14505 291 14561 329
rect 14591 342 14753 379
tri 14591 326 14607 342 ne
rect 14607 326 14753 342
tri 14667 296 14697 326 ne
rect 14505 257 14515 291
rect 14549 257 14561 291
rect 14505 223 14561 257
rect 14505 189 14515 223
rect 14549 189 14561 223
tri 14591 280 14607 296 se
rect 14607 280 14651 296
tri 14651 280 14667 296 sw
rect 14591 247 14667 280
rect 14591 213 14612 247
rect 14646 213 14667 247
rect 14591 211 14667 213
tri 14591 195 14607 211 ne
rect 14607 195 14651 211
tri 14651 195 14667 211 nw
rect 14697 291 14753 326
rect 14697 257 14709 291
rect 14743 257 14753 291
rect 14697 223 14753 257
rect 14505 165 14561 189
tri 14561 165 14591 195 sw
tri 14667 165 14697 195 se
rect 14697 189 14709 223
rect 14743 189 14753 223
rect 14697 165 14753 189
rect 14505 153 14753 165
rect 14505 119 14515 153
rect 14549 119 14612 153
rect 14646 119 14709 153
rect 14743 119 14753 153
rect 14505 103 14753 119
rect 14986 361 15042 377
rect 14986 327 14996 361
rect 15030 327 15042 361
rect 14986 289 15042 327
rect 15072 361 15236 377
rect 15072 332 15093 361
tri 15072 316 15088 332 ne
rect 15088 327 15093 332
rect 15127 327 15190 361
rect 15224 327 15236 361
rect 15088 316 15236 327
rect 15266 340 15428 377
tri 15266 324 15282 340 ne
rect 15282 324 15428 340
rect 14986 255 14996 289
rect 15030 255 15042 289
tri 15148 286 15178 316 ne
rect 15178 289 15236 316
tri 15342 294 15372 324 ne
rect 14986 221 15042 255
rect 14986 187 14996 221
rect 15030 187 15042 221
rect 14986 155 15042 187
tri 15072 270 15088 286 se
rect 15088 270 15132 286
tri 15132 270 15148 286 sw
rect 15072 236 15148 270
rect 15072 202 15093 236
rect 15127 202 15148 236
rect 15072 201 15148 202
tri 15072 185 15088 201 ne
rect 15088 185 15132 201
tri 15132 185 15148 201 nw
rect 15178 255 15190 289
rect 15224 255 15236 289
rect 15178 221 15236 255
rect 15178 187 15190 221
rect 15224 187 15236 221
tri 15266 278 15282 294 se
rect 15282 278 15326 294
tri 15326 278 15342 294 sw
rect 15266 245 15342 278
rect 15266 211 15287 245
rect 15321 211 15342 245
rect 15266 209 15342 211
tri 15266 193 15282 209 ne
rect 15282 193 15326 209
tri 15326 193 15342 209 nw
rect 15372 289 15428 324
rect 15372 255 15384 289
rect 15418 255 15428 289
rect 15372 221 15428 255
tri 15042 155 15072 185 sw
tri 15148 155 15178 185 se
rect 15178 163 15236 187
tri 15236 163 15266 193 sw
tri 15342 163 15372 193 se
rect 15372 187 15384 221
rect 15418 187 15428 221
rect 15372 163 15428 187
rect 15178 155 15428 163
rect 14986 151 15428 155
rect 14986 117 14996 151
rect 15030 117 15190 151
rect 15224 117 15287 151
rect 15321 117 15384 151
rect 15418 117 15428 151
rect 14986 101 15428 117
rect 15652 361 15708 377
rect 15652 327 15662 361
rect 15696 327 15708 361
rect 15652 289 15708 327
rect 15738 361 15902 377
rect 15738 332 15759 361
tri 15738 316 15754 332 ne
rect 15754 327 15759 332
rect 15793 327 15856 361
rect 15890 327 15902 361
rect 15754 316 15902 327
rect 15932 361 16092 377
rect 15932 340 16050 361
tri 15932 324 15948 340 ne
rect 15948 327 16050 340
rect 16084 327 16092 361
rect 15948 324 16092 327
rect 15652 255 15662 289
rect 15696 255 15708 289
tri 15814 286 15844 316 ne
rect 15844 289 15902 316
tri 16008 294 16038 324 ne
rect 15652 221 15708 255
rect 15652 187 15662 221
rect 15696 187 15708 221
rect 15652 155 15708 187
tri 15738 270 15754 286 se
rect 15754 270 15798 286
tri 15798 270 15814 286 sw
rect 15738 236 15814 270
rect 15738 202 15759 236
rect 15793 202 15814 236
rect 15738 201 15814 202
tri 15738 185 15754 201 ne
rect 15754 185 15798 201
tri 15798 185 15814 201 nw
rect 15844 255 15856 289
rect 15890 255 15902 289
rect 15844 221 15902 255
rect 15844 187 15856 221
rect 15890 187 15902 221
tri 15932 278 15948 294 se
rect 15948 278 15992 294
tri 15992 278 16008 294 sw
rect 15932 245 16008 278
rect 15932 211 15952 245
rect 15986 211 16008 245
rect 15932 209 16008 211
tri 15932 193 15948 209 ne
rect 15948 193 15992 209
tri 15992 193 16008 209 nw
rect 16038 289 16092 324
rect 16038 255 16050 289
rect 16084 255 16092 289
rect 16038 221 16092 255
tri 15708 155 15738 185 sw
tri 15814 155 15844 185 se
rect 15844 163 15902 187
tri 15902 163 15932 193 sw
tri 16008 163 16038 193 se
rect 16038 187 16050 221
rect 16084 187 16092 221
rect 16038 163 16092 187
rect 15844 155 16092 163
rect 15652 151 16092 155
rect 15652 117 15662 151
rect 15696 117 15856 151
rect 15890 117 15952 151
rect 15986 117 16050 151
rect 16084 117 16092 151
rect 15652 101 16092 117
rect 16318 361 16374 377
rect 16318 327 16328 361
rect 16362 327 16374 361
rect 16318 289 16374 327
rect 16404 361 16674 377
rect 16404 332 16425 361
tri 16404 316 16420 332 ne
rect 16420 327 16425 332
rect 16459 327 16522 361
rect 16556 340 16674 361
rect 16556 327 16658 340
rect 16420 324 16658 327
tri 16658 324 16674 340 nw
rect 16704 361 16760 377
rect 16704 327 16716 361
rect 16750 327 16760 361
rect 16420 316 16568 324
rect 16318 255 16328 289
rect 16362 255 16374 289
tri 16480 286 16510 316 ne
rect 16510 289 16568 316
tri 16568 294 16598 324 nw
rect 16318 221 16374 255
rect 16318 187 16328 221
rect 16362 187 16374 221
rect 16318 155 16374 187
tri 16404 270 16420 286 se
rect 16420 270 16464 286
tri 16464 270 16480 286 sw
rect 16404 236 16480 270
rect 16404 202 16425 236
rect 16459 202 16480 236
rect 16404 201 16480 202
tri 16404 185 16420 201 ne
rect 16420 185 16464 201
tri 16464 185 16480 201 nw
rect 16510 255 16522 289
rect 16556 255 16568 289
rect 16510 221 16568 255
rect 16510 187 16522 221
rect 16556 187 16568 221
tri 16598 278 16614 294 se
rect 16614 278 16658 294
tri 16658 278 16674 294 sw
rect 16598 245 16674 278
rect 16598 211 16619 245
rect 16653 211 16674 245
rect 16598 209 16674 211
tri 16598 193 16614 209 ne
rect 16614 193 16658 209
tri 16658 193 16674 209 nw
rect 16704 289 16760 327
rect 16704 255 16716 289
rect 16750 255 16760 289
rect 16704 221 16760 255
tri 16374 155 16404 185 sw
tri 16480 155 16510 185 se
rect 16510 163 16568 187
tri 16568 163 16598 193 sw
tri 16674 163 16704 193 se
rect 16704 187 16716 221
rect 16750 187 16760 221
rect 16704 163 16760 187
rect 16510 155 16760 163
rect 16318 151 16760 155
rect 16318 117 16328 151
rect 16362 117 16522 151
rect 16556 117 16619 151
rect 16653 117 16716 151
rect 16750 117 16760 151
rect 16318 101 16760 117
rect 16984 361 17040 377
rect 16984 327 16994 361
rect 17028 327 17040 361
rect 16984 289 17040 327
rect 17070 361 17234 377
rect 17070 332 17091 361
tri 17070 316 17086 332 ne
rect 17086 327 17091 332
rect 17125 327 17188 361
rect 17222 327 17234 361
rect 17086 316 17234 327
rect 17264 340 17426 377
tri 17264 324 17280 340 ne
rect 17280 324 17426 340
rect 16984 255 16994 289
rect 17028 255 17040 289
tri 17146 286 17176 316 ne
rect 17176 289 17234 316
tri 17340 294 17370 324 ne
rect 16984 221 17040 255
rect 16984 187 16994 221
rect 17028 187 17040 221
rect 16984 155 17040 187
tri 17070 270 17086 286 se
rect 17086 270 17130 286
tri 17130 270 17146 286 sw
rect 17070 236 17146 270
rect 17070 202 17091 236
rect 17125 202 17146 236
rect 17070 201 17146 202
tri 17070 185 17086 201 ne
rect 17086 185 17130 201
tri 17130 185 17146 201 nw
rect 17176 255 17188 289
rect 17222 255 17234 289
tri 17265 279 17280 294 se
rect 17280 279 17324 294
tri 17324 279 17339 294 sw
rect 17370 289 17426 324
rect 17176 221 17234 255
rect 17176 187 17188 221
rect 17222 187 17234 221
rect 17264 245 17340 279
rect 17264 211 17285 245
rect 17319 211 17340 245
rect 17264 209 17340 211
tri 17264 193 17280 209 ne
rect 17280 193 17324 209
tri 17324 193 17340 209 nw
rect 17370 255 17382 289
rect 17416 255 17426 289
rect 17370 221 17426 255
tri 17040 155 17070 185 sw
tri 17146 155 17176 185 se
rect 17176 163 17234 187
tri 17234 163 17264 193 sw
tri 17340 163 17370 193 se
rect 17370 187 17382 221
rect 17416 187 17426 221
rect 17370 163 17426 187
rect 17176 155 17426 163
rect 16984 151 17426 155
rect 16984 117 16994 151
rect 17028 117 17188 151
rect 17222 117 17285 151
rect 17319 117 17382 151
rect 17416 117 17426 151
rect 16984 101 17426 117
rect 17637 361 17693 377
rect 17637 327 17647 361
rect 17681 327 17693 361
rect 17637 289 17693 327
rect 17723 361 17883 377
rect 17723 340 17841 361
tri 17723 324 17739 340 ne
rect 17739 327 17841 340
rect 17875 327 17883 361
rect 17739 324 17883 327
tri 17799 294 17829 324 ne
rect 17637 255 17647 289
rect 17681 255 17693 289
rect 17637 221 17693 255
rect 17637 187 17647 221
rect 17681 187 17693 221
tri 17723 278 17739 294 se
rect 17739 278 17783 294
tri 17783 278 17799 294 sw
rect 17723 245 17799 278
rect 17723 211 17743 245
rect 17777 211 17799 245
rect 17723 209 17799 211
tri 17723 193 17739 209 ne
rect 17739 193 17783 209
tri 17783 193 17799 209 nw
rect 17829 289 17883 324
rect 17829 255 17841 289
rect 17875 255 17883 289
rect 17829 221 17883 255
rect 17637 163 17693 187
tri 17693 163 17723 193 sw
tri 17799 163 17829 193 se
rect 17829 187 17841 221
rect 17875 187 17883 221
rect 17829 163 17883 187
rect 17637 151 17883 163
rect 17637 117 17647 151
rect 17681 117 17743 151
rect 17777 117 17841 151
rect 17875 117 17883 151
rect 17637 101 17883 117
<< pdiff >>
rect 191 1412 247 1450
rect 191 1378 201 1412
rect 235 1378 247 1412
rect 191 1344 247 1378
rect 191 1310 201 1344
rect 235 1310 247 1344
rect 191 1276 247 1310
rect 191 1242 201 1276
rect 235 1242 247 1276
rect 191 1208 247 1242
rect 191 1174 201 1208
rect 235 1174 247 1208
rect 191 1139 247 1174
rect 191 1105 201 1139
rect 235 1105 247 1139
rect 191 1050 247 1105
rect 277 1412 335 1450
rect 277 1378 289 1412
rect 323 1378 335 1412
rect 277 1344 335 1378
rect 277 1310 289 1344
rect 323 1310 335 1344
rect 277 1276 335 1310
rect 277 1242 289 1276
rect 323 1242 335 1276
rect 277 1208 335 1242
rect 277 1174 289 1208
rect 323 1174 335 1208
rect 277 1139 335 1174
rect 277 1105 289 1139
rect 323 1105 335 1139
rect 277 1050 335 1105
rect 365 1412 423 1450
rect 365 1378 377 1412
rect 411 1378 423 1412
rect 365 1344 423 1378
rect 365 1310 377 1344
rect 411 1310 423 1344
rect 365 1276 423 1310
rect 365 1242 377 1276
rect 411 1242 423 1276
rect 365 1208 423 1242
rect 365 1174 377 1208
rect 411 1174 423 1208
rect 365 1050 423 1174
rect 453 1412 511 1450
rect 453 1378 465 1412
rect 499 1378 511 1412
rect 453 1344 511 1378
rect 453 1310 465 1344
rect 499 1310 511 1344
rect 453 1276 511 1310
rect 453 1242 465 1276
rect 499 1242 511 1276
rect 453 1208 511 1242
rect 453 1174 465 1208
rect 499 1174 511 1208
rect 453 1139 511 1174
rect 453 1105 465 1139
rect 499 1105 511 1139
rect 453 1050 511 1105
rect 541 1412 599 1450
rect 541 1378 553 1412
rect 587 1378 599 1412
rect 541 1344 599 1378
rect 541 1310 553 1344
rect 587 1310 599 1344
rect 541 1276 599 1310
rect 541 1242 553 1276
rect 587 1242 599 1276
rect 541 1208 599 1242
rect 541 1174 553 1208
rect 587 1174 599 1208
rect 541 1050 599 1174
rect 629 1412 687 1450
rect 629 1378 641 1412
rect 675 1378 687 1412
rect 629 1344 687 1378
rect 629 1310 641 1344
rect 675 1310 687 1344
rect 629 1276 687 1310
rect 629 1242 641 1276
rect 675 1242 687 1276
rect 629 1208 687 1242
rect 629 1174 641 1208
rect 675 1174 687 1208
rect 629 1139 687 1174
rect 629 1105 641 1139
rect 675 1105 687 1139
rect 629 1050 687 1105
rect 717 1412 771 1450
rect 717 1378 729 1412
rect 763 1378 771 1412
rect 717 1344 771 1378
rect 717 1310 729 1344
rect 763 1310 771 1344
rect 717 1276 771 1310
rect 717 1242 729 1276
rect 763 1242 771 1276
rect 717 1208 771 1242
rect 717 1174 729 1208
rect 763 1174 771 1208
rect 717 1050 771 1174
rect 1153 1412 1209 1450
rect 1153 1378 1163 1412
rect 1197 1378 1209 1412
rect 1153 1344 1209 1378
rect 1153 1310 1163 1344
rect 1197 1310 1209 1344
rect 1153 1276 1209 1310
rect 1153 1242 1163 1276
rect 1197 1242 1209 1276
rect 1153 1208 1209 1242
rect 1153 1174 1163 1208
rect 1197 1174 1209 1208
rect 1153 1139 1209 1174
rect 1153 1105 1163 1139
rect 1197 1105 1209 1139
rect 1153 1050 1209 1105
rect 1239 1412 1297 1450
rect 1239 1378 1251 1412
rect 1285 1378 1297 1412
rect 1239 1344 1297 1378
rect 1239 1310 1251 1344
rect 1285 1310 1297 1344
rect 1239 1276 1297 1310
rect 1239 1242 1251 1276
rect 1285 1242 1297 1276
rect 1239 1208 1297 1242
rect 1239 1174 1251 1208
rect 1285 1174 1297 1208
rect 1239 1139 1297 1174
rect 1239 1105 1251 1139
rect 1285 1105 1297 1139
rect 1239 1050 1297 1105
rect 1327 1412 1385 1450
rect 1327 1378 1339 1412
rect 1373 1378 1385 1412
rect 1327 1344 1385 1378
rect 1327 1310 1339 1344
rect 1373 1310 1385 1344
rect 1327 1276 1385 1310
rect 1327 1242 1339 1276
rect 1373 1242 1385 1276
rect 1327 1208 1385 1242
rect 1327 1174 1339 1208
rect 1373 1174 1385 1208
rect 1327 1050 1385 1174
rect 1415 1412 1473 1450
rect 1415 1378 1427 1412
rect 1461 1378 1473 1412
rect 1415 1344 1473 1378
rect 1415 1310 1427 1344
rect 1461 1310 1473 1344
rect 1415 1276 1473 1310
rect 1415 1242 1427 1276
rect 1461 1242 1473 1276
rect 1415 1208 1473 1242
rect 1415 1174 1427 1208
rect 1461 1174 1473 1208
rect 1415 1139 1473 1174
rect 1415 1105 1427 1139
rect 1461 1105 1473 1139
rect 1415 1050 1473 1105
rect 1503 1412 1561 1450
rect 1503 1378 1515 1412
rect 1549 1378 1561 1412
rect 1503 1344 1561 1378
rect 1503 1310 1515 1344
rect 1549 1310 1561 1344
rect 1503 1276 1561 1310
rect 1503 1242 1515 1276
rect 1549 1242 1561 1276
rect 1503 1208 1561 1242
rect 1503 1174 1515 1208
rect 1549 1174 1561 1208
rect 1503 1050 1561 1174
rect 1591 1412 1649 1450
rect 1591 1378 1603 1412
rect 1637 1378 1649 1412
rect 1591 1344 1649 1378
rect 1591 1310 1603 1344
rect 1637 1310 1649 1344
rect 1591 1276 1649 1310
rect 1591 1242 1603 1276
rect 1637 1242 1649 1276
rect 1591 1208 1649 1242
rect 1591 1174 1603 1208
rect 1637 1174 1649 1208
rect 1591 1139 1649 1174
rect 1591 1105 1603 1139
rect 1637 1105 1649 1139
rect 1591 1050 1649 1105
rect 1679 1412 1733 1450
rect 1679 1378 1691 1412
rect 1725 1378 1733 1412
rect 1679 1344 1733 1378
rect 1679 1310 1691 1344
rect 1725 1310 1733 1344
rect 1679 1276 1733 1310
rect 1679 1242 1691 1276
rect 1725 1242 1733 1276
rect 1679 1208 1733 1242
rect 1679 1174 1691 1208
rect 1725 1174 1733 1208
rect 1679 1050 1733 1174
rect 2055 1412 2111 1450
rect 2055 1378 2065 1412
rect 2099 1378 2111 1412
rect 2055 1344 2111 1378
rect 2055 1310 2065 1344
rect 2099 1310 2111 1344
rect 2055 1276 2111 1310
rect 2055 1242 2065 1276
rect 2099 1242 2111 1276
rect 2055 1208 2111 1242
rect 2055 1174 2065 1208
rect 2099 1174 2111 1208
rect 2055 1139 2111 1174
rect 2055 1105 2065 1139
rect 2099 1105 2111 1139
rect 2055 1050 2111 1105
rect 2141 1412 2199 1450
rect 2141 1378 2153 1412
rect 2187 1378 2199 1412
rect 2141 1344 2199 1378
rect 2141 1310 2153 1344
rect 2187 1310 2199 1344
rect 2141 1276 2199 1310
rect 2141 1242 2153 1276
rect 2187 1242 2199 1276
rect 2141 1208 2199 1242
rect 2141 1174 2153 1208
rect 2187 1174 2199 1208
rect 2141 1139 2199 1174
rect 2141 1105 2153 1139
rect 2187 1105 2199 1139
rect 2141 1050 2199 1105
rect 2229 1412 2287 1450
rect 2229 1378 2241 1412
rect 2275 1378 2287 1412
rect 2229 1344 2287 1378
rect 2229 1310 2241 1344
rect 2275 1310 2287 1344
rect 2229 1276 2287 1310
rect 2229 1242 2241 1276
rect 2275 1242 2287 1276
rect 2229 1208 2287 1242
rect 2229 1174 2241 1208
rect 2275 1174 2287 1208
rect 2229 1050 2287 1174
rect 2317 1412 2375 1450
rect 2317 1378 2329 1412
rect 2363 1378 2375 1412
rect 2317 1344 2375 1378
rect 2317 1310 2329 1344
rect 2363 1310 2375 1344
rect 2317 1276 2375 1310
rect 2317 1242 2329 1276
rect 2363 1242 2375 1276
rect 2317 1208 2375 1242
rect 2317 1174 2329 1208
rect 2363 1174 2375 1208
rect 2317 1139 2375 1174
rect 2317 1105 2329 1139
rect 2363 1105 2375 1139
rect 2317 1050 2375 1105
rect 2405 1412 2459 1450
rect 2405 1378 2417 1412
rect 2451 1378 2459 1412
rect 2405 1344 2459 1378
rect 2405 1310 2417 1344
rect 2451 1310 2459 1344
rect 2405 1276 2459 1310
rect 2405 1242 2417 1276
rect 2451 1242 2459 1276
rect 2405 1208 2459 1242
rect 2405 1174 2417 1208
rect 2451 1174 2459 1208
rect 2405 1050 2459 1174
rect 2781 1412 2837 1450
rect 2781 1378 2791 1412
rect 2825 1378 2837 1412
rect 2781 1344 2837 1378
rect 2781 1310 2791 1344
rect 2825 1310 2837 1344
rect 2781 1276 2837 1310
rect 2781 1242 2791 1276
rect 2825 1242 2837 1276
rect 2781 1208 2837 1242
rect 2781 1174 2791 1208
rect 2825 1174 2837 1208
rect 2781 1139 2837 1174
rect 2781 1105 2791 1139
rect 2825 1105 2837 1139
rect 2781 1050 2837 1105
rect 2867 1412 2925 1450
rect 2867 1378 2879 1412
rect 2913 1378 2925 1412
rect 2867 1344 2925 1378
rect 2867 1310 2879 1344
rect 2913 1310 2925 1344
rect 2867 1276 2925 1310
rect 2867 1242 2879 1276
rect 2913 1242 2925 1276
rect 2867 1208 2925 1242
rect 2867 1174 2879 1208
rect 2913 1174 2925 1208
rect 2867 1139 2925 1174
rect 2867 1105 2879 1139
rect 2913 1105 2925 1139
rect 2867 1050 2925 1105
rect 2955 1412 3013 1450
rect 2955 1378 2967 1412
rect 3001 1378 3013 1412
rect 2955 1344 3013 1378
rect 2955 1310 2967 1344
rect 3001 1310 3013 1344
rect 2955 1276 3013 1310
rect 2955 1242 2967 1276
rect 3001 1242 3013 1276
rect 2955 1208 3013 1242
rect 2955 1174 2967 1208
rect 3001 1174 3013 1208
rect 2955 1050 3013 1174
rect 3043 1412 3101 1450
rect 3043 1378 3055 1412
rect 3089 1378 3101 1412
rect 3043 1344 3101 1378
rect 3043 1310 3055 1344
rect 3089 1310 3101 1344
rect 3043 1276 3101 1310
rect 3043 1242 3055 1276
rect 3089 1242 3101 1276
rect 3043 1208 3101 1242
rect 3043 1174 3055 1208
rect 3089 1174 3101 1208
rect 3043 1139 3101 1174
rect 3043 1105 3055 1139
rect 3089 1105 3101 1139
rect 3043 1050 3101 1105
rect 3131 1412 3189 1450
rect 3131 1378 3143 1412
rect 3177 1378 3189 1412
rect 3131 1344 3189 1378
rect 3131 1310 3143 1344
rect 3177 1310 3189 1344
rect 3131 1276 3189 1310
rect 3131 1242 3143 1276
rect 3177 1242 3189 1276
rect 3131 1208 3189 1242
rect 3131 1174 3143 1208
rect 3177 1174 3189 1208
rect 3131 1050 3189 1174
rect 3219 1412 3277 1450
rect 3219 1378 3231 1412
rect 3265 1378 3277 1412
rect 3219 1344 3277 1378
rect 3219 1310 3231 1344
rect 3265 1310 3277 1344
rect 3219 1276 3277 1310
rect 3219 1242 3231 1276
rect 3265 1242 3277 1276
rect 3219 1208 3277 1242
rect 3219 1174 3231 1208
rect 3265 1174 3277 1208
rect 3219 1139 3277 1174
rect 3219 1105 3231 1139
rect 3265 1105 3277 1139
rect 3219 1050 3277 1105
rect 3307 1412 3361 1450
rect 3307 1378 3319 1412
rect 3353 1378 3361 1412
rect 3307 1344 3361 1378
rect 3307 1310 3319 1344
rect 3353 1310 3361 1344
rect 3307 1276 3361 1310
rect 3307 1242 3319 1276
rect 3353 1242 3361 1276
rect 3307 1208 3361 1242
rect 3307 1174 3319 1208
rect 3353 1174 3361 1208
rect 3307 1050 3361 1174
rect 3743 1412 3799 1450
rect 3743 1378 3753 1412
rect 3787 1378 3799 1412
rect 3743 1344 3799 1378
rect 3743 1310 3753 1344
rect 3787 1310 3799 1344
rect 3743 1276 3799 1310
rect 3743 1242 3753 1276
rect 3787 1242 3799 1276
rect 3743 1208 3799 1242
rect 3743 1174 3753 1208
rect 3787 1174 3799 1208
rect 3743 1139 3799 1174
rect 3743 1105 3753 1139
rect 3787 1105 3799 1139
rect 3743 1050 3799 1105
rect 3829 1412 3887 1450
rect 3829 1378 3841 1412
rect 3875 1378 3887 1412
rect 3829 1344 3887 1378
rect 3829 1310 3841 1344
rect 3875 1310 3887 1344
rect 3829 1276 3887 1310
rect 3829 1242 3841 1276
rect 3875 1242 3887 1276
rect 3829 1208 3887 1242
rect 3829 1174 3841 1208
rect 3875 1174 3887 1208
rect 3829 1139 3887 1174
rect 3829 1105 3841 1139
rect 3875 1105 3887 1139
rect 3829 1050 3887 1105
rect 3917 1412 3975 1450
rect 3917 1378 3929 1412
rect 3963 1378 3975 1412
rect 3917 1344 3975 1378
rect 3917 1310 3929 1344
rect 3963 1310 3975 1344
rect 3917 1276 3975 1310
rect 3917 1242 3929 1276
rect 3963 1242 3975 1276
rect 3917 1208 3975 1242
rect 3917 1174 3929 1208
rect 3963 1174 3975 1208
rect 3917 1050 3975 1174
rect 4005 1412 4063 1450
rect 4005 1378 4017 1412
rect 4051 1378 4063 1412
rect 4005 1344 4063 1378
rect 4005 1310 4017 1344
rect 4051 1310 4063 1344
rect 4005 1276 4063 1310
rect 4005 1242 4017 1276
rect 4051 1242 4063 1276
rect 4005 1208 4063 1242
rect 4005 1174 4017 1208
rect 4051 1174 4063 1208
rect 4005 1139 4063 1174
rect 4005 1105 4017 1139
rect 4051 1105 4063 1139
rect 4005 1050 4063 1105
rect 4093 1412 4151 1450
rect 4093 1378 4105 1412
rect 4139 1378 4151 1412
rect 4093 1344 4151 1378
rect 4093 1310 4105 1344
rect 4139 1310 4151 1344
rect 4093 1276 4151 1310
rect 4093 1242 4105 1276
rect 4139 1242 4151 1276
rect 4093 1208 4151 1242
rect 4093 1174 4105 1208
rect 4139 1174 4151 1208
rect 4093 1050 4151 1174
rect 4181 1412 4239 1450
rect 4181 1378 4193 1412
rect 4227 1378 4239 1412
rect 4181 1344 4239 1378
rect 4181 1310 4193 1344
rect 4227 1310 4239 1344
rect 4181 1276 4239 1310
rect 4181 1242 4193 1276
rect 4227 1242 4239 1276
rect 4181 1208 4239 1242
rect 4181 1174 4193 1208
rect 4227 1174 4239 1208
rect 4181 1139 4239 1174
rect 4181 1105 4193 1139
rect 4227 1105 4239 1139
rect 4181 1050 4239 1105
rect 4269 1412 4323 1450
rect 4269 1378 4281 1412
rect 4315 1378 4323 1412
rect 4269 1344 4323 1378
rect 4269 1310 4281 1344
rect 4315 1310 4323 1344
rect 4269 1276 4323 1310
rect 4269 1242 4281 1276
rect 4315 1242 4323 1276
rect 4269 1208 4323 1242
rect 4269 1174 4281 1208
rect 4315 1174 4323 1208
rect 4269 1050 4323 1174
rect 4645 1412 4701 1450
rect 4645 1378 4655 1412
rect 4689 1378 4701 1412
rect 4645 1344 4701 1378
rect 4645 1310 4655 1344
rect 4689 1310 4701 1344
rect 4645 1276 4701 1310
rect 4645 1242 4655 1276
rect 4689 1242 4701 1276
rect 4645 1208 4701 1242
rect 4645 1174 4655 1208
rect 4689 1174 4701 1208
rect 4645 1139 4701 1174
rect 4645 1105 4655 1139
rect 4689 1105 4701 1139
rect 4645 1050 4701 1105
rect 4731 1412 4789 1450
rect 4731 1378 4743 1412
rect 4777 1378 4789 1412
rect 4731 1344 4789 1378
rect 4731 1310 4743 1344
rect 4777 1310 4789 1344
rect 4731 1276 4789 1310
rect 4731 1242 4743 1276
rect 4777 1242 4789 1276
rect 4731 1208 4789 1242
rect 4731 1174 4743 1208
rect 4777 1174 4789 1208
rect 4731 1139 4789 1174
rect 4731 1105 4743 1139
rect 4777 1105 4789 1139
rect 4731 1050 4789 1105
rect 4819 1412 4877 1450
rect 4819 1378 4831 1412
rect 4865 1378 4877 1412
rect 4819 1344 4877 1378
rect 4819 1310 4831 1344
rect 4865 1310 4877 1344
rect 4819 1276 4877 1310
rect 4819 1242 4831 1276
rect 4865 1242 4877 1276
rect 4819 1208 4877 1242
rect 4819 1174 4831 1208
rect 4865 1174 4877 1208
rect 4819 1050 4877 1174
rect 4907 1412 4965 1450
rect 4907 1378 4919 1412
rect 4953 1378 4965 1412
rect 4907 1344 4965 1378
rect 4907 1310 4919 1344
rect 4953 1310 4965 1344
rect 4907 1276 4965 1310
rect 4907 1242 4919 1276
rect 4953 1242 4965 1276
rect 4907 1208 4965 1242
rect 4907 1174 4919 1208
rect 4953 1174 4965 1208
rect 4907 1139 4965 1174
rect 4907 1105 4919 1139
rect 4953 1105 4965 1139
rect 4907 1050 4965 1105
rect 4995 1412 5049 1450
rect 4995 1378 5007 1412
rect 5041 1378 5049 1412
rect 4995 1344 5049 1378
rect 4995 1310 5007 1344
rect 5041 1310 5049 1344
rect 4995 1276 5049 1310
rect 4995 1242 5007 1276
rect 5041 1242 5049 1276
rect 4995 1208 5049 1242
rect 4995 1174 5007 1208
rect 5041 1174 5049 1208
rect 4995 1050 5049 1174
rect 5371 1412 5427 1450
rect 5371 1378 5381 1412
rect 5415 1378 5427 1412
rect 5371 1344 5427 1378
rect 5371 1310 5381 1344
rect 5415 1310 5427 1344
rect 5371 1276 5427 1310
rect 5371 1242 5381 1276
rect 5415 1242 5427 1276
rect 5371 1208 5427 1242
rect 5371 1174 5381 1208
rect 5415 1174 5427 1208
rect 5371 1139 5427 1174
rect 5371 1105 5381 1139
rect 5415 1105 5427 1139
rect 5371 1050 5427 1105
rect 5457 1412 5515 1450
rect 5457 1378 5469 1412
rect 5503 1378 5515 1412
rect 5457 1344 5515 1378
rect 5457 1310 5469 1344
rect 5503 1310 5515 1344
rect 5457 1276 5515 1310
rect 5457 1242 5469 1276
rect 5503 1242 5515 1276
rect 5457 1208 5515 1242
rect 5457 1174 5469 1208
rect 5503 1174 5515 1208
rect 5457 1139 5515 1174
rect 5457 1105 5469 1139
rect 5503 1105 5515 1139
rect 5457 1050 5515 1105
rect 5545 1412 5603 1450
rect 5545 1378 5557 1412
rect 5591 1378 5603 1412
rect 5545 1344 5603 1378
rect 5545 1310 5557 1344
rect 5591 1310 5603 1344
rect 5545 1276 5603 1310
rect 5545 1242 5557 1276
rect 5591 1242 5603 1276
rect 5545 1208 5603 1242
rect 5545 1174 5557 1208
rect 5591 1174 5603 1208
rect 5545 1050 5603 1174
rect 5633 1412 5691 1450
rect 5633 1378 5645 1412
rect 5679 1378 5691 1412
rect 5633 1344 5691 1378
rect 5633 1310 5645 1344
rect 5679 1310 5691 1344
rect 5633 1276 5691 1310
rect 5633 1242 5645 1276
rect 5679 1242 5691 1276
rect 5633 1208 5691 1242
rect 5633 1174 5645 1208
rect 5679 1174 5691 1208
rect 5633 1139 5691 1174
rect 5633 1105 5645 1139
rect 5679 1105 5691 1139
rect 5633 1050 5691 1105
rect 5721 1412 5779 1450
rect 5721 1378 5733 1412
rect 5767 1378 5779 1412
rect 5721 1344 5779 1378
rect 5721 1310 5733 1344
rect 5767 1310 5779 1344
rect 5721 1276 5779 1310
rect 5721 1242 5733 1276
rect 5767 1242 5779 1276
rect 5721 1208 5779 1242
rect 5721 1174 5733 1208
rect 5767 1174 5779 1208
rect 5721 1050 5779 1174
rect 5809 1412 5867 1450
rect 5809 1378 5821 1412
rect 5855 1378 5867 1412
rect 5809 1344 5867 1378
rect 5809 1310 5821 1344
rect 5855 1310 5867 1344
rect 5809 1276 5867 1310
rect 5809 1242 5821 1276
rect 5855 1242 5867 1276
rect 5809 1208 5867 1242
rect 5809 1174 5821 1208
rect 5855 1174 5867 1208
rect 5809 1139 5867 1174
rect 5809 1105 5821 1139
rect 5855 1105 5867 1139
rect 5809 1050 5867 1105
rect 5897 1412 5951 1450
rect 5897 1378 5909 1412
rect 5943 1378 5951 1412
rect 5897 1344 5951 1378
rect 5897 1310 5909 1344
rect 5943 1310 5951 1344
rect 5897 1276 5951 1310
rect 5897 1242 5909 1276
rect 5943 1242 5951 1276
rect 5897 1208 5951 1242
rect 5897 1174 5909 1208
rect 5943 1174 5951 1208
rect 5897 1050 5951 1174
rect 6333 1412 6389 1450
rect 6333 1378 6343 1412
rect 6377 1378 6389 1412
rect 6333 1344 6389 1378
rect 6333 1310 6343 1344
rect 6377 1310 6389 1344
rect 6333 1276 6389 1310
rect 6333 1242 6343 1276
rect 6377 1242 6389 1276
rect 6333 1208 6389 1242
rect 6333 1174 6343 1208
rect 6377 1174 6389 1208
rect 6333 1139 6389 1174
rect 6333 1105 6343 1139
rect 6377 1105 6389 1139
rect 6333 1050 6389 1105
rect 6419 1412 6477 1450
rect 6419 1378 6431 1412
rect 6465 1378 6477 1412
rect 6419 1344 6477 1378
rect 6419 1310 6431 1344
rect 6465 1310 6477 1344
rect 6419 1276 6477 1310
rect 6419 1242 6431 1276
rect 6465 1242 6477 1276
rect 6419 1208 6477 1242
rect 6419 1174 6431 1208
rect 6465 1174 6477 1208
rect 6419 1139 6477 1174
rect 6419 1105 6431 1139
rect 6465 1105 6477 1139
rect 6419 1050 6477 1105
rect 6507 1412 6565 1450
rect 6507 1378 6519 1412
rect 6553 1378 6565 1412
rect 6507 1344 6565 1378
rect 6507 1310 6519 1344
rect 6553 1310 6565 1344
rect 6507 1276 6565 1310
rect 6507 1242 6519 1276
rect 6553 1242 6565 1276
rect 6507 1208 6565 1242
rect 6507 1174 6519 1208
rect 6553 1174 6565 1208
rect 6507 1050 6565 1174
rect 6595 1412 6653 1450
rect 6595 1378 6607 1412
rect 6641 1378 6653 1412
rect 6595 1344 6653 1378
rect 6595 1310 6607 1344
rect 6641 1310 6653 1344
rect 6595 1276 6653 1310
rect 6595 1242 6607 1276
rect 6641 1242 6653 1276
rect 6595 1208 6653 1242
rect 6595 1174 6607 1208
rect 6641 1174 6653 1208
rect 6595 1139 6653 1174
rect 6595 1105 6607 1139
rect 6641 1105 6653 1139
rect 6595 1050 6653 1105
rect 6683 1412 6741 1450
rect 6683 1378 6695 1412
rect 6729 1378 6741 1412
rect 6683 1344 6741 1378
rect 6683 1310 6695 1344
rect 6729 1310 6741 1344
rect 6683 1276 6741 1310
rect 6683 1242 6695 1276
rect 6729 1242 6741 1276
rect 6683 1208 6741 1242
rect 6683 1174 6695 1208
rect 6729 1174 6741 1208
rect 6683 1050 6741 1174
rect 6771 1412 6829 1450
rect 6771 1378 6783 1412
rect 6817 1378 6829 1412
rect 6771 1344 6829 1378
rect 6771 1310 6783 1344
rect 6817 1310 6829 1344
rect 6771 1276 6829 1310
rect 6771 1242 6783 1276
rect 6817 1242 6829 1276
rect 6771 1208 6829 1242
rect 6771 1174 6783 1208
rect 6817 1174 6829 1208
rect 6771 1139 6829 1174
rect 6771 1105 6783 1139
rect 6817 1105 6829 1139
rect 6771 1050 6829 1105
rect 6859 1412 6913 1450
rect 6859 1378 6871 1412
rect 6905 1378 6913 1412
rect 6859 1344 6913 1378
rect 6859 1310 6871 1344
rect 6905 1310 6913 1344
rect 6859 1276 6913 1310
rect 6859 1242 6871 1276
rect 6905 1242 6913 1276
rect 6859 1208 6913 1242
rect 6859 1174 6871 1208
rect 6905 1174 6913 1208
rect 6859 1050 6913 1174
rect 7235 1412 7291 1450
rect 7235 1378 7245 1412
rect 7279 1378 7291 1412
rect 7235 1344 7291 1378
rect 7235 1310 7245 1344
rect 7279 1310 7291 1344
rect 7235 1276 7291 1310
rect 7235 1242 7245 1276
rect 7279 1242 7291 1276
rect 7235 1208 7291 1242
rect 7235 1174 7245 1208
rect 7279 1174 7291 1208
rect 7235 1139 7291 1174
rect 7235 1105 7245 1139
rect 7279 1105 7291 1139
rect 7235 1050 7291 1105
rect 7321 1412 7379 1450
rect 7321 1378 7333 1412
rect 7367 1378 7379 1412
rect 7321 1344 7379 1378
rect 7321 1310 7333 1344
rect 7367 1310 7379 1344
rect 7321 1276 7379 1310
rect 7321 1242 7333 1276
rect 7367 1242 7379 1276
rect 7321 1208 7379 1242
rect 7321 1174 7333 1208
rect 7367 1174 7379 1208
rect 7321 1139 7379 1174
rect 7321 1105 7333 1139
rect 7367 1105 7379 1139
rect 7321 1050 7379 1105
rect 7409 1412 7467 1450
rect 7409 1378 7421 1412
rect 7455 1378 7467 1412
rect 7409 1344 7467 1378
rect 7409 1310 7421 1344
rect 7455 1310 7467 1344
rect 7409 1276 7467 1310
rect 7409 1242 7421 1276
rect 7455 1242 7467 1276
rect 7409 1208 7467 1242
rect 7409 1174 7421 1208
rect 7455 1174 7467 1208
rect 7409 1050 7467 1174
rect 7497 1412 7555 1450
rect 7497 1378 7509 1412
rect 7543 1378 7555 1412
rect 7497 1344 7555 1378
rect 7497 1310 7509 1344
rect 7543 1310 7555 1344
rect 7497 1276 7555 1310
rect 7497 1242 7509 1276
rect 7543 1242 7555 1276
rect 7497 1208 7555 1242
rect 7497 1174 7509 1208
rect 7543 1174 7555 1208
rect 7497 1139 7555 1174
rect 7497 1105 7509 1139
rect 7543 1105 7555 1139
rect 7497 1050 7555 1105
rect 7585 1412 7639 1450
rect 7585 1378 7597 1412
rect 7631 1378 7639 1412
rect 7585 1344 7639 1378
rect 7585 1310 7597 1344
rect 7631 1310 7639 1344
rect 7585 1276 7639 1310
rect 7585 1242 7597 1276
rect 7631 1242 7639 1276
rect 7585 1208 7639 1242
rect 7585 1174 7597 1208
rect 7631 1174 7639 1208
rect 7585 1050 7639 1174
rect 7961 1412 8017 1450
rect 7961 1378 7971 1412
rect 8005 1378 8017 1412
rect 7961 1344 8017 1378
rect 7961 1310 7971 1344
rect 8005 1310 8017 1344
rect 7961 1276 8017 1310
rect 7961 1242 7971 1276
rect 8005 1242 8017 1276
rect 7961 1208 8017 1242
rect 7961 1174 7971 1208
rect 8005 1174 8017 1208
rect 7961 1139 8017 1174
rect 7961 1105 7971 1139
rect 8005 1105 8017 1139
rect 7961 1050 8017 1105
rect 8047 1412 8105 1450
rect 8047 1378 8059 1412
rect 8093 1378 8105 1412
rect 8047 1344 8105 1378
rect 8047 1310 8059 1344
rect 8093 1310 8105 1344
rect 8047 1276 8105 1310
rect 8047 1242 8059 1276
rect 8093 1242 8105 1276
rect 8047 1208 8105 1242
rect 8047 1174 8059 1208
rect 8093 1174 8105 1208
rect 8047 1139 8105 1174
rect 8047 1105 8059 1139
rect 8093 1105 8105 1139
rect 8047 1050 8105 1105
rect 8135 1412 8193 1450
rect 8135 1378 8147 1412
rect 8181 1378 8193 1412
rect 8135 1344 8193 1378
rect 8135 1310 8147 1344
rect 8181 1310 8193 1344
rect 8135 1276 8193 1310
rect 8135 1242 8147 1276
rect 8181 1242 8193 1276
rect 8135 1208 8193 1242
rect 8135 1174 8147 1208
rect 8181 1174 8193 1208
rect 8135 1050 8193 1174
rect 8223 1412 8281 1450
rect 8223 1378 8235 1412
rect 8269 1378 8281 1412
rect 8223 1344 8281 1378
rect 8223 1310 8235 1344
rect 8269 1310 8281 1344
rect 8223 1276 8281 1310
rect 8223 1242 8235 1276
rect 8269 1242 8281 1276
rect 8223 1208 8281 1242
rect 8223 1174 8235 1208
rect 8269 1174 8281 1208
rect 8223 1139 8281 1174
rect 8223 1105 8235 1139
rect 8269 1105 8281 1139
rect 8223 1050 8281 1105
rect 8311 1412 8369 1450
rect 8311 1378 8323 1412
rect 8357 1378 8369 1412
rect 8311 1344 8369 1378
rect 8311 1310 8323 1344
rect 8357 1310 8369 1344
rect 8311 1276 8369 1310
rect 8311 1242 8323 1276
rect 8357 1242 8369 1276
rect 8311 1208 8369 1242
rect 8311 1174 8323 1208
rect 8357 1174 8369 1208
rect 8311 1050 8369 1174
rect 8399 1412 8457 1450
rect 8399 1378 8411 1412
rect 8445 1378 8457 1412
rect 8399 1344 8457 1378
rect 8399 1310 8411 1344
rect 8445 1310 8457 1344
rect 8399 1276 8457 1310
rect 8399 1242 8411 1276
rect 8445 1242 8457 1276
rect 8399 1208 8457 1242
rect 8399 1174 8411 1208
rect 8445 1174 8457 1208
rect 8399 1139 8457 1174
rect 8399 1105 8411 1139
rect 8445 1105 8457 1139
rect 8399 1050 8457 1105
rect 8487 1412 8541 1450
rect 8487 1378 8499 1412
rect 8533 1378 8541 1412
rect 8487 1344 8541 1378
rect 8487 1310 8499 1344
rect 8533 1310 8541 1344
rect 8487 1276 8541 1310
rect 8487 1242 8499 1276
rect 8533 1242 8541 1276
rect 8487 1208 8541 1242
rect 8487 1174 8499 1208
rect 8533 1174 8541 1208
rect 8487 1050 8541 1174
rect 8923 1412 8979 1450
rect 8923 1378 8933 1412
rect 8967 1378 8979 1412
rect 8923 1344 8979 1378
rect 8923 1310 8933 1344
rect 8967 1310 8979 1344
rect 8923 1276 8979 1310
rect 8923 1242 8933 1276
rect 8967 1242 8979 1276
rect 8923 1208 8979 1242
rect 8923 1174 8933 1208
rect 8967 1174 8979 1208
rect 8923 1139 8979 1174
rect 8923 1105 8933 1139
rect 8967 1105 8979 1139
rect 8923 1050 8979 1105
rect 9009 1412 9067 1450
rect 9009 1378 9021 1412
rect 9055 1378 9067 1412
rect 9009 1344 9067 1378
rect 9009 1310 9021 1344
rect 9055 1310 9067 1344
rect 9009 1276 9067 1310
rect 9009 1242 9021 1276
rect 9055 1242 9067 1276
rect 9009 1208 9067 1242
rect 9009 1174 9021 1208
rect 9055 1174 9067 1208
rect 9009 1139 9067 1174
rect 9009 1105 9021 1139
rect 9055 1105 9067 1139
rect 9009 1050 9067 1105
rect 9097 1412 9155 1450
rect 9097 1378 9109 1412
rect 9143 1378 9155 1412
rect 9097 1344 9155 1378
rect 9097 1310 9109 1344
rect 9143 1310 9155 1344
rect 9097 1276 9155 1310
rect 9097 1242 9109 1276
rect 9143 1242 9155 1276
rect 9097 1208 9155 1242
rect 9097 1174 9109 1208
rect 9143 1174 9155 1208
rect 9097 1050 9155 1174
rect 9185 1412 9243 1450
rect 9185 1378 9197 1412
rect 9231 1378 9243 1412
rect 9185 1344 9243 1378
rect 9185 1310 9197 1344
rect 9231 1310 9243 1344
rect 9185 1276 9243 1310
rect 9185 1242 9197 1276
rect 9231 1242 9243 1276
rect 9185 1208 9243 1242
rect 9185 1174 9197 1208
rect 9231 1174 9243 1208
rect 9185 1139 9243 1174
rect 9185 1105 9197 1139
rect 9231 1105 9243 1139
rect 9185 1050 9243 1105
rect 9273 1412 9331 1450
rect 9273 1378 9285 1412
rect 9319 1378 9331 1412
rect 9273 1344 9331 1378
rect 9273 1310 9285 1344
rect 9319 1310 9331 1344
rect 9273 1276 9331 1310
rect 9273 1242 9285 1276
rect 9319 1242 9331 1276
rect 9273 1208 9331 1242
rect 9273 1174 9285 1208
rect 9319 1174 9331 1208
rect 9273 1050 9331 1174
rect 9361 1412 9419 1450
rect 9361 1378 9373 1412
rect 9407 1378 9419 1412
rect 9361 1344 9419 1378
rect 9361 1310 9373 1344
rect 9407 1310 9419 1344
rect 9361 1276 9419 1310
rect 9361 1242 9373 1276
rect 9407 1242 9419 1276
rect 9361 1208 9419 1242
rect 9361 1174 9373 1208
rect 9407 1174 9419 1208
rect 9361 1139 9419 1174
rect 9361 1105 9373 1139
rect 9407 1105 9419 1139
rect 9361 1050 9419 1105
rect 9449 1412 9503 1450
rect 9449 1378 9461 1412
rect 9495 1378 9503 1412
rect 9449 1344 9503 1378
rect 9449 1310 9461 1344
rect 9495 1310 9503 1344
rect 9449 1276 9503 1310
rect 9449 1242 9461 1276
rect 9495 1242 9503 1276
rect 9449 1208 9503 1242
rect 9449 1174 9461 1208
rect 9495 1174 9503 1208
rect 9449 1050 9503 1174
rect 9825 1412 9881 1450
rect 9825 1378 9835 1412
rect 9869 1378 9881 1412
rect 9825 1344 9881 1378
rect 9825 1310 9835 1344
rect 9869 1310 9881 1344
rect 9825 1276 9881 1310
rect 9825 1242 9835 1276
rect 9869 1242 9881 1276
rect 9825 1208 9881 1242
rect 9825 1174 9835 1208
rect 9869 1174 9881 1208
rect 9825 1139 9881 1174
rect 9825 1105 9835 1139
rect 9869 1105 9881 1139
rect 9825 1050 9881 1105
rect 9911 1412 9969 1450
rect 9911 1378 9923 1412
rect 9957 1378 9969 1412
rect 9911 1344 9969 1378
rect 9911 1310 9923 1344
rect 9957 1310 9969 1344
rect 9911 1276 9969 1310
rect 9911 1242 9923 1276
rect 9957 1242 9969 1276
rect 9911 1208 9969 1242
rect 9911 1174 9923 1208
rect 9957 1174 9969 1208
rect 9911 1139 9969 1174
rect 9911 1105 9923 1139
rect 9957 1105 9969 1139
rect 9911 1050 9969 1105
rect 9999 1412 10057 1450
rect 9999 1378 10011 1412
rect 10045 1378 10057 1412
rect 9999 1344 10057 1378
rect 9999 1310 10011 1344
rect 10045 1310 10057 1344
rect 9999 1276 10057 1310
rect 9999 1242 10011 1276
rect 10045 1242 10057 1276
rect 9999 1208 10057 1242
rect 9999 1174 10011 1208
rect 10045 1174 10057 1208
rect 9999 1050 10057 1174
rect 10087 1412 10145 1450
rect 10087 1378 10099 1412
rect 10133 1378 10145 1412
rect 10087 1344 10145 1378
rect 10087 1310 10099 1344
rect 10133 1310 10145 1344
rect 10087 1276 10145 1310
rect 10087 1242 10099 1276
rect 10133 1242 10145 1276
rect 10087 1208 10145 1242
rect 10087 1174 10099 1208
rect 10133 1174 10145 1208
rect 10087 1139 10145 1174
rect 10087 1105 10099 1139
rect 10133 1105 10145 1139
rect 10087 1050 10145 1105
rect 10175 1412 10229 1450
rect 10175 1378 10187 1412
rect 10221 1378 10229 1412
rect 10175 1344 10229 1378
rect 10175 1310 10187 1344
rect 10221 1310 10229 1344
rect 10175 1276 10229 1310
rect 10175 1242 10187 1276
rect 10221 1242 10229 1276
rect 10175 1208 10229 1242
rect 10175 1174 10187 1208
rect 10221 1174 10229 1208
rect 10175 1050 10229 1174
rect 10551 1412 10607 1450
rect 10551 1378 10561 1412
rect 10595 1378 10607 1412
rect 10551 1344 10607 1378
rect 10551 1310 10561 1344
rect 10595 1310 10607 1344
rect 10551 1276 10607 1310
rect 10551 1242 10561 1276
rect 10595 1242 10607 1276
rect 10551 1208 10607 1242
rect 10551 1174 10561 1208
rect 10595 1174 10607 1208
rect 10551 1139 10607 1174
rect 10551 1105 10561 1139
rect 10595 1105 10607 1139
rect 10551 1050 10607 1105
rect 10637 1412 10695 1450
rect 10637 1378 10649 1412
rect 10683 1378 10695 1412
rect 10637 1344 10695 1378
rect 10637 1310 10649 1344
rect 10683 1310 10695 1344
rect 10637 1276 10695 1310
rect 10637 1242 10649 1276
rect 10683 1242 10695 1276
rect 10637 1208 10695 1242
rect 10637 1174 10649 1208
rect 10683 1174 10695 1208
rect 10637 1139 10695 1174
rect 10637 1105 10649 1139
rect 10683 1105 10695 1139
rect 10637 1050 10695 1105
rect 10725 1412 10783 1450
rect 10725 1378 10737 1412
rect 10771 1378 10783 1412
rect 10725 1344 10783 1378
rect 10725 1310 10737 1344
rect 10771 1310 10783 1344
rect 10725 1276 10783 1310
rect 10725 1242 10737 1276
rect 10771 1242 10783 1276
rect 10725 1208 10783 1242
rect 10725 1174 10737 1208
rect 10771 1174 10783 1208
rect 10725 1050 10783 1174
rect 10813 1412 10871 1450
rect 10813 1378 10825 1412
rect 10859 1378 10871 1412
rect 10813 1344 10871 1378
rect 10813 1310 10825 1344
rect 10859 1310 10871 1344
rect 10813 1276 10871 1310
rect 10813 1242 10825 1276
rect 10859 1242 10871 1276
rect 10813 1208 10871 1242
rect 10813 1174 10825 1208
rect 10859 1174 10871 1208
rect 10813 1139 10871 1174
rect 10813 1105 10825 1139
rect 10859 1105 10871 1139
rect 10813 1050 10871 1105
rect 10901 1412 10959 1450
rect 10901 1378 10913 1412
rect 10947 1378 10959 1412
rect 10901 1344 10959 1378
rect 10901 1310 10913 1344
rect 10947 1310 10959 1344
rect 10901 1276 10959 1310
rect 10901 1242 10913 1276
rect 10947 1242 10959 1276
rect 10901 1208 10959 1242
rect 10901 1174 10913 1208
rect 10947 1174 10959 1208
rect 10901 1050 10959 1174
rect 10989 1412 11047 1450
rect 10989 1378 11001 1412
rect 11035 1378 11047 1412
rect 10989 1344 11047 1378
rect 10989 1310 11001 1344
rect 11035 1310 11047 1344
rect 10989 1276 11047 1310
rect 10989 1242 11001 1276
rect 11035 1242 11047 1276
rect 10989 1208 11047 1242
rect 10989 1174 11001 1208
rect 11035 1174 11047 1208
rect 10989 1139 11047 1174
rect 10989 1105 11001 1139
rect 11035 1105 11047 1139
rect 10989 1050 11047 1105
rect 11077 1412 11131 1450
rect 11077 1378 11089 1412
rect 11123 1378 11131 1412
rect 11077 1344 11131 1378
rect 11077 1310 11089 1344
rect 11123 1310 11131 1344
rect 11077 1276 11131 1310
rect 11077 1242 11089 1276
rect 11123 1242 11131 1276
rect 11077 1208 11131 1242
rect 11077 1174 11089 1208
rect 11123 1174 11131 1208
rect 11077 1050 11131 1174
rect 11513 1412 11569 1450
rect 11513 1378 11523 1412
rect 11557 1378 11569 1412
rect 11513 1344 11569 1378
rect 11513 1310 11523 1344
rect 11557 1310 11569 1344
rect 11513 1276 11569 1310
rect 11513 1242 11523 1276
rect 11557 1242 11569 1276
rect 11513 1208 11569 1242
rect 11513 1174 11523 1208
rect 11557 1174 11569 1208
rect 11513 1139 11569 1174
rect 11513 1105 11523 1139
rect 11557 1105 11569 1139
rect 11513 1050 11569 1105
rect 11599 1412 11657 1450
rect 11599 1378 11611 1412
rect 11645 1378 11657 1412
rect 11599 1344 11657 1378
rect 11599 1310 11611 1344
rect 11645 1310 11657 1344
rect 11599 1276 11657 1310
rect 11599 1242 11611 1276
rect 11645 1242 11657 1276
rect 11599 1208 11657 1242
rect 11599 1174 11611 1208
rect 11645 1174 11657 1208
rect 11599 1139 11657 1174
rect 11599 1105 11611 1139
rect 11645 1105 11657 1139
rect 11599 1050 11657 1105
rect 11687 1412 11745 1450
rect 11687 1378 11699 1412
rect 11733 1378 11745 1412
rect 11687 1344 11745 1378
rect 11687 1310 11699 1344
rect 11733 1310 11745 1344
rect 11687 1276 11745 1310
rect 11687 1242 11699 1276
rect 11733 1242 11745 1276
rect 11687 1208 11745 1242
rect 11687 1174 11699 1208
rect 11733 1174 11745 1208
rect 11687 1050 11745 1174
rect 11775 1412 11833 1450
rect 11775 1378 11787 1412
rect 11821 1378 11833 1412
rect 11775 1344 11833 1378
rect 11775 1310 11787 1344
rect 11821 1310 11833 1344
rect 11775 1276 11833 1310
rect 11775 1242 11787 1276
rect 11821 1242 11833 1276
rect 11775 1208 11833 1242
rect 11775 1174 11787 1208
rect 11821 1174 11833 1208
rect 11775 1139 11833 1174
rect 11775 1105 11787 1139
rect 11821 1105 11833 1139
rect 11775 1050 11833 1105
rect 11863 1412 11921 1450
rect 11863 1378 11875 1412
rect 11909 1378 11921 1412
rect 11863 1344 11921 1378
rect 11863 1310 11875 1344
rect 11909 1310 11921 1344
rect 11863 1276 11921 1310
rect 11863 1242 11875 1276
rect 11909 1242 11921 1276
rect 11863 1208 11921 1242
rect 11863 1174 11875 1208
rect 11909 1174 11921 1208
rect 11863 1050 11921 1174
rect 11951 1412 12009 1450
rect 11951 1378 11963 1412
rect 11997 1378 12009 1412
rect 11951 1344 12009 1378
rect 11951 1310 11963 1344
rect 11997 1310 12009 1344
rect 11951 1276 12009 1310
rect 11951 1242 11963 1276
rect 11997 1242 12009 1276
rect 11951 1208 12009 1242
rect 11951 1174 11963 1208
rect 11997 1174 12009 1208
rect 11951 1139 12009 1174
rect 11951 1105 11963 1139
rect 11997 1105 12009 1139
rect 11951 1050 12009 1105
rect 12039 1412 12093 1450
rect 12039 1378 12051 1412
rect 12085 1378 12093 1412
rect 12039 1344 12093 1378
rect 12039 1310 12051 1344
rect 12085 1310 12093 1344
rect 12039 1276 12093 1310
rect 12039 1242 12051 1276
rect 12085 1242 12093 1276
rect 12039 1208 12093 1242
rect 12039 1174 12051 1208
rect 12085 1174 12093 1208
rect 12039 1050 12093 1174
rect 12415 1412 12471 1450
rect 12415 1378 12425 1412
rect 12459 1378 12471 1412
rect 12415 1344 12471 1378
rect 12415 1310 12425 1344
rect 12459 1310 12471 1344
rect 12415 1276 12471 1310
rect 12415 1242 12425 1276
rect 12459 1242 12471 1276
rect 12415 1208 12471 1242
rect 12415 1174 12425 1208
rect 12459 1174 12471 1208
rect 12415 1139 12471 1174
rect 12415 1105 12425 1139
rect 12459 1105 12471 1139
rect 12415 1050 12471 1105
rect 12501 1412 12559 1450
rect 12501 1378 12513 1412
rect 12547 1378 12559 1412
rect 12501 1344 12559 1378
rect 12501 1310 12513 1344
rect 12547 1310 12559 1344
rect 12501 1276 12559 1310
rect 12501 1242 12513 1276
rect 12547 1242 12559 1276
rect 12501 1208 12559 1242
rect 12501 1174 12513 1208
rect 12547 1174 12559 1208
rect 12501 1139 12559 1174
rect 12501 1105 12513 1139
rect 12547 1105 12559 1139
rect 12501 1050 12559 1105
rect 12589 1412 12647 1450
rect 12589 1378 12601 1412
rect 12635 1378 12647 1412
rect 12589 1344 12647 1378
rect 12589 1310 12601 1344
rect 12635 1310 12647 1344
rect 12589 1276 12647 1310
rect 12589 1242 12601 1276
rect 12635 1242 12647 1276
rect 12589 1208 12647 1242
rect 12589 1174 12601 1208
rect 12635 1174 12647 1208
rect 12589 1050 12647 1174
rect 12677 1412 12735 1450
rect 12677 1378 12689 1412
rect 12723 1378 12735 1412
rect 12677 1344 12735 1378
rect 12677 1310 12689 1344
rect 12723 1310 12735 1344
rect 12677 1276 12735 1310
rect 12677 1242 12689 1276
rect 12723 1242 12735 1276
rect 12677 1208 12735 1242
rect 12677 1174 12689 1208
rect 12723 1174 12735 1208
rect 12677 1139 12735 1174
rect 12677 1105 12689 1139
rect 12723 1105 12735 1139
rect 12677 1050 12735 1105
rect 12765 1412 12819 1450
rect 12765 1378 12777 1412
rect 12811 1378 12819 1412
rect 12765 1344 12819 1378
rect 12765 1310 12777 1344
rect 12811 1310 12819 1344
rect 12765 1276 12819 1310
rect 12765 1242 12777 1276
rect 12811 1242 12819 1276
rect 12765 1208 12819 1242
rect 12765 1174 12777 1208
rect 12811 1174 12819 1208
rect 12765 1050 12819 1174
rect 13141 1412 13197 1450
rect 13141 1378 13151 1412
rect 13185 1378 13197 1412
rect 13141 1344 13197 1378
rect 13141 1310 13151 1344
rect 13185 1310 13197 1344
rect 13141 1276 13197 1310
rect 13141 1242 13151 1276
rect 13185 1242 13197 1276
rect 13141 1208 13197 1242
rect 13141 1174 13151 1208
rect 13185 1174 13197 1208
rect 13141 1139 13197 1174
rect 13141 1105 13151 1139
rect 13185 1105 13197 1139
rect 13141 1050 13197 1105
rect 13227 1412 13285 1450
rect 13227 1378 13239 1412
rect 13273 1378 13285 1412
rect 13227 1344 13285 1378
rect 13227 1310 13239 1344
rect 13273 1310 13285 1344
rect 13227 1276 13285 1310
rect 13227 1242 13239 1276
rect 13273 1242 13285 1276
rect 13227 1208 13285 1242
rect 13227 1174 13239 1208
rect 13273 1174 13285 1208
rect 13227 1139 13285 1174
rect 13227 1105 13239 1139
rect 13273 1105 13285 1139
rect 13227 1050 13285 1105
rect 13315 1412 13373 1450
rect 13315 1378 13327 1412
rect 13361 1378 13373 1412
rect 13315 1344 13373 1378
rect 13315 1310 13327 1344
rect 13361 1310 13373 1344
rect 13315 1276 13373 1310
rect 13315 1242 13327 1276
rect 13361 1242 13373 1276
rect 13315 1208 13373 1242
rect 13315 1174 13327 1208
rect 13361 1174 13373 1208
rect 13315 1050 13373 1174
rect 13403 1412 13461 1450
rect 13403 1378 13415 1412
rect 13449 1378 13461 1412
rect 13403 1344 13461 1378
rect 13403 1310 13415 1344
rect 13449 1310 13461 1344
rect 13403 1276 13461 1310
rect 13403 1242 13415 1276
rect 13449 1242 13461 1276
rect 13403 1208 13461 1242
rect 13403 1174 13415 1208
rect 13449 1174 13461 1208
rect 13403 1139 13461 1174
rect 13403 1105 13415 1139
rect 13449 1105 13461 1139
rect 13403 1050 13461 1105
rect 13491 1412 13549 1450
rect 13491 1378 13503 1412
rect 13537 1378 13549 1412
rect 13491 1344 13549 1378
rect 13491 1310 13503 1344
rect 13537 1310 13549 1344
rect 13491 1276 13549 1310
rect 13491 1242 13503 1276
rect 13537 1242 13549 1276
rect 13491 1208 13549 1242
rect 13491 1174 13503 1208
rect 13537 1174 13549 1208
rect 13491 1050 13549 1174
rect 13579 1412 13637 1450
rect 13579 1378 13591 1412
rect 13625 1378 13637 1412
rect 13579 1344 13637 1378
rect 13579 1310 13591 1344
rect 13625 1310 13637 1344
rect 13579 1276 13637 1310
rect 13579 1242 13591 1276
rect 13625 1242 13637 1276
rect 13579 1208 13637 1242
rect 13579 1174 13591 1208
rect 13625 1174 13637 1208
rect 13579 1139 13637 1174
rect 13579 1105 13591 1139
rect 13625 1105 13637 1139
rect 13579 1050 13637 1105
rect 13667 1412 13721 1450
rect 13667 1378 13679 1412
rect 13713 1378 13721 1412
rect 13667 1344 13721 1378
rect 13667 1310 13679 1344
rect 13713 1310 13721 1344
rect 13667 1276 13721 1310
rect 13667 1242 13679 1276
rect 13713 1242 13721 1276
rect 13667 1208 13721 1242
rect 13667 1174 13679 1208
rect 13713 1174 13721 1208
rect 13667 1050 13721 1174
rect 14103 1412 14159 1450
rect 14103 1378 14113 1412
rect 14147 1378 14159 1412
rect 14103 1344 14159 1378
rect 14103 1310 14113 1344
rect 14147 1310 14159 1344
rect 14103 1276 14159 1310
rect 14103 1242 14113 1276
rect 14147 1242 14159 1276
rect 14103 1208 14159 1242
rect 14103 1174 14113 1208
rect 14147 1174 14159 1208
rect 14103 1139 14159 1174
rect 14103 1105 14113 1139
rect 14147 1105 14159 1139
rect 14103 1050 14159 1105
rect 14189 1412 14247 1450
rect 14189 1378 14201 1412
rect 14235 1378 14247 1412
rect 14189 1344 14247 1378
rect 14189 1310 14201 1344
rect 14235 1310 14247 1344
rect 14189 1276 14247 1310
rect 14189 1242 14201 1276
rect 14235 1242 14247 1276
rect 14189 1208 14247 1242
rect 14189 1174 14201 1208
rect 14235 1174 14247 1208
rect 14189 1139 14247 1174
rect 14189 1105 14201 1139
rect 14235 1105 14247 1139
rect 14189 1050 14247 1105
rect 14277 1412 14335 1450
rect 14277 1378 14289 1412
rect 14323 1378 14335 1412
rect 14277 1344 14335 1378
rect 14277 1310 14289 1344
rect 14323 1310 14335 1344
rect 14277 1276 14335 1310
rect 14277 1242 14289 1276
rect 14323 1242 14335 1276
rect 14277 1208 14335 1242
rect 14277 1174 14289 1208
rect 14323 1174 14335 1208
rect 14277 1050 14335 1174
rect 14365 1412 14423 1450
rect 14365 1378 14377 1412
rect 14411 1378 14423 1412
rect 14365 1344 14423 1378
rect 14365 1310 14377 1344
rect 14411 1310 14423 1344
rect 14365 1276 14423 1310
rect 14365 1242 14377 1276
rect 14411 1242 14423 1276
rect 14365 1208 14423 1242
rect 14365 1174 14377 1208
rect 14411 1174 14423 1208
rect 14365 1139 14423 1174
rect 14365 1105 14377 1139
rect 14411 1105 14423 1139
rect 14365 1050 14423 1105
rect 14453 1412 14511 1450
rect 14453 1378 14465 1412
rect 14499 1378 14511 1412
rect 14453 1344 14511 1378
rect 14453 1310 14465 1344
rect 14499 1310 14511 1344
rect 14453 1276 14511 1310
rect 14453 1242 14465 1276
rect 14499 1242 14511 1276
rect 14453 1208 14511 1242
rect 14453 1174 14465 1208
rect 14499 1174 14511 1208
rect 14453 1050 14511 1174
rect 14541 1412 14599 1450
rect 14541 1378 14553 1412
rect 14587 1378 14599 1412
rect 14541 1344 14599 1378
rect 14541 1310 14553 1344
rect 14587 1310 14599 1344
rect 14541 1276 14599 1310
rect 14541 1242 14553 1276
rect 14587 1242 14599 1276
rect 14541 1208 14599 1242
rect 14541 1174 14553 1208
rect 14587 1174 14599 1208
rect 14541 1139 14599 1174
rect 14541 1105 14553 1139
rect 14587 1105 14599 1139
rect 14541 1050 14599 1105
rect 14629 1412 14683 1450
rect 14629 1378 14641 1412
rect 14675 1378 14683 1412
rect 14629 1344 14683 1378
rect 14629 1310 14641 1344
rect 14675 1310 14683 1344
rect 14629 1276 14683 1310
rect 14629 1242 14641 1276
rect 14675 1242 14683 1276
rect 14629 1208 14683 1242
rect 14629 1174 14641 1208
rect 14675 1174 14683 1208
rect 14629 1050 14683 1174
rect 15005 1412 15061 1450
rect 15005 1378 15015 1412
rect 15049 1378 15061 1412
rect 15005 1344 15061 1378
rect 15005 1310 15015 1344
rect 15049 1310 15061 1344
rect 15005 1276 15061 1310
rect 15005 1242 15015 1276
rect 15049 1242 15061 1276
rect 15005 1208 15061 1242
rect 15005 1174 15015 1208
rect 15049 1174 15061 1208
rect 15005 1139 15061 1174
rect 15005 1105 15015 1139
rect 15049 1105 15061 1139
rect 15005 1050 15061 1105
rect 15091 1412 15149 1450
rect 15091 1378 15103 1412
rect 15137 1378 15149 1412
rect 15091 1344 15149 1378
rect 15091 1310 15103 1344
rect 15137 1310 15149 1344
rect 15091 1276 15149 1310
rect 15091 1242 15103 1276
rect 15137 1242 15149 1276
rect 15091 1208 15149 1242
rect 15091 1174 15103 1208
rect 15137 1174 15149 1208
rect 15091 1139 15149 1174
rect 15091 1105 15103 1139
rect 15137 1105 15149 1139
rect 15091 1050 15149 1105
rect 15179 1412 15237 1450
rect 15179 1378 15191 1412
rect 15225 1378 15237 1412
rect 15179 1344 15237 1378
rect 15179 1310 15191 1344
rect 15225 1310 15237 1344
rect 15179 1276 15237 1310
rect 15179 1242 15191 1276
rect 15225 1242 15237 1276
rect 15179 1208 15237 1242
rect 15179 1174 15191 1208
rect 15225 1174 15237 1208
rect 15179 1050 15237 1174
rect 15267 1412 15325 1450
rect 15267 1378 15279 1412
rect 15313 1378 15325 1412
rect 15267 1344 15325 1378
rect 15267 1310 15279 1344
rect 15313 1310 15325 1344
rect 15267 1276 15325 1310
rect 15267 1242 15279 1276
rect 15313 1242 15325 1276
rect 15267 1208 15325 1242
rect 15267 1174 15279 1208
rect 15313 1174 15325 1208
rect 15267 1139 15325 1174
rect 15267 1105 15279 1139
rect 15313 1105 15325 1139
rect 15267 1050 15325 1105
rect 15355 1412 15409 1450
rect 15355 1378 15367 1412
rect 15401 1378 15409 1412
rect 15355 1344 15409 1378
rect 15355 1310 15367 1344
rect 15401 1310 15409 1344
rect 15355 1276 15409 1310
rect 15355 1242 15367 1276
rect 15401 1242 15409 1276
rect 15355 1208 15409 1242
rect 15355 1174 15367 1208
rect 15401 1174 15409 1208
rect 15355 1050 15409 1174
rect 15671 1411 15727 1451
rect 15671 1377 15681 1411
rect 15715 1377 15727 1411
rect 15671 1343 15727 1377
rect 15671 1309 15681 1343
rect 15715 1309 15727 1343
rect 15671 1275 15727 1309
rect 15671 1241 15681 1275
rect 15715 1241 15727 1275
rect 15671 1207 15727 1241
rect 15671 1173 15681 1207
rect 15715 1173 15727 1207
rect 15671 1139 15727 1173
rect 15671 1105 15681 1139
rect 15715 1105 15727 1139
rect 15671 1051 15727 1105
rect 15757 1411 15815 1451
rect 15757 1377 15769 1411
rect 15803 1377 15815 1411
rect 15757 1343 15815 1377
rect 15757 1309 15769 1343
rect 15803 1309 15815 1343
rect 15757 1275 15815 1309
rect 15757 1241 15769 1275
rect 15803 1241 15815 1275
rect 15757 1207 15815 1241
rect 15757 1173 15769 1207
rect 15803 1173 15815 1207
rect 15757 1139 15815 1173
rect 15757 1105 15769 1139
rect 15803 1105 15815 1139
rect 15757 1051 15815 1105
rect 15845 1411 15903 1451
rect 15845 1377 15857 1411
rect 15891 1377 15903 1411
rect 15845 1343 15903 1377
rect 15845 1309 15857 1343
rect 15891 1309 15903 1343
rect 15845 1275 15903 1309
rect 15845 1241 15857 1275
rect 15891 1241 15903 1275
rect 15845 1207 15903 1241
rect 15845 1173 15857 1207
rect 15891 1173 15903 1207
rect 15845 1051 15903 1173
rect 15933 1411 15991 1451
rect 15933 1377 15945 1411
rect 15979 1377 15991 1411
rect 15933 1343 15991 1377
rect 15933 1309 15945 1343
rect 15979 1309 15991 1343
rect 15933 1275 15991 1309
rect 15933 1241 15945 1275
rect 15979 1241 15991 1275
rect 15933 1207 15991 1241
rect 15933 1173 15945 1207
rect 15979 1173 15991 1207
rect 15933 1051 15991 1173
rect 16021 1411 16075 1451
rect 16021 1377 16033 1411
rect 16067 1377 16075 1411
rect 16021 1343 16075 1377
rect 16021 1309 16033 1343
rect 16067 1309 16075 1343
rect 16021 1275 16075 1309
rect 16021 1241 16033 1275
rect 16067 1241 16075 1275
rect 16021 1207 16075 1241
rect 16021 1173 16033 1207
rect 16067 1173 16075 1207
rect 16021 1139 16075 1173
rect 16021 1105 16033 1139
rect 16067 1105 16075 1139
rect 16021 1051 16075 1105
rect 16337 1411 16391 1451
rect 16337 1377 16345 1411
rect 16379 1377 16391 1411
rect 16337 1343 16391 1377
rect 16337 1309 16345 1343
rect 16379 1309 16391 1343
rect 16337 1275 16391 1309
rect 16337 1241 16345 1275
rect 16379 1241 16391 1275
rect 16337 1207 16391 1241
rect 16337 1173 16345 1207
rect 16379 1173 16391 1207
rect 16337 1051 16391 1173
rect 16421 1343 16479 1451
rect 16421 1309 16433 1343
rect 16467 1309 16479 1343
rect 16421 1275 16479 1309
rect 16421 1241 16433 1275
rect 16467 1241 16479 1275
rect 16421 1207 16479 1241
rect 16421 1173 16433 1207
rect 16467 1173 16479 1207
rect 16421 1139 16479 1173
rect 16421 1105 16433 1139
rect 16467 1105 16479 1139
rect 16421 1051 16479 1105
rect 16509 1411 16567 1451
rect 16509 1377 16521 1411
rect 16555 1377 16567 1411
rect 16509 1343 16567 1377
rect 16509 1309 16521 1343
rect 16555 1309 16567 1343
rect 16509 1275 16567 1309
rect 16509 1241 16521 1275
rect 16555 1241 16567 1275
rect 16509 1207 16567 1241
rect 16509 1173 16521 1207
rect 16555 1173 16567 1207
rect 16509 1051 16567 1173
rect 16597 1343 16655 1451
rect 16597 1309 16609 1343
rect 16643 1309 16655 1343
rect 16597 1275 16655 1309
rect 16597 1241 16609 1275
rect 16643 1241 16655 1275
rect 16597 1207 16655 1241
rect 16597 1173 16609 1207
rect 16643 1173 16655 1207
rect 16597 1051 16655 1173
rect 16685 1411 16741 1451
rect 16685 1377 16697 1411
rect 16731 1377 16741 1411
rect 16685 1343 16741 1377
rect 16685 1309 16697 1343
rect 16731 1309 16741 1343
rect 16685 1275 16741 1309
rect 16685 1241 16697 1275
rect 16731 1241 16741 1275
rect 16685 1207 16741 1241
rect 16685 1173 16697 1207
rect 16731 1173 16741 1207
rect 16685 1051 16741 1173
rect 17003 1411 17059 1451
rect 17003 1377 17013 1411
rect 17047 1377 17059 1411
rect 17003 1343 17059 1377
rect 17003 1309 17013 1343
rect 17047 1309 17059 1343
rect 17003 1275 17059 1309
rect 17003 1241 17013 1275
rect 17047 1241 17059 1275
rect 17003 1207 17059 1241
rect 17003 1173 17013 1207
rect 17047 1173 17059 1207
rect 17003 1051 17059 1173
rect 17089 1343 17147 1451
rect 17089 1309 17101 1343
rect 17135 1309 17147 1343
rect 17089 1275 17147 1309
rect 17089 1241 17101 1275
rect 17135 1241 17147 1275
rect 17089 1207 17147 1241
rect 17089 1173 17101 1207
rect 17135 1173 17147 1207
rect 17089 1139 17147 1173
rect 17089 1105 17101 1139
rect 17135 1105 17147 1139
rect 17089 1051 17147 1105
rect 17177 1411 17235 1451
rect 17177 1377 17189 1411
rect 17223 1377 17235 1411
rect 17177 1343 17235 1377
rect 17177 1309 17189 1343
rect 17223 1309 17235 1343
rect 17177 1275 17235 1309
rect 17177 1241 17189 1275
rect 17223 1241 17235 1275
rect 17177 1207 17235 1241
rect 17177 1173 17189 1207
rect 17223 1173 17235 1207
rect 17177 1051 17235 1173
rect 17265 1343 17323 1451
rect 17265 1309 17277 1343
rect 17311 1309 17323 1343
rect 17265 1275 17323 1309
rect 17265 1241 17277 1275
rect 17311 1241 17323 1275
rect 17265 1207 17323 1241
rect 17265 1173 17277 1207
rect 17311 1173 17323 1207
rect 17265 1139 17323 1173
rect 17265 1105 17277 1139
rect 17311 1105 17323 1139
rect 17265 1051 17323 1105
rect 17353 1411 17407 1451
rect 17353 1377 17365 1411
rect 17399 1377 17407 1411
rect 17353 1343 17407 1377
rect 17353 1309 17365 1343
rect 17399 1309 17407 1343
rect 17353 1275 17407 1309
rect 17353 1241 17365 1275
rect 17399 1241 17407 1275
rect 17353 1207 17407 1241
rect 17353 1173 17365 1207
rect 17399 1173 17407 1207
rect 17353 1051 17407 1173
rect 17645 1412 17701 1450
rect 17645 1378 17655 1412
rect 17689 1378 17701 1412
rect 17645 1344 17701 1378
rect 17645 1310 17655 1344
rect 17689 1310 17701 1344
rect 17645 1276 17701 1310
rect 17645 1242 17655 1276
rect 17689 1242 17701 1276
rect 17645 1208 17701 1242
rect 17645 1174 17655 1208
rect 17689 1174 17701 1208
rect 17645 1139 17701 1174
rect 17645 1105 17655 1139
rect 17689 1105 17701 1139
rect 17645 1050 17701 1105
rect 17731 1412 17789 1450
rect 17731 1378 17743 1412
rect 17777 1378 17789 1412
rect 17731 1344 17789 1378
rect 17731 1310 17743 1344
rect 17777 1310 17789 1344
rect 17731 1276 17789 1310
rect 17731 1242 17743 1276
rect 17777 1242 17789 1276
rect 17731 1208 17789 1242
rect 17731 1174 17743 1208
rect 17777 1174 17789 1208
rect 17731 1139 17789 1174
rect 17731 1105 17743 1139
rect 17777 1105 17789 1139
rect 17731 1050 17789 1105
rect 17819 1412 17873 1450
rect 17819 1378 17831 1412
rect 17865 1378 17873 1412
rect 17819 1344 17873 1378
rect 17819 1310 17831 1344
rect 17865 1310 17873 1344
rect 17819 1276 17873 1310
rect 17819 1242 17831 1276
rect 17865 1242 17873 1276
rect 17819 1208 17873 1242
rect 17819 1174 17831 1208
rect 17865 1174 17873 1208
rect 17819 1139 17873 1174
rect 17819 1105 17831 1139
rect 17865 1105 17873 1139
rect 17819 1050 17873 1105
<< ndiffc >>
rect 101 329 135 363
rect 198 329 232 363
rect 295 329 329 363
rect 392 329 426 363
rect 489 329 523 363
rect 101 257 135 291
rect 101 189 135 223
rect 198 204 232 238
rect 295 257 329 291
rect 295 189 329 223
rect 393 210 427 244
rect 101 119 135 153
rect 295 119 329 153
rect 392 119 426 153
rect 489 119 523 153
rect 603 329 637 363
rect 603 257 637 291
rect 603 189 637 223
rect 700 213 734 247
rect 797 257 831 291
rect 797 189 831 223
rect 603 119 637 153
rect 700 119 734 153
rect 797 119 831 153
rect 1063 329 1097 363
rect 1160 329 1194 363
rect 1257 329 1291 363
rect 1354 329 1388 363
rect 1451 329 1485 363
rect 1063 257 1097 291
rect 1063 189 1097 223
rect 1160 204 1194 238
rect 1257 257 1291 291
rect 1257 189 1291 223
rect 1355 210 1389 244
rect 1063 119 1097 153
rect 1257 119 1291 153
rect 1354 119 1388 153
rect 1451 119 1485 153
rect 1565 329 1599 363
rect 1565 257 1599 291
rect 1565 189 1599 223
rect 1662 213 1696 247
rect 1759 257 1793 291
rect 1759 189 1793 223
rect 1565 119 1599 153
rect 1662 119 1696 153
rect 1759 119 1793 153
rect 2046 327 2080 361
rect 2143 327 2177 361
rect 2240 327 2274 361
rect 2046 255 2080 289
rect 2046 187 2080 221
rect 2143 202 2177 236
rect 2240 255 2274 289
rect 2240 187 2274 221
rect 2337 211 2371 245
rect 2434 255 2468 289
rect 2434 187 2468 221
rect 2046 117 2080 151
rect 2240 117 2274 151
rect 2337 117 2371 151
rect 2434 117 2468 151
rect 2691 329 2725 363
rect 2788 329 2822 363
rect 2885 329 2919 363
rect 2982 329 3016 363
rect 3079 329 3113 363
rect 2691 257 2725 291
rect 2691 189 2725 223
rect 2788 204 2822 238
rect 2885 257 2919 291
rect 2885 189 2919 223
rect 2983 210 3017 244
rect 2691 119 2725 153
rect 2885 119 2919 153
rect 2982 119 3016 153
rect 3079 119 3113 153
rect 3193 329 3227 363
rect 3193 257 3227 291
rect 3193 189 3227 223
rect 3290 213 3324 247
rect 3387 257 3421 291
rect 3387 189 3421 223
rect 3193 119 3227 153
rect 3290 119 3324 153
rect 3387 119 3421 153
rect 3653 329 3687 363
rect 3750 329 3784 363
rect 3847 329 3881 363
rect 3944 329 3978 363
rect 4041 329 4075 363
rect 3653 257 3687 291
rect 3653 189 3687 223
rect 3750 204 3784 238
rect 3847 257 3881 291
rect 3847 189 3881 223
rect 3945 210 3979 244
rect 3653 119 3687 153
rect 3847 119 3881 153
rect 3944 119 3978 153
rect 4041 119 4075 153
rect 4155 329 4189 363
rect 4155 257 4189 291
rect 4155 189 4189 223
rect 4252 213 4286 247
rect 4349 257 4383 291
rect 4349 189 4383 223
rect 4155 119 4189 153
rect 4252 119 4286 153
rect 4349 119 4383 153
rect 4636 327 4670 361
rect 4733 327 4767 361
rect 4830 327 4864 361
rect 4636 255 4670 289
rect 4636 187 4670 221
rect 4733 202 4767 236
rect 4830 255 4864 289
rect 4830 187 4864 221
rect 4927 211 4961 245
rect 5024 255 5058 289
rect 5024 187 5058 221
rect 4636 117 4670 151
rect 4830 117 4864 151
rect 4927 117 4961 151
rect 5024 117 5058 151
rect 5281 329 5315 363
rect 5378 329 5412 363
rect 5475 329 5509 363
rect 5572 329 5606 363
rect 5669 329 5703 363
rect 5281 257 5315 291
rect 5281 189 5315 223
rect 5378 204 5412 238
rect 5475 257 5509 291
rect 5475 189 5509 223
rect 5573 210 5607 244
rect 5281 119 5315 153
rect 5475 119 5509 153
rect 5572 119 5606 153
rect 5669 119 5703 153
rect 5783 329 5817 363
rect 5783 257 5817 291
rect 5783 189 5817 223
rect 5880 213 5914 247
rect 5977 257 6011 291
rect 5977 189 6011 223
rect 5783 119 5817 153
rect 5880 119 5914 153
rect 5977 119 6011 153
rect 6243 329 6277 363
rect 6340 329 6374 363
rect 6437 329 6471 363
rect 6534 329 6568 363
rect 6631 329 6665 363
rect 6243 257 6277 291
rect 6243 189 6277 223
rect 6340 204 6374 238
rect 6437 257 6471 291
rect 6437 189 6471 223
rect 6535 210 6569 244
rect 6243 119 6277 153
rect 6437 119 6471 153
rect 6534 119 6568 153
rect 6631 119 6665 153
rect 6745 329 6779 363
rect 6745 257 6779 291
rect 6745 189 6779 223
rect 6842 213 6876 247
rect 6939 257 6973 291
rect 6939 189 6973 223
rect 6745 119 6779 153
rect 6842 119 6876 153
rect 6939 119 6973 153
rect 7226 327 7260 361
rect 7323 327 7357 361
rect 7420 327 7454 361
rect 7226 255 7260 289
rect 7226 187 7260 221
rect 7323 202 7357 236
rect 7420 255 7454 289
rect 7420 187 7454 221
rect 7517 211 7551 245
rect 7614 255 7648 289
rect 7614 187 7648 221
rect 7226 117 7260 151
rect 7420 117 7454 151
rect 7517 117 7551 151
rect 7614 117 7648 151
rect 7871 329 7905 363
rect 7968 329 8002 363
rect 8065 329 8099 363
rect 8162 329 8196 363
rect 8259 329 8293 363
rect 7871 257 7905 291
rect 7871 189 7905 223
rect 7968 204 8002 238
rect 8065 257 8099 291
rect 8065 189 8099 223
rect 8163 210 8197 244
rect 7871 119 7905 153
rect 8065 119 8099 153
rect 8162 119 8196 153
rect 8259 119 8293 153
rect 8373 329 8407 363
rect 8373 257 8407 291
rect 8373 189 8407 223
rect 8470 213 8504 247
rect 8567 257 8601 291
rect 8567 189 8601 223
rect 8373 119 8407 153
rect 8470 119 8504 153
rect 8567 119 8601 153
rect 8833 329 8867 363
rect 8930 329 8964 363
rect 9027 329 9061 363
rect 9124 329 9158 363
rect 9221 329 9255 363
rect 8833 257 8867 291
rect 8833 189 8867 223
rect 8930 204 8964 238
rect 9027 257 9061 291
rect 9027 189 9061 223
rect 9125 210 9159 244
rect 8833 119 8867 153
rect 9027 119 9061 153
rect 9124 119 9158 153
rect 9221 119 9255 153
rect 9335 329 9369 363
rect 9335 257 9369 291
rect 9335 189 9369 223
rect 9432 213 9466 247
rect 9529 257 9563 291
rect 9529 189 9563 223
rect 9335 119 9369 153
rect 9432 119 9466 153
rect 9529 119 9563 153
rect 9816 327 9850 361
rect 9913 327 9947 361
rect 10010 327 10044 361
rect 9816 255 9850 289
rect 9816 187 9850 221
rect 9913 202 9947 236
rect 10010 255 10044 289
rect 10010 187 10044 221
rect 10107 211 10141 245
rect 10204 255 10238 289
rect 10204 187 10238 221
rect 9816 117 9850 151
rect 10010 117 10044 151
rect 10107 117 10141 151
rect 10204 117 10238 151
rect 10461 329 10495 363
rect 10558 329 10592 363
rect 10655 329 10689 363
rect 10752 329 10786 363
rect 10849 329 10883 363
rect 10461 257 10495 291
rect 10461 189 10495 223
rect 10558 204 10592 238
rect 10655 257 10689 291
rect 10655 189 10689 223
rect 10753 210 10787 244
rect 10461 119 10495 153
rect 10655 119 10689 153
rect 10752 119 10786 153
rect 10849 119 10883 153
rect 10963 329 10997 363
rect 10963 257 10997 291
rect 10963 189 10997 223
rect 11060 213 11094 247
rect 11157 257 11191 291
rect 11157 189 11191 223
rect 10963 119 10997 153
rect 11060 119 11094 153
rect 11157 119 11191 153
rect 11423 329 11457 363
rect 11520 329 11554 363
rect 11617 329 11651 363
rect 11714 329 11748 363
rect 11811 329 11845 363
rect 11423 257 11457 291
rect 11423 189 11457 223
rect 11520 204 11554 238
rect 11617 257 11651 291
rect 11617 189 11651 223
rect 11715 210 11749 244
rect 11423 119 11457 153
rect 11617 119 11651 153
rect 11714 119 11748 153
rect 11811 119 11845 153
rect 11925 329 11959 363
rect 11925 257 11959 291
rect 11925 189 11959 223
rect 12022 213 12056 247
rect 12119 257 12153 291
rect 12119 189 12153 223
rect 11925 119 11959 153
rect 12022 119 12056 153
rect 12119 119 12153 153
rect 12406 327 12440 361
rect 12503 327 12537 361
rect 12600 327 12634 361
rect 12406 255 12440 289
rect 12406 187 12440 221
rect 12503 202 12537 236
rect 12600 255 12634 289
rect 12600 187 12634 221
rect 12697 211 12731 245
rect 12794 255 12828 289
rect 12794 187 12828 221
rect 12406 117 12440 151
rect 12600 117 12634 151
rect 12697 117 12731 151
rect 12794 117 12828 151
rect 13051 329 13085 363
rect 13148 329 13182 363
rect 13245 329 13279 363
rect 13342 329 13376 363
rect 13439 329 13473 363
rect 13051 257 13085 291
rect 13051 189 13085 223
rect 13148 204 13182 238
rect 13245 257 13279 291
rect 13245 189 13279 223
rect 13343 210 13377 244
rect 13051 119 13085 153
rect 13245 119 13279 153
rect 13342 119 13376 153
rect 13439 119 13473 153
rect 13553 329 13587 363
rect 13553 257 13587 291
rect 13553 189 13587 223
rect 13650 213 13684 247
rect 13747 257 13781 291
rect 13747 189 13781 223
rect 13553 119 13587 153
rect 13650 119 13684 153
rect 13747 119 13781 153
rect 14013 329 14047 363
rect 14110 329 14144 363
rect 14207 329 14241 363
rect 14304 329 14338 363
rect 14401 329 14435 363
rect 14013 257 14047 291
rect 14013 189 14047 223
rect 14110 204 14144 238
rect 14207 257 14241 291
rect 14207 189 14241 223
rect 14305 210 14339 244
rect 14013 119 14047 153
rect 14207 119 14241 153
rect 14304 119 14338 153
rect 14401 119 14435 153
rect 14515 329 14549 363
rect 14515 257 14549 291
rect 14515 189 14549 223
rect 14612 213 14646 247
rect 14709 257 14743 291
rect 14709 189 14743 223
rect 14515 119 14549 153
rect 14612 119 14646 153
rect 14709 119 14743 153
rect 14996 327 15030 361
rect 15093 327 15127 361
rect 15190 327 15224 361
rect 14996 255 15030 289
rect 14996 187 15030 221
rect 15093 202 15127 236
rect 15190 255 15224 289
rect 15190 187 15224 221
rect 15287 211 15321 245
rect 15384 255 15418 289
rect 15384 187 15418 221
rect 14996 117 15030 151
rect 15190 117 15224 151
rect 15287 117 15321 151
rect 15384 117 15418 151
rect 15662 327 15696 361
rect 15759 327 15793 361
rect 15856 327 15890 361
rect 16050 327 16084 361
rect 15662 255 15696 289
rect 15662 187 15696 221
rect 15759 202 15793 236
rect 15856 255 15890 289
rect 15856 187 15890 221
rect 15952 211 15986 245
rect 16050 255 16084 289
rect 16050 187 16084 221
rect 15662 117 15696 151
rect 15856 117 15890 151
rect 15952 117 15986 151
rect 16050 117 16084 151
rect 16328 327 16362 361
rect 16425 327 16459 361
rect 16522 327 16556 361
rect 16716 327 16750 361
rect 16328 255 16362 289
rect 16328 187 16362 221
rect 16425 202 16459 236
rect 16522 255 16556 289
rect 16522 187 16556 221
rect 16619 211 16653 245
rect 16716 255 16750 289
rect 16716 187 16750 221
rect 16328 117 16362 151
rect 16522 117 16556 151
rect 16619 117 16653 151
rect 16716 117 16750 151
rect 16994 327 17028 361
rect 17091 327 17125 361
rect 17188 327 17222 361
rect 16994 255 17028 289
rect 16994 187 17028 221
rect 17091 202 17125 236
rect 17188 255 17222 289
rect 17188 187 17222 221
rect 17285 211 17319 245
rect 17382 255 17416 289
rect 17382 187 17416 221
rect 16994 117 17028 151
rect 17188 117 17222 151
rect 17285 117 17319 151
rect 17382 117 17416 151
rect 17647 327 17681 361
rect 17841 327 17875 361
rect 17647 255 17681 289
rect 17647 187 17681 221
rect 17743 211 17777 245
rect 17841 255 17875 289
rect 17841 187 17875 221
rect 17647 117 17681 151
rect 17743 117 17777 151
rect 17841 117 17875 151
<< pdiffc >>
rect 201 1378 235 1412
rect 201 1310 235 1344
rect 201 1242 235 1276
rect 201 1174 235 1208
rect 201 1105 235 1139
rect 289 1378 323 1412
rect 289 1310 323 1344
rect 289 1242 323 1276
rect 289 1174 323 1208
rect 289 1105 323 1139
rect 377 1378 411 1412
rect 377 1310 411 1344
rect 377 1242 411 1276
rect 377 1174 411 1208
rect 465 1378 499 1412
rect 465 1310 499 1344
rect 465 1242 499 1276
rect 465 1174 499 1208
rect 465 1105 499 1139
rect 553 1378 587 1412
rect 553 1310 587 1344
rect 553 1242 587 1276
rect 553 1174 587 1208
rect 641 1378 675 1412
rect 641 1310 675 1344
rect 641 1242 675 1276
rect 641 1174 675 1208
rect 641 1105 675 1139
rect 729 1378 763 1412
rect 729 1310 763 1344
rect 729 1242 763 1276
rect 729 1174 763 1208
rect 1163 1378 1197 1412
rect 1163 1310 1197 1344
rect 1163 1242 1197 1276
rect 1163 1174 1197 1208
rect 1163 1105 1197 1139
rect 1251 1378 1285 1412
rect 1251 1310 1285 1344
rect 1251 1242 1285 1276
rect 1251 1174 1285 1208
rect 1251 1105 1285 1139
rect 1339 1378 1373 1412
rect 1339 1310 1373 1344
rect 1339 1242 1373 1276
rect 1339 1174 1373 1208
rect 1427 1378 1461 1412
rect 1427 1310 1461 1344
rect 1427 1242 1461 1276
rect 1427 1174 1461 1208
rect 1427 1105 1461 1139
rect 1515 1378 1549 1412
rect 1515 1310 1549 1344
rect 1515 1242 1549 1276
rect 1515 1174 1549 1208
rect 1603 1378 1637 1412
rect 1603 1310 1637 1344
rect 1603 1242 1637 1276
rect 1603 1174 1637 1208
rect 1603 1105 1637 1139
rect 1691 1378 1725 1412
rect 1691 1310 1725 1344
rect 1691 1242 1725 1276
rect 1691 1174 1725 1208
rect 2065 1378 2099 1412
rect 2065 1310 2099 1344
rect 2065 1242 2099 1276
rect 2065 1174 2099 1208
rect 2065 1105 2099 1139
rect 2153 1378 2187 1412
rect 2153 1310 2187 1344
rect 2153 1242 2187 1276
rect 2153 1174 2187 1208
rect 2153 1105 2187 1139
rect 2241 1378 2275 1412
rect 2241 1310 2275 1344
rect 2241 1242 2275 1276
rect 2241 1174 2275 1208
rect 2329 1378 2363 1412
rect 2329 1310 2363 1344
rect 2329 1242 2363 1276
rect 2329 1174 2363 1208
rect 2329 1105 2363 1139
rect 2417 1378 2451 1412
rect 2417 1310 2451 1344
rect 2417 1242 2451 1276
rect 2417 1174 2451 1208
rect 2791 1378 2825 1412
rect 2791 1310 2825 1344
rect 2791 1242 2825 1276
rect 2791 1174 2825 1208
rect 2791 1105 2825 1139
rect 2879 1378 2913 1412
rect 2879 1310 2913 1344
rect 2879 1242 2913 1276
rect 2879 1174 2913 1208
rect 2879 1105 2913 1139
rect 2967 1378 3001 1412
rect 2967 1310 3001 1344
rect 2967 1242 3001 1276
rect 2967 1174 3001 1208
rect 3055 1378 3089 1412
rect 3055 1310 3089 1344
rect 3055 1242 3089 1276
rect 3055 1174 3089 1208
rect 3055 1105 3089 1139
rect 3143 1378 3177 1412
rect 3143 1310 3177 1344
rect 3143 1242 3177 1276
rect 3143 1174 3177 1208
rect 3231 1378 3265 1412
rect 3231 1310 3265 1344
rect 3231 1242 3265 1276
rect 3231 1174 3265 1208
rect 3231 1105 3265 1139
rect 3319 1378 3353 1412
rect 3319 1310 3353 1344
rect 3319 1242 3353 1276
rect 3319 1174 3353 1208
rect 3753 1378 3787 1412
rect 3753 1310 3787 1344
rect 3753 1242 3787 1276
rect 3753 1174 3787 1208
rect 3753 1105 3787 1139
rect 3841 1378 3875 1412
rect 3841 1310 3875 1344
rect 3841 1242 3875 1276
rect 3841 1174 3875 1208
rect 3841 1105 3875 1139
rect 3929 1378 3963 1412
rect 3929 1310 3963 1344
rect 3929 1242 3963 1276
rect 3929 1174 3963 1208
rect 4017 1378 4051 1412
rect 4017 1310 4051 1344
rect 4017 1242 4051 1276
rect 4017 1174 4051 1208
rect 4017 1105 4051 1139
rect 4105 1378 4139 1412
rect 4105 1310 4139 1344
rect 4105 1242 4139 1276
rect 4105 1174 4139 1208
rect 4193 1378 4227 1412
rect 4193 1310 4227 1344
rect 4193 1242 4227 1276
rect 4193 1174 4227 1208
rect 4193 1105 4227 1139
rect 4281 1378 4315 1412
rect 4281 1310 4315 1344
rect 4281 1242 4315 1276
rect 4281 1174 4315 1208
rect 4655 1378 4689 1412
rect 4655 1310 4689 1344
rect 4655 1242 4689 1276
rect 4655 1174 4689 1208
rect 4655 1105 4689 1139
rect 4743 1378 4777 1412
rect 4743 1310 4777 1344
rect 4743 1242 4777 1276
rect 4743 1174 4777 1208
rect 4743 1105 4777 1139
rect 4831 1378 4865 1412
rect 4831 1310 4865 1344
rect 4831 1242 4865 1276
rect 4831 1174 4865 1208
rect 4919 1378 4953 1412
rect 4919 1310 4953 1344
rect 4919 1242 4953 1276
rect 4919 1174 4953 1208
rect 4919 1105 4953 1139
rect 5007 1378 5041 1412
rect 5007 1310 5041 1344
rect 5007 1242 5041 1276
rect 5007 1174 5041 1208
rect 5381 1378 5415 1412
rect 5381 1310 5415 1344
rect 5381 1242 5415 1276
rect 5381 1174 5415 1208
rect 5381 1105 5415 1139
rect 5469 1378 5503 1412
rect 5469 1310 5503 1344
rect 5469 1242 5503 1276
rect 5469 1174 5503 1208
rect 5469 1105 5503 1139
rect 5557 1378 5591 1412
rect 5557 1310 5591 1344
rect 5557 1242 5591 1276
rect 5557 1174 5591 1208
rect 5645 1378 5679 1412
rect 5645 1310 5679 1344
rect 5645 1242 5679 1276
rect 5645 1174 5679 1208
rect 5645 1105 5679 1139
rect 5733 1378 5767 1412
rect 5733 1310 5767 1344
rect 5733 1242 5767 1276
rect 5733 1174 5767 1208
rect 5821 1378 5855 1412
rect 5821 1310 5855 1344
rect 5821 1242 5855 1276
rect 5821 1174 5855 1208
rect 5821 1105 5855 1139
rect 5909 1378 5943 1412
rect 5909 1310 5943 1344
rect 5909 1242 5943 1276
rect 5909 1174 5943 1208
rect 6343 1378 6377 1412
rect 6343 1310 6377 1344
rect 6343 1242 6377 1276
rect 6343 1174 6377 1208
rect 6343 1105 6377 1139
rect 6431 1378 6465 1412
rect 6431 1310 6465 1344
rect 6431 1242 6465 1276
rect 6431 1174 6465 1208
rect 6431 1105 6465 1139
rect 6519 1378 6553 1412
rect 6519 1310 6553 1344
rect 6519 1242 6553 1276
rect 6519 1174 6553 1208
rect 6607 1378 6641 1412
rect 6607 1310 6641 1344
rect 6607 1242 6641 1276
rect 6607 1174 6641 1208
rect 6607 1105 6641 1139
rect 6695 1378 6729 1412
rect 6695 1310 6729 1344
rect 6695 1242 6729 1276
rect 6695 1174 6729 1208
rect 6783 1378 6817 1412
rect 6783 1310 6817 1344
rect 6783 1242 6817 1276
rect 6783 1174 6817 1208
rect 6783 1105 6817 1139
rect 6871 1378 6905 1412
rect 6871 1310 6905 1344
rect 6871 1242 6905 1276
rect 6871 1174 6905 1208
rect 7245 1378 7279 1412
rect 7245 1310 7279 1344
rect 7245 1242 7279 1276
rect 7245 1174 7279 1208
rect 7245 1105 7279 1139
rect 7333 1378 7367 1412
rect 7333 1310 7367 1344
rect 7333 1242 7367 1276
rect 7333 1174 7367 1208
rect 7333 1105 7367 1139
rect 7421 1378 7455 1412
rect 7421 1310 7455 1344
rect 7421 1242 7455 1276
rect 7421 1174 7455 1208
rect 7509 1378 7543 1412
rect 7509 1310 7543 1344
rect 7509 1242 7543 1276
rect 7509 1174 7543 1208
rect 7509 1105 7543 1139
rect 7597 1378 7631 1412
rect 7597 1310 7631 1344
rect 7597 1242 7631 1276
rect 7597 1174 7631 1208
rect 7971 1378 8005 1412
rect 7971 1310 8005 1344
rect 7971 1242 8005 1276
rect 7971 1174 8005 1208
rect 7971 1105 8005 1139
rect 8059 1378 8093 1412
rect 8059 1310 8093 1344
rect 8059 1242 8093 1276
rect 8059 1174 8093 1208
rect 8059 1105 8093 1139
rect 8147 1378 8181 1412
rect 8147 1310 8181 1344
rect 8147 1242 8181 1276
rect 8147 1174 8181 1208
rect 8235 1378 8269 1412
rect 8235 1310 8269 1344
rect 8235 1242 8269 1276
rect 8235 1174 8269 1208
rect 8235 1105 8269 1139
rect 8323 1378 8357 1412
rect 8323 1310 8357 1344
rect 8323 1242 8357 1276
rect 8323 1174 8357 1208
rect 8411 1378 8445 1412
rect 8411 1310 8445 1344
rect 8411 1242 8445 1276
rect 8411 1174 8445 1208
rect 8411 1105 8445 1139
rect 8499 1378 8533 1412
rect 8499 1310 8533 1344
rect 8499 1242 8533 1276
rect 8499 1174 8533 1208
rect 8933 1378 8967 1412
rect 8933 1310 8967 1344
rect 8933 1242 8967 1276
rect 8933 1174 8967 1208
rect 8933 1105 8967 1139
rect 9021 1378 9055 1412
rect 9021 1310 9055 1344
rect 9021 1242 9055 1276
rect 9021 1174 9055 1208
rect 9021 1105 9055 1139
rect 9109 1378 9143 1412
rect 9109 1310 9143 1344
rect 9109 1242 9143 1276
rect 9109 1174 9143 1208
rect 9197 1378 9231 1412
rect 9197 1310 9231 1344
rect 9197 1242 9231 1276
rect 9197 1174 9231 1208
rect 9197 1105 9231 1139
rect 9285 1378 9319 1412
rect 9285 1310 9319 1344
rect 9285 1242 9319 1276
rect 9285 1174 9319 1208
rect 9373 1378 9407 1412
rect 9373 1310 9407 1344
rect 9373 1242 9407 1276
rect 9373 1174 9407 1208
rect 9373 1105 9407 1139
rect 9461 1378 9495 1412
rect 9461 1310 9495 1344
rect 9461 1242 9495 1276
rect 9461 1174 9495 1208
rect 9835 1378 9869 1412
rect 9835 1310 9869 1344
rect 9835 1242 9869 1276
rect 9835 1174 9869 1208
rect 9835 1105 9869 1139
rect 9923 1378 9957 1412
rect 9923 1310 9957 1344
rect 9923 1242 9957 1276
rect 9923 1174 9957 1208
rect 9923 1105 9957 1139
rect 10011 1378 10045 1412
rect 10011 1310 10045 1344
rect 10011 1242 10045 1276
rect 10011 1174 10045 1208
rect 10099 1378 10133 1412
rect 10099 1310 10133 1344
rect 10099 1242 10133 1276
rect 10099 1174 10133 1208
rect 10099 1105 10133 1139
rect 10187 1378 10221 1412
rect 10187 1310 10221 1344
rect 10187 1242 10221 1276
rect 10187 1174 10221 1208
rect 10561 1378 10595 1412
rect 10561 1310 10595 1344
rect 10561 1242 10595 1276
rect 10561 1174 10595 1208
rect 10561 1105 10595 1139
rect 10649 1378 10683 1412
rect 10649 1310 10683 1344
rect 10649 1242 10683 1276
rect 10649 1174 10683 1208
rect 10649 1105 10683 1139
rect 10737 1378 10771 1412
rect 10737 1310 10771 1344
rect 10737 1242 10771 1276
rect 10737 1174 10771 1208
rect 10825 1378 10859 1412
rect 10825 1310 10859 1344
rect 10825 1242 10859 1276
rect 10825 1174 10859 1208
rect 10825 1105 10859 1139
rect 10913 1378 10947 1412
rect 10913 1310 10947 1344
rect 10913 1242 10947 1276
rect 10913 1174 10947 1208
rect 11001 1378 11035 1412
rect 11001 1310 11035 1344
rect 11001 1242 11035 1276
rect 11001 1174 11035 1208
rect 11001 1105 11035 1139
rect 11089 1378 11123 1412
rect 11089 1310 11123 1344
rect 11089 1242 11123 1276
rect 11089 1174 11123 1208
rect 11523 1378 11557 1412
rect 11523 1310 11557 1344
rect 11523 1242 11557 1276
rect 11523 1174 11557 1208
rect 11523 1105 11557 1139
rect 11611 1378 11645 1412
rect 11611 1310 11645 1344
rect 11611 1242 11645 1276
rect 11611 1174 11645 1208
rect 11611 1105 11645 1139
rect 11699 1378 11733 1412
rect 11699 1310 11733 1344
rect 11699 1242 11733 1276
rect 11699 1174 11733 1208
rect 11787 1378 11821 1412
rect 11787 1310 11821 1344
rect 11787 1242 11821 1276
rect 11787 1174 11821 1208
rect 11787 1105 11821 1139
rect 11875 1378 11909 1412
rect 11875 1310 11909 1344
rect 11875 1242 11909 1276
rect 11875 1174 11909 1208
rect 11963 1378 11997 1412
rect 11963 1310 11997 1344
rect 11963 1242 11997 1276
rect 11963 1174 11997 1208
rect 11963 1105 11997 1139
rect 12051 1378 12085 1412
rect 12051 1310 12085 1344
rect 12051 1242 12085 1276
rect 12051 1174 12085 1208
rect 12425 1378 12459 1412
rect 12425 1310 12459 1344
rect 12425 1242 12459 1276
rect 12425 1174 12459 1208
rect 12425 1105 12459 1139
rect 12513 1378 12547 1412
rect 12513 1310 12547 1344
rect 12513 1242 12547 1276
rect 12513 1174 12547 1208
rect 12513 1105 12547 1139
rect 12601 1378 12635 1412
rect 12601 1310 12635 1344
rect 12601 1242 12635 1276
rect 12601 1174 12635 1208
rect 12689 1378 12723 1412
rect 12689 1310 12723 1344
rect 12689 1242 12723 1276
rect 12689 1174 12723 1208
rect 12689 1105 12723 1139
rect 12777 1378 12811 1412
rect 12777 1310 12811 1344
rect 12777 1242 12811 1276
rect 12777 1174 12811 1208
rect 13151 1378 13185 1412
rect 13151 1310 13185 1344
rect 13151 1242 13185 1276
rect 13151 1174 13185 1208
rect 13151 1105 13185 1139
rect 13239 1378 13273 1412
rect 13239 1310 13273 1344
rect 13239 1242 13273 1276
rect 13239 1174 13273 1208
rect 13239 1105 13273 1139
rect 13327 1378 13361 1412
rect 13327 1310 13361 1344
rect 13327 1242 13361 1276
rect 13327 1174 13361 1208
rect 13415 1378 13449 1412
rect 13415 1310 13449 1344
rect 13415 1242 13449 1276
rect 13415 1174 13449 1208
rect 13415 1105 13449 1139
rect 13503 1378 13537 1412
rect 13503 1310 13537 1344
rect 13503 1242 13537 1276
rect 13503 1174 13537 1208
rect 13591 1378 13625 1412
rect 13591 1310 13625 1344
rect 13591 1242 13625 1276
rect 13591 1174 13625 1208
rect 13591 1105 13625 1139
rect 13679 1378 13713 1412
rect 13679 1310 13713 1344
rect 13679 1242 13713 1276
rect 13679 1174 13713 1208
rect 14113 1378 14147 1412
rect 14113 1310 14147 1344
rect 14113 1242 14147 1276
rect 14113 1174 14147 1208
rect 14113 1105 14147 1139
rect 14201 1378 14235 1412
rect 14201 1310 14235 1344
rect 14201 1242 14235 1276
rect 14201 1174 14235 1208
rect 14201 1105 14235 1139
rect 14289 1378 14323 1412
rect 14289 1310 14323 1344
rect 14289 1242 14323 1276
rect 14289 1174 14323 1208
rect 14377 1378 14411 1412
rect 14377 1310 14411 1344
rect 14377 1242 14411 1276
rect 14377 1174 14411 1208
rect 14377 1105 14411 1139
rect 14465 1378 14499 1412
rect 14465 1310 14499 1344
rect 14465 1242 14499 1276
rect 14465 1174 14499 1208
rect 14553 1378 14587 1412
rect 14553 1310 14587 1344
rect 14553 1242 14587 1276
rect 14553 1174 14587 1208
rect 14553 1105 14587 1139
rect 14641 1378 14675 1412
rect 14641 1310 14675 1344
rect 14641 1242 14675 1276
rect 14641 1174 14675 1208
rect 15015 1378 15049 1412
rect 15015 1310 15049 1344
rect 15015 1242 15049 1276
rect 15015 1174 15049 1208
rect 15015 1105 15049 1139
rect 15103 1378 15137 1412
rect 15103 1310 15137 1344
rect 15103 1242 15137 1276
rect 15103 1174 15137 1208
rect 15103 1105 15137 1139
rect 15191 1378 15225 1412
rect 15191 1310 15225 1344
rect 15191 1242 15225 1276
rect 15191 1174 15225 1208
rect 15279 1378 15313 1412
rect 15279 1310 15313 1344
rect 15279 1242 15313 1276
rect 15279 1174 15313 1208
rect 15279 1105 15313 1139
rect 15367 1378 15401 1412
rect 15367 1310 15401 1344
rect 15367 1242 15401 1276
rect 15367 1174 15401 1208
rect 15681 1377 15715 1411
rect 15681 1309 15715 1343
rect 15681 1241 15715 1275
rect 15681 1173 15715 1207
rect 15681 1105 15715 1139
rect 15769 1377 15803 1411
rect 15769 1309 15803 1343
rect 15769 1241 15803 1275
rect 15769 1173 15803 1207
rect 15769 1105 15803 1139
rect 15857 1377 15891 1411
rect 15857 1309 15891 1343
rect 15857 1241 15891 1275
rect 15857 1173 15891 1207
rect 15945 1377 15979 1411
rect 15945 1309 15979 1343
rect 15945 1241 15979 1275
rect 15945 1173 15979 1207
rect 16033 1377 16067 1411
rect 16033 1309 16067 1343
rect 16033 1241 16067 1275
rect 16033 1173 16067 1207
rect 16033 1105 16067 1139
rect 16345 1377 16379 1411
rect 16345 1309 16379 1343
rect 16345 1241 16379 1275
rect 16345 1173 16379 1207
rect 16433 1309 16467 1343
rect 16433 1241 16467 1275
rect 16433 1173 16467 1207
rect 16433 1105 16467 1139
rect 16521 1377 16555 1411
rect 16521 1309 16555 1343
rect 16521 1241 16555 1275
rect 16521 1173 16555 1207
rect 16609 1309 16643 1343
rect 16609 1241 16643 1275
rect 16609 1173 16643 1207
rect 16697 1377 16731 1411
rect 16697 1309 16731 1343
rect 16697 1241 16731 1275
rect 16697 1173 16731 1207
rect 17013 1377 17047 1411
rect 17013 1309 17047 1343
rect 17013 1241 17047 1275
rect 17013 1173 17047 1207
rect 17101 1309 17135 1343
rect 17101 1241 17135 1275
rect 17101 1173 17135 1207
rect 17101 1105 17135 1139
rect 17189 1377 17223 1411
rect 17189 1309 17223 1343
rect 17189 1241 17223 1275
rect 17189 1173 17223 1207
rect 17277 1309 17311 1343
rect 17277 1241 17311 1275
rect 17277 1173 17311 1207
rect 17277 1105 17311 1139
rect 17365 1377 17399 1411
rect 17365 1309 17399 1343
rect 17365 1241 17399 1275
rect 17365 1173 17399 1207
rect 17655 1378 17689 1412
rect 17655 1310 17689 1344
rect 17655 1242 17689 1276
rect 17655 1174 17689 1208
rect 17655 1105 17689 1139
rect 17743 1378 17777 1412
rect 17743 1310 17777 1344
rect 17743 1242 17777 1276
rect 17743 1174 17777 1208
rect 17743 1105 17777 1139
rect 17831 1378 17865 1412
rect 17831 1310 17865 1344
rect 17831 1242 17865 1276
rect 17831 1174 17865 1208
rect 17831 1105 17865 1139
<< psubdiff >>
rect -31 546 18013 572
rect -31 512 -17 546
rect 17 512 945 546
rect 979 512 1907 546
rect 1941 512 2573 546
rect 2607 512 3535 546
rect 3569 512 4497 546
rect 4531 512 5163 546
rect 5197 512 6125 546
rect 6159 512 7087 546
rect 7121 512 7753 546
rect 7787 512 8715 546
rect 8749 512 9677 546
rect 9711 512 10343 546
rect 10377 512 11305 546
rect 11339 512 12267 546
rect 12301 512 12933 546
rect 12967 512 13895 546
rect 13929 512 14857 546
rect 14891 512 15523 546
rect 15557 512 16189 546
rect 16223 512 16855 546
rect 16889 512 17521 546
rect 17555 512 17965 546
rect 17999 512 18013 546
rect -31 510 18013 512
rect -31 474 31 510
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect -31 368 -17 402
rect 17 368 31 402
rect 931 474 993 510
rect 931 440 945 474
rect 979 440 993 474
rect 931 402 993 440
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect 931 368 945 402
rect 979 368 993 402
rect 1893 474 1955 510
rect 1893 440 1907 474
rect 1941 440 1955 474
rect 1893 402 1955 440
rect 931 330 993 368
rect 931 296 945 330
rect 979 296 993 330
rect 931 258 993 296
rect 931 224 945 258
rect 979 224 993 258
rect 931 186 993 224
rect 931 152 945 186
rect 979 152 993 186
rect 931 114 993 152
rect -31 47 31 80
rect 931 80 945 114
rect 979 80 993 114
rect 1893 368 1907 402
rect 1941 368 1955 402
rect 2559 474 2621 510
rect 2559 440 2573 474
rect 2607 440 2621 474
rect 2559 402 2621 440
rect 1893 330 1955 368
rect 1893 296 1907 330
rect 1941 296 1955 330
rect 1893 258 1955 296
rect 1893 224 1907 258
rect 1941 224 1955 258
rect 1893 186 1955 224
rect 1893 152 1907 186
rect 1941 152 1955 186
rect 1893 114 1955 152
rect 931 47 993 80
rect 1893 80 1907 114
rect 1941 80 1955 114
rect 2559 368 2573 402
rect 2607 368 2621 402
rect 3521 474 3583 510
rect 3521 440 3535 474
rect 3569 440 3583 474
rect 3521 402 3583 440
rect 2559 330 2621 368
rect 2559 296 2573 330
rect 2607 296 2621 330
rect 2559 258 2621 296
rect 2559 224 2573 258
rect 2607 224 2621 258
rect 2559 186 2621 224
rect 2559 152 2573 186
rect 2607 152 2621 186
rect 2559 114 2621 152
rect 1893 47 1955 80
rect 2559 80 2573 114
rect 2607 80 2621 114
rect 3521 368 3535 402
rect 3569 368 3583 402
rect 4483 474 4545 510
rect 4483 440 4497 474
rect 4531 440 4545 474
rect 4483 402 4545 440
rect 3521 330 3583 368
rect 3521 296 3535 330
rect 3569 296 3583 330
rect 3521 258 3583 296
rect 3521 224 3535 258
rect 3569 224 3583 258
rect 3521 186 3583 224
rect 3521 152 3535 186
rect 3569 152 3583 186
rect 3521 114 3583 152
rect 2559 47 2621 80
rect 3521 80 3535 114
rect 3569 80 3583 114
rect 4483 368 4497 402
rect 4531 368 4545 402
rect 5149 474 5211 510
rect 5149 440 5163 474
rect 5197 440 5211 474
rect 5149 402 5211 440
rect 4483 330 4545 368
rect 4483 296 4497 330
rect 4531 296 4545 330
rect 4483 258 4545 296
rect 4483 224 4497 258
rect 4531 224 4545 258
rect 4483 186 4545 224
rect 4483 152 4497 186
rect 4531 152 4545 186
rect 4483 114 4545 152
rect 3521 47 3583 80
rect 4483 80 4497 114
rect 4531 80 4545 114
rect 5149 368 5163 402
rect 5197 368 5211 402
rect 6111 474 6173 510
rect 6111 440 6125 474
rect 6159 440 6173 474
rect 6111 402 6173 440
rect 5149 330 5211 368
rect 5149 296 5163 330
rect 5197 296 5211 330
rect 5149 258 5211 296
rect 5149 224 5163 258
rect 5197 224 5211 258
rect 5149 186 5211 224
rect 5149 152 5163 186
rect 5197 152 5211 186
rect 5149 114 5211 152
rect 4483 47 4545 80
rect 5149 80 5163 114
rect 5197 80 5211 114
rect 6111 368 6125 402
rect 6159 368 6173 402
rect 7073 474 7135 510
rect 7073 440 7087 474
rect 7121 440 7135 474
rect 7073 402 7135 440
rect 6111 330 6173 368
rect 6111 296 6125 330
rect 6159 296 6173 330
rect 6111 258 6173 296
rect 6111 224 6125 258
rect 6159 224 6173 258
rect 6111 186 6173 224
rect 6111 152 6125 186
rect 6159 152 6173 186
rect 6111 114 6173 152
rect 5149 47 5211 80
rect 6111 80 6125 114
rect 6159 80 6173 114
rect 7073 368 7087 402
rect 7121 368 7135 402
rect 7739 474 7801 510
rect 7739 440 7753 474
rect 7787 440 7801 474
rect 7739 402 7801 440
rect 7073 330 7135 368
rect 7073 296 7087 330
rect 7121 296 7135 330
rect 7073 258 7135 296
rect 7073 224 7087 258
rect 7121 224 7135 258
rect 7073 186 7135 224
rect 7073 152 7087 186
rect 7121 152 7135 186
rect 7073 114 7135 152
rect 6111 47 6173 80
rect 7073 80 7087 114
rect 7121 80 7135 114
rect 7739 368 7753 402
rect 7787 368 7801 402
rect 8701 474 8763 510
rect 8701 440 8715 474
rect 8749 440 8763 474
rect 8701 402 8763 440
rect 7739 330 7801 368
rect 7739 296 7753 330
rect 7787 296 7801 330
rect 7739 258 7801 296
rect 7739 224 7753 258
rect 7787 224 7801 258
rect 7739 186 7801 224
rect 7739 152 7753 186
rect 7787 152 7801 186
rect 7739 114 7801 152
rect 7073 47 7135 80
rect 7739 80 7753 114
rect 7787 80 7801 114
rect 8701 368 8715 402
rect 8749 368 8763 402
rect 9663 474 9725 510
rect 9663 440 9677 474
rect 9711 440 9725 474
rect 9663 402 9725 440
rect 8701 330 8763 368
rect 8701 296 8715 330
rect 8749 296 8763 330
rect 8701 258 8763 296
rect 8701 224 8715 258
rect 8749 224 8763 258
rect 8701 186 8763 224
rect 8701 152 8715 186
rect 8749 152 8763 186
rect 8701 114 8763 152
rect 7739 47 7801 80
rect 8701 80 8715 114
rect 8749 80 8763 114
rect 9663 368 9677 402
rect 9711 368 9725 402
rect 10329 474 10391 510
rect 10329 440 10343 474
rect 10377 440 10391 474
rect 10329 402 10391 440
rect 9663 330 9725 368
rect 9663 296 9677 330
rect 9711 296 9725 330
rect 9663 258 9725 296
rect 9663 224 9677 258
rect 9711 224 9725 258
rect 9663 186 9725 224
rect 9663 152 9677 186
rect 9711 152 9725 186
rect 9663 114 9725 152
rect 8701 47 8763 80
rect 9663 80 9677 114
rect 9711 80 9725 114
rect 10329 368 10343 402
rect 10377 368 10391 402
rect 11291 474 11353 510
rect 11291 440 11305 474
rect 11339 440 11353 474
rect 11291 402 11353 440
rect 10329 330 10391 368
rect 10329 296 10343 330
rect 10377 296 10391 330
rect 10329 258 10391 296
rect 10329 224 10343 258
rect 10377 224 10391 258
rect 10329 186 10391 224
rect 10329 152 10343 186
rect 10377 152 10391 186
rect 10329 114 10391 152
rect 9663 47 9725 80
rect 10329 80 10343 114
rect 10377 80 10391 114
rect 11291 368 11305 402
rect 11339 368 11353 402
rect 12253 474 12315 510
rect 12253 440 12267 474
rect 12301 440 12315 474
rect 12253 402 12315 440
rect 11291 330 11353 368
rect 11291 296 11305 330
rect 11339 296 11353 330
rect 11291 258 11353 296
rect 11291 224 11305 258
rect 11339 224 11353 258
rect 11291 186 11353 224
rect 11291 152 11305 186
rect 11339 152 11353 186
rect 11291 114 11353 152
rect 10329 47 10391 80
rect 11291 80 11305 114
rect 11339 80 11353 114
rect 12253 368 12267 402
rect 12301 368 12315 402
rect 12919 474 12981 510
rect 12919 440 12933 474
rect 12967 440 12981 474
rect 12919 402 12981 440
rect 12253 330 12315 368
rect 12253 296 12267 330
rect 12301 296 12315 330
rect 12253 258 12315 296
rect 12253 224 12267 258
rect 12301 224 12315 258
rect 12253 186 12315 224
rect 12253 152 12267 186
rect 12301 152 12315 186
rect 12253 114 12315 152
rect 11291 47 11353 80
rect 12253 80 12267 114
rect 12301 80 12315 114
rect 12919 368 12933 402
rect 12967 368 12981 402
rect 13881 474 13943 510
rect 13881 440 13895 474
rect 13929 440 13943 474
rect 13881 402 13943 440
rect 12919 330 12981 368
rect 12919 296 12933 330
rect 12967 296 12981 330
rect 12919 258 12981 296
rect 12919 224 12933 258
rect 12967 224 12981 258
rect 12919 186 12981 224
rect 12919 152 12933 186
rect 12967 152 12981 186
rect 12919 114 12981 152
rect 12253 47 12315 80
rect 12919 80 12933 114
rect 12967 80 12981 114
rect 13881 368 13895 402
rect 13929 368 13943 402
rect 14843 474 14905 510
rect 14843 440 14857 474
rect 14891 440 14905 474
rect 14843 402 14905 440
rect 13881 330 13943 368
rect 13881 296 13895 330
rect 13929 296 13943 330
rect 13881 258 13943 296
rect 13881 224 13895 258
rect 13929 224 13943 258
rect 13881 186 13943 224
rect 13881 152 13895 186
rect 13929 152 13943 186
rect 13881 114 13943 152
rect 12919 47 12981 80
rect 13881 80 13895 114
rect 13929 80 13943 114
rect 14843 368 14857 402
rect 14891 368 14905 402
rect 15509 474 15571 510
rect 15509 440 15523 474
rect 15557 440 15571 474
rect 15509 402 15571 440
rect 16175 474 16237 510
rect 16175 440 16189 474
rect 16223 440 16237 474
rect 14843 330 14905 368
rect 14843 296 14857 330
rect 14891 296 14905 330
rect 14843 258 14905 296
rect 14843 224 14857 258
rect 14891 224 14905 258
rect 14843 186 14905 224
rect 14843 152 14857 186
rect 14891 152 14905 186
rect 14843 114 14905 152
rect 13881 47 13943 80
rect 14843 80 14857 114
rect 14891 80 14905 114
rect 15509 368 15523 402
rect 15557 368 15571 402
rect 16175 402 16237 440
rect 15509 330 15571 368
rect 15509 296 15523 330
rect 15557 296 15571 330
rect 15509 258 15571 296
rect 15509 224 15523 258
rect 15557 224 15571 258
rect 15509 186 15571 224
rect 15509 152 15523 186
rect 15557 152 15571 186
rect 15509 114 15571 152
rect 14843 47 14905 80
rect 15509 80 15523 114
rect 15557 80 15571 114
rect 16175 368 16189 402
rect 16223 368 16237 402
rect 16841 474 16903 510
rect 16841 440 16855 474
rect 16889 440 16903 474
rect 16841 402 16903 440
rect 17507 474 17569 510
rect 17507 440 17521 474
rect 17555 440 17569 474
rect 16175 330 16237 368
rect 16175 296 16189 330
rect 16223 296 16237 330
rect 16175 258 16237 296
rect 16175 224 16189 258
rect 16223 224 16237 258
rect 16175 186 16237 224
rect 16175 152 16189 186
rect 16223 152 16237 186
rect 16175 114 16237 152
rect 15509 47 15571 80
rect 16175 80 16189 114
rect 16223 80 16237 114
rect 16841 368 16855 402
rect 16889 368 16903 402
rect 17507 402 17569 440
rect 17951 474 18013 510
rect 16841 330 16903 368
rect 16841 296 16855 330
rect 16889 296 16903 330
rect 16841 258 16903 296
rect 16841 224 16855 258
rect 16889 224 16903 258
rect 16841 186 16903 224
rect 16841 152 16855 186
rect 16889 152 16903 186
rect 16841 114 16903 152
rect 16175 47 16237 80
rect 16841 80 16855 114
rect 16889 80 16903 114
rect 17507 368 17521 402
rect 17555 368 17569 402
rect 17951 440 17965 474
rect 17999 440 18013 474
rect 17951 402 18013 440
rect 17507 330 17569 368
rect 17507 296 17521 330
rect 17555 296 17569 330
rect 17507 258 17569 296
rect 17507 224 17521 258
rect 17555 224 17569 258
rect 17507 186 17569 224
rect 17507 152 17521 186
rect 17555 152 17569 186
rect 17507 114 17569 152
rect 16841 47 16903 80
rect 17507 80 17521 114
rect 17555 80 17569 114
rect 17951 368 17965 402
rect 17999 368 18013 402
rect 17951 330 18013 368
rect 17951 296 17965 330
rect 17999 296 18013 330
rect 17951 258 18013 296
rect 17951 224 17965 258
rect 17999 224 18013 258
rect 17951 186 18013 224
rect 17951 152 17965 186
rect 17999 152 18013 186
rect 17951 114 18013 152
rect 17507 47 17569 80
rect 17951 80 17965 114
rect 17999 80 18013 114
rect 17951 47 18013 80
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 343 47
rect 377 13 415 47
rect 449 13 513 47
rect 547 13 585 47
rect 619 13 657 47
rect 691 13 729 47
rect 763 13 801 47
rect 835 13 873 47
rect 907 13 1017 47
rect 1051 13 1089 47
rect 1123 13 1161 47
rect 1195 13 1233 47
rect 1267 13 1305 47
rect 1339 13 1377 47
rect 1411 13 1475 47
rect 1509 13 1547 47
rect 1581 13 1619 47
rect 1653 13 1691 47
rect 1725 13 1763 47
rect 1797 13 1835 47
rect 1869 13 1979 47
rect 2013 13 2051 47
rect 2085 13 2123 47
rect 2157 13 2195 47
rect 2229 13 2285 47
rect 2319 13 2357 47
rect 2391 13 2429 47
rect 2463 13 2501 47
rect 2535 13 2645 47
rect 2679 13 2717 47
rect 2751 13 2789 47
rect 2823 13 2861 47
rect 2895 13 2933 47
rect 2967 13 3005 47
rect 3039 13 3103 47
rect 3137 13 3175 47
rect 3209 13 3247 47
rect 3281 13 3319 47
rect 3353 13 3391 47
rect 3425 13 3463 47
rect 3497 13 3607 47
rect 3641 13 3679 47
rect 3713 13 3751 47
rect 3785 13 3823 47
rect 3857 13 3895 47
rect 3929 13 3967 47
rect 4001 13 4065 47
rect 4099 13 4137 47
rect 4171 13 4209 47
rect 4243 13 4281 47
rect 4315 13 4353 47
rect 4387 13 4425 47
rect 4459 13 4569 47
rect 4603 13 4641 47
rect 4675 13 4713 47
rect 4747 13 4785 47
rect 4819 13 4875 47
rect 4909 13 4947 47
rect 4981 13 5019 47
rect 5053 13 5091 47
rect 5125 13 5235 47
rect 5269 13 5307 47
rect 5341 13 5379 47
rect 5413 13 5451 47
rect 5485 13 5523 47
rect 5557 13 5595 47
rect 5629 13 5693 47
rect 5727 13 5765 47
rect 5799 13 5837 47
rect 5871 13 5909 47
rect 5943 13 5981 47
rect 6015 13 6053 47
rect 6087 13 6197 47
rect 6231 13 6269 47
rect 6303 13 6341 47
rect 6375 13 6413 47
rect 6447 13 6485 47
rect 6519 13 6557 47
rect 6591 13 6655 47
rect 6689 13 6727 47
rect 6761 13 6799 47
rect 6833 13 6871 47
rect 6905 13 6943 47
rect 6977 13 7015 47
rect 7049 13 7159 47
rect 7193 13 7231 47
rect 7265 13 7303 47
rect 7337 13 7375 47
rect 7409 13 7465 47
rect 7499 13 7537 47
rect 7571 13 7609 47
rect 7643 13 7681 47
rect 7715 13 7825 47
rect 7859 13 7897 47
rect 7931 13 7969 47
rect 8003 13 8041 47
rect 8075 13 8113 47
rect 8147 13 8185 47
rect 8219 13 8283 47
rect 8317 13 8355 47
rect 8389 13 8427 47
rect 8461 13 8499 47
rect 8533 13 8571 47
rect 8605 13 8643 47
rect 8677 13 8787 47
rect 8821 13 8859 47
rect 8893 13 8931 47
rect 8965 13 9003 47
rect 9037 13 9075 47
rect 9109 13 9147 47
rect 9181 13 9245 47
rect 9279 13 9317 47
rect 9351 13 9389 47
rect 9423 13 9461 47
rect 9495 13 9533 47
rect 9567 13 9605 47
rect 9639 13 9749 47
rect 9783 13 9821 47
rect 9855 13 9893 47
rect 9927 13 9965 47
rect 9999 13 10055 47
rect 10089 13 10127 47
rect 10161 13 10199 47
rect 10233 13 10271 47
rect 10305 13 10415 47
rect 10449 13 10487 47
rect 10521 13 10559 47
rect 10593 13 10631 47
rect 10665 13 10703 47
rect 10737 13 10775 47
rect 10809 13 10873 47
rect 10907 13 10945 47
rect 10979 13 11017 47
rect 11051 13 11089 47
rect 11123 13 11161 47
rect 11195 13 11233 47
rect 11267 13 11377 47
rect 11411 13 11449 47
rect 11483 13 11521 47
rect 11555 13 11593 47
rect 11627 13 11665 47
rect 11699 13 11737 47
rect 11771 13 11835 47
rect 11869 13 11907 47
rect 11941 13 11979 47
rect 12013 13 12051 47
rect 12085 13 12123 47
rect 12157 13 12195 47
rect 12229 13 12339 47
rect 12373 13 12411 47
rect 12445 13 12483 47
rect 12517 13 12555 47
rect 12589 13 12645 47
rect 12679 13 12717 47
rect 12751 13 12789 47
rect 12823 13 12861 47
rect 12895 13 13005 47
rect 13039 13 13077 47
rect 13111 13 13149 47
rect 13183 13 13221 47
rect 13255 13 13293 47
rect 13327 13 13365 47
rect 13399 13 13463 47
rect 13497 13 13535 47
rect 13569 13 13607 47
rect 13641 13 13679 47
rect 13713 13 13751 47
rect 13785 13 13823 47
rect 13857 13 13967 47
rect 14001 13 14039 47
rect 14073 13 14111 47
rect 14145 13 14183 47
rect 14217 13 14255 47
rect 14289 13 14327 47
rect 14361 13 14425 47
rect 14459 13 14497 47
rect 14531 13 14569 47
rect 14603 13 14641 47
rect 14675 13 14713 47
rect 14747 13 14785 47
rect 14819 13 14929 47
rect 14963 13 15001 47
rect 15035 13 15073 47
rect 15107 13 15145 47
rect 15179 13 15235 47
rect 15269 13 15307 47
rect 15341 13 15379 47
rect 15413 13 15451 47
rect 15485 13 15595 47
rect 15629 13 15667 47
rect 15701 13 15739 47
rect 15773 13 15811 47
rect 15845 13 15901 47
rect 15935 13 15973 47
rect 16007 13 16045 47
rect 16079 13 16117 47
rect 16151 13 16261 47
rect 16295 13 16333 47
rect 16367 13 16405 47
rect 16439 13 16477 47
rect 16511 13 16567 47
rect 16601 13 16639 47
rect 16673 13 16711 47
rect 16745 13 16783 47
rect 16817 13 16927 47
rect 16961 13 16999 47
rect 17033 13 17071 47
rect 17105 13 17143 47
rect 17177 13 17233 47
rect 17267 13 17305 47
rect 17339 13 17377 47
rect 17411 13 17449 47
rect 17483 13 17593 47
rect 17627 13 17665 47
rect 17699 13 17743 47
rect 17777 13 17821 47
rect 17855 13 17893 47
rect 17927 13 18013 47
rect -31 11 31 13
rect 931 11 993 13
rect 1893 11 1955 13
rect 2559 11 2621 13
rect 3521 11 3583 13
rect 4483 11 4545 13
rect 5149 11 5211 13
rect 6111 11 6173 13
rect 7073 11 7135 13
rect 7739 11 7801 13
rect 8701 11 8763 13
rect 9663 11 9725 13
rect 10329 11 10391 13
rect 11291 11 11353 13
rect 12253 11 12315 13
rect 12919 11 12981 13
rect 13881 11 13943 13
rect 14843 11 14905 13
rect 15509 11 15571 13
rect 16175 11 16237 13
rect 16841 11 16903 13
rect 17507 11 17569 13
rect 17951 11 18013 13
<< nsubdiff >>
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 343 1539
rect 377 1505 415 1539
rect 449 1505 513 1539
rect 547 1505 585 1539
rect 619 1505 657 1539
rect 691 1505 729 1539
rect 763 1505 801 1539
rect 835 1505 873 1539
rect 907 1505 1017 1539
rect 1051 1505 1089 1539
rect 1123 1505 1161 1539
rect 1195 1505 1233 1539
rect 1267 1505 1305 1539
rect 1339 1505 1377 1539
rect 1411 1505 1475 1539
rect 1509 1505 1547 1539
rect 1581 1505 1619 1539
rect 1653 1505 1691 1539
rect 1725 1505 1763 1539
rect 1797 1505 1835 1539
rect 1869 1505 1979 1539
rect 2013 1505 2051 1539
rect 2085 1505 2123 1539
rect 2157 1505 2195 1539
rect 2229 1505 2285 1539
rect 2319 1505 2357 1539
rect 2391 1505 2429 1539
rect 2463 1505 2501 1539
rect 2535 1505 2645 1539
rect 2679 1505 2717 1539
rect 2751 1505 2789 1539
rect 2823 1505 2861 1539
rect 2895 1505 2933 1539
rect 2967 1505 3005 1539
rect 3039 1505 3103 1539
rect 3137 1505 3175 1539
rect 3209 1505 3247 1539
rect 3281 1505 3319 1539
rect 3353 1505 3391 1539
rect 3425 1505 3463 1539
rect 3497 1505 3607 1539
rect 3641 1505 3679 1539
rect 3713 1505 3751 1539
rect 3785 1505 3823 1539
rect 3857 1505 3895 1539
rect 3929 1505 3967 1539
rect 4001 1505 4065 1539
rect 4099 1505 4137 1539
rect 4171 1505 4209 1539
rect 4243 1505 4281 1539
rect 4315 1505 4353 1539
rect 4387 1505 4425 1539
rect 4459 1505 4569 1539
rect 4603 1505 4641 1539
rect 4675 1505 4713 1539
rect 4747 1505 4785 1539
rect 4819 1505 4875 1539
rect 4909 1505 4947 1539
rect 4981 1505 5019 1539
rect 5053 1505 5091 1539
rect 5125 1505 5235 1539
rect 5269 1505 5307 1539
rect 5341 1505 5379 1539
rect 5413 1505 5451 1539
rect 5485 1505 5523 1539
rect 5557 1505 5595 1539
rect 5629 1505 5693 1539
rect 5727 1505 5765 1539
rect 5799 1505 5837 1539
rect 5871 1505 5909 1539
rect 5943 1505 5981 1539
rect 6015 1505 6053 1539
rect 6087 1505 6197 1539
rect 6231 1505 6269 1539
rect 6303 1505 6341 1539
rect 6375 1505 6413 1539
rect 6447 1505 6485 1539
rect 6519 1505 6557 1539
rect 6591 1505 6655 1539
rect 6689 1505 6727 1539
rect 6761 1505 6799 1539
rect 6833 1505 6871 1539
rect 6905 1505 6943 1539
rect 6977 1505 7015 1539
rect 7049 1505 7159 1539
rect 7193 1505 7231 1539
rect 7265 1505 7303 1539
rect 7337 1505 7375 1539
rect 7409 1505 7465 1539
rect 7499 1505 7537 1539
rect 7571 1505 7609 1539
rect 7643 1505 7681 1539
rect 7715 1505 7825 1539
rect 7859 1505 7897 1539
rect 7931 1505 7969 1539
rect 8003 1505 8041 1539
rect 8075 1505 8113 1539
rect 8147 1505 8185 1539
rect 8219 1505 8283 1539
rect 8317 1505 8355 1539
rect 8389 1505 8427 1539
rect 8461 1505 8499 1539
rect 8533 1505 8571 1539
rect 8605 1505 8643 1539
rect 8677 1505 8787 1539
rect 8821 1505 8859 1539
rect 8893 1505 8931 1539
rect 8965 1505 9003 1539
rect 9037 1505 9075 1539
rect 9109 1505 9147 1539
rect 9181 1505 9245 1539
rect 9279 1505 9317 1539
rect 9351 1505 9389 1539
rect 9423 1505 9461 1539
rect 9495 1505 9533 1539
rect 9567 1505 9605 1539
rect 9639 1505 9749 1539
rect 9783 1505 9821 1539
rect 9855 1505 9893 1539
rect 9927 1505 9965 1539
rect 9999 1505 10055 1539
rect 10089 1505 10127 1539
rect 10161 1505 10199 1539
rect 10233 1505 10271 1539
rect 10305 1505 10415 1539
rect 10449 1505 10487 1539
rect 10521 1505 10559 1539
rect 10593 1505 10631 1539
rect 10665 1505 10703 1539
rect 10737 1505 10775 1539
rect 10809 1505 10873 1539
rect 10907 1505 10945 1539
rect 10979 1505 11017 1539
rect 11051 1505 11089 1539
rect 11123 1505 11161 1539
rect 11195 1505 11233 1539
rect 11267 1505 11377 1539
rect 11411 1505 11449 1539
rect 11483 1505 11521 1539
rect 11555 1505 11593 1539
rect 11627 1505 11665 1539
rect 11699 1505 11737 1539
rect 11771 1505 11835 1539
rect 11869 1505 11907 1539
rect 11941 1505 11979 1539
rect 12013 1505 12051 1539
rect 12085 1505 12123 1539
rect 12157 1505 12195 1539
rect 12229 1505 12339 1539
rect 12373 1505 12411 1539
rect 12445 1505 12483 1539
rect 12517 1505 12555 1539
rect 12589 1505 12645 1539
rect 12679 1505 12717 1539
rect 12751 1505 12789 1539
rect 12823 1505 12861 1539
rect 12895 1505 13005 1539
rect 13039 1505 13077 1539
rect 13111 1505 13149 1539
rect 13183 1505 13221 1539
rect 13255 1505 13293 1539
rect 13327 1505 13365 1539
rect 13399 1505 13463 1539
rect 13497 1505 13535 1539
rect 13569 1505 13607 1539
rect 13641 1505 13679 1539
rect 13713 1505 13751 1539
rect 13785 1505 13823 1539
rect 13857 1505 13967 1539
rect 14001 1505 14039 1539
rect 14073 1505 14111 1539
rect 14145 1505 14183 1539
rect 14217 1505 14255 1539
rect 14289 1505 14327 1539
rect 14361 1505 14425 1539
rect 14459 1505 14497 1539
rect 14531 1505 14569 1539
rect 14603 1505 14641 1539
rect 14675 1505 14713 1539
rect 14747 1505 14785 1539
rect 14819 1505 14929 1539
rect 14963 1505 15001 1539
rect 15035 1505 15073 1539
rect 15107 1505 15145 1539
rect 15179 1505 15235 1539
rect 15269 1505 15307 1539
rect 15341 1505 15379 1539
rect 15413 1505 15451 1539
rect 15485 1505 15595 1539
rect 15629 1505 15667 1539
rect 15701 1505 15739 1539
rect 15773 1505 15811 1539
rect 15845 1505 15901 1539
rect 15935 1505 15973 1539
rect 16007 1505 16045 1539
rect 16079 1505 16117 1539
rect 16151 1505 16261 1539
rect 16295 1505 16333 1539
rect 16367 1505 16405 1539
rect 16439 1505 16477 1539
rect 16511 1505 16567 1539
rect 16601 1505 16639 1539
rect 16673 1505 16711 1539
rect 16745 1505 16783 1539
rect 16817 1505 16927 1539
rect 16961 1505 16999 1539
rect 17033 1505 17071 1539
rect 17105 1505 17143 1539
rect 17177 1505 17233 1539
rect 17267 1505 17305 1539
rect 17339 1505 17377 1539
rect 17411 1505 17449 1539
rect 17483 1505 17593 1539
rect 17627 1505 17665 1539
rect 17699 1505 17743 1539
rect 17777 1505 17821 1539
rect 17855 1505 17893 1539
rect 17927 1505 18013 1539
rect -31 1470 31 1505
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect 931 1470 993 1505
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect -31 1038 31 1076
rect 931 1436 945 1470
rect 979 1436 993 1470
rect 1893 1470 1955 1505
rect 931 1398 993 1436
rect 931 1364 945 1398
rect 979 1364 993 1398
rect 931 1326 993 1364
rect 931 1292 945 1326
rect 979 1292 993 1326
rect 931 1254 993 1292
rect 931 1220 945 1254
rect 979 1220 993 1254
rect 931 1182 993 1220
rect 931 1148 945 1182
rect 979 1148 993 1182
rect 931 1110 993 1148
rect 931 1076 945 1110
rect 979 1076 993 1110
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect 931 1038 993 1076
rect 1893 1436 1907 1470
rect 1941 1436 1955 1470
rect 2559 1470 2621 1505
rect 1893 1398 1955 1436
rect 1893 1364 1907 1398
rect 1941 1364 1955 1398
rect 1893 1326 1955 1364
rect 1893 1292 1907 1326
rect 1941 1292 1955 1326
rect 1893 1254 1955 1292
rect 1893 1220 1907 1254
rect 1941 1220 1955 1254
rect 1893 1182 1955 1220
rect 1893 1148 1907 1182
rect 1941 1148 1955 1182
rect 1893 1110 1955 1148
rect 1893 1076 1907 1110
rect 1941 1076 1955 1110
rect 931 1004 945 1038
rect 979 1004 993 1038
rect 931 966 993 1004
rect -31 930 31 932
rect 931 932 945 966
rect 979 932 993 966
rect 1893 1038 1955 1076
rect 2559 1436 2573 1470
rect 2607 1436 2621 1470
rect 3521 1470 3583 1505
rect 2559 1398 2621 1436
rect 2559 1364 2573 1398
rect 2607 1364 2621 1398
rect 2559 1326 2621 1364
rect 2559 1292 2573 1326
rect 2607 1292 2621 1326
rect 2559 1254 2621 1292
rect 2559 1220 2573 1254
rect 2607 1220 2621 1254
rect 2559 1182 2621 1220
rect 2559 1148 2573 1182
rect 2607 1148 2621 1182
rect 2559 1110 2621 1148
rect 2559 1076 2573 1110
rect 2607 1076 2621 1110
rect 1893 1004 1907 1038
rect 1941 1004 1955 1038
rect 1893 966 1955 1004
rect 931 930 993 932
rect 1893 932 1907 966
rect 1941 932 1955 966
rect 2559 1038 2621 1076
rect 3521 1436 3535 1470
rect 3569 1436 3583 1470
rect 4483 1470 4545 1505
rect 3521 1398 3583 1436
rect 3521 1364 3535 1398
rect 3569 1364 3583 1398
rect 3521 1326 3583 1364
rect 3521 1292 3535 1326
rect 3569 1292 3583 1326
rect 3521 1254 3583 1292
rect 3521 1220 3535 1254
rect 3569 1220 3583 1254
rect 3521 1182 3583 1220
rect 3521 1148 3535 1182
rect 3569 1148 3583 1182
rect 3521 1110 3583 1148
rect 3521 1076 3535 1110
rect 3569 1076 3583 1110
rect 2559 1004 2573 1038
rect 2607 1004 2621 1038
rect 2559 966 2621 1004
rect 1893 930 1955 932
rect 2559 932 2573 966
rect 2607 932 2621 966
rect 3521 1038 3583 1076
rect 4483 1436 4497 1470
rect 4531 1436 4545 1470
rect 5149 1470 5211 1505
rect 4483 1398 4545 1436
rect 4483 1364 4497 1398
rect 4531 1364 4545 1398
rect 4483 1326 4545 1364
rect 4483 1292 4497 1326
rect 4531 1292 4545 1326
rect 4483 1254 4545 1292
rect 4483 1220 4497 1254
rect 4531 1220 4545 1254
rect 4483 1182 4545 1220
rect 4483 1148 4497 1182
rect 4531 1148 4545 1182
rect 4483 1110 4545 1148
rect 4483 1076 4497 1110
rect 4531 1076 4545 1110
rect 3521 1004 3535 1038
rect 3569 1004 3583 1038
rect 3521 966 3583 1004
rect 2559 930 2621 932
rect 3521 932 3535 966
rect 3569 932 3583 966
rect 4483 1038 4545 1076
rect 5149 1436 5163 1470
rect 5197 1436 5211 1470
rect 6111 1470 6173 1505
rect 5149 1398 5211 1436
rect 5149 1364 5163 1398
rect 5197 1364 5211 1398
rect 5149 1326 5211 1364
rect 5149 1292 5163 1326
rect 5197 1292 5211 1326
rect 5149 1254 5211 1292
rect 5149 1220 5163 1254
rect 5197 1220 5211 1254
rect 5149 1182 5211 1220
rect 5149 1148 5163 1182
rect 5197 1148 5211 1182
rect 5149 1110 5211 1148
rect 5149 1076 5163 1110
rect 5197 1076 5211 1110
rect 4483 1004 4497 1038
rect 4531 1004 4545 1038
rect 4483 966 4545 1004
rect 3521 930 3583 932
rect 4483 932 4497 966
rect 4531 932 4545 966
rect 5149 1038 5211 1076
rect 6111 1436 6125 1470
rect 6159 1436 6173 1470
rect 7073 1470 7135 1505
rect 6111 1398 6173 1436
rect 6111 1364 6125 1398
rect 6159 1364 6173 1398
rect 6111 1326 6173 1364
rect 6111 1292 6125 1326
rect 6159 1292 6173 1326
rect 6111 1254 6173 1292
rect 6111 1220 6125 1254
rect 6159 1220 6173 1254
rect 6111 1182 6173 1220
rect 6111 1148 6125 1182
rect 6159 1148 6173 1182
rect 6111 1110 6173 1148
rect 6111 1076 6125 1110
rect 6159 1076 6173 1110
rect 5149 1004 5163 1038
rect 5197 1004 5211 1038
rect 5149 966 5211 1004
rect 4483 930 4545 932
rect 5149 932 5163 966
rect 5197 932 5211 966
rect 6111 1038 6173 1076
rect 7073 1436 7087 1470
rect 7121 1436 7135 1470
rect 7739 1470 7801 1505
rect 7073 1398 7135 1436
rect 7073 1364 7087 1398
rect 7121 1364 7135 1398
rect 7073 1326 7135 1364
rect 7073 1292 7087 1326
rect 7121 1292 7135 1326
rect 7073 1254 7135 1292
rect 7073 1220 7087 1254
rect 7121 1220 7135 1254
rect 7073 1182 7135 1220
rect 7073 1148 7087 1182
rect 7121 1148 7135 1182
rect 7073 1110 7135 1148
rect 7073 1076 7087 1110
rect 7121 1076 7135 1110
rect 6111 1004 6125 1038
rect 6159 1004 6173 1038
rect 6111 966 6173 1004
rect 5149 930 5211 932
rect 6111 932 6125 966
rect 6159 932 6173 966
rect 7073 1038 7135 1076
rect 7739 1436 7753 1470
rect 7787 1436 7801 1470
rect 8701 1470 8763 1505
rect 7739 1398 7801 1436
rect 7739 1364 7753 1398
rect 7787 1364 7801 1398
rect 7739 1326 7801 1364
rect 7739 1292 7753 1326
rect 7787 1292 7801 1326
rect 7739 1254 7801 1292
rect 7739 1220 7753 1254
rect 7787 1220 7801 1254
rect 7739 1182 7801 1220
rect 7739 1148 7753 1182
rect 7787 1148 7801 1182
rect 7739 1110 7801 1148
rect 7739 1076 7753 1110
rect 7787 1076 7801 1110
rect 7073 1004 7087 1038
rect 7121 1004 7135 1038
rect 7073 966 7135 1004
rect 6111 930 6173 932
rect 7073 932 7087 966
rect 7121 932 7135 966
rect 7739 1038 7801 1076
rect 8701 1436 8715 1470
rect 8749 1436 8763 1470
rect 9663 1470 9725 1505
rect 8701 1398 8763 1436
rect 8701 1364 8715 1398
rect 8749 1364 8763 1398
rect 8701 1326 8763 1364
rect 8701 1292 8715 1326
rect 8749 1292 8763 1326
rect 8701 1254 8763 1292
rect 8701 1220 8715 1254
rect 8749 1220 8763 1254
rect 8701 1182 8763 1220
rect 8701 1148 8715 1182
rect 8749 1148 8763 1182
rect 8701 1110 8763 1148
rect 8701 1076 8715 1110
rect 8749 1076 8763 1110
rect 7739 1004 7753 1038
rect 7787 1004 7801 1038
rect 7739 966 7801 1004
rect 7073 930 7135 932
rect 7739 932 7753 966
rect 7787 932 7801 966
rect 8701 1038 8763 1076
rect 9663 1436 9677 1470
rect 9711 1436 9725 1470
rect 10329 1470 10391 1505
rect 9663 1398 9725 1436
rect 9663 1364 9677 1398
rect 9711 1364 9725 1398
rect 9663 1326 9725 1364
rect 9663 1292 9677 1326
rect 9711 1292 9725 1326
rect 9663 1254 9725 1292
rect 9663 1220 9677 1254
rect 9711 1220 9725 1254
rect 9663 1182 9725 1220
rect 9663 1148 9677 1182
rect 9711 1148 9725 1182
rect 9663 1110 9725 1148
rect 9663 1076 9677 1110
rect 9711 1076 9725 1110
rect 8701 1004 8715 1038
rect 8749 1004 8763 1038
rect 8701 966 8763 1004
rect 7739 930 7801 932
rect 8701 932 8715 966
rect 8749 932 8763 966
rect 9663 1038 9725 1076
rect 10329 1436 10343 1470
rect 10377 1436 10391 1470
rect 11291 1470 11353 1505
rect 10329 1398 10391 1436
rect 10329 1364 10343 1398
rect 10377 1364 10391 1398
rect 10329 1326 10391 1364
rect 10329 1292 10343 1326
rect 10377 1292 10391 1326
rect 10329 1254 10391 1292
rect 10329 1220 10343 1254
rect 10377 1220 10391 1254
rect 10329 1182 10391 1220
rect 10329 1148 10343 1182
rect 10377 1148 10391 1182
rect 10329 1110 10391 1148
rect 10329 1076 10343 1110
rect 10377 1076 10391 1110
rect 9663 1004 9677 1038
rect 9711 1004 9725 1038
rect 9663 966 9725 1004
rect 8701 930 8763 932
rect 9663 932 9677 966
rect 9711 932 9725 966
rect 10329 1038 10391 1076
rect 11291 1436 11305 1470
rect 11339 1436 11353 1470
rect 12253 1470 12315 1505
rect 11291 1398 11353 1436
rect 11291 1364 11305 1398
rect 11339 1364 11353 1398
rect 11291 1326 11353 1364
rect 11291 1292 11305 1326
rect 11339 1292 11353 1326
rect 11291 1254 11353 1292
rect 11291 1220 11305 1254
rect 11339 1220 11353 1254
rect 11291 1182 11353 1220
rect 11291 1148 11305 1182
rect 11339 1148 11353 1182
rect 11291 1110 11353 1148
rect 11291 1076 11305 1110
rect 11339 1076 11353 1110
rect 10329 1004 10343 1038
rect 10377 1004 10391 1038
rect 10329 966 10391 1004
rect 9663 930 9725 932
rect 10329 932 10343 966
rect 10377 932 10391 966
rect 11291 1038 11353 1076
rect 12253 1436 12267 1470
rect 12301 1436 12315 1470
rect 12919 1470 12981 1505
rect 12253 1398 12315 1436
rect 12253 1364 12267 1398
rect 12301 1364 12315 1398
rect 12253 1326 12315 1364
rect 12253 1292 12267 1326
rect 12301 1292 12315 1326
rect 12253 1254 12315 1292
rect 12253 1220 12267 1254
rect 12301 1220 12315 1254
rect 12253 1182 12315 1220
rect 12253 1148 12267 1182
rect 12301 1148 12315 1182
rect 12253 1110 12315 1148
rect 12253 1076 12267 1110
rect 12301 1076 12315 1110
rect 11291 1004 11305 1038
rect 11339 1004 11353 1038
rect 11291 966 11353 1004
rect 10329 930 10391 932
rect 11291 932 11305 966
rect 11339 932 11353 966
rect 12253 1038 12315 1076
rect 12919 1436 12933 1470
rect 12967 1436 12981 1470
rect 13881 1470 13943 1505
rect 12919 1398 12981 1436
rect 12919 1364 12933 1398
rect 12967 1364 12981 1398
rect 12919 1326 12981 1364
rect 12919 1292 12933 1326
rect 12967 1292 12981 1326
rect 12919 1254 12981 1292
rect 12919 1220 12933 1254
rect 12967 1220 12981 1254
rect 12919 1182 12981 1220
rect 12919 1148 12933 1182
rect 12967 1148 12981 1182
rect 12919 1110 12981 1148
rect 12919 1076 12933 1110
rect 12967 1076 12981 1110
rect 12253 1004 12267 1038
rect 12301 1004 12315 1038
rect 12253 966 12315 1004
rect 11291 930 11353 932
rect 12253 932 12267 966
rect 12301 932 12315 966
rect 12919 1038 12981 1076
rect 13881 1436 13895 1470
rect 13929 1436 13943 1470
rect 14843 1470 14905 1505
rect 13881 1398 13943 1436
rect 13881 1364 13895 1398
rect 13929 1364 13943 1398
rect 13881 1326 13943 1364
rect 13881 1292 13895 1326
rect 13929 1292 13943 1326
rect 13881 1254 13943 1292
rect 13881 1220 13895 1254
rect 13929 1220 13943 1254
rect 13881 1182 13943 1220
rect 13881 1148 13895 1182
rect 13929 1148 13943 1182
rect 13881 1110 13943 1148
rect 13881 1076 13895 1110
rect 13929 1076 13943 1110
rect 12919 1004 12933 1038
rect 12967 1004 12981 1038
rect 12919 966 12981 1004
rect 12253 930 12315 932
rect 12919 932 12933 966
rect 12967 932 12981 966
rect 13881 1038 13943 1076
rect 14843 1436 14857 1470
rect 14891 1436 14905 1470
rect 15509 1470 15571 1505
rect 14843 1398 14905 1436
rect 14843 1364 14857 1398
rect 14891 1364 14905 1398
rect 14843 1326 14905 1364
rect 14843 1292 14857 1326
rect 14891 1292 14905 1326
rect 14843 1254 14905 1292
rect 14843 1220 14857 1254
rect 14891 1220 14905 1254
rect 14843 1182 14905 1220
rect 14843 1148 14857 1182
rect 14891 1148 14905 1182
rect 14843 1110 14905 1148
rect 14843 1076 14857 1110
rect 14891 1076 14905 1110
rect 13881 1004 13895 1038
rect 13929 1004 13943 1038
rect 13881 966 13943 1004
rect 12919 930 12981 932
rect 13881 932 13895 966
rect 13929 932 13943 966
rect 14843 1038 14905 1076
rect 15509 1436 15523 1470
rect 15557 1436 15571 1470
rect 16175 1470 16237 1505
rect 15509 1398 15571 1436
rect 15509 1364 15523 1398
rect 15557 1364 15571 1398
rect 15509 1326 15571 1364
rect 15509 1292 15523 1326
rect 15557 1292 15571 1326
rect 15509 1254 15571 1292
rect 15509 1220 15523 1254
rect 15557 1220 15571 1254
rect 15509 1182 15571 1220
rect 15509 1148 15523 1182
rect 15557 1148 15571 1182
rect 15509 1110 15571 1148
rect 15509 1076 15523 1110
rect 15557 1076 15571 1110
rect 14843 1004 14857 1038
rect 14891 1004 14905 1038
rect 14843 966 14905 1004
rect 13881 930 13943 932
rect 14843 932 14857 966
rect 14891 932 14905 966
rect 15509 1038 15571 1076
rect 16175 1436 16189 1470
rect 16223 1436 16237 1470
rect 16841 1470 16903 1505
rect 16175 1398 16237 1436
rect 16175 1364 16189 1398
rect 16223 1364 16237 1398
rect 16175 1326 16237 1364
rect 16175 1292 16189 1326
rect 16223 1292 16237 1326
rect 16175 1254 16237 1292
rect 16175 1220 16189 1254
rect 16223 1220 16237 1254
rect 16175 1182 16237 1220
rect 16175 1148 16189 1182
rect 16223 1148 16237 1182
rect 16175 1110 16237 1148
rect 16175 1076 16189 1110
rect 16223 1076 16237 1110
rect 15509 1004 15523 1038
rect 15557 1004 15571 1038
rect 15509 966 15571 1004
rect 14843 930 14905 932
rect 15509 932 15523 966
rect 15557 932 15571 966
rect 16175 1038 16237 1076
rect 16841 1436 16855 1470
rect 16889 1436 16903 1470
rect 17507 1470 17569 1505
rect 16841 1398 16903 1436
rect 16841 1364 16855 1398
rect 16889 1364 16903 1398
rect 16841 1326 16903 1364
rect 16841 1292 16855 1326
rect 16889 1292 16903 1326
rect 16841 1254 16903 1292
rect 16841 1220 16855 1254
rect 16889 1220 16903 1254
rect 16841 1182 16903 1220
rect 16841 1148 16855 1182
rect 16889 1148 16903 1182
rect 16841 1110 16903 1148
rect 16841 1076 16855 1110
rect 16889 1076 16903 1110
rect 16175 1004 16189 1038
rect 16223 1004 16237 1038
rect 16175 966 16237 1004
rect 15509 930 15571 932
rect 16175 932 16189 966
rect 16223 932 16237 966
rect 16841 1038 16903 1076
rect 17507 1436 17521 1470
rect 17555 1436 17569 1470
rect 17951 1470 18013 1505
rect 17507 1398 17569 1436
rect 17507 1364 17521 1398
rect 17555 1364 17569 1398
rect 17507 1326 17569 1364
rect 17507 1292 17521 1326
rect 17555 1292 17569 1326
rect 17507 1254 17569 1292
rect 17507 1220 17521 1254
rect 17555 1220 17569 1254
rect 17507 1182 17569 1220
rect 17507 1148 17521 1182
rect 17555 1148 17569 1182
rect 17507 1110 17569 1148
rect 17507 1076 17521 1110
rect 17555 1076 17569 1110
rect 16841 1004 16855 1038
rect 16889 1004 16903 1038
rect 16841 966 16903 1004
rect 16175 930 16237 932
rect 16841 932 16855 966
rect 16889 932 16903 966
rect 17507 1038 17569 1076
rect 17951 1436 17965 1470
rect 17999 1436 18013 1470
rect 17951 1398 18013 1436
rect 17951 1364 17965 1398
rect 17999 1364 18013 1398
rect 17951 1326 18013 1364
rect 17951 1292 17965 1326
rect 17999 1292 18013 1326
rect 17951 1254 18013 1292
rect 17951 1220 17965 1254
rect 17999 1220 18013 1254
rect 17951 1182 18013 1220
rect 17951 1148 17965 1182
rect 17999 1148 18013 1182
rect 17951 1110 18013 1148
rect 17951 1076 17965 1110
rect 17999 1076 18013 1110
rect 17507 1004 17521 1038
rect 17555 1004 17569 1038
rect 17507 966 17569 1004
rect 16841 930 16903 932
rect 17507 932 17521 966
rect 17555 932 17569 966
rect 17951 1038 18013 1076
rect 17951 1004 17965 1038
rect 17999 1004 18013 1038
rect 17951 966 18013 1004
rect 17507 930 17569 932
rect 17951 932 17965 966
rect 17999 932 18013 966
rect 17951 930 18013 932
rect -31 868 18013 930
<< psubdiffcont >>
rect -17 512 17 546
rect 945 512 979 546
rect 1907 512 1941 546
rect 2573 512 2607 546
rect 3535 512 3569 546
rect 4497 512 4531 546
rect 5163 512 5197 546
rect 6125 512 6159 546
rect 7087 512 7121 546
rect 7753 512 7787 546
rect 8715 512 8749 546
rect 9677 512 9711 546
rect 10343 512 10377 546
rect 11305 512 11339 546
rect 12267 512 12301 546
rect 12933 512 12967 546
rect 13895 512 13929 546
rect 14857 512 14891 546
rect 15523 512 15557 546
rect 16189 512 16223 546
rect 16855 512 16889 546
rect 17521 512 17555 546
rect 17965 512 17999 546
rect -17 440 17 474
rect -17 368 17 402
rect 945 440 979 474
rect -17 296 17 330
rect -17 224 17 258
rect -17 152 17 186
rect -17 80 17 114
rect 945 368 979 402
rect 1907 440 1941 474
rect 945 296 979 330
rect 945 224 979 258
rect 945 152 979 186
rect 945 80 979 114
rect 1907 368 1941 402
rect 2573 440 2607 474
rect 1907 296 1941 330
rect 1907 224 1941 258
rect 1907 152 1941 186
rect 1907 80 1941 114
rect 2573 368 2607 402
rect 3535 440 3569 474
rect 2573 296 2607 330
rect 2573 224 2607 258
rect 2573 152 2607 186
rect 2573 80 2607 114
rect 3535 368 3569 402
rect 4497 440 4531 474
rect 3535 296 3569 330
rect 3535 224 3569 258
rect 3535 152 3569 186
rect 3535 80 3569 114
rect 4497 368 4531 402
rect 5163 440 5197 474
rect 4497 296 4531 330
rect 4497 224 4531 258
rect 4497 152 4531 186
rect 4497 80 4531 114
rect 5163 368 5197 402
rect 6125 440 6159 474
rect 5163 296 5197 330
rect 5163 224 5197 258
rect 5163 152 5197 186
rect 5163 80 5197 114
rect 6125 368 6159 402
rect 7087 440 7121 474
rect 6125 296 6159 330
rect 6125 224 6159 258
rect 6125 152 6159 186
rect 6125 80 6159 114
rect 7087 368 7121 402
rect 7753 440 7787 474
rect 7087 296 7121 330
rect 7087 224 7121 258
rect 7087 152 7121 186
rect 7087 80 7121 114
rect 7753 368 7787 402
rect 8715 440 8749 474
rect 7753 296 7787 330
rect 7753 224 7787 258
rect 7753 152 7787 186
rect 7753 80 7787 114
rect 8715 368 8749 402
rect 9677 440 9711 474
rect 8715 296 8749 330
rect 8715 224 8749 258
rect 8715 152 8749 186
rect 8715 80 8749 114
rect 9677 368 9711 402
rect 10343 440 10377 474
rect 9677 296 9711 330
rect 9677 224 9711 258
rect 9677 152 9711 186
rect 9677 80 9711 114
rect 10343 368 10377 402
rect 11305 440 11339 474
rect 10343 296 10377 330
rect 10343 224 10377 258
rect 10343 152 10377 186
rect 10343 80 10377 114
rect 11305 368 11339 402
rect 12267 440 12301 474
rect 11305 296 11339 330
rect 11305 224 11339 258
rect 11305 152 11339 186
rect 11305 80 11339 114
rect 12267 368 12301 402
rect 12933 440 12967 474
rect 12267 296 12301 330
rect 12267 224 12301 258
rect 12267 152 12301 186
rect 12267 80 12301 114
rect 12933 368 12967 402
rect 13895 440 13929 474
rect 12933 296 12967 330
rect 12933 224 12967 258
rect 12933 152 12967 186
rect 12933 80 12967 114
rect 13895 368 13929 402
rect 14857 440 14891 474
rect 13895 296 13929 330
rect 13895 224 13929 258
rect 13895 152 13929 186
rect 13895 80 13929 114
rect 14857 368 14891 402
rect 15523 440 15557 474
rect 16189 440 16223 474
rect 14857 296 14891 330
rect 14857 224 14891 258
rect 14857 152 14891 186
rect 14857 80 14891 114
rect 15523 368 15557 402
rect 15523 296 15557 330
rect 15523 224 15557 258
rect 15523 152 15557 186
rect 15523 80 15557 114
rect 16189 368 16223 402
rect 16855 440 16889 474
rect 17521 440 17555 474
rect 16189 296 16223 330
rect 16189 224 16223 258
rect 16189 152 16223 186
rect 16189 80 16223 114
rect 16855 368 16889 402
rect 16855 296 16889 330
rect 16855 224 16889 258
rect 16855 152 16889 186
rect 16855 80 16889 114
rect 17521 368 17555 402
rect 17965 440 17999 474
rect 17521 296 17555 330
rect 17521 224 17555 258
rect 17521 152 17555 186
rect 17521 80 17555 114
rect 17965 368 17999 402
rect 17965 296 17999 330
rect 17965 224 17999 258
rect 17965 152 17999 186
rect 17965 80 17999 114
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 343 13 377 47
rect 415 13 449 47
rect 513 13 547 47
rect 585 13 619 47
rect 657 13 691 47
rect 729 13 763 47
rect 801 13 835 47
rect 873 13 907 47
rect 1017 13 1051 47
rect 1089 13 1123 47
rect 1161 13 1195 47
rect 1233 13 1267 47
rect 1305 13 1339 47
rect 1377 13 1411 47
rect 1475 13 1509 47
rect 1547 13 1581 47
rect 1619 13 1653 47
rect 1691 13 1725 47
rect 1763 13 1797 47
rect 1835 13 1869 47
rect 1979 13 2013 47
rect 2051 13 2085 47
rect 2123 13 2157 47
rect 2195 13 2229 47
rect 2285 13 2319 47
rect 2357 13 2391 47
rect 2429 13 2463 47
rect 2501 13 2535 47
rect 2645 13 2679 47
rect 2717 13 2751 47
rect 2789 13 2823 47
rect 2861 13 2895 47
rect 2933 13 2967 47
rect 3005 13 3039 47
rect 3103 13 3137 47
rect 3175 13 3209 47
rect 3247 13 3281 47
rect 3319 13 3353 47
rect 3391 13 3425 47
rect 3463 13 3497 47
rect 3607 13 3641 47
rect 3679 13 3713 47
rect 3751 13 3785 47
rect 3823 13 3857 47
rect 3895 13 3929 47
rect 3967 13 4001 47
rect 4065 13 4099 47
rect 4137 13 4171 47
rect 4209 13 4243 47
rect 4281 13 4315 47
rect 4353 13 4387 47
rect 4425 13 4459 47
rect 4569 13 4603 47
rect 4641 13 4675 47
rect 4713 13 4747 47
rect 4785 13 4819 47
rect 4875 13 4909 47
rect 4947 13 4981 47
rect 5019 13 5053 47
rect 5091 13 5125 47
rect 5235 13 5269 47
rect 5307 13 5341 47
rect 5379 13 5413 47
rect 5451 13 5485 47
rect 5523 13 5557 47
rect 5595 13 5629 47
rect 5693 13 5727 47
rect 5765 13 5799 47
rect 5837 13 5871 47
rect 5909 13 5943 47
rect 5981 13 6015 47
rect 6053 13 6087 47
rect 6197 13 6231 47
rect 6269 13 6303 47
rect 6341 13 6375 47
rect 6413 13 6447 47
rect 6485 13 6519 47
rect 6557 13 6591 47
rect 6655 13 6689 47
rect 6727 13 6761 47
rect 6799 13 6833 47
rect 6871 13 6905 47
rect 6943 13 6977 47
rect 7015 13 7049 47
rect 7159 13 7193 47
rect 7231 13 7265 47
rect 7303 13 7337 47
rect 7375 13 7409 47
rect 7465 13 7499 47
rect 7537 13 7571 47
rect 7609 13 7643 47
rect 7681 13 7715 47
rect 7825 13 7859 47
rect 7897 13 7931 47
rect 7969 13 8003 47
rect 8041 13 8075 47
rect 8113 13 8147 47
rect 8185 13 8219 47
rect 8283 13 8317 47
rect 8355 13 8389 47
rect 8427 13 8461 47
rect 8499 13 8533 47
rect 8571 13 8605 47
rect 8643 13 8677 47
rect 8787 13 8821 47
rect 8859 13 8893 47
rect 8931 13 8965 47
rect 9003 13 9037 47
rect 9075 13 9109 47
rect 9147 13 9181 47
rect 9245 13 9279 47
rect 9317 13 9351 47
rect 9389 13 9423 47
rect 9461 13 9495 47
rect 9533 13 9567 47
rect 9605 13 9639 47
rect 9749 13 9783 47
rect 9821 13 9855 47
rect 9893 13 9927 47
rect 9965 13 9999 47
rect 10055 13 10089 47
rect 10127 13 10161 47
rect 10199 13 10233 47
rect 10271 13 10305 47
rect 10415 13 10449 47
rect 10487 13 10521 47
rect 10559 13 10593 47
rect 10631 13 10665 47
rect 10703 13 10737 47
rect 10775 13 10809 47
rect 10873 13 10907 47
rect 10945 13 10979 47
rect 11017 13 11051 47
rect 11089 13 11123 47
rect 11161 13 11195 47
rect 11233 13 11267 47
rect 11377 13 11411 47
rect 11449 13 11483 47
rect 11521 13 11555 47
rect 11593 13 11627 47
rect 11665 13 11699 47
rect 11737 13 11771 47
rect 11835 13 11869 47
rect 11907 13 11941 47
rect 11979 13 12013 47
rect 12051 13 12085 47
rect 12123 13 12157 47
rect 12195 13 12229 47
rect 12339 13 12373 47
rect 12411 13 12445 47
rect 12483 13 12517 47
rect 12555 13 12589 47
rect 12645 13 12679 47
rect 12717 13 12751 47
rect 12789 13 12823 47
rect 12861 13 12895 47
rect 13005 13 13039 47
rect 13077 13 13111 47
rect 13149 13 13183 47
rect 13221 13 13255 47
rect 13293 13 13327 47
rect 13365 13 13399 47
rect 13463 13 13497 47
rect 13535 13 13569 47
rect 13607 13 13641 47
rect 13679 13 13713 47
rect 13751 13 13785 47
rect 13823 13 13857 47
rect 13967 13 14001 47
rect 14039 13 14073 47
rect 14111 13 14145 47
rect 14183 13 14217 47
rect 14255 13 14289 47
rect 14327 13 14361 47
rect 14425 13 14459 47
rect 14497 13 14531 47
rect 14569 13 14603 47
rect 14641 13 14675 47
rect 14713 13 14747 47
rect 14785 13 14819 47
rect 14929 13 14963 47
rect 15001 13 15035 47
rect 15073 13 15107 47
rect 15145 13 15179 47
rect 15235 13 15269 47
rect 15307 13 15341 47
rect 15379 13 15413 47
rect 15451 13 15485 47
rect 15595 13 15629 47
rect 15667 13 15701 47
rect 15739 13 15773 47
rect 15811 13 15845 47
rect 15901 13 15935 47
rect 15973 13 16007 47
rect 16045 13 16079 47
rect 16117 13 16151 47
rect 16261 13 16295 47
rect 16333 13 16367 47
rect 16405 13 16439 47
rect 16477 13 16511 47
rect 16567 13 16601 47
rect 16639 13 16673 47
rect 16711 13 16745 47
rect 16783 13 16817 47
rect 16927 13 16961 47
rect 16999 13 17033 47
rect 17071 13 17105 47
rect 17143 13 17177 47
rect 17233 13 17267 47
rect 17305 13 17339 47
rect 17377 13 17411 47
rect 17449 13 17483 47
rect 17593 13 17627 47
rect 17665 13 17699 47
rect 17743 13 17777 47
rect 17821 13 17855 47
rect 17893 13 17927 47
<< nsubdiffcont >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 343 1505 377 1539
rect 415 1505 449 1539
rect 513 1505 547 1539
rect 585 1505 619 1539
rect 657 1505 691 1539
rect 729 1505 763 1539
rect 801 1505 835 1539
rect 873 1505 907 1539
rect 1017 1505 1051 1539
rect 1089 1505 1123 1539
rect 1161 1505 1195 1539
rect 1233 1505 1267 1539
rect 1305 1505 1339 1539
rect 1377 1505 1411 1539
rect 1475 1505 1509 1539
rect 1547 1505 1581 1539
rect 1619 1505 1653 1539
rect 1691 1505 1725 1539
rect 1763 1505 1797 1539
rect 1835 1505 1869 1539
rect 1979 1505 2013 1539
rect 2051 1505 2085 1539
rect 2123 1505 2157 1539
rect 2195 1505 2229 1539
rect 2285 1505 2319 1539
rect 2357 1505 2391 1539
rect 2429 1505 2463 1539
rect 2501 1505 2535 1539
rect 2645 1505 2679 1539
rect 2717 1505 2751 1539
rect 2789 1505 2823 1539
rect 2861 1505 2895 1539
rect 2933 1505 2967 1539
rect 3005 1505 3039 1539
rect 3103 1505 3137 1539
rect 3175 1505 3209 1539
rect 3247 1505 3281 1539
rect 3319 1505 3353 1539
rect 3391 1505 3425 1539
rect 3463 1505 3497 1539
rect 3607 1505 3641 1539
rect 3679 1505 3713 1539
rect 3751 1505 3785 1539
rect 3823 1505 3857 1539
rect 3895 1505 3929 1539
rect 3967 1505 4001 1539
rect 4065 1505 4099 1539
rect 4137 1505 4171 1539
rect 4209 1505 4243 1539
rect 4281 1505 4315 1539
rect 4353 1505 4387 1539
rect 4425 1505 4459 1539
rect 4569 1505 4603 1539
rect 4641 1505 4675 1539
rect 4713 1505 4747 1539
rect 4785 1505 4819 1539
rect 4875 1505 4909 1539
rect 4947 1505 4981 1539
rect 5019 1505 5053 1539
rect 5091 1505 5125 1539
rect 5235 1505 5269 1539
rect 5307 1505 5341 1539
rect 5379 1505 5413 1539
rect 5451 1505 5485 1539
rect 5523 1505 5557 1539
rect 5595 1505 5629 1539
rect 5693 1505 5727 1539
rect 5765 1505 5799 1539
rect 5837 1505 5871 1539
rect 5909 1505 5943 1539
rect 5981 1505 6015 1539
rect 6053 1505 6087 1539
rect 6197 1505 6231 1539
rect 6269 1505 6303 1539
rect 6341 1505 6375 1539
rect 6413 1505 6447 1539
rect 6485 1505 6519 1539
rect 6557 1505 6591 1539
rect 6655 1505 6689 1539
rect 6727 1505 6761 1539
rect 6799 1505 6833 1539
rect 6871 1505 6905 1539
rect 6943 1505 6977 1539
rect 7015 1505 7049 1539
rect 7159 1505 7193 1539
rect 7231 1505 7265 1539
rect 7303 1505 7337 1539
rect 7375 1505 7409 1539
rect 7465 1505 7499 1539
rect 7537 1505 7571 1539
rect 7609 1505 7643 1539
rect 7681 1505 7715 1539
rect 7825 1505 7859 1539
rect 7897 1505 7931 1539
rect 7969 1505 8003 1539
rect 8041 1505 8075 1539
rect 8113 1505 8147 1539
rect 8185 1505 8219 1539
rect 8283 1505 8317 1539
rect 8355 1505 8389 1539
rect 8427 1505 8461 1539
rect 8499 1505 8533 1539
rect 8571 1505 8605 1539
rect 8643 1505 8677 1539
rect 8787 1505 8821 1539
rect 8859 1505 8893 1539
rect 8931 1505 8965 1539
rect 9003 1505 9037 1539
rect 9075 1505 9109 1539
rect 9147 1505 9181 1539
rect 9245 1505 9279 1539
rect 9317 1505 9351 1539
rect 9389 1505 9423 1539
rect 9461 1505 9495 1539
rect 9533 1505 9567 1539
rect 9605 1505 9639 1539
rect 9749 1505 9783 1539
rect 9821 1505 9855 1539
rect 9893 1505 9927 1539
rect 9965 1505 9999 1539
rect 10055 1505 10089 1539
rect 10127 1505 10161 1539
rect 10199 1505 10233 1539
rect 10271 1505 10305 1539
rect 10415 1505 10449 1539
rect 10487 1505 10521 1539
rect 10559 1505 10593 1539
rect 10631 1505 10665 1539
rect 10703 1505 10737 1539
rect 10775 1505 10809 1539
rect 10873 1505 10907 1539
rect 10945 1505 10979 1539
rect 11017 1505 11051 1539
rect 11089 1505 11123 1539
rect 11161 1505 11195 1539
rect 11233 1505 11267 1539
rect 11377 1505 11411 1539
rect 11449 1505 11483 1539
rect 11521 1505 11555 1539
rect 11593 1505 11627 1539
rect 11665 1505 11699 1539
rect 11737 1505 11771 1539
rect 11835 1505 11869 1539
rect 11907 1505 11941 1539
rect 11979 1505 12013 1539
rect 12051 1505 12085 1539
rect 12123 1505 12157 1539
rect 12195 1505 12229 1539
rect 12339 1505 12373 1539
rect 12411 1505 12445 1539
rect 12483 1505 12517 1539
rect 12555 1505 12589 1539
rect 12645 1505 12679 1539
rect 12717 1505 12751 1539
rect 12789 1505 12823 1539
rect 12861 1505 12895 1539
rect 13005 1505 13039 1539
rect 13077 1505 13111 1539
rect 13149 1505 13183 1539
rect 13221 1505 13255 1539
rect 13293 1505 13327 1539
rect 13365 1505 13399 1539
rect 13463 1505 13497 1539
rect 13535 1505 13569 1539
rect 13607 1505 13641 1539
rect 13679 1505 13713 1539
rect 13751 1505 13785 1539
rect 13823 1505 13857 1539
rect 13967 1505 14001 1539
rect 14039 1505 14073 1539
rect 14111 1505 14145 1539
rect 14183 1505 14217 1539
rect 14255 1505 14289 1539
rect 14327 1505 14361 1539
rect 14425 1505 14459 1539
rect 14497 1505 14531 1539
rect 14569 1505 14603 1539
rect 14641 1505 14675 1539
rect 14713 1505 14747 1539
rect 14785 1505 14819 1539
rect 14929 1505 14963 1539
rect 15001 1505 15035 1539
rect 15073 1505 15107 1539
rect 15145 1505 15179 1539
rect 15235 1505 15269 1539
rect 15307 1505 15341 1539
rect 15379 1505 15413 1539
rect 15451 1505 15485 1539
rect 15595 1505 15629 1539
rect 15667 1505 15701 1539
rect 15739 1505 15773 1539
rect 15811 1505 15845 1539
rect 15901 1505 15935 1539
rect 15973 1505 16007 1539
rect 16045 1505 16079 1539
rect 16117 1505 16151 1539
rect 16261 1505 16295 1539
rect 16333 1505 16367 1539
rect 16405 1505 16439 1539
rect 16477 1505 16511 1539
rect 16567 1505 16601 1539
rect 16639 1505 16673 1539
rect 16711 1505 16745 1539
rect 16783 1505 16817 1539
rect 16927 1505 16961 1539
rect 16999 1505 17033 1539
rect 17071 1505 17105 1539
rect 17143 1505 17177 1539
rect 17233 1505 17267 1539
rect 17305 1505 17339 1539
rect 17377 1505 17411 1539
rect 17449 1505 17483 1539
rect 17593 1505 17627 1539
rect 17665 1505 17699 1539
rect 17743 1505 17777 1539
rect 17821 1505 17855 1539
rect 17893 1505 17927 1539
rect -17 1436 17 1470
rect -17 1364 17 1398
rect -17 1292 17 1326
rect -17 1220 17 1254
rect -17 1148 17 1182
rect -17 1076 17 1110
rect 945 1436 979 1470
rect 945 1364 979 1398
rect 945 1292 979 1326
rect 945 1220 979 1254
rect 945 1148 979 1182
rect 945 1076 979 1110
rect -17 1004 17 1038
rect -17 932 17 966
rect 1907 1436 1941 1470
rect 1907 1364 1941 1398
rect 1907 1292 1941 1326
rect 1907 1220 1941 1254
rect 1907 1148 1941 1182
rect 1907 1076 1941 1110
rect 945 1004 979 1038
rect 945 932 979 966
rect 2573 1436 2607 1470
rect 2573 1364 2607 1398
rect 2573 1292 2607 1326
rect 2573 1220 2607 1254
rect 2573 1148 2607 1182
rect 2573 1076 2607 1110
rect 1907 1004 1941 1038
rect 1907 932 1941 966
rect 3535 1436 3569 1470
rect 3535 1364 3569 1398
rect 3535 1292 3569 1326
rect 3535 1220 3569 1254
rect 3535 1148 3569 1182
rect 3535 1076 3569 1110
rect 2573 1004 2607 1038
rect 2573 932 2607 966
rect 4497 1436 4531 1470
rect 4497 1364 4531 1398
rect 4497 1292 4531 1326
rect 4497 1220 4531 1254
rect 4497 1148 4531 1182
rect 4497 1076 4531 1110
rect 3535 1004 3569 1038
rect 3535 932 3569 966
rect 5163 1436 5197 1470
rect 5163 1364 5197 1398
rect 5163 1292 5197 1326
rect 5163 1220 5197 1254
rect 5163 1148 5197 1182
rect 5163 1076 5197 1110
rect 4497 1004 4531 1038
rect 4497 932 4531 966
rect 6125 1436 6159 1470
rect 6125 1364 6159 1398
rect 6125 1292 6159 1326
rect 6125 1220 6159 1254
rect 6125 1148 6159 1182
rect 6125 1076 6159 1110
rect 5163 1004 5197 1038
rect 5163 932 5197 966
rect 7087 1436 7121 1470
rect 7087 1364 7121 1398
rect 7087 1292 7121 1326
rect 7087 1220 7121 1254
rect 7087 1148 7121 1182
rect 7087 1076 7121 1110
rect 6125 1004 6159 1038
rect 6125 932 6159 966
rect 7753 1436 7787 1470
rect 7753 1364 7787 1398
rect 7753 1292 7787 1326
rect 7753 1220 7787 1254
rect 7753 1148 7787 1182
rect 7753 1076 7787 1110
rect 7087 1004 7121 1038
rect 7087 932 7121 966
rect 8715 1436 8749 1470
rect 8715 1364 8749 1398
rect 8715 1292 8749 1326
rect 8715 1220 8749 1254
rect 8715 1148 8749 1182
rect 8715 1076 8749 1110
rect 7753 1004 7787 1038
rect 7753 932 7787 966
rect 9677 1436 9711 1470
rect 9677 1364 9711 1398
rect 9677 1292 9711 1326
rect 9677 1220 9711 1254
rect 9677 1148 9711 1182
rect 9677 1076 9711 1110
rect 8715 1004 8749 1038
rect 8715 932 8749 966
rect 10343 1436 10377 1470
rect 10343 1364 10377 1398
rect 10343 1292 10377 1326
rect 10343 1220 10377 1254
rect 10343 1148 10377 1182
rect 10343 1076 10377 1110
rect 9677 1004 9711 1038
rect 9677 932 9711 966
rect 11305 1436 11339 1470
rect 11305 1364 11339 1398
rect 11305 1292 11339 1326
rect 11305 1220 11339 1254
rect 11305 1148 11339 1182
rect 11305 1076 11339 1110
rect 10343 1004 10377 1038
rect 10343 932 10377 966
rect 12267 1436 12301 1470
rect 12267 1364 12301 1398
rect 12267 1292 12301 1326
rect 12267 1220 12301 1254
rect 12267 1148 12301 1182
rect 12267 1076 12301 1110
rect 11305 1004 11339 1038
rect 11305 932 11339 966
rect 12933 1436 12967 1470
rect 12933 1364 12967 1398
rect 12933 1292 12967 1326
rect 12933 1220 12967 1254
rect 12933 1148 12967 1182
rect 12933 1076 12967 1110
rect 12267 1004 12301 1038
rect 12267 932 12301 966
rect 13895 1436 13929 1470
rect 13895 1364 13929 1398
rect 13895 1292 13929 1326
rect 13895 1220 13929 1254
rect 13895 1148 13929 1182
rect 13895 1076 13929 1110
rect 12933 1004 12967 1038
rect 12933 932 12967 966
rect 14857 1436 14891 1470
rect 14857 1364 14891 1398
rect 14857 1292 14891 1326
rect 14857 1220 14891 1254
rect 14857 1148 14891 1182
rect 14857 1076 14891 1110
rect 13895 1004 13929 1038
rect 13895 932 13929 966
rect 15523 1436 15557 1470
rect 15523 1364 15557 1398
rect 15523 1292 15557 1326
rect 15523 1220 15557 1254
rect 15523 1148 15557 1182
rect 15523 1076 15557 1110
rect 14857 1004 14891 1038
rect 14857 932 14891 966
rect 16189 1436 16223 1470
rect 16189 1364 16223 1398
rect 16189 1292 16223 1326
rect 16189 1220 16223 1254
rect 16189 1148 16223 1182
rect 16189 1076 16223 1110
rect 15523 1004 15557 1038
rect 15523 932 15557 966
rect 16855 1436 16889 1470
rect 16855 1364 16889 1398
rect 16855 1292 16889 1326
rect 16855 1220 16889 1254
rect 16855 1148 16889 1182
rect 16855 1076 16889 1110
rect 16189 1004 16223 1038
rect 16189 932 16223 966
rect 17521 1436 17555 1470
rect 17521 1364 17555 1398
rect 17521 1292 17555 1326
rect 17521 1220 17555 1254
rect 17521 1148 17555 1182
rect 17521 1076 17555 1110
rect 16855 1004 16889 1038
rect 16855 932 16889 966
rect 17965 1436 17999 1470
rect 17965 1364 17999 1398
rect 17965 1292 17999 1326
rect 17965 1220 17999 1254
rect 17965 1148 17999 1182
rect 17965 1076 17999 1110
rect 17521 1004 17555 1038
rect 17521 932 17555 966
rect 17965 1004 17999 1038
rect 17965 932 17999 966
<< poly >>
rect 247 1450 277 1476
rect 335 1450 365 1476
rect 423 1450 453 1476
rect 511 1450 541 1476
rect 599 1450 629 1476
rect 687 1450 717 1476
rect 1209 1450 1239 1476
rect 1297 1450 1327 1476
rect 1385 1450 1415 1476
rect 1473 1450 1503 1476
rect 1561 1450 1591 1476
rect 1649 1450 1679 1476
rect 247 1019 277 1050
rect 335 1019 365 1050
rect 423 1019 453 1050
rect 511 1019 541 1050
rect 195 1003 365 1019
rect 195 969 205 1003
rect 239 989 365 1003
rect 417 1003 541 1019
rect 239 969 249 989
rect 195 953 249 969
rect 417 969 427 1003
rect 461 989 541 1003
rect 599 1019 629 1050
rect 687 1019 717 1050
rect 599 1003 717 1019
rect 599 989 649 1003
rect 461 969 471 989
rect 417 953 471 969
rect 639 969 649 989
rect 683 989 717 1003
rect 2111 1450 2141 1476
rect 2199 1450 2229 1476
rect 2287 1450 2317 1476
rect 2375 1450 2405 1476
rect 1209 1019 1239 1050
rect 1297 1019 1327 1050
rect 1385 1019 1415 1050
rect 1473 1019 1503 1050
rect 683 969 693 989
rect 639 953 693 969
rect 1157 1003 1327 1019
rect 1157 969 1167 1003
rect 1201 989 1327 1003
rect 1379 1003 1503 1019
rect 1201 969 1211 989
rect 1157 953 1211 969
rect 1379 969 1389 1003
rect 1423 989 1503 1003
rect 1561 1019 1591 1050
rect 1649 1019 1679 1050
rect 1561 1003 1679 1019
rect 1561 989 1611 1003
rect 1423 969 1433 989
rect 1379 953 1433 969
rect 1601 969 1611 989
rect 1645 989 1679 1003
rect 2837 1450 2867 1476
rect 2925 1450 2955 1476
rect 3013 1450 3043 1476
rect 3101 1450 3131 1476
rect 3189 1450 3219 1476
rect 3277 1450 3307 1476
rect 1645 969 1655 989
rect 1601 953 1655 969
rect 2111 1019 2141 1050
rect 2199 1019 2229 1050
rect 2287 1019 2317 1050
rect 2375 1019 2405 1050
rect 2111 1003 2229 1019
rect 2111 989 2129 1003
rect 2119 969 2129 989
rect 2163 989 2229 1003
rect 2273 1003 2405 1019
rect 2163 969 2173 989
rect 2119 953 2173 969
rect 2273 969 2283 1003
rect 2317 989 2405 1003
rect 3799 1450 3829 1476
rect 3887 1450 3917 1476
rect 3975 1450 4005 1476
rect 4063 1450 4093 1476
rect 4151 1450 4181 1476
rect 4239 1450 4269 1476
rect 2837 1019 2867 1050
rect 2925 1019 2955 1050
rect 3013 1019 3043 1050
rect 3101 1019 3131 1050
rect 2317 969 2327 989
rect 2273 953 2327 969
rect 2785 1003 2955 1019
rect 2785 969 2795 1003
rect 2829 989 2955 1003
rect 3007 1003 3131 1019
rect 2829 969 2839 989
rect 2785 953 2839 969
rect 3007 969 3017 1003
rect 3051 989 3131 1003
rect 3189 1019 3219 1050
rect 3277 1019 3307 1050
rect 3189 1003 3307 1019
rect 3189 989 3239 1003
rect 3051 969 3061 989
rect 3007 953 3061 969
rect 3229 969 3239 989
rect 3273 989 3307 1003
rect 4701 1450 4731 1476
rect 4789 1450 4819 1476
rect 4877 1450 4907 1476
rect 4965 1450 4995 1476
rect 3799 1019 3829 1050
rect 3887 1019 3917 1050
rect 3975 1019 4005 1050
rect 4063 1019 4093 1050
rect 3273 969 3283 989
rect 3229 953 3283 969
rect 3747 1003 3917 1019
rect 3747 969 3757 1003
rect 3791 989 3917 1003
rect 3969 1003 4093 1019
rect 3791 969 3801 989
rect 3747 953 3801 969
rect 3969 969 3979 1003
rect 4013 989 4093 1003
rect 4151 1019 4181 1050
rect 4239 1019 4269 1050
rect 4151 1003 4269 1019
rect 4151 989 4201 1003
rect 4013 969 4023 989
rect 3969 953 4023 969
rect 4191 969 4201 989
rect 4235 989 4269 1003
rect 5427 1450 5457 1476
rect 5515 1450 5545 1476
rect 5603 1450 5633 1476
rect 5691 1450 5721 1476
rect 5779 1450 5809 1476
rect 5867 1450 5897 1476
rect 4235 969 4245 989
rect 4191 953 4245 969
rect 4701 1019 4731 1050
rect 4789 1019 4819 1050
rect 4877 1019 4907 1050
rect 4965 1019 4995 1050
rect 4701 1003 4819 1019
rect 4701 989 4719 1003
rect 4709 969 4719 989
rect 4753 989 4819 1003
rect 4863 1003 4995 1019
rect 4753 969 4763 989
rect 4709 953 4763 969
rect 4863 969 4873 1003
rect 4907 989 4995 1003
rect 6389 1450 6419 1476
rect 6477 1450 6507 1476
rect 6565 1450 6595 1476
rect 6653 1450 6683 1476
rect 6741 1450 6771 1476
rect 6829 1450 6859 1476
rect 5427 1019 5457 1050
rect 5515 1019 5545 1050
rect 5603 1019 5633 1050
rect 5691 1019 5721 1050
rect 4907 969 4917 989
rect 4863 953 4917 969
rect 5375 1003 5545 1019
rect 5375 969 5385 1003
rect 5419 989 5545 1003
rect 5597 1003 5721 1019
rect 5419 969 5429 989
rect 5375 953 5429 969
rect 5597 969 5607 1003
rect 5641 989 5721 1003
rect 5779 1019 5809 1050
rect 5867 1019 5897 1050
rect 5779 1003 5897 1019
rect 5779 989 5829 1003
rect 5641 969 5651 989
rect 5597 953 5651 969
rect 5819 969 5829 989
rect 5863 989 5897 1003
rect 7291 1450 7321 1476
rect 7379 1450 7409 1476
rect 7467 1450 7497 1476
rect 7555 1450 7585 1476
rect 6389 1019 6419 1050
rect 6477 1019 6507 1050
rect 6565 1019 6595 1050
rect 6653 1019 6683 1050
rect 5863 969 5873 989
rect 5819 953 5873 969
rect 6337 1003 6507 1019
rect 6337 969 6347 1003
rect 6381 989 6507 1003
rect 6559 1003 6683 1019
rect 6381 969 6391 989
rect 6337 953 6391 969
rect 6559 969 6569 1003
rect 6603 989 6683 1003
rect 6741 1019 6771 1050
rect 6829 1019 6859 1050
rect 6741 1003 6859 1019
rect 6741 989 6791 1003
rect 6603 969 6613 989
rect 6559 953 6613 969
rect 6781 969 6791 989
rect 6825 989 6859 1003
rect 8017 1450 8047 1476
rect 8105 1450 8135 1476
rect 8193 1450 8223 1476
rect 8281 1450 8311 1476
rect 8369 1450 8399 1476
rect 8457 1450 8487 1476
rect 6825 969 6835 989
rect 6781 953 6835 969
rect 7291 1019 7321 1050
rect 7379 1019 7409 1050
rect 7467 1019 7497 1050
rect 7555 1019 7585 1050
rect 7291 1003 7409 1019
rect 7291 989 7309 1003
rect 7299 969 7309 989
rect 7343 989 7409 1003
rect 7453 1003 7585 1019
rect 7343 969 7353 989
rect 7299 953 7353 969
rect 7453 969 7463 1003
rect 7497 989 7585 1003
rect 8979 1450 9009 1476
rect 9067 1450 9097 1476
rect 9155 1450 9185 1476
rect 9243 1450 9273 1476
rect 9331 1450 9361 1476
rect 9419 1450 9449 1476
rect 8017 1019 8047 1050
rect 8105 1019 8135 1050
rect 8193 1019 8223 1050
rect 8281 1019 8311 1050
rect 7497 969 7507 989
rect 7453 953 7507 969
rect 7965 1003 8135 1019
rect 7965 969 7975 1003
rect 8009 989 8135 1003
rect 8187 1003 8311 1019
rect 8009 969 8019 989
rect 7965 953 8019 969
rect 8187 969 8197 1003
rect 8231 989 8311 1003
rect 8369 1019 8399 1050
rect 8457 1019 8487 1050
rect 8369 1003 8487 1019
rect 8369 989 8419 1003
rect 8231 969 8241 989
rect 8187 953 8241 969
rect 8409 969 8419 989
rect 8453 989 8487 1003
rect 9881 1450 9911 1476
rect 9969 1450 9999 1476
rect 10057 1450 10087 1476
rect 10145 1450 10175 1476
rect 8979 1019 9009 1050
rect 9067 1019 9097 1050
rect 9155 1019 9185 1050
rect 9243 1019 9273 1050
rect 8453 969 8463 989
rect 8409 953 8463 969
rect 8927 1003 9097 1019
rect 8927 969 8937 1003
rect 8971 989 9097 1003
rect 9149 1003 9273 1019
rect 8971 969 8981 989
rect 8927 953 8981 969
rect 9149 969 9159 1003
rect 9193 989 9273 1003
rect 9331 1019 9361 1050
rect 9419 1019 9449 1050
rect 9331 1003 9449 1019
rect 9331 989 9381 1003
rect 9193 969 9203 989
rect 9149 953 9203 969
rect 9371 969 9381 989
rect 9415 989 9449 1003
rect 10607 1450 10637 1476
rect 10695 1450 10725 1476
rect 10783 1450 10813 1476
rect 10871 1450 10901 1476
rect 10959 1450 10989 1476
rect 11047 1450 11077 1476
rect 9415 969 9425 989
rect 9371 953 9425 969
rect 9881 1019 9911 1050
rect 9969 1019 9999 1050
rect 10057 1019 10087 1050
rect 10145 1019 10175 1050
rect 9881 1003 9999 1019
rect 9881 989 9899 1003
rect 9889 969 9899 989
rect 9933 989 9999 1003
rect 10043 1003 10175 1019
rect 9933 969 9943 989
rect 9889 953 9943 969
rect 10043 969 10053 1003
rect 10087 989 10175 1003
rect 11569 1450 11599 1476
rect 11657 1450 11687 1476
rect 11745 1450 11775 1476
rect 11833 1450 11863 1476
rect 11921 1450 11951 1476
rect 12009 1450 12039 1476
rect 10607 1019 10637 1050
rect 10695 1019 10725 1050
rect 10783 1019 10813 1050
rect 10871 1019 10901 1050
rect 10087 969 10097 989
rect 10043 953 10097 969
rect 10555 1003 10725 1019
rect 10555 969 10565 1003
rect 10599 989 10725 1003
rect 10777 1003 10901 1019
rect 10599 969 10609 989
rect 10555 953 10609 969
rect 10777 969 10787 1003
rect 10821 989 10901 1003
rect 10959 1019 10989 1050
rect 11047 1019 11077 1050
rect 10959 1003 11077 1019
rect 10959 989 11009 1003
rect 10821 969 10831 989
rect 10777 953 10831 969
rect 10999 969 11009 989
rect 11043 989 11077 1003
rect 12471 1450 12501 1476
rect 12559 1450 12589 1476
rect 12647 1450 12677 1476
rect 12735 1450 12765 1476
rect 11569 1019 11599 1050
rect 11657 1019 11687 1050
rect 11745 1019 11775 1050
rect 11833 1019 11863 1050
rect 11043 969 11053 989
rect 10999 953 11053 969
rect 11517 1003 11687 1019
rect 11517 969 11527 1003
rect 11561 989 11687 1003
rect 11739 1003 11863 1019
rect 11561 969 11571 989
rect 11517 953 11571 969
rect 11739 969 11749 1003
rect 11783 989 11863 1003
rect 11921 1019 11951 1050
rect 12009 1019 12039 1050
rect 11921 1003 12039 1019
rect 11921 989 11971 1003
rect 11783 969 11793 989
rect 11739 953 11793 969
rect 11961 969 11971 989
rect 12005 989 12039 1003
rect 13197 1450 13227 1476
rect 13285 1450 13315 1476
rect 13373 1450 13403 1476
rect 13461 1450 13491 1476
rect 13549 1450 13579 1476
rect 13637 1450 13667 1476
rect 12005 969 12015 989
rect 11961 953 12015 969
rect 12471 1019 12501 1050
rect 12559 1019 12589 1050
rect 12647 1019 12677 1050
rect 12735 1019 12765 1050
rect 12471 1003 12589 1019
rect 12471 989 12489 1003
rect 12479 969 12489 989
rect 12523 989 12589 1003
rect 12633 1003 12765 1019
rect 12523 969 12533 989
rect 12479 953 12533 969
rect 12633 969 12643 1003
rect 12677 989 12765 1003
rect 14159 1450 14189 1476
rect 14247 1450 14277 1476
rect 14335 1450 14365 1476
rect 14423 1450 14453 1476
rect 14511 1450 14541 1476
rect 14599 1450 14629 1476
rect 13197 1019 13227 1050
rect 13285 1019 13315 1050
rect 13373 1019 13403 1050
rect 13461 1019 13491 1050
rect 12677 969 12687 989
rect 12633 953 12687 969
rect 13145 1003 13315 1019
rect 13145 969 13155 1003
rect 13189 989 13315 1003
rect 13367 1003 13491 1019
rect 13189 969 13199 989
rect 13145 953 13199 969
rect 13367 969 13377 1003
rect 13411 989 13491 1003
rect 13549 1019 13579 1050
rect 13637 1019 13667 1050
rect 13549 1003 13667 1019
rect 13549 989 13599 1003
rect 13411 969 13421 989
rect 13367 953 13421 969
rect 13589 969 13599 989
rect 13633 989 13667 1003
rect 15061 1450 15091 1476
rect 15149 1450 15179 1476
rect 15237 1450 15267 1476
rect 15325 1450 15355 1476
rect 14159 1019 14189 1050
rect 14247 1019 14277 1050
rect 14335 1019 14365 1050
rect 14423 1019 14453 1050
rect 13633 969 13643 989
rect 13589 953 13643 969
rect 14107 1003 14277 1019
rect 14107 969 14117 1003
rect 14151 989 14277 1003
rect 14329 1003 14453 1019
rect 14151 969 14161 989
rect 14107 953 14161 969
rect 14329 969 14339 1003
rect 14373 989 14453 1003
rect 14511 1019 14541 1050
rect 14599 1019 14629 1050
rect 14511 1003 14629 1019
rect 14511 989 14561 1003
rect 14373 969 14383 989
rect 14329 953 14383 969
rect 14551 969 14561 989
rect 14595 989 14629 1003
rect 15727 1451 15757 1477
rect 15815 1451 15845 1477
rect 15903 1451 15933 1477
rect 15991 1451 16021 1477
rect 14595 969 14605 989
rect 14551 953 14605 969
rect 15061 1019 15091 1050
rect 15149 1019 15179 1050
rect 15237 1019 15267 1050
rect 15325 1019 15355 1050
rect 15061 1003 15179 1019
rect 15061 989 15079 1003
rect 15069 969 15079 989
rect 15113 989 15179 1003
rect 15223 1003 15355 1019
rect 15113 969 15123 989
rect 15069 953 15123 969
rect 15223 969 15233 1003
rect 15267 989 15355 1003
rect 16391 1451 16421 1477
rect 16479 1451 16509 1477
rect 16567 1451 16597 1477
rect 16655 1451 16685 1477
rect 15727 1020 15757 1051
rect 15815 1020 15845 1051
rect 15903 1020 15933 1051
rect 15991 1020 16021 1051
rect 15267 969 15277 989
rect 15223 953 15277 969
rect 15661 1004 15845 1020
rect 15661 970 15671 1004
rect 15705 990 15845 1004
rect 15891 1004 16021 1020
rect 15705 970 15715 990
rect 15661 954 15715 970
rect 15891 970 15901 1004
rect 15935 990 16021 1004
rect 17059 1451 17089 1477
rect 17147 1451 17177 1477
rect 17235 1451 17265 1477
rect 17323 1451 17353 1477
rect 15935 970 15945 990
rect 15891 954 15945 970
rect 16391 1020 16421 1051
rect 16479 1020 16509 1051
rect 16391 1004 16509 1020
rect 16391 990 16411 1004
rect 16401 970 16411 990
rect 16445 990 16509 1004
rect 16567 1020 16597 1051
rect 16655 1020 16685 1051
rect 17701 1450 17731 1476
rect 17789 1450 17819 1476
rect 16567 1004 16751 1020
rect 16567 990 16707 1004
rect 16445 970 16455 990
rect 16401 954 16455 970
rect 16697 970 16707 990
rect 16741 970 16751 1004
rect 16697 954 16751 970
rect 17059 1020 17089 1051
rect 17147 1020 17177 1051
rect 17235 1020 17265 1051
rect 17323 1020 17353 1051
rect 16993 1004 17177 1020
rect 16993 970 17003 1004
rect 17037 990 17177 1004
rect 17219 1004 17353 1020
rect 17037 970 17047 990
rect 16993 954 17047 970
rect 17219 970 17229 1004
rect 17263 990 17353 1004
rect 17701 1019 17731 1050
rect 17789 1019 17819 1050
rect 17263 970 17273 990
rect 17219 954 17273 970
rect 17659 1003 17819 1019
rect 17659 969 17669 1003
rect 17703 989 17819 1003
rect 17703 969 17713 989
rect 17659 953 17713 969
rect 195 461 249 477
rect 195 441 205 461
rect 147 427 205 441
rect 239 427 249 461
rect 147 411 249 427
rect 417 461 471 477
rect 417 427 427 461
rect 461 441 471 461
rect 639 461 693 477
rect 461 427 477 441
rect 417 411 477 427
rect 639 427 649 461
rect 683 427 693 461
rect 639 411 693 427
rect 1157 461 1211 477
rect 1157 441 1167 461
rect 147 379 177 411
rect 447 379 477 411
rect 649 379 679 411
rect 1109 427 1167 441
rect 1201 427 1211 461
rect 1109 411 1211 427
rect 1379 461 1433 477
rect 1379 427 1389 461
rect 1423 441 1433 461
rect 1601 461 1655 477
rect 1423 427 1439 441
rect 1379 411 1439 427
rect 1601 427 1611 461
rect 1645 427 1655 461
rect 1601 411 1655 427
rect 2119 461 2173 477
rect 2119 441 2129 461
rect 1109 379 1139 411
rect 1409 379 1439 411
rect 1611 379 1641 411
rect 2092 427 2129 441
rect 2163 427 2173 461
rect 2092 411 2173 427
rect 2267 461 2321 477
rect 2267 427 2277 461
rect 2311 427 2321 461
rect 2267 411 2321 427
rect 2785 461 2839 477
rect 2785 441 2795 461
rect 2092 377 2122 411
rect 2286 377 2316 411
rect 2737 427 2795 441
rect 2829 427 2839 461
rect 2737 411 2839 427
rect 3007 461 3061 477
rect 3007 427 3017 461
rect 3051 441 3061 461
rect 3229 461 3283 477
rect 3051 427 3067 441
rect 3007 411 3067 427
rect 3229 427 3239 461
rect 3273 427 3283 461
rect 3229 411 3283 427
rect 3747 461 3801 477
rect 3747 441 3757 461
rect 2737 379 2767 411
rect 3037 379 3067 411
rect 3239 379 3269 411
rect 3699 427 3757 441
rect 3791 427 3801 461
rect 3699 411 3801 427
rect 3969 461 4023 477
rect 3969 427 3979 461
rect 4013 441 4023 461
rect 4191 461 4245 477
rect 4013 427 4029 441
rect 3969 411 4029 427
rect 4191 427 4201 461
rect 4235 427 4245 461
rect 4191 411 4245 427
rect 4709 461 4763 477
rect 4709 441 4719 461
rect 3699 379 3729 411
rect 3999 379 4029 411
rect 4201 379 4231 411
rect 4682 427 4719 441
rect 4753 427 4763 461
rect 4682 411 4763 427
rect 4857 461 4911 477
rect 4857 427 4867 461
rect 4901 427 4911 461
rect 4857 411 4911 427
rect 5375 461 5429 477
rect 5375 441 5385 461
rect 4682 377 4712 411
rect 4876 377 4906 411
rect 5327 427 5385 441
rect 5419 427 5429 461
rect 5327 411 5429 427
rect 5597 461 5651 477
rect 5597 427 5607 461
rect 5641 441 5651 461
rect 5819 461 5873 477
rect 5641 427 5657 441
rect 5597 411 5657 427
rect 5819 427 5829 461
rect 5863 427 5873 461
rect 5819 411 5873 427
rect 6337 461 6391 477
rect 6337 441 6347 461
rect 5327 379 5357 411
rect 5627 379 5657 411
rect 5829 379 5859 411
rect 6289 427 6347 441
rect 6381 427 6391 461
rect 6289 411 6391 427
rect 6559 461 6613 477
rect 6559 427 6569 461
rect 6603 441 6613 461
rect 6781 461 6835 477
rect 6603 427 6619 441
rect 6559 411 6619 427
rect 6781 427 6791 461
rect 6825 427 6835 461
rect 6781 411 6835 427
rect 7299 461 7353 477
rect 7299 441 7309 461
rect 6289 379 6319 411
rect 6589 379 6619 411
rect 6791 379 6821 411
rect 7272 427 7309 441
rect 7343 427 7353 461
rect 7272 411 7353 427
rect 7447 461 7501 477
rect 7447 427 7457 461
rect 7491 427 7501 461
rect 7447 411 7501 427
rect 7965 461 8019 477
rect 7965 441 7975 461
rect 7272 377 7302 411
rect 7466 377 7496 411
rect 7917 427 7975 441
rect 8009 427 8019 461
rect 7917 411 8019 427
rect 8187 461 8241 477
rect 8187 427 8197 461
rect 8231 441 8241 461
rect 8409 461 8463 477
rect 8231 427 8247 441
rect 8187 411 8247 427
rect 8409 427 8419 461
rect 8453 427 8463 461
rect 8409 411 8463 427
rect 8927 461 8981 477
rect 8927 441 8937 461
rect 7917 379 7947 411
rect 8217 379 8247 411
rect 8419 379 8449 411
rect 8879 427 8937 441
rect 8971 427 8981 461
rect 8879 411 8981 427
rect 9149 461 9203 477
rect 9149 427 9159 461
rect 9193 441 9203 461
rect 9371 461 9425 477
rect 9193 427 9209 441
rect 9149 411 9209 427
rect 9371 427 9381 461
rect 9415 427 9425 461
rect 9371 411 9425 427
rect 9889 461 9943 477
rect 9889 441 9899 461
rect 8879 379 8909 411
rect 9179 379 9209 411
rect 9381 379 9411 411
rect 9862 427 9899 441
rect 9933 427 9943 461
rect 9862 411 9943 427
rect 10037 461 10091 477
rect 10037 427 10047 461
rect 10081 427 10091 461
rect 10037 411 10091 427
rect 10555 461 10609 477
rect 10555 441 10565 461
rect 9862 377 9892 411
rect 10056 377 10086 411
rect 10507 427 10565 441
rect 10599 427 10609 461
rect 10507 411 10609 427
rect 10777 461 10831 477
rect 10777 427 10787 461
rect 10821 441 10831 461
rect 10999 461 11053 477
rect 10821 427 10837 441
rect 10777 411 10837 427
rect 10999 427 11009 461
rect 11043 427 11053 461
rect 10999 411 11053 427
rect 11517 461 11571 477
rect 11517 441 11527 461
rect 10507 379 10537 411
rect 10807 379 10837 411
rect 11009 379 11039 411
rect 11469 427 11527 441
rect 11561 427 11571 461
rect 11469 411 11571 427
rect 11739 461 11793 477
rect 11739 427 11749 461
rect 11783 441 11793 461
rect 11961 461 12015 477
rect 11783 427 11799 441
rect 11739 411 11799 427
rect 11961 427 11971 461
rect 12005 427 12015 461
rect 11961 411 12015 427
rect 12479 461 12533 477
rect 12479 441 12489 461
rect 11469 379 11499 411
rect 11769 379 11799 411
rect 11971 379 12001 411
rect 12452 427 12489 441
rect 12523 427 12533 461
rect 12452 411 12533 427
rect 12627 461 12681 477
rect 12627 427 12637 461
rect 12671 427 12681 461
rect 12627 411 12681 427
rect 13145 461 13199 477
rect 13145 441 13155 461
rect 12452 377 12482 411
rect 12646 377 12676 411
rect 13097 427 13155 441
rect 13189 427 13199 461
rect 13097 411 13199 427
rect 13367 461 13421 477
rect 13367 427 13377 461
rect 13411 441 13421 461
rect 13589 461 13643 477
rect 13411 427 13427 441
rect 13367 411 13427 427
rect 13589 427 13599 461
rect 13633 427 13643 461
rect 13589 411 13643 427
rect 14107 461 14161 477
rect 14107 441 14117 461
rect 13097 379 13127 411
rect 13397 379 13427 411
rect 13599 379 13629 411
rect 14059 427 14117 441
rect 14151 427 14161 461
rect 14059 411 14161 427
rect 14329 461 14383 477
rect 14329 427 14339 461
rect 14373 441 14383 461
rect 14551 461 14605 477
rect 14373 427 14389 441
rect 14329 411 14389 427
rect 14551 427 14561 461
rect 14595 427 14605 461
rect 14551 411 14605 427
rect 15069 461 15123 477
rect 15069 441 15079 461
rect 14059 379 14089 411
rect 14359 379 14389 411
rect 14561 379 14591 411
rect 15042 427 15079 441
rect 15113 427 15123 461
rect 15042 411 15123 427
rect 15217 461 15271 477
rect 15217 427 15227 461
rect 15261 427 15271 461
rect 15217 411 15271 427
rect 15042 377 15072 411
rect 15236 377 15266 411
rect 15661 461 15715 477
rect 15661 427 15671 461
rect 15705 441 15715 461
rect 15883 461 15937 477
rect 15705 427 15738 441
rect 15661 411 15738 427
rect 15883 427 15893 461
rect 15927 427 15937 461
rect 15883 411 15937 427
rect 16401 461 16455 477
rect 16401 441 16411 461
rect 15708 377 15738 411
rect 15902 377 15932 411
rect 16374 427 16411 441
rect 16445 427 16455 461
rect 16697 461 16751 477
rect 16697 441 16707 461
rect 16374 411 16455 427
rect 16674 427 16707 441
rect 16741 427 16751 461
rect 16674 411 16751 427
rect 16374 377 16404 411
rect 16674 377 16704 411
rect 16993 461 17047 477
rect 16993 427 17003 461
rect 17037 441 17047 461
rect 17215 461 17269 477
rect 17037 427 17070 441
rect 16993 411 17070 427
rect 17215 427 17225 461
rect 17259 427 17269 461
rect 17215 411 17269 427
rect 17040 377 17070 411
rect 17234 377 17264 411
rect 17659 461 17713 477
rect 17659 427 17669 461
rect 17703 441 17713 461
rect 17703 427 17723 441
rect 17659 411 17723 427
rect 17693 377 17723 411
<< polycont >>
rect 205 969 239 1003
rect 427 969 461 1003
rect 649 969 683 1003
rect 1167 969 1201 1003
rect 1389 969 1423 1003
rect 1611 969 1645 1003
rect 2129 969 2163 1003
rect 2283 969 2317 1003
rect 2795 969 2829 1003
rect 3017 969 3051 1003
rect 3239 969 3273 1003
rect 3757 969 3791 1003
rect 3979 969 4013 1003
rect 4201 969 4235 1003
rect 4719 969 4753 1003
rect 4873 969 4907 1003
rect 5385 969 5419 1003
rect 5607 969 5641 1003
rect 5829 969 5863 1003
rect 6347 969 6381 1003
rect 6569 969 6603 1003
rect 6791 969 6825 1003
rect 7309 969 7343 1003
rect 7463 969 7497 1003
rect 7975 969 8009 1003
rect 8197 969 8231 1003
rect 8419 969 8453 1003
rect 8937 969 8971 1003
rect 9159 969 9193 1003
rect 9381 969 9415 1003
rect 9899 969 9933 1003
rect 10053 969 10087 1003
rect 10565 969 10599 1003
rect 10787 969 10821 1003
rect 11009 969 11043 1003
rect 11527 969 11561 1003
rect 11749 969 11783 1003
rect 11971 969 12005 1003
rect 12489 969 12523 1003
rect 12643 969 12677 1003
rect 13155 969 13189 1003
rect 13377 969 13411 1003
rect 13599 969 13633 1003
rect 14117 969 14151 1003
rect 14339 969 14373 1003
rect 14561 969 14595 1003
rect 15079 969 15113 1003
rect 15233 969 15267 1003
rect 15671 970 15705 1004
rect 15901 970 15935 1004
rect 16411 970 16445 1004
rect 16707 970 16741 1004
rect 17003 970 17037 1004
rect 17229 970 17263 1004
rect 17669 969 17703 1003
rect 205 427 239 461
rect 427 427 461 461
rect 649 427 683 461
rect 1167 427 1201 461
rect 1389 427 1423 461
rect 1611 427 1645 461
rect 2129 427 2163 461
rect 2277 427 2311 461
rect 2795 427 2829 461
rect 3017 427 3051 461
rect 3239 427 3273 461
rect 3757 427 3791 461
rect 3979 427 4013 461
rect 4201 427 4235 461
rect 4719 427 4753 461
rect 4867 427 4901 461
rect 5385 427 5419 461
rect 5607 427 5641 461
rect 5829 427 5863 461
rect 6347 427 6381 461
rect 6569 427 6603 461
rect 6791 427 6825 461
rect 7309 427 7343 461
rect 7457 427 7491 461
rect 7975 427 8009 461
rect 8197 427 8231 461
rect 8419 427 8453 461
rect 8937 427 8971 461
rect 9159 427 9193 461
rect 9381 427 9415 461
rect 9899 427 9933 461
rect 10047 427 10081 461
rect 10565 427 10599 461
rect 10787 427 10821 461
rect 11009 427 11043 461
rect 11527 427 11561 461
rect 11749 427 11783 461
rect 11971 427 12005 461
rect 12489 427 12523 461
rect 12637 427 12671 461
rect 13155 427 13189 461
rect 13377 427 13411 461
rect 13599 427 13633 461
rect 14117 427 14151 461
rect 14339 427 14373 461
rect 14561 427 14595 461
rect 15079 427 15113 461
rect 15227 427 15261 461
rect 15671 427 15705 461
rect 15893 427 15927 461
rect 16411 427 16445 461
rect 16707 427 16741 461
rect 17003 427 17037 461
rect 17225 427 17259 461
rect 17669 427 17703 461
<< locali >>
rect -31 1539 18013 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 343 1539
rect 377 1505 415 1539
rect 449 1505 513 1539
rect 547 1505 585 1539
rect 619 1505 657 1539
rect 691 1505 729 1539
rect 763 1505 801 1539
rect 835 1505 873 1539
rect 907 1505 1017 1539
rect 1051 1505 1089 1539
rect 1123 1505 1161 1539
rect 1195 1505 1233 1539
rect 1267 1505 1305 1539
rect 1339 1505 1377 1539
rect 1411 1505 1475 1539
rect 1509 1505 1547 1539
rect 1581 1505 1619 1539
rect 1653 1505 1691 1539
rect 1725 1505 1763 1539
rect 1797 1505 1835 1539
rect 1869 1505 1979 1539
rect 2013 1505 2051 1539
rect 2085 1505 2123 1539
rect 2157 1505 2195 1539
rect 2229 1505 2285 1539
rect 2319 1505 2357 1539
rect 2391 1505 2429 1539
rect 2463 1505 2501 1539
rect 2535 1505 2645 1539
rect 2679 1505 2717 1539
rect 2751 1505 2789 1539
rect 2823 1505 2861 1539
rect 2895 1505 2933 1539
rect 2967 1505 3005 1539
rect 3039 1505 3103 1539
rect 3137 1505 3175 1539
rect 3209 1505 3247 1539
rect 3281 1505 3319 1539
rect 3353 1505 3391 1539
rect 3425 1505 3463 1539
rect 3497 1505 3607 1539
rect 3641 1505 3679 1539
rect 3713 1505 3751 1539
rect 3785 1505 3823 1539
rect 3857 1505 3895 1539
rect 3929 1505 3967 1539
rect 4001 1505 4065 1539
rect 4099 1505 4137 1539
rect 4171 1505 4209 1539
rect 4243 1505 4281 1539
rect 4315 1505 4353 1539
rect 4387 1505 4425 1539
rect 4459 1505 4569 1539
rect 4603 1505 4641 1539
rect 4675 1505 4713 1539
rect 4747 1505 4785 1539
rect 4819 1505 4875 1539
rect 4909 1505 4947 1539
rect 4981 1505 5019 1539
rect 5053 1505 5091 1539
rect 5125 1505 5235 1539
rect 5269 1505 5307 1539
rect 5341 1505 5379 1539
rect 5413 1505 5451 1539
rect 5485 1505 5523 1539
rect 5557 1505 5595 1539
rect 5629 1505 5693 1539
rect 5727 1505 5765 1539
rect 5799 1505 5837 1539
rect 5871 1505 5909 1539
rect 5943 1505 5981 1539
rect 6015 1505 6053 1539
rect 6087 1505 6197 1539
rect 6231 1505 6269 1539
rect 6303 1505 6341 1539
rect 6375 1505 6413 1539
rect 6447 1505 6485 1539
rect 6519 1505 6557 1539
rect 6591 1505 6655 1539
rect 6689 1505 6727 1539
rect 6761 1505 6799 1539
rect 6833 1505 6871 1539
rect 6905 1505 6943 1539
rect 6977 1505 7015 1539
rect 7049 1505 7159 1539
rect 7193 1505 7231 1539
rect 7265 1505 7303 1539
rect 7337 1505 7375 1539
rect 7409 1505 7465 1539
rect 7499 1505 7537 1539
rect 7571 1505 7609 1539
rect 7643 1505 7681 1539
rect 7715 1505 7825 1539
rect 7859 1505 7897 1539
rect 7931 1505 7969 1539
rect 8003 1505 8041 1539
rect 8075 1505 8113 1539
rect 8147 1505 8185 1539
rect 8219 1505 8283 1539
rect 8317 1505 8355 1539
rect 8389 1505 8427 1539
rect 8461 1505 8499 1539
rect 8533 1505 8571 1539
rect 8605 1505 8643 1539
rect 8677 1505 8787 1539
rect 8821 1505 8859 1539
rect 8893 1505 8931 1539
rect 8965 1505 9003 1539
rect 9037 1505 9075 1539
rect 9109 1505 9147 1539
rect 9181 1505 9245 1539
rect 9279 1505 9317 1539
rect 9351 1505 9389 1539
rect 9423 1505 9461 1539
rect 9495 1505 9533 1539
rect 9567 1505 9605 1539
rect 9639 1505 9749 1539
rect 9783 1505 9821 1539
rect 9855 1505 9893 1539
rect 9927 1505 9965 1539
rect 9999 1505 10055 1539
rect 10089 1505 10127 1539
rect 10161 1505 10199 1539
rect 10233 1505 10271 1539
rect 10305 1505 10415 1539
rect 10449 1505 10487 1539
rect 10521 1505 10559 1539
rect 10593 1505 10631 1539
rect 10665 1505 10703 1539
rect 10737 1505 10775 1539
rect 10809 1505 10873 1539
rect 10907 1505 10945 1539
rect 10979 1505 11017 1539
rect 11051 1505 11089 1539
rect 11123 1505 11161 1539
rect 11195 1505 11233 1539
rect 11267 1505 11377 1539
rect 11411 1505 11449 1539
rect 11483 1505 11521 1539
rect 11555 1505 11593 1539
rect 11627 1505 11665 1539
rect 11699 1505 11737 1539
rect 11771 1505 11835 1539
rect 11869 1505 11907 1539
rect 11941 1505 11979 1539
rect 12013 1505 12051 1539
rect 12085 1505 12123 1539
rect 12157 1505 12195 1539
rect 12229 1505 12339 1539
rect 12373 1505 12411 1539
rect 12445 1505 12483 1539
rect 12517 1505 12555 1539
rect 12589 1505 12645 1539
rect 12679 1505 12717 1539
rect 12751 1505 12789 1539
rect 12823 1505 12861 1539
rect 12895 1505 13005 1539
rect 13039 1505 13077 1539
rect 13111 1505 13149 1539
rect 13183 1505 13221 1539
rect 13255 1505 13293 1539
rect 13327 1505 13365 1539
rect 13399 1505 13463 1539
rect 13497 1505 13535 1539
rect 13569 1505 13607 1539
rect 13641 1505 13679 1539
rect 13713 1505 13751 1539
rect 13785 1505 13823 1539
rect 13857 1505 13967 1539
rect 14001 1505 14039 1539
rect 14073 1505 14111 1539
rect 14145 1505 14183 1539
rect 14217 1505 14255 1539
rect 14289 1505 14327 1539
rect 14361 1505 14425 1539
rect 14459 1505 14497 1539
rect 14531 1505 14569 1539
rect 14603 1505 14641 1539
rect 14675 1505 14713 1539
rect 14747 1505 14785 1539
rect 14819 1505 14929 1539
rect 14963 1505 15001 1539
rect 15035 1505 15073 1539
rect 15107 1505 15145 1539
rect 15179 1505 15235 1539
rect 15269 1505 15307 1539
rect 15341 1505 15379 1539
rect 15413 1505 15451 1539
rect 15485 1505 15595 1539
rect 15629 1505 15667 1539
rect 15701 1505 15739 1539
rect 15773 1505 15811 1539
rect 15845 1505 15901 1539
rect 15935 1505 15973 1539
rect 16007 1505 16045 1539
rect 16079 1505 16117 1539
rect 16151 1505 16261 1539
rect 16295 1505 16333 1539
rect 16367 1505 16405 1539
rect 16439 1505 16477 1539
rect 16511 1505 16567 1539
rect 16601 1505 16639 1539
rect 16673 1505 16711 1539
rect 16745 1505 16783 1539
rect 16817 1505 16927 1539
rect 16961 1505 16999 1539
rect 17033 1505 17071 1539
rect 17105 1505 17143 1539
rect 17177 1505 17233 1539
rect 17267 1505 17305 1539
rect 17339 1505 17377 1539
rect 17411 1505 17449 1539
rect 17483 1505 17593 1539
rect 17627 1505 17665 1539
rect 17699 1505 17743 1539
rect 17777 1505 17821 1539
rect 17855 1505 17893 1539
rect 17927 1505 18013 1539
rect -31 1492 18013 1505
rect -31 1470 31 1492
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect 201 1412 235 1492
rect 201 1344 235 1378
rect 201 1276 235 1310
rect 201 1208 235 1242
rect 201 1139 235 1174
rect 201 1089 235 1105
rect 289 1412 323 1450
rect 289 1344 323 1378
rect 289 1276 323 1310
rect 289 1208 323 1242
rect 289 1139 323 1174
rect 377 1412 411 1492
rect 377 1344 411 1378
rect 377 1276 411 1310
rect 377 1208 411 1242
rect 377 1157 411 1174
rect 465 1412 499 1450
rect 465 1344 499 1378
rect 465 1276 499 1310
rect 465 1208 499 1242
rect 289 1094 323 1105
rect 465 1139 499 1174
rect 553 1412 587 1492
rect 553 1344 587 1378
rect 553 1276 587 1310
rect 553 1208 587 1242
rect 553 1157 587 1174
rect 641 1412 675 1450
rect 641 1344 675 1378
rect 641 1276 675 1310
rect 641 1208 675 1242
rect 465 1094 499 1105
rect 641 1139 675 1174
rect 729 1412 763 1492
rect 729 1344 763 1378
rect 729 1276 763 1310
rect 729 1208 763 1242
rect 729 1157 763 1174
rect 931 1470 993 1492
rect 931 1436 945 1470
rect 979 1436 993 1470
rect 931 1398 993 1436
rect 931 1364 945 1398
rect 979 1364 993 1398
rect 931 1326 993 1364
rect 931 1292 945 1326
rect 979 1292 993 1326
rect 931 1254 993 1292
rect 931 1220 945 1254
rect 979 1220 993 1254
rect 931 1182 993 1220
rect 641 1094 675 1105
rect 931 1148 945 1182
rect 979 1148 993 1182
rect 931 1110 993 1148
rect -31 1038 31 1076
rect 289 1060 831 1094
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect -31 868 31 932
rect 205 1003 239 1019
rect 205 757 239 969
rect -31 546 31 572
rect -31 512 -17 546
rect 17 512 31 546
rect -31 474 31 512
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect 205 461 239 723
rect 205 411 239 427
rect 427 1003 461 1019
rect 427 831 461 969
rect 427 461 461 797
rect 427 411 461 427
rect 649 1003 683 1019
rect 649 609 683 969
rect 649 461 683 575
rect 649 411 683 427
rect 797 905 831 1060
rect -31 368 -17 402
rect 17 368 31 402
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect 101 363 135 379
rect 295 363 329 379
rect 489 363 523 379
rect 135 329 198 363
rect 232 329 295 363
rect 329 329 392 363
rect 426 329 489 363
rect 101 291 135 329
rect 101 223 135 257
rect 295 291 329 329
rect 489 313 523 329
rect 603 363 637 379
rect 797 378 831 871
rect 931 1076 945 1110
rect 979 1076 993 1110
rect 1163 1412 1197 1492
rect 1163 1344 1197 1378
rect 1163 1276 1197 1310
rect 1163 1208 1197 1242
rect 1163 1139 1197 1174
rect 1163 1089 1197 1105
rect 1251 1412 1285 1450
rect 1251 1344 1285 1378
rect 1251 1276 1285 1310
rect 1251 1208 1285 1242
rect 1251 1139 1285 1174
rect 1339 1412 1373 1492
rect 1339 1344 1373 1378
rect 1339 1276 1373 1310
rect 1339 1208 1373 1242
rect 1339 1157 1373 1174
rect 1427 1412 1461 1450
rect 1427 1344 1461 1378
rect 1427 1276 1461 1310
rect 1427 1208 1461 1242
rect 1251 1094 1285 1105
rect 1427 1139 1461 1174
rect 1515 1412 1549 1492
rect 1515 1344 1549 1378
rect 1515 1276 1549 1310
rect 1515 1208 1549 1242
rect 1515 1157 1549 1174
rect 1603 1412 1637 1450
rect 1603 1344 1637 1378
rect 1603 1276 1637 1310
rect 1603 1208 1637 1242
rect 1427 1094 1461 1105
rect 1603 1139 1637 1174
rect 1691 1412 1725 1492
rect 1691 1344 1725 1378
rect 1691 1276 1725 1310
rect 1691 1208 1725 1242
rect 1691 1157 1725 1174
rect 1893 1470 1955 1492
rect 1893 1436 1907 1470
rect 1941 1436 1955 1470
rect 1893 1398 1955 1436
rect 1893 1364 1907 1398
rect 1941 1364 1955 1398
rect 1893 1326 1955 1364
rect 1893 1292 1907 1326
rect 1941 1292 1955 1326
rect 1893 1254 1955 1292
rect 1893 1220 1907 1254
rect 1941 1220 1955 1254
rect 1893 1182 1955 1220
rect 1603 1094 1637 1105
rect 1893 1148 1907 1182
rect 1941 1148 1955 1182
rect 1893 1110 1955 1148
rect 931 1038 993 1076
rect 1251 1060 1793 1094
rect 931 1004 945 1038
rect 979 1004 993 1038
rect 931 966 993 1004
rect 931 932 945 966
rect 979 932 993 966
rect 931 868 993 932
rect 1167 1003 1201 1019
rect 1167 905 1201 969
rect 603 291 637 329
rect 101 153 135 189
rect 101 103 135 119
rect 198 238 232 254
rect -31 62 31 80
rect 198 62 232 204
rect 295 223 329 257
rect 393 244 427 260
rect 603 244 637 257
rect 427 223 637 244
rect 427 210 603 223
rect 393 194 427 210
rect 295 153 329 189
rect 700 344 831 378
rect 931 546 993 572
rect 931 512 945 546
rect 979 512 993 546
rect 931 474 993 512
rect 931 440 945 474
rect 979 440 993 474
rect 931 402 993 440
rect 1167 461 1201 871
rect 1167 411 1201 427
rect 1389 1003 1423 1019
rect 1389 461 1423 969
rect 1389 411 1423 427
rect 1611 1003 1645 1019
rect 1611 683 1645 969
rect 1611 461 1645 649
rect 1611 411 1645 427
rect 1759 609 1793 1060
rect 1893 1076 1907 1110
rect 1941 1076 1955 1110
rect 1893 1038 1955 1076
rect 2065 1412 2099 1492
rect 2065 1344 2099 1378
rect 2065 1276 2099 1310
rect 2065 1208 2099 1242
rect 2065 1139 2099 1174
rect 2065 1073 2099 1105
rect 2153 1412 2187 1450
rect 2153 1344 2187 1378
rect 2153 1276 2187 1310
rect 2153 1208 2187 1242
rect 2153 1139 2187 1174
rect 2241 1412 2275 1492
rect 2241 1344 2275 1378
rect 2241 1276 2275 1310
rect 2241 1208 2275 1242
rect 2241 1157 2275 1174
rect 2329 1412 2363 1450
rect 2329 1344 2363 1378
rect 2329 1276 2363 1310
rect 2329 1208 2363 1242
rect 2153 1103 2187 1105
rect 2329 1139 2363 1174
rect 2417 1412 2451 1492
rect 2417 1344 2451 1378
rect 2417 1276 2451 1310
rect 2417 1208 2451 1242
rect 2417 1157 2451 1174
rect 2559 1470 2621 1492
rect 2559 1436 2573 1470
rect 2607 1436 2621 1470
rect 2559 1398 2621 1436
rect 2559 1364 2573 1398
rect 2607 1364 2621 1398
rect 2559 1326 2621 1364
rect 2559 1292 2573 1326
rect 2607 1292 2621 1326
rect 2559 1254 2621 1292
rect 2559 1220 2573 1254
rect 2607 1220 2621 1254
rect 2559 1182 2621 1220
rect 2329 1103 2363 1105
rect 2559 1148 2573 1182
rect 2607 1148 2621 1182
rect 2559 1110 2621 1148
rect 2153 1069 2459 1103
rect 1893 1004 1907 1038
rect 1941 1004 1955 1038
rect 1893 966 1955 1004
rect 1893 932 1907 966
rect 1941 932 1955 966
rect 1893 868 1955 932
rect 2129 1003 2163 1019
rect 2283 1003 2317 1019
rect 931 368 945 402
rect 979 368 993 402
rect 700 247 734 344
rect 931 330 993 368
rect 700 197 734 213
rect 797 291 831 307
rect 797 223 831 257
rect 489 153 523 169
rect 329 119 392 153
rect 426 119 489 153
rect 295 103 329 119
rect 489 103 523 119
rect 603 153 637 189
rect 797 153 831 189
rect 637 119 700 153
rect 734 119 797 153
rect 603 103 637 119
rect 797 103 831 119
rect 931 296 945 330
rect 979 296 993 330
rect 931 258 993 296
rect 931 224 945 258
rect 979 224 993 258
rect 931 186 993 224
rect 931 152 945 186
rect 979 152 993 186
rect 931 114 993 152
rect 931 80 945 114
rect 979 80 993 114
rect 1063 363 1097 379
rect 1257 363 1291 379
rect 1451 363 1485 379
rect 1097 329 1160 363
rect 1194 329 1257 363
rect 1291 329 1354 363
rect 1388 329 1451 363
rect 1063 291 1097 329
rect 1063 223 1097 257
rect 1257 291 1291 329
rect 1451 313 1485 329
rect 1565 363 1599 379
rect 1759 378 1793 575
rect 2129 609 2163 969
rect 1565 291 1599 329
rect 1063 153 1097 189
rect 1063 103 1097 119
rect 1160 238 1194 254
rect 931 62 993 80
rect 1160 62 1194 204
rect 1257 223 1291 257
rect 1355 244 1389 260
rect 1565 244 1599 257
rect 1389 223 1599 244
rect 1389 210 1565 223
rect 1355 194 1389 210
rect 1257 153 1291 189
rect 1662 344 1793 378
rect 1893 546 1955 572
rect 1893 512 1907 546
rect 1941 512 1955 546
rect 1893 474 1955 512
rect 1893 440 1907 474
rect 1941 440 1955 474
rect 1893 402 1955 440
rect 2129 461 2163 575
rect 2129 411 2163 427
rect 2277 969 2283 988
rect 2277 953 2317 969
rect 2277 757 2311 953
rect 2277 461 2311 723
rect 2277 411 2311 427
rect 2425 609 2459 1069
rect 2559 1076 2573 1110
rect 2607 1076 2621 1110
rect 2791 1412 2825 1492
rect 2791 1344 2825 1378
rect 2791 1276 2825 1310
rect 2791 1208 2825 1242
rect 2791 1139 2825 1174
rect 2791 1089 2825 1105
rect 2879 1412 2913 1450
rect 2879 1344 2913 1378
rect 2879 1276 2913 1310
rect 2879 1208 2913 1242
rect 2879 1139 2913 1174
rect 2967 1412 3001 1492
rect 2967 1344 3001 1378
rect 2967 1276 3001 1310
rect 2967 1208 3001 1242
rect 2967 1157 3001 1174
rect 3055 1412 3089 1450
rect 3055 1344 3089 1378
rect 3055 1276 3089 1310
rect 3055 1208 3089 1242
rect 2879 1094 2913 1105
rect 3055 1139 3089 1174
rect 3143 1412 3177 1492
rect 3143 1344 3177 1378
rect 3143 1276 3177 1310
rect 3143 1208 3177 1242
rect 3143 1157 3177 1174
rect 3231 1412 3265 1450
rect 3231 1344 3265 1378
rect 3231 1276 3265 1310
rect 3231 1208 3265 1242
rect 3055 1094 3089 1105
rect 3231 1139 3265 1174
rect 3319 1412 3353 1492
rect 3319 1344 3353 1378
rect 3319 1276 3353 1310
rect 3319 1208 3353 1242
rect 3319 1157 3353 1174
rect 3521 1470 3583 1492
rect 3521 1436 3535 1470
rect 3569 1436 3583 1470
rect 3521 1398 3583 1436
rect 3521 1364 3535 1398
rect 3569 1364 3583 1398
rect 3521 1326 3583 1364
rect 3521 1292 3535 1326
rect 3569 1292 3583 1326
rect 3521 1254 3583 1292
rect 3521 1220 3535 1254
rect 3569 1220 3583 1254
rect 3521 1182 3583 1220
rect 3231 1094 3265 1105
rect 3521 1148 3535 1182
rect 3569 1148 3583 1182
rect 3521 1110 3583 1148
rect 2559 1038 2621 1076
rect 2879 1060 3421 1094
rect 2559 1004 2573 1038
rect 2607 1004 2621 1038
rect 2559 966 2621 1004
rect 2559 932 2573 966
rect 2607 932 2621 966
rect 2559 868 2621 932
rect 2795 1003 2829 1019
rect 1893 368 1907 402
rect 1941 368 1955 402
rect 1662 247 1696 344
rect 1893 330 1955 368
rect 1662 197 1696 213
rect 1759 291 1793 307
rect 1759 223 1793 257
rect 1451 153 1485 169
rect 1291 119 1354 153
rect 1388 119 1451 153
rect 1257 103 1291 119
rect 1451 103 1485 119
rect 1565 153 1599 189
rect 1759 153 1793 189
rect 1599 119 1662 153
rect 1696 119 1759 153
rect 1565 103 1599 119
rect 1759 103 1793 119
rect 1893 296 1907 330
rect 1941 296 1955 330
rect 1893 258 1955 296
rect 1893 224 1907 258
rect 1941 224 1955 258
rect 1893 186 1955 224
rect 1893 152 1907 186
rect 1941 152 1955 186
rect 1893 114 1955 152
rect 1893 80 1907 114
rect 1941 80 1955 114
rect 2046 361 2080 377
rect 2240 361 2274 377
rect 2425 376 2459 575
rect 2795 609 2829 969
rect 2080 327 2143 361
rect 2177 327 2240 361
rect 2046 289 2080 327
rect 2046 221 2080 255
rect 2240 289 2274 327
rect 2046 151 2080 187
rect 2046 101 2080 117
rect 2143 236 2177 252
rect 1893 62 1955 80
rect 2143 62 2177 202
rect 2240 221 2274 255
rect 2337 342 2459 376
rect 2559 546 2621 572
rect 2559 512 2573 546
rect 2607 512 2621 546
rect 2559 474 2621 512
rect 2559 440 2573 474
rect 2607 440 2621 474
rect 2559 402 2621 440
rect 2795 461 2829 575
rect 2795 411 2829 427
rect 3017 1003 3051 1019
rect 3017 831 3051 969
rect 3017 461 3051 797
rect 3017 411 3051 427
rect 3239 1003 3273 1019
rect 3239 683 3273 969
rect 3239 461 3273 649
rect 3239 411 3273 427
rect 3387 757 3421 1060
rect 3521 1076 3535 1110
rect 3569 1076 3583 1110
rect 3753 1412 3787 1492
rect 3753 1344 3787 1378
rect 3753 1276 3787 1310
rect 3753 1208 3787 1242
rect 3753 1139 3787 1174
rect 3753 1089 3787 1105
rect 3841 1412 3875 1450
rect 3841 1344 3875 1378
rect 3841 1276 3875 1310
rect 3841 1208 3875 1242
rect 3841 1139 3875 1174
rect 3929 1412 3963 1492
rect 3929 1344 3963 1378
rect 3929 1276 3963 1310
rect 3929 1208 3963 1242
rect 3929 1157 3963 1174
rect 4017 1412 4051 1450
rect 4017 1344 4051 1378
rect 4017 1276 4051 1310
rect 4017 1208 4051 1242
rect 3841 1094 3875 1105
rect 4017 1139 4051 1174
rect 4105 1412 4139 1492
rect 4105 1344 4139 1378
rect 4105 1276 4139 1310
rect 4105 1208 4139 1242
rect 4105 1157 4139 1174
rect 4193 1412 4227 1450
rect 4193 1344 4227 1378
rect 4193 1276 4227 1310
rect 4193 1208 4227 1242
rect 4017 1094 4051 1105
rect 4193 1139 4227 1174
rect 4281 1412 4315 1492
rect 4281 1344 4315 1378
rect 4281 1276 4315 1310
rect 4281 1208 4315 1242
rect 4281 1157 4315 1174
rect 4483 1470 4545 1492
rect 4483 1436 4497 1470
rect 4531 1436 4545 1470
rect 4483 1398 4545 1436
rect 4483 1364 4497 1398
rect 4531 1364 4545 1398
rect 4483 1326 4545 1364
rect 4483 1292 4497 1326
rect 4531 1292 4545 1326
rect 4483 1254 4545 1292
rect 4483 1220 4497 1254
rect 4531 1220 4545 1254
rect 4483 1182 4545 1220
rect 4193 1094 4227 1105
rect 4483 1148 4497 1182
rect 4531 1148 4545 1182
rect 4483 1110 4545 1148
rect 3521 1038 3583 1076
rect 3841 1060 4383 1094
rect 3521 1004 3535 1038
rect 3569 1004 3583 1038
rect 3521 966 3583 1004
rect 3521 932 3535 966
rect 3569 932 3583 966
rect 3521 868 3583 932
rect 3757 1003 3791 1019
rect 3757 905 3791 969
rect 2559 368 2573 402
rect 2607 368 2621 402
rect 2337 245 2371 342
rect 2559 330 2621 368
rect 2337 195 2371 211
rect 2434 289 2468 305
rect 2434 221 2468 255
rect 2240 151 2274 187
rect 2434 151 2468 187
rect 2274 117 2337 151
rect 2371 117 2434 151
rect 2240 101 2274 117
rect 2434 101 2468 117
rect 2559 296 2573 330
rect 2607 296 2621 330
rect 2559 258 2621 296
rect 2559 224 2573 258
rect 2607 224 2621 258
rect 2559 186 2621 224
rect 2559 152 2573 186
rect 2607 152 2621 186
rect 2559 114 2621 152
rect 2559 80 2573 114
rect 2607 80 2621 114
rect 2691 363 2725 379
rect 2885 363 2919 379
rect 3079 363 3113 379
rect 2725 329 2788 363
rect 2822 329 2885 363
rect 2919 329 2982 363
rect 3016 329 3079 363
rect 2691 291 2725 329
rect 2691 223 2725 257
rect 2885 291 2919 329
rect 3079 313 3113 329
rect 3193 363 3227 379
rect 3387 378 3421 723
rect 3193 291 3227 329
rect 2691 153 2725 189
rect 2691 103 2725 119
rect 2788 238 2822 254
rect 2559 62 2621 80
rect 2788 62 2822 204
rect 2885 223 2919 257
rect 2983 244 3017 260
rect 3193 244 3227 257
rect 3017 223 3227 244
rect 3017 210 3193 223
rect 2983 194 3017 210
rect 2885 153 2919 189
rect 3290 344 3421 378
rect 3521 546 3583 572
rect 3521 512 3535 546
rect 3569 512 3583 546
rect 3521 474 3583 512
rect 3521 440 3535 474
rect 3569 440 3583 474
rect 3521 402 3583 440
rect 3757 461 3791 871
rect 3757 411 3791 427
rect 3979 1003 4013 1019
rect 3979 683 4013 969
rect 3979 461 4013 649
rect 3979 411 4013 427
rect 4201 1003 4235 1019
rect 4201 461 4235 945
rect 4201 411 4235 427
rect 4349 905 4383 1060
rect 3521 368 3535 402
rect 3569 368 3583 402
rect 3290 247 3324 344
rect 3521 330 3583 368
rect 3290 197 3324 213
rect 3387 291 3421 307
rect 3387 223 3421 257
rect 3079 153 3113 169
rect 2919 119 2982 153
rect 3016 119 3079 153
rect 2885 103 2919 119
rect 3079 103 3113 119
rect 3193 153 3227 189
rect 3387 153 3421 189
rect 3227 119 3290 153
rect 3324 119 3387 153
rect 3193 103 3227 119
rect 3387 103 3421 119
rect 3521 296 3535 330
rect 3569 296 3583 330
rect 3521 258 3583 296
rect 3521 224 3535 258
rect 3569 224 3583 258
rect 3521 186 3583 224
rect 3521 152 3535 186
rect 3569 152 3583 186
rect 3521 114 3583 152
rect 3521 80 3535 114
rect 3569 80 3583 114
rect 3653 363 3687 379
rect 3847 363 3881 379
rect 4041 363 4075 379
rect 3687 329 3750 363
rect 3784 329 3847 363
rect 3881 329 3944 363
rect 3978 329 4041 363
rect 3653 291 3687 329
rect 3653 223 3687 257
rect 3847 291 3881 329
rect 4041 313 4075 329
rect 4155 363 4189 379
rect 4349 378 4383 871
rect 4483 1076 4497 1110
rect 4531 1076 4545 1110
rect 4483 1038 4545 1076
rect 4655 1412 4689 1492
rect 4655 1344 4689 1378
rect 4655 1276 4689 1310
rect 4655 1208 4689 1242
rect 4655 1139 4689 1174
rect 4655 1073 4689 1105
rect 4743 1412 4777 1450
rect 4743 1344 4777 1378
rect 4743 1276 4777 1310
rect 4743 1208 4777 1242
rect 4743 1139 4777 1174
rect 4831 1412 4865 1492
rect 4831 1344 4865 1378
rect 4831 1276 4865 1310
rect 4831 1208 4865 1242
rect 4831 1157 4865 1174
rect 4919 1412 4953 1450
rect 4919 1344 4953 1378
rect 4919 1276 4953 1310
rect 4919 1208 4953 1242
rect 4743 1103 4777 1105
rect 4919 1139 4953 1174
rect 5007 1412 5041 1492
rect 5007 1344 5041 1378
rect 5007 1276 5041 1310
rect 5007 1208 5041 1242
rect 5007 1157 5041 1174
rect 5149 1470 5211 1492
rect 5149 1436 5163 1470
rect 5197 1436 5211 1470
rect 5149 1398 5211 1436
rect 5149 1364 5163 1398
rect 5197 1364 5211 1398
rect 5149 1326 5211 1364
rect 5149 1292 5163 1326
rect 5197 1292 5211 1326
rect 5149 1254 5211 1292
rect 5149 1220 5163 1254
rect 5197 1220 5211 1254
rect 5149 1182 5211 1220
rect 4919 1103 4953 1105
rect 5149 1148 5163 1182
rect 5197 1148 5211 1182
rect 5149 1110 5211 1148
rect 4743 1069 5049 1103
rect 4483 1004 4497 1038
rect 4531 1004 4545 1038
rect 4483 966 4545 1004
rect 4483 932 4497 966
rect 4531 932 4545 966
rect 4483 868 4545 932
rect 4719 1003 4753 1019
rect 4873 1003 4907 1019
rect 4719 905 4753 969
rect 4155 291 4189 329
rect 3653 153 3687 189
rect 3653 103 3687 119
rect 3750 238 3784 254
rect 3521 62 3583 80
rect 3750 62 3784 204
rect 3847 223 3881 257
rect 3945 244 3979 260
rect 4155 244 4189 257
rect 3979 223 4189 244
rect 3979 210 4155 223
rect 3945 194 3979 210
rect 3847 153 3881 189
rect 4252 344 4383 378
rect 4483 546 4545 572
rect 4483 512 4497 546
rect 4531 512 4545 546
rect 4483 474 4545 512
rect 4483 440 4497 474
rect 4531 440 4545 474
rect 4483 402 4545 440
rect 4719 461 4753 871
rect 4719 411 4753 427
rect 4867 969 4873 988
rect 4867 953 4907 969
rect 5015 979 5049 1069
rect 4867 757 4901 953
rect 4867 461 4901 723
rect 4867 411 4901 427
rect 4483 368 4497 402
rect 4531 368 4545 402
rect 4252 247 4286 344
rect 4483 330 4545 368
rect 4252 197 4286 213
rect 4349 291 4383 307
rect 4349 223 4383 257
rect 4041 153 4075 169
rect 3881 119 3944 153
rect 3978 119 4041 153
rect 3847 103 3881 119
rect 4041 103 4075 119
rect 4155 153 4189 189
rect 4349 153 4383 189
rect 4189 119 4252 153
rect 4286 119 4349 153
rect 4155 103 4189 119
rect 4349 103 4383 119
rect 4483 296 4497 330
rect 4531 296 4545 330
rect 4483 258 4545 296
rect 4483 224 4497 258
rect 4531 224 4545 258
rect 4483 186 4545 224
rect 4483 152 4497 186
rect 4531 152 4545 186
rect 4483 114 4545 152
rect 4483 80 4497 114
rect 4531 80 4545 114
rect 4636 361 4670 377
rect 4830 361 4864 377
rect 5015 376 5049 945
rect 5149 1076 5163 1110
rect 5197 1076 5211 1110
rect 5381 1412 5415 1492
rect 5381 1344 5415 1378
rect 5381 1276 5415 1310
rect 5381 1208 5415 1242
rect 5381 1139 5415 1174
rect 5381 1089 5415 1105
rect 5469 1412 5503 1450
rect 5469 1344 5503 1378
rect 5469 1276 5503 1310
rect 5469 1208 5503 1242
rect 5469 1139 5503 1174
rect 5557 1412 5591 1492
rect 5557 1344 5591 1378
rect 5557 1276 5591 1310
rect 5557 1208 5591 1242
rect 5557 1157 5591 1174
rect 5645 1412 5679 1450
rect 5645 1344 5679 1378
rect 5645 1276 5679 1310
rect 5645 1208 5679 1242
rect 5469 1094 5503 1105
rect 5645 1139 5679 1174
rect 5733 1412 5767 1492
rect 5733 1344 5767 1378
rect 5733 1276 5767 1310
rect 5733 1208 5767 1242
rect 5733 1157 5767 1174
rect 5821 1412 5855 1450
rect 5821 1344 5855 1378
rect 5821 1276 5855 1310
rect 5821 1208 5855 1242
rect 5645 1094 5679 1105
rect 5821 1139 5855 1174
rect 5909 1412 5943 1492
rect 5909 1344 5943 1378
rect 5909 1276 5943 1310
rect 5909 1208 5943 1242
rect 5909 1157 5943 1174
rect 6111 1470 6173 1492
rect 6111 1436 6125 1470
rect 6159 1436 6173 1470
rect 6111 1398 6173 1436
rect 6111 1364 6125 1398
rect 6159 1364 6173 1398
rect 6111 1326 6173 1364
rect 6111 1292 6125 1326
rect 6159 1292 6173 1326
rect 6111 1254 6173 1292
rect 6111 1220 6125 1254
rect 6159 1220 6173 1254
rect 6111 1182 6173 1220
rect 5821 1094 5855 1105
rect 6111 1148 6125 1182
rect 6159 1148 6173 1182
rect 6111 1110 6173 1148
rect 5149 1038 5211 1076
rect 5469 1060 6011 1094
rect 5149 1004 5163 1038
rect 5197 1004 5211 1038
rect 5149 966 5211 1004
rect 5149 932 5163 966
rect 5197 932 5211 966
rect 5149 868 5211 932
rect 5385 1003 5419 1019
rect 5385 757 5419 969
rect 4670 327 4733 361
rect 4767 327 4830 361
rect 4636 289 4670 327
rect 4636 221 4670 255
rect 4830 289 4864 327
rect 4636 151 4670 187
rect 4636 101 4670 117
rect 4733 236 4767 252
rect 4483 62 4545 80
rect 4733 62 4767 202
rect 4830 221 4864 255
rect 4927 342 5049 376
rect 5149 546 5211 572
rect 5149 512 5163 546
rect 5197 512 5211 546
rect 5149 474 5211 512
rect 5149 440 5163 474
rect 5197 440 5211 474
rect 5149 402 5211 440
rect 5385 461 5419 723
rect 5385 411 5419 427
rect 5607 1003 5641 1019
rect 5607 831 5641 969
rect 5607 461 5641 797
rect 5607 411 5641 427
rect 5829 1003 5863 1019
rect 5829 609 5863 969
rect 5829 461 5863 575
rect 5829 411 5863 427
rect 5977 905 6011 1060
rect 5149 368 5163 402
rect 5197 368 5211 402
rect 4927 245 4961 342
rect 5149 330 5211 368
rect 4927 195 4961 211
rect 5024 289 5058 305
rect 5024 221 5058 255
rect 4830 151 4864 187
rect 5024 151 5058 187
rect 4864 117 4927 151
rect 4961 117 5024 151
rect 4830 101 4864 117
rect 5024 101 5058 117
rect 5149 296 5163 330
rect 5197 296 5211 330
rect 5149 258 5211 296
rect 5149 224 5163 258
rect 5197 224 5211 258
rect 5149 186 5211 224
rect 5149 152 5163 186
rect 5197 152 5211 186
rect 5149 114 5211 152
rect 5149 80 5163 114
rect 5197 80 5211 114
rect 5281 363 5315 379
rect 5475 363 5509 379
rect 5669 363 5703 379
rect 5315 329 5378 363
rect 5412 329 5475 363
rect 5509 329 5572 363
rect 5606 329 5669 363
rect 5281 291 5315 329
rect 5281 223 5315 257
rect 5475 291 5509 329
rect 5669 313 5703 329
rect 5783 363 5817 379
rect 5977 378 6011 871
rect 6111 1076 6125 1110
rect 6159 1076 6173 1110
rect 6343 1412 6377 1492
rect 6343 1344 6377 1378
rect 6343 1276 6377 1310
rect 6343 1208 6377 1242
rect 6343 1139 6377 1174
rect 6343 1089 6377 1105
rect 6431 1412 6465 1450
rect 6431 1344 6465 1378
rect 6431 1276 6465 1310
rect 6431 1208 6465 1242
rect 6431 1139 6465 1174
rect 6519 1412 6553 1492
rect 6519 1344 6553 1378
rect 6519 1276 6553 1310
rect 6519 1208 6553 1242
rect 6519 1157 6553 1174
rect 6607 1412 6641 1450
rect 6607 1344 6641 1378
rect 6607 1276 6641 1310
rect 6607 1208 6641 1242
rect 6431 1094 6465 1105
rect 6607 1139 6641 1174
rect 6695 1412 6729 1492
rect 6695 1344 6729 1378
rect 6695 1276 6729 1310
rect 6695 1208 6729 1242
rect 6695 1157 6729 1174
rect 6783 1412 6817 1450
rect 6783 1344 6817 1378
rect 6783 1276 6817 1310
rect 6783 1208 6817 1242
rect 6607 1094 6641 1105
rect 6783 1139 6817 1174
rect 6871 1412 6905 1492
rect 6871 1344 6905 1378
rect 6871 1276 6905 1310
rect 6871 1208 6905 1242
rect 6871 1157 6905 1174
rect 7073 1470 7135 1492
rect 7073 1436 7087 1470
rect 7121 1436 7135 1470
rect 7073 1398 7135 1436
rect 7073 1364 7087 1398
rect 7121 1364 7135 1398
rect 7073 1326 7135 1364
rect 7073 1292 7087 1326
rect 7121 1292 7135 1326
rect 7073 1254 7135 1292
rect 7073 1220 7087 1254
rect 7121 1220 7135 1254
rect 7073 1182 7135 1220
rect 6783 1094 6817 1105
rect 7073 1148 7087 1182
rect 7121 1148 7135 1182
rect 7073 1110 7135 1148
rect 6111 1038 6173 1076
rect 6431 1060 6973 1094
rect 6111 1004 6125 1038
rect 6159 1004 6173 1038
rect 6111 966 6173 1004
rect 6111 932 6125 966
rect 6159 932 6173 966
rect 6111 868 6173 932
rect 6347 1003 6381 1019
rect 6347 905 6381 969
rect 5783 291 5817 329
rect 5281 153 5315 189
rect 5281 103 5315 119
rect 5378 238 5412 254
rect 5149 62 5211 80
rect 5378 62 5412 204
rect 5475 223 5509 257
rect 5573 244 5607 260
rect 5783 244 5817 257
rect 5607 223 5817 244
rect 5607 210 5783 223
rect 5573 194 5607 210
rect 5475 153 5509 189
rect 5880 344 6011 378
rect 6111 546 6173 572
rect 6111 512 6125 546
rect 6159 512 6173 546
rect 6111 474 6173 512
rect 6111 440 6125 474
rect 6159 440 6173 474
rect 6111 402 6173 440
rect 6347 461 6381 871
rect 6347 411 6381 427
rect 6569 1003 6603 1019
rect 6569 461 6603 969
rect 6569 411 6603 427
rect 6791 1003 6825 1019
rect 6791 683 6825 969
rect 6791 461 6825 649
rect 6791 411 6825 427
rect 6939 609 6973 1060
rect 7073 1076 7087 1110
rect 7121 1076 7135 1110
rect 7073 1038 7135 1076
rect 7245 1412 7279 1492
rect 7245 1344 7279 1378
rect 7245 1276 7279 1310
rect 7245 1208 7279 1242
rect 7245 1139 7279 1174
rect 7245 1073 7279 1105
rect 7333 1412 7367 1450
rect 7333 1344 7367 1378
rect 7333 1276 7367 1310
rect 7333 1208 7367 1242
rect 7333 1139 7367 1174
rect 7421 1412 7455 1492
rect 7421 1344 7455 1378
rect 7421 1276 7455 1310
rect 7421 1208 7455 1242
rect 7421 1157 7455 1174
rect 7509 1412 7543 1450
rect 7509 1344 7543 1378
rect 7509 1276 7543 1310
rect 7509 1208 7543 1242
rect 7333 1103 7367 1105
rect 7509 1139 7543 1174
rect 7597 1412 7631 1492
rect 7597 1344 7631 1378
rect 7597 1276 7631 1310
rect 7597 1208 7631 1242
rect 7597 1157 7631 1174
rect 7739 1470 7801 1492
rect 7739 1436 7753 1470
rect 7787 1436 7801 1470
rect 7739 1398 7801 1436
rect 7739 1364 7753 1398
rect 7787 1364 7801 1398
rect 7739 1326 7801 1364
rect 7739 1292 7753 1326
rect 7787 1292 7801 1326
rect 7739 1254 7801 1292
rect 7739 1220 7753 1254
rect 7787 1220 7801 1254
rect 7739 1182 7801 1220
rect 7509 1103 7543 1105
rect 7739 1148 7753 1182
rect 7787 1148 7801 1182
rect 7739 1110 7801 1148
rect 7333 1069 7639 1103
rect 7073 1004 7087 1038
rect 7121 1004 7135 1038
rect 7073 966 7135 1004
rect 7073 932 7087 966
rect 7121 932 7135 966
rect 7073 868 7135 932
rect 7309 1003 7343 1019
rect 7463 1003 7497 1019
rect 6111 368 6125 402
rect 6159 368 6173 402
rect 5880 247 5914 344
rect 6111 330 6173 368
rect 5880 197 5914 213
rect 5977 291 6011 307
rect 5977 223 6011 257
rect 5669 153 5703 169
rect 5509 119 5572 153
rect 5606 119 5669 153
rect 5475 103 5509 119
rect 5669 103 5703 119
rect 5783 153 5817 189
rect 5977 153 6011 189
rect 5817 119 5880 153
rect 5914 119 5977 153
rect 5783 103 5817 119
rect 5977 103 6011 119
rect 6111 296 6125 330
rect 6159 296 6173 330
rect 6111 258 6173 296
rect 6111 224 6125 258
rect 6159 224 6173 258
rect 6111 186 6173 224
rect 6111 152 6125 186
rect 6159 152 6173 186
rect 6111 114 6173 152
rect 6111 80 6125 114
rect 6159 80 6173 114
rect 6243 363 6277 379
rect 6437 363 6471 379
rect 6631 363 6665 379
rect 6277 329 6340 363
rect 6374 329 6437 363
rect 6471 329 6534 363
rect 6568 329 6631 363
rect 6243 291 6277 329
rect 6243 223 6277 257
rect 6437 291 6471 329
rect 6631 313 6665 329
rect 6745 363 6779 379
rect 6939 378 6973 575
rect 7309 609 7343 969
rect 6745 291 6779 329
rect 6243 153 6277 189
rect 6243 103 6277 119
rect 6340 238 6374 254
rect 6111 62 6173 80
rect 6340 62 6374 204
rect 6437 223 6471 257
rect 6535 244 6569 260
rect 6745 244 6779 257
rect 6569 223 6779 244
rect 6569 210 6745 223
rect 6535 194 6569 210
rect 6437 153 6471 189
rect 6842 344 6973 378
rect 7073 546 7135 572
rect 7073 512 7087 546
rect 7121 512 7135 546
rect 7073 474 7135 512
rect 7073 440 7087 474
rect 7121 440 7135 474
rect 7073 402 7135 440
rect 7309 461 7343 575
rect 7309 411 7343 427
rect 7457 969 7463 988
rect 7457 953 7497 969
rect 7457 757 7491 953
rect 7457 461 7491 723
rect 7457 411 7491 427
rect 7605 609 7639 1069
rect 7739 1076 7753 1110
rect 7787 1076 7801 1110
rect 7971 1412 8005 1492
rect 7971 1344 8005 1378
rect 7971 1276 8005 1310
rect 7971 1208 8005 1242
rect 7971 1139 8005 1174
rect 7971 1089 8005 1105
rect 8059 1412 8093 1450
rect 8059 1344 8093 1378
rect 8059 1276 8093 1310
rect 8059 1208 8093 1242
rect 8059 1139 8093 1174
rect 8147 1412 8181 1492
rect 8147 1344 8181 1378
rect 8147 1276 8181 1310
rect 8147 1208 8181 1242
rect 8147 1157 8181 1174
rect 8235 1412 8269 1450
rect 8235 1344 8269 1378
rect 8235 1276 8269 1310
rect 8235 1208 8269 1242
rect 8059 1094 8093 1105
rect 8235 1139 8269 1174
rect 8323 1412 8357 1492
rect 8323 1344 8357 1378
rect 8323 1276 8357 1310
rect 8323 1208 8357 1242
rect 8323 1157 8357 1174
rect 8411 1412 8445 1450
rect 8411 1344 8445 1378
rect 8411 1276 8445 1310
rect 8411 1208 8445 1242
rect 8235 1094 8269 1105
rect 8411 1139 8445 1174
rect 8499 1412 8533 1492
rect 8499 1344 8533 1378
rect 8499 1276 8533 1310
rect 8499 1208 8533 1242
rect 8499 1157 8533 1174
rect 8701 1470 8763 1492
rect 8701 1436 8715 1470
rect 8749 1436 8763 1470
rect 8701 1398 8763 1436
rect 8701 1364 8715 1398
rect 8749 1364 8763 1398
rect 8701 1326 8763 1364
rect 8701 1292 8715 1326
rect 8749 1292 8763 1326
rect 8701 1254 8763 1292
rect 8701 1220 8715 1254
rect 8749 1220 8763 1254
rect 8701 1182 8763 1220
rect 8411 1094 8445 1105
rect 8701 1148 8715 1182
rect 8749 1148 8763 1182
rect 8701 1110 8763 1148
rect 7739 1038 7801 1076
rect 8059 1060 8601 1094
rect 7739 1004 7753 1038
rect 7787 1004 7801 1038
rect 7739 966 7801 1004
rect 7739 932 7753 966
rect 7787 932 7801 966
rect 7739 868 7801 932
rect 7975 1003 8009 1019
rect 7073 368 7087 402
rect 7121 368 7135 402
rect 6842 247 6876 344
rect 7073 330 7135 368
rect 6842 197 6876 213
rect 6939 291 6973 307
rect 6939 223 6973 257
rect 6631 153 6665 169
rect 6471 119 6534 153
rect 6568 119 6631 153
rect 6437 103 6471 119
rect 6631 103 6665 119
rect 6745 153 6779 189
rect 6939 153 6973 189
rect 6779 119 6842 153
rect 6876 119 6939 153
rect 6745 103 6779 119
rect 6939 103 6973 119
rect 7073 296 7087 330
rect 7121 296 7135 330
rect 7073 258 7135 296
rect 7073 224 7087 258
rect 7121 224 7135 258
rect 7073 186 7135 224
rect 7073 152 7087 186
rect 7121 152 7135 186
rect 7073 114 7135 152
rect 7073 80 7087 114
rect 7121 80 7135 114
rect 7226 361 7260 377
rect 7420 361 7454 377
rect 7605 376 7639 575
rect 7975 609 8009 969
rect 7260 327 7323 361
rect 7357 327 7420 361
rect 7226 289 7260 327
rect 7226 221 7260 255
rect 7420 289 7454 327
rect 7226 151 7260 187
rect 7226 101 7260 117
rect 7323 236 7357 252
rect 7073 62 7135 80
rect 7323 62 7357 202
rect 7420 221 7454 255
rect 7517 342 7639 376
rect 7739 546 7801 572
rect 7739 512 7753 546
rect 7787 512 7801 546
rect 7739 474 7801 512
rect 7739 440 7753 474
rect 7787 440 7801 474
rect 7739 402 7801 440
rect 7975 461 8009 575
rect 7975 411 8009 427
rect 8197 1003 8231 1019
rect 8197 831 8231 969
rect 8197 461 8231 797
rect 8197 411 8231 427
rect 8419 1003 8453 1019
rect 8419 683 8453 969
rect 8419 461 8453 649
rect 8419 411 8453 427
rect 8567 757 8601 1060
rect 8701 1076 8715 1110
rect 8749 1076 8763 1110
rect 8933 1412 8967 1492
rect 8933 1344 8967 1378
rect 8933 1276 8967 1310
rect 8933 1208 8967 1242
rect 8933 1139 8967 1174
rect 8933 1089 8967 1105
rect 9021 1412 9055 1450
rect 9021 1344 9055 1378
rect 9021 1276 9055 1310
rect 9021 1208 9055 1242
rect 9021 1139 9055 1174
rect 9109 1412 9143 1492
rect 9109 1344 9143 1378
rect 9109 1276 9143 1310
rect 9109 1208 9143 1242
rect 9109 1157 9143 1174
rect 9197 1412 9231 1450
rect 9197 1344 9231 1378
rect 9197 1276 9231 1310
rect 9197 1208 9231 1242
rect 9021 1094 9055 1105
rect 9197 1139 9231 1174
rect 9285 1412 9319 1492
rect 9285 1344 9319 1378
rect 9285 1276 9319 1310
rect 9285 1208 9319 1242
rect 9285 1157 9319 1174
rect 9373 1412 9407 1450
rect 9373 1344 9407 1378
rect 9373 1276 9407 1310
rect 9373 1208 9407 1242
rect 9197 1094 9231 1105
rect 9373 1139 9407 1174
rect 9461 1412 9495 1492
rect 9461 1344 9495 1378
rect 9461 1276 9495 1310
rect 9461 1208 9495 1242
rect 9461 1157 9495 1174
rect 9663 1470 9725 1492
rect 9663 1436 9677 1470
rect 9711 1436 9725 1470
rect 9663 1398 9725 1436
rect 9663 1364 9677 1398
rect 9711 1364 9725 1398
rect 9663 1326 9725 1364
rect 9663 1292 9677 1326
rect 9711 1292 9725 1326
rect 9663 1254 9725 1292
rect 9663 1220 9677 1254
rect 9711 1220 9725 1254
rect 9663 1182 9725 1220
rect 9373 1094 9407 1105
rect 9663 1148 9677 1182
rect 9711 1148 9725 1182
rect 9663 1110 9725 1148
rect 8701 1038 8763 1076
rect 9021 1060 9563 1094
rect 8701 1004 8715 1038
rect 8749 1004 8763 1038
rect 8701 966 8763 1004
rect 8701 932 8715 966
rect 8749 932 8763 966
rect 8701 868 8763 932
rect 8937 1003 8971 1019
rect 8937 905 8971 969
rect 7739 368 7753 402
rect 7787 368 7801 402
rect 7517 245 7551 342
rect 7739 330 7801 368
rect 7517 195 7551 211
rect 7614 289 7648 305
rect 7614 221 7648 255
rect 7420 151 7454 187
rect 7614 151 7648 187
rect 7454 117 7517 151
rect 7551 117 7614 151
rect 7420 101 7454 117
rect 7614 101 7648 117
rect 7739 296 7753 330
rect 7787 296 7801 330
rect 7739 258 7801 296
rect 7739 224 7753 258
rect 7787 224 7801 258
rect 7739 186 7801 224
rect 7739 152 7753 186
rect 7787 152 7801 186
rect 7739 114 7801 152
rect 7739 80 7753 114
rect 7787 80 7801 114
rect 7871 363 7905 379
rect 8065 363 8099 379
rect 8259 363 8293 379
rect 7905 329 7968 363
rect 8002 329 8065 363
rect 8099 329 8162 363
rect 8196 329 8259 363
rect 7871 291 7905 329
rect 7871 223 7905 257
rect 8065 291 8099 329
rect 8259 313 8293 329
rect 8373 363 8407 379
rect 8567 378 8601 723
rect 8373 291 8407 329
rect 7871 153 7905 189
rect 7871 103 7905 119
rect 7968 238 8002 254
rect 7739 62 7801 80
rect 7968 62 8002 204
rect 8065 223 8099 257
rect 8163 244 8197 260
rect 8373 244 8407 257
rect 8197 223 8407 244
rect 8197 210 8373 223
rect 8163 194 8197 210
rect 8065 153 8099 189
rect 8470 344 8601 378
rect 8701 546 8763 572
rect 8701 512 8715 546
rect 8749 512 8763 546
rect 8701 474 8763 512
rect 8701 440 8715 474
rect 8749 440 8763 474
rect 8701 402 8763 440
rect 8937 461 8971 871
rect 8937 411 8971 427
rect 9159 1003 9193 1019
rect 9159 683 9193 969
rect 9159 461 9193 649
rect 9159 411 9193 427
rect 9381 1003 9415 1019
rect 9381 535 9415 969
rect 9381 461 9415 501
rect 9381 411 9415 427
rect 9529 905 9563 1060
rect 8701 368 8715 402
rect 8749 368 8763 402
rect 8470 247 8504 344
rect 8701 330 8763 368
rect 8470 197 8504 213
rect 8567 291 8601 307
rect 8567 223 8601 257
rect 8259 153 8293 169
rect 8099 119 8162 153
rect 8196 119 8259 153
rect 8065 103 8099 119
rect 8259 103 8293 119
rect 8373 153 8407 189
rect 8567 153 8601 189
rect 8407 119 8470 153
rect 8504 119 8567 153
rect 8373 103 8407 119
rect 8567 103 8601 119
rect 8701 296 8715 330
rect 8749 296 8763 330
rect 8701 258 8763 296
rect 8701 224 8715 258
rect 8749 224 8763 258
rect 8701 186 8763 224
rect 8701 152 8715 186
rect 8749 152 8763 186
rect 8701 114 8763 152
rect 8701 80 8715 114
rect 8749 80 8763 114
rect 8833 363 8867 379
rect 9027 363 9061 379
rect 9221 363 9255 379
rect 8867 329 8930 363
rect 8964 329 9027 363
rect 9061 329 9124 363
rect 9158 329 9221 363
rect 8833 291 8867 329
rect 8833 223 8867 257
rect 9027 291 9061 329
rect 9221 313 9255 329
rect 9335 363 9369 379
rect 9529 378 9563 871
rect 9663 1076 9677 1110
rect 9711 1076 9725 1110
rect 9663 1038 9725 1076
rect 9835 1412 9869 1492
rect 9835 1344 9869 1378
rect 9835 1276 9869 1310
rect 9835 1208 9869 1242
rect 9835 1139 9869 1174
rect 9835 1073 9869 1105
rect 9923 1412 9957 1450
rect 9923 1344 9957 1378
rect 9923 1276 9957 1310
rect 9923 1208 9957 1242
rect 9923 1139 9957 1174
rect 10011 1412 10045 1492
rect 10011 1344 10045 1378
rect 10011 1276 10045 1310
rect 10011 1208 10045 1242
rect 10011 1157 10045 1174
rect 10099 1412 10133 1450
rect 10099 1344 10133 1378
rect 10099 1276 10133 1310
rect 10099 1208 10133 1242
rect 9923 1103 9957 1105
rect 10099 1139 10133 1174
rect 10187 1412 10221 1492
rect 10187 1344 10221 1378
rect 10187 1276 10221 1310
rect 10187 1208 10221 1242
rect 10187 1157 10221 1174
rect 10329 1470 10391 1492
rect 10329 1436 10343 1470
rect 10377 1436 10391 1470
rect 10329 1398 10391 1436
rect 10329 1364 10343 1398
rect 10377 1364 10391 1398
rect 10329 1326 10391 1364
rect 10329 1292 10343 1326
rect 10377 1292 10391 1326
rect 10329 1254 10391 1292
rect 10329 1220 10343 1254
rect 10377 1220 10391 1254
rect 10329 1182 10391 1220
rect 10099 1103 10133 1105
rect 10329 1148 10343 1182
rect 10377 1148 10391 1182
rect 10329 1110 10391 1148
rect 9923 1069 10229 1103
rect 9663 1004 9677 1038
rect 9711 1004 9725 1038
rect 9663 966 9725 1004
rect 9663 932 9677 966
rect 9711 932 9725 966
rect 9663 868 9725 932
rect 9899 1003 9933 1019
rect 10053 1003 10087 1019
rect 9899 905 9933 969
rect 9335 291 9369 329
rect 8833 153 8867 189
rect 8833 103 8867 119
rect 8930 238 8964 254
rect 8701 62 8763 80
rect 8930 62 8964 204
rect 9027 223 9061 257
rect 9125 244 9159 260
rect 9335 244 9369 257
rect 9159 223 9369 244
rect 9159 210 9335 223
rect 9125 194 9159 210
rect 9027 153 9061 189
rect 9432 344 9563 378
rect 9663 546 9725 572
rect 9663 512 9677 546
rect 9711 512 9725 546
rect 9663 474 9725 512
rect 9663 440 9677 474
rect 9711 440 9725 474
rect 9663 402 9725 440
rect 9899 461 9933 871
rect 9899 411 9933 427
rect 10047 969 10053 988
rect 10047 953 10087 969
rect 10047 757 10081 953
rect 10047 461 10081 723
rect 10047 411 10081 427
rect 10195 535 10229 1069
rect 10329 1076 10343 1110
rect 10377 1076 10391 1110
rect 10561 1412 10595 1492
rect 10561 1344 10595 1378
rect 10561 1276 10595 1310
rect 10561 1208 10595 1242
rect 10561 1139 10595 1174
rect 10561 1089 10595 1105
rect 10649 1412 10683 1450
rect 10649 1344 10683 1378
rect 10649 1276 10683 1310
rect 10649 1208 10683 1242
rect 10649 1139 10683 1174
rect 10737 1412 10771 1492
rect 10737 1344 10771 1378
rect 10737 1276 10771 1310
rect 10737 1208 10771 1242
rect 10737 1157 10771 1174
rect 10825 1412 10859 1450
rect 10825 1344 10859 1378
rect 10825 1276 10859 1310
rect 10825 1208 10859 1242
rect 10649 1094 10683 1105
rect 10825 1139 10859 1174
rect 10913 1412 10947 1492
rect 10913 1344 10947 1378
rect 10913 1276 10947 1310
rect 10913 1208 10947 1242
rect 10913 1157 10947 1174
rect 11001 1412 11035 1450
rect 11001 1344 11035 1378
rect 11001 1276 11035 1310
rect 11001 1208 11035 1242
rect 10825 1094 10859 1105
rect 11001 1139 11035 1174
rect 11089 1412 11123 1492
rect 11089 1344 11123 1378
rect 11089 1276 11123 1310
rect 11089 1208 11123 1242
rect 11089 1157 11123 1174
rect 11291 1470 11353 1492
rect 11291 1436 11305 1470
rect 11339 1436 11353 1470
rect 11291 1398 11353 1436
rect 11291 1364 11305 1398
rect 11339 1364 11353 1398
rect 11291 1326 11353 1364
rect 11291 1292 11305 1326
rect 11339 1292 11353 1326
rect 11291 1254 11353 1292
rect 11291 1220 11305 1254
rect 11339 1220 11353 1254
rect 11291 1182 11353 1220
rect 11001 1094 11035 1105
rect 11291 1148 11305 1182
rect 11339 1148 11353 1182
rect 11291 1110 11353 1148
rect 10329 1038 10391 1076
rect 10649 1060 11191 1094
rect 10329 1004 10343 1038
rect 10377 1004 10391 1038
rect 10329 966 10391 1004
rect 10329 932 10343 966
rect 10377 932 10391 966
rect 10329 868 10391 932
rect 10565 1003 10599 1019
rect 10565 757 10599 969
rect 9663 368 9677 402
rect 9711 368 9725 402
rect 9432 247 9466 344
rect 9663 330 9725 368
rect 9432 197 9466 213
rect 9529 291 9563 307
rect 9529 223 9563 257
rect 9221 153 9255 169
rect 9061 119 9124 153
rect 9158 119 9221 153
rect 9027 103 9061 119
rect 9221 103 9255 119
rect 9335 153 9369 189
rect 9529 153 9563 189
rect 9369 119 9432 153
rect 9466 119 9529 153
rect 9335 103 9369 119
rect 9529 103 9563 119
rect 9663 296 9677 330
rect 9711 296 9725 330
rect 9663 258 9725 296
rect 9663 224 9677 258
rect 9711 224 9725 258
rect 9663 186 9725 224
rect 9663 152 9677 186
rect 9711 152 9725 186
rect 9663 114 9725 152
rect 9663 80 9677 114
rect 9711 80 9725 114
rect 9816 361 9850 377
rect 10010 361 10044 377
rect 10195 376 10229 501
rect 9850 327 9913 361
rect 9947 327 10010 361
rect 9816 289 9850 327
rect 9816 221 9850 255
rect 10010 289 10044 327
rect 9816 151 9850 187
rect 9816 101 9850 117
rect 9913 236 9947 252
rect 9663 62 9725 80
rect 9913 62 9947 202
rect 10010 221 10044 255
rect 10107 342 10229 376
rect 10329 546 10391 572
rect 10329 512 10343 546
rect 10377 512 10391 546
rect 10329 474 10391 512
rect 10329 440 10343 474
rect 10377 440 10391 474
rect 10329 402 10391 440
rect 10565 461 10599 723
rect 10565 411 10599 427
rect 10787 1003 10821 1019
rect 10787 831 10821 969
rect 10787 461 10821 797
rect 10787 411 10821 427
rect 11009 1003 11043 1019
rect 11009 609 11043 969
rect 11009 461 11043 575
rect 11009 411 11043 427
rect 11157 905 11191 1060
rect 10329 368 10343 402
rect 10377 368 10391 402
rect 10107 245 10141 342
rect 10329 330 10391 368
rect 10107 195 10141 211
rect 10204 289 10238 305
rect 10204 221 10238 255
rect 10010 151 10044 187
rect 10204 151 10238 187
rect 10044 117 10107 151
rect 10141 117 10204 151
rect 10010 101 10044 117
rect 10204 101 10238 117
rect 10329 296 10343 330
rect 10377 296 10391 330
rect 10329 258 10391 296
rect 10329 224 10343 258
rect 10377 224 10391 258
rect 10329 186 10391 224
rect 10329 152 10343 186
rect 10377 152 10391 186
rect 10329 114 10391 152
rect 10329 80 10343 114
rect 10377 80 10391 114
rect 10461 363 10495 379
rect 10655 363 10689 379
rect 10849 363 10883 379
rect 10495 329 10558 363
rect 10592 329 10655 363
rect 10689 329 10752 363
rect 10786 329 10849 363
rect 10461 291 10495 329
rect 10461 223 10495 257
rect 10655 291 10689 329
rect 10849 313 10883 329
rect 10963 363 10997 379
rect 11157 378 11191 871
rect 11291 1076 11305 1110
rect 11339 1076 11353 1110
rect 11523 1412 11557 1492
rect 11523 1344 11557 1378
rect 11523 1276 11557 1310
rect 11523 1208 11557 1242
rect 11523 1139 11557 1174
rect 11523 1089 11557 1105
rect 11611 1412 11645 1450
rect 11611 1344 11645 1378
rect 11611 1276 11645 1310
rect 11611 1208 11645 1242
rect 11611 1139 11645 1174
rect 11699 1412 11733 1492
rect 11699 1344 11733 1378
rect 11699 1276 11733 1310
rect 11699 1208 11733 1242
rect 11699 1157 11733 1174
rect 11787 1412 11821 1450
rect 11787 1344 11821 1378
rect 11787 1276 11821 1310
rect 11787 1208 11821 1242
rect 11611 1094 11645 1105
rect 11787 1139 11821 1174
rect 11875 1412 11909 1492
rect 11875 1344 11909 1378
rect 11875 1276 11909 1310
rect 11875 1208 11909 1242
rect 11875 1157 11909 1174
rect 11963 1412 11997 1450
rect 11963 1344 11997 1378
rect 11963 1276 11997 1310
rect 11963 1208 11997 1242
rect 11787 1094 11821 1105
rect 11963 1139 11997 1174
rect 12051 1412 12085 1492
rect 12051 1344 12085 1378
rect 12051 1276 12085 1310
rect 12051 1208 12085 1242
rect 12051 1157 12085 1174
rect 12253 1470 12315 1492
rect 12253 1436 12267 1470
rect 12301 1436 12315 1470
rect 12253 1398 12315 1436
rect 12253 1364 12267 1398
rect 12301 1364 12315 1398
rect 12253 1326 12315 1364
rect 12253 1292 12267 1326
rect 12301 1292 12315 1326
rect 12253 1254 12315 1292
rect 12253 1220 12267 1254
rect 12301 1220 12315 1254
rect 12253 1182 12315 1220
rect 11963 1094 11997 1105
rect 12253 1148 12267 1182
rect 12301 1148 12315 1182
rect 12253 1110 12315 1148
rect 11291 1038 11353 1076
rect 11611 1060 12153 1094
rect 11291 1004 11305 1038
rect 11339 1004 11353 1038
rect 11291 966 11353 1004
rect 11291 932 11305 966
rect 11339 932 11353 966
rect 11291 868 11353 932
rect 11527 1003 11561 1019
rect 11527 905 11561 969
rect 10963 291 10997 329
rect 10461 153 10495 189
rect 10461 103 10495 119
rect 10558 238 10592 254
rect 10329 62 10391 80
rect 10558 62 10592 204
rect 10655 223 10689 257
rect 10753 244 10787 260
rect 10963 244 10997 257
rect 10787 223 10997 244
rect 10787 210 10963 223
rect 10753 194 10787 210
rect 10655 153 10689 189
rect 11060 344 11191 378
rect 11291 546 11353 572
rect 11291 512 11305 546
rect 11339 512 11353 546
rect 11291 474 11353 512
rect 11291 440 11305 474
rect 11339 440 11353 474
rect 11291 402 11353 440
rect 11527 461 11561 871
rect 11527 411 11561 427
rect 11749 1003 11783 1019
rect 11749 461 11783 969
rect 11749 411 11783 427
rect 11971 1003 12005 1019
rect 11971 683 12005 969
rect 11971 461 12005 649
rect 11971 411 12005 427
rect 12119 609 12153 1060
rect 12253 1076 12267 1110
rect 12301 1076 12315 1110
rect 12253 1038 12315 1076
rect 12425 1412 12459 1492
rect 12425 1344 12459 1378
rect 12425 1276 12459 1310
rect 12425 1208 12459 1242
rect 12425 1139 12459 1174
rect 12425 1073 12459 1105
rect 12513 1412 12547 1450
rect 12513 1344 12547 1378
rect 12513 1276 12547 1310
rect 12513 1208 12547 1242
rect 12513 1139 12547 1174
rect 12601 1412 12635 1492
rect 12601 1344 12635 1378
rect 12601 1276 12635 1310
rect 12601 1208 12635 1242
rect 12601 1157 12635 1174
rect 12689 1412 12723 1450
rect 12689 1344 12723 1378
rect 12689 1276 12723 1310
rect 12689 1208 12723 1242
rect 12513 1103 12547 1105
rect 12689 1139 12723 1174
rect 12777 1412 12811 1492
rect 12777 1344 12811 1378
rect 12777 1276 12811 1310
rect 12777 1208 12811 1242
rect 12777 1157 12811 1174
rect 12919 1470 12981 1492
rect 12919 1436 12933 1470
rect 12967 1436 12981 1470
rect 12919 1398 12981 1436
rect 12919 1364 12933 1398
rect 12967 1364 12981 1398
rect 12919 1326 12981 1364
rect 12919 1292 12933 1326
rect 12967 1292 12981 1326
rect 12919 1254 12981 1292
rect 12919 1220 12933 1254
rect 12967 1220 12981 1254
rect 12919 1182 12981 1220
rect 12689 1103 12723 1105
rect 12919 1148 12933 1182
rect 12967 1148 12981 1182
rect 12919 1110 12981 1148
rect 12513 1069 12819 1103
rect 12253 1004 12267 1038
rect 12301 1004 12315 1038
rect 12253 966 12315 1004
rect 12253 932 12267 966
rect 12301 932 12315 966
rect 12253 868 12315 932
rect 12489 1003 12523 1019
rect 12643 1003 12677 1019
rect 11291 368 11305 402
rect 11339 368 11353 402
rect 11060 247 11094 344
rect 11291 330 11353 368
rect 11060 197 11094 213
rect 11157 291 11191 307
rect 11157 223 11191 257
rect 10849 153 10883 169
rect 10689 119 10752 153
rect 10786 119 10849 153
rect 10655 103 10689 119
rect 10849 103 10883 119
rect 10963 153 10997 189
rect 11157 153 11191 189
rect 10997 119 11060 153
rect 11094 119 11157 153
rect 10963 103 10997 119
rect 11157 103 11191 119
rect 11291 296 11305 330
rect 11339 296 11353 330
rect 11291 258 11353 296
rect 11291 224 11305 258
rect 11339 224 11353 258
rect 11291 186 11353 224
rect 11291 152 11305 186
rect 11339 152 11353 186
rect 11291 114 11353 152
rect 11291 80 11305 114
rect 11339 80 11353 114
rect 11423 363 11457 379
rect 11617 363 11651 379
rect 11811 363 11845 379
rect 11457 329 11520 363
rect 11554 329 11617 363
rect 11651 329 11714 363
rect 11748 329 11811 363
rect 11423 291 11457 329
rect 11423 223 11457 257
rect 11617 291 11651 329
rect 11811 313 11845 329
rect 11925 363 11959 379
rect 12119 378 12153 575
rect 12489 609 12523 969
rect 11925 291 11959 329
rect 11423 153 11457 189
rect 11423 103 11457 119
rect 11520 238 11554 254
rect 11291 62 11353 80
rect 11520 62 11554 204
rect 11617 223 11651 257
rect 11715 244 11749 260
rect 11925 244 11959 257
rect 11749 223 11959 244
rect 11749 210 11925 223
rect 11715 194 11749 210
rect 11617 153 11651 189
rect 12022 344 12153 378
rect 12253 546 12315 572
rect 12253 512 12267 546
rect 12301 512 12315 546
rect 12253 474 12315 512
rect 12253 440 12267 474
rect 12301 440 12315 474
rect 12253 402 12315 440
rect 12489 461 12523 575
rect 12489 411 12523 427
rect 12637 969 12643 988
rect 12637 953 12677 969
rect 12637 757 12671 953
rect 12637 461 12671 723
rect 12637 411 12671 427
rect 12785 609 12819 1069
rect 12919 1076 12933 1110
rect 12967 1076 12981 1110
rect 13151 1412 13185 1492
rect 13151 1344 13185 1378
rect 13151 1276 13185 1310
rect 13151 1208 13185 1242
rect 13151 1139 13185 1174
rect 13151 1089 13185 1105
rect 13239 1412 13273 1450
rect 13239 1344 13273 1378
rect 13239 1276 13273 1310
rect 13239 1208 13273 1242
rect 13239 1139 13273 1174
rect 13327 1412 13361 1492
rect 13327 1344 13361 1378
rect 13327 1276 13361 1310
rect 13327 1208 13361 1242
rect 13327 1157 13361 1174
rect 13415 1412 13449 1450
rect 13415 1344 13449 1378
rect 13415 1276 13449 1310
rect 13415 1208 13449 1242
rect 13239 1094 13273 1105
rect 13415 1139 13449 1174
rect 13503 1412 13537 1492
rect 13503 1344 13537 1378
rect 13503 1276 13537 1310
rect 13503 1208 13537 1242
rect 13503 1157 13537 1174
rect 13591 1412 13625 1450
rect 13591 1344 13625 1378
rect 13591 1276 13625 1310
rect 13591 1208 13625 1242
rect 13415 1094 13449 1105
rect 13591 1139 13625 1174
rect 13679 1412 13713 1492
rect 13679 1344 13713 1378
rect 13679 1276 13713 1310
rect 13679 1208 13713 1242
rect 13679 1157 13713 1174
rect 13881 1470 13943 1492
rect 13881 1436 13895 1470
rect 13929 1436 13943 1470
rect 13881 1398 13943 1436
rect 13881 1364 13895 1398
rect 13929 1364 13943 1398
rect 13881 1326 13943 1364
rect 13881 1292 13895 1326
rect 13929 1292 13943 1326
rect 13881 1254 13943 1292
rect 13881 1220 13895 1254
rect 13929 1220 13943 1254
rect 13881 1182 13943 1220
rect 13591 1094 13625 1105
rect 13881 1148 13895 1182
rect 13929 1148 13943 1182
rect 13881 1110 13943 1148
rect 12919 1038 12981 1076
rect 13239 1060 13781 1094
rect 12919 1004 12933 1038
rect 12967 1004 12981 1038
rect 12919 966 12981 1004
rect 12919 932 12933 966
rect 12967 932 12981 966
rect 12919 868 12981 932
rect 13155 1003 13189 1019
rect 12253 368 12267 402
rect 12301 368 12315 402
rect 12022 247 12056 344
rect 12253 330 12315 368
rect 12022 197 12056 213
rect 12119 291 12153 307
rect 12119 223 12153 257
rect 11811 153 11845 169
rect 11651 119 11714 153
rect 11748 119 11811 153
rect 11617 103 11651 119
rect 11811 103 11845 119
rect 11925 153 11959 189
rect 12119 153 12153 189
rect 11959 119 12022 153
rect 12056 119 12119 153
rect 11925 103 11959 119
rect 12119 103 12153 119
rect 12253 296 12267 330
rect 12301 296 12315 330
rect 12253 258 12315 296
rect 12253 224 12267 258
rect 12301 224 12315 258
rect 12253 186 12315 224
rect 12253 152 12267 186
rect 12301 152 12315 186
rect 12253 114 12315 152
rect 12253 80 12267 114
rect 12301 80 12315 114
rect 12406 361 12440 377
rect 12600 361 12634 377
rect 12785 376 12819 575
rect 13155 609 13189 969
rect 12440 327 12503 361
rect 12537 327 12600 361
rect 12406 289 12440 327
rect 12406 221 12440 255
rect 12600 289 12634 327
rect 12406 151 12440 187
rect 12406 101 12440 117
rect 12503 236 12537 252
rect 12253 62 12315 80
rect 12503 62 12537 202
rect 12600 221 12634 255
rect 12697 342 12819 376
rect 12919 546 12981 572
rect 12919 512 12933 546
rect 12967 512 12981 546
rect 12919 474 12981 512
rect 12919 440 12933 474
rect 12967 440 12981 474
rect 12919 402 12981 440
rect 13155 461 13189 575
rect 13155 411 13189 427
rect 13377 1003 13411 1019
rect 13377 831 13411 969
rect 13377 461 13411 797
rect 13377 411 13411 427
rect 13599 1003 13633 1019
rect 13599 683 13633 969
rect 13599 461 13633 649
rect 13599 411 13633 427
rect 13747 757 13781 1060
rect 13881 1076 13895 1110
rect 13929 1076 13943 1110
rect 14113 1412 14147 1492
rect 14113 1344 14147 1378
rect 14113 1276 14147 1310
rect 14113 1208 14147 1242
rect 14113 1139 14147 1174
rect 14113 1089 14147 1105
rect 14201 1412 14235 1450
rect 14201 1344 14235 1378
rect 14201 1276 14235 1310
rect 14201 1208 14235 1242
rect 14201 1139 14235 1174
rect 14289 1412 14323 1492
rect 14289 1344 14323 1378
rect 14289 1276 14323 1310
rect 14289 1208 14323 1242
rect 14289 1157 14323 1174
rect 14377 1412 14411 1450
rect 14377 1344 14411 1378
rect 14377 1276 14411 1310
rect 14377 1208 14411 1242
rect 14201 1094 14235 1105
rect 14377 1139 14411 1174
rect 14465 1412 14499 1492
rect 14465 1344 14499 1378
rect 14465 1276 14499 1310
rect 14465 1208 14499 1242
rect 14465 1157 14499 1174
rect 14553 1412 14587 1450
rect 14553 1344 14587 1378
rect 14553 1276 14587 1310
rect 14553 1208 14587 1242
rect 14377 1094 14411 1105
rect 14553 1139 14587 1174
rect 14641 1412 14675 1492
rect 14641 1344 14675 1378
rect 14641 1276 14675 1310
rect 14641 1208 14675 1242
rect 14641 1157 14675 1174
rect 14843 1470 14905 1492
rect 14843 1436 14857 1470
rect 14891 1436 14905 1470
rect 14843 1398 14905 1436
rect 14843 1364 14857 1398
rect 14891 1364 14905 1398
rect 14843 1326 14905 1364
rect 14843 1292 14857 1326
rect 14891 1292 14905 1326
rect 14843 1254 14905 1292
rect 14843 1220 14857 1254
rect 14891 1220 14905 1254
rect 14843 1182 14905 1220
rect 14553 1094 14587 1105
rect 14843 1148 14857 1182
rect 14891 1148 14905 1182
rect 14843 1110 14905 1148
rect 13881 1038 13943 1076
rect 14201 1060 14743 1094
rect 13881 1004 13895 1038
rect 13929 1004 13943 1038
rect 13881 966 13943 1004
rect 13881 932 13895 966
rect 13929 932 13943 966
rect 13881 868 13943 932
rect 14117 1003 14151 1019
rect 14117 905 14151 969
rect 12919 368 12933 402
rect 12967 368 12981 402
rect 12697 245 12731 342
rect 12919 330 12981 368
rect 12697 195 12731 211
rect 12794 289 12828 305
rect 12794 221 12828 255
rect 12600 151 12634 187
rect 12794 151 12828 187
rect 12634 117 12697 151
rect 12731 117 12794 151
rect 12600 101 12634 117
rect 12794 101 12828 117
rect 12919 296 12933 330
rect 12967 296 12981 330
rect 12919 258 12981 296
rect 12919 224 12933 258
rect 12967 224 12981 258
rect 12919 186 12981 224
rect 12919 152 12933 186
rect 12967 152 12981 186
rect 12919 114 12981 152
rect 12919 80 12933 114
rect 12967 80 12981 114
rect 13051 363 13085 379
rect 13245 363 13279 379
rect 13439 363 13473 379
rect 13085 329 13148 363
rect 13182 329 13245 363
rect 13279 329 13342 363
rect 13376 329 13439 363
rect 13051 291 13085 329
rect 13051 223 13085 257
rect 13245 291 13279 329
rect 13439 313 13473 329
rect 13553 363 13587 379
rect 13747 378 13781 723
rect 13553 291 13587 329
rect 13051 153 13085 189
rect 13051 103 13085 119
rect 13148 238 13182 254
rect 12919 62 12981 80
rect 13148 62 13182 204
rect 13245 223 13279 257
rect 13343 244 13377 260
rect 13553 244 13587 257
rect 13377 223 13587 244
rect 13377 210 13553 223
rect 13343 194 13377 210
rect 13245 153 13279 189
rect 13650 344 13781 378
rect 13881 546 13943 572
rect 13881 512 13895 546
rect 13929 512 13943 546
rect 13881 474 13943 512
rect 13881 440 13895 474
rect 13929 440 13943 474
rect 13881 402 13943 440
rect 14117 461 14151 871
rect 14117 411 14151 427
rect 14339 1003 14373 1019
rect 14339 683 14373 969
rect 14339 461 14373 649
rect 14339 411 14373 427
rect 14561 1003 14595 1019
rect 14561 461 14595 969
rect 14561 411 14595 427
rect 14709 905 14743 1060
rect 13881 368 13895 402
rect 13929 368 13943 402
rect 13650 247 13684 344
rect 13881 330 13943 368
rect 13650 197 13684 213
rect 13747 291 13781 307
rect 13747 223 13781 257
rect 13439 153 13473 169
rect 13279 119 13342 153
rect 13376 119 13439 153
rect 13245 103 13279 119
rect 13439 103 13473 119
rect 13553 153 13587 189
rect 13747 153 13781 189
rect 13587 119 13650 153
rect 13684 119 13747 153
rect 13553 103 13587 119
rect 13747 103 13781 119
rect 13881 296 13895 330
rect 13929 296 13943 330
rect 13881 258 13943 296
rect 13881 224 13895 258
rect 13929 224 13943 258
rect 13881 186 13943 224
rect 13881 152 13895 186
rect 13929 152 13943 186
rect 13881 114 13943 152
rect 13881 80 13895 114
rect 13929 80 13943 114
rect 14013 363 14047 379
rect 14207 363 14241 379
rect 14401 363 14435 379
rect 14047 329 14110 363
rect 14144 329 14207 363
rect 14241 329 14304 363
rect 14338 329 14401 363
rect 14013 291 14047 329
rect 14013 223 14047 257
rect 14207 291 14241 329
rect 14401 313 14435 329
rect 14515 363 14549 379
rect 14709 378 14743 871
rect 14843 1076 14857 1110
rect 14891 1076 14905 1110
rect 14843 1038 14905 1076
rect 15015 1412 15049 1492
rect 15015 1344 15049 1378
rect 15015 1276 15049 1310
rect 15015 1208 15049 1242
rect 15015 1139 15049 1174
rect 15015 1073 15049 1105
rect 15103 1412 15137 1450
rect 15103 1344 15137 1378
rect 15103 1276 15137 1310
rect 15103 1208 15137 1242
rect 15103 1139 15137 1174
rect 15191 1412 15225 1492
rect 15191 1344 15225 1378
rect 15191 1276 15225 1310
rect 15191 1208 15225 1242
rect 15191 1157 15225 1174
rect 15279 1412 15313 1450
rect 15279 1344 15313 1378
rect 15279 1276 15313 1310
rect 15279 1208 15313 1242
rect 15103 1103 15137 1105
rect 15279 1139 15313 1174
rect 15367 1412 15401 1492
rect 15367 1344 15401 1378
rect 15367 1276 15401 1310
rect 15367 1208 15401 1242
rect 15367 1157 15401 1174
rect 15509 1470 15571 1492
rect 15509 1436 15523 1470
rect 15557 1436 15571 1470
rect 15509 1398 15571 1436
rect 15509 1364 15523 1398
rect 15557 1364 15571 1398
rect 15509 1326 15571 1364
rect 15509 1292 15523 1326
rect 15557 1292 15571 1326
rect 15509 1254 15571 1292
rect 15509 1220 15523 1254
rect 15557 1220 15571 1254
rect 15509 1182 15571 1220
rect 15279 1103 15313 1105
rect 15509 1148 15523 1182
rect 15557 1148 15571 1182
rect 15509 1110 15571 1148
rect 15103 1069 15409 1103
rect 14843 1004 14857 1038
rect 14891 1004 14905 1038
rect 14843 966 14905 1004
rect 14843 932 14857 966
rect 14891 932 14905 966
rect 14843 868 14905 932
rect 15079 1003 15113 1019
rect 15233 1003 15267 1019
rect 15079 905 15113 969
rect 14515 291 14549 329
rect 14013 153 14047 189
rect 14013 103 14047 119
rect 14110 238 14144 254
rect 13881 62 13943 80
rect 14110 62 14144 204
rect 14207 223 14241 257
rect 14305 244 14339 260
rect 14515 244 14549 257
rect 14339 223 14549 244
rect 14339 210 14515 223
rect 14305 194 14339 210
rect 14207 153 14241 189
rect 14612 344 14743 378
rect 14843 546 14905 572
rect 14843 512 14857 546
rect 14891 512 14905 546
rect 14843 474 14905 512
rect 14843 440 14857 474
rect 14891 440 14905 474
rect 14843 402 14905 440
rect 15079 461 15113 871
rect 15079 411 15113 427
rect 15227 969 15233 988
rect 15227 953 15267 969
rect 15227 757 15261 953
rect 15227 461 15261 723
rect 15227 411 15261 427
rect 15375 757 15409 1069
rect 15509 1076 15523 1110
rect 15557 1076 15571 1110
rect 15509 1038 15571 1076
rect 15681 1411 15715 1492
rect 15681 1343 15715 1377
rect 15681 1275 15715 1309
rect 15681 1207 15715 1241
rect 15681 1139 15715 1173
rect 15681 1071 15715 1105
rect 15769 1411 15805 1445
rect 15857 1411 15891 1492
rect 15769 1343 15803 1377
rect 15769 1275 15803 1309
rect 15769 1207 15803 1241
rect 15769 1139 15803 1173
rect 15857 1343 15891 1377
rect 15857 1275 15891 1309
rect 15857 1207 15891 1241
rect 15857 1157 15891 1173
rect 15945 1411 15979 1445
rect 15945 1343 15979 1377
rect 15945 1275 15979 1309
rect 15945 1207 15979 1241
rect 15945 1105 15979 1173
rect 15769 1071 15945 1105
rect 16033 1411 16067 1492
rect 16033 1343 16067 1377
rect 16033 1275 16067 1309
rect 16033 1207 16067 1241
rect 16033 1139 16067 1173
rect 16033 1071 16067 1105
rect 16175 1470 16237 1492
rect 16175 1436 16189 1470
rect 16223 1436 16237 1470
rect 16841 1470 16903 1492
rect 16175 1398 16237 1436
rect 16175 1364 16189 1398
rect 16223 1364 16237 1398
rect 16175 1326 16237 1364
rect 16175 1292 16189 1326
rect 16223 1292 16237 1326
rect 16175 1254 16237 1292
rect 16175 1220 16189 1254
rect 16223 1220 16237 1254
rect 16175 1182 16237 1220
rect 16175 1148 16189 1182
rect 16223 1148 16237 1182
rect 16175 1110 16237 1148
rect 16175 1076 16189 1110
rect 16223 1076 16237 1110
rect 15945 1055 15979 1071
rect 15509 1004 15523 1038
rect 15557 1004 15571 1038
rect 16175 1038 16237 1076
rect 16345 1411 16731 1445
rect 16345 1343 16379 1377
rect 16345 1275 16379 1309
rect 16345 1207 16379 1241
rect 16345 1105 16379 1173
rect 16433 1343 16467 1359
rect 16433 1275 16467 1309
rect 16433 1207 16467 1241
rect 16433 1139 16467 1173
rect 16521 1343 16555 1377
rect 16521 1275 16555 1309
rect 16521 1207 16555 1241
rect 16521 1157 16555 1173
rect 16609 1343 16643 1359
rect 16609 1275 16643 1309
rect 16609 1207 16643 1241
rect 16609 1105 16643 1173
rect 16697 1343 16731 1377
rect 16697 1275 16731 1309
rect 16697 1207 16731 1241
rect 16697 1121 16731 1173
rect 16841 1436 16855 1470
rect 16889 1436 16903 1470
rect 17507 1470 17569 1492
rect 16841 1398 16903 1436
rect 16841 1364 16855 1398
rect 16889 1364 16903 1398
rect 16841 1326 16903 1364
rect 16841 1292 16855 1326
rect 16889 1292 16903 1326
rect 16841 1254 16903 1292
rect 16841 1220 16855 1254
rect 16889 1220 16903 1254
rect 16841 1182 16903 1220
rect 16841 1148 16855 1182
rect 16889 1148 16903 1182
rect 16433 1071 16609 1105
rect 16345 1055 16379 1071
rect 16609 1055 16643 1071
rect 16841 1110 16903 1148
rect 16841 1076 16855 1110
rect 16889 1076 16903 1110
rect 15509 966 15571 1004
rect 15509 932 15523 966
rect 15557 932 15571 966
rect 15509 868 15571 932
rect 15671 1004 15705 1020
rect 15901 1004 15935 1020
rect 15671 905 15705 970
rect 14843 368 14857 402
rect 14891 368 14905 402
rect 14612 247 14646 344
rect 14843 330 14905 368
rect 14612 197 14646 213
rect 14709 291 14743 307
rect 14709 223 14743 257
rect 14401 153 14435 169
rect 14241 119 14304 153
rect 14338 119 14401 153
rect 14207 103 14241 119
rect 14401 103 14435 119
rect 14515 153 14549 189
rect 14709 153 14743 189
rect 14549 119 14612 153
rect 14646 119 14709 153
rect 14515 103 14549 119
rect 14709 103 14743 119
rect 14843 296 14857 330
rect 14891 296 14905 330
rect 14843 258 14905 296
rect 14843 224 14857 258
rect 14891 224 14905 258
rect 14843 186 14905 224
rect 14843 152 14857 186
rect 14891 152 14905 186
rect 14843 114 14905 152
rect 14843 80 14857 114
rect 14891 80 14905 114
rect 14996 361 15030 377
rect 15190 361 15224 377
rect 15375 376 15409 723
rect 15030 327 15093 361
rect 15127 327 15190 361
rect 14996 289 15030 327
rect 14996 221 15030 255
rect 15190 289 15224 327
rect 14996 151 15030 187
rect 14996 101 15030 117
rect 15093 236 15127 252
rect 14843 62 14905 80
rect 15093 62 15127 202
rect 15190 221 15224 255
rect 15287 342 15409 376
rect 15509 546 15571 572
rect 15509 512 15523 546
rect 15557 512 15571 546
rect 15509 474 15571 512
rect 15509 440 15523 474
rect 15557 440 15571 474
rect 15509 402 15571 440
rect 15671 535 15705 871
rect 15671 461 15705 501
rect 15671 411 15705 427
rect 15893 979 15901 995
rect 15927 954 15935 970
rect 16175 1004 16189 1038
rect 16223 1004 16237 1038
rect 16841 1038 16903 1076
rect 17013 1411 17399 1445
rect 17013 1343 17047 1377
rect 17013 1275 17047 1309
rect 17013 1207 17047 1241
rect 17013 1105 17047 1173
rect 17101 1343 17135 1359
rect 17101 1275 17135 1309
rect 17101 1207 17135 1241
rect 17101 1139 17135 1173
rect 17189 1343 17223 1377
rect 17189 1275 17223 1309
rect 17189 1207 17223 1241
rect 17189 1157 17223 1173
rect 17277 1343 17311 1359
rect 17277 1275 17311 1309
rect 17277 1207 17311 1241
rect 17277 1139 17311 1173
rect 17365 1343 17399 1377
rect 17365 1275 17399 1309
rect 17365 1207 17399 1241
rect 17365 1157 17399 1173
rect 17507 1436 17521 1470
rect 17555 1436 17569 1470
rect 17507 1398 17569 1436
rect 17507 1364 17521 1398
rect 17555 1364 17569 1398
rect 17507 1326 17569 1364
rect 17507 1292 17521 1326
rect 17555 1292 17569 1326
rect 17507 1254 17569 1292
rect 17507 1220 17521 1254
rect 17555 1220 17569 1254
rect 17507 1182 17569 1220
rect 17507 1148 17521 1182
rect 17555 1148 17569 1182
rect 17507 1110 17569 1148
rect 17101 1071 17407 1105
rect 17013 1055 17047 1071
rect 16175 966 16237 1004
rect 15893 831 15927 945
rect 16175 932 16189 966
rect 16223 932 16237 966
rect 16175 868 16237 932
rect 16411 1004 16445 1020
rect 16411 905 16445 970
rect 16411 847 16445 871
rect 16707 1004 16741 1020
rect 16707 905 16741 970
rect 15893 461 15927 797
rect 16707 757 16741 871
rect 16841 1004 16855 1038
rect 16889 1004 16903 1038
rect 16841 966 16903 1004
rect 16841 932 16855 966
rect 16889 932 16903 966
rect 16841 868 16903 932
rect 17003 1004 17037 1020
rect 17003 905 17037 970
rect 17003 847 17037 871
rect 17225 1004 17263 1020
rect 17225 970 17229 1004
rect 17225 954 17263 970
rect 15893 411 15927 427
rect 16175 546 16237 572
rect 16175 512 16189 546
rect 16223 512 16237 546
rect 16175 474 16237 512
rect 16175 440 16189 474
rect 16223 440 16237 474
rect 15509 368 15523 402
rect 15557 368 15571 402
rect 16175 402 16237 440
rect 16411 535 16445 551
rect 16411 461 16445 501
rect 16411 411 16445 427
rect 16707 535 16741 723
rect 17225 831 17259 954
rect 16707 461 16741 501
rect 16707 411 16741 427
rect 16841 546 16903 572
rect 16841 512 16855 546
rect 16889 512 16903 546
rect 16841 474 16903 512
rect 16841 440 16855 474
rect 16889 440 16903 474
rect 15287 245 15321 342
rect 15509 330 15571 368
rect 15287 195 15321 211
rect 15384 289 15418 305
rect 15384 221 15418 255
rect 15190 151 15224 187
rect 15384 151 15418 187
rect 15224 117 15287 151
rect 15321 117 15384 151
rect 15190 101 15224 117
rect 15384 101 15418 117
rect 15509 296 15523 330
rect 15557 296 15571 330
rect 15509 258 15571 296
rect 15509 224 15523 258
rect 15557 224 15571 258
rect 15509 186 15571 224
rect 15509 152 15523 186
rect 15557 152 15571 186
rect 15509 114 15571 152
rect 15509 80 15523 114
rect 15557 80 15571 114
rect 15662 361 15696 377
rect 15856 361 15890 377
rect 15696 327 15759 361
rect 15793 327 15856 361
rect 15662 289 15696 327
rect 15662 221 15696 255
rect 15856 289 15890 327
rect 16050 361 16084 377
rect 15953 281 15987 297
rect 15662 151 15696 187
rect 15662 101 15696 117
rect 15759 236 15793 252
rect 15509 62 15571 80
rect 15759 62 15793 202
rect 15856 221 15890 255
rect 15952 247 15953 262
rect 15952 245 15987 247
rect 15986 231 15987 245
rect 16050 289 16084 327
rect 15952 195 15986 211
rect 16050 221 16084 255
rect 15856 151 15890 187
rect 16050 151 16084 187
rect 15890 117 15952 151
rect 15986 117 16050 151
rect 15856 101 15890 117
rect 16050 101 16084 117
rect 16175 368 16189 402
rect 16223 368 16237 402
rect 16841 402 16903 440
rect 17003 535 17037 551
rect 17003 461 17037 501
rect 17003 411 17037 427
rect 17225 461 17259 797
rect 17225 411 17259 427
rect 17373 831 17407 1071
rect 17507 1076 17521 1110
rect 17555 1076 17569 1110
rect 17655 1412 17689 1492
rect 17655 1344 17689 1378
rect 17655 1276 17689 1310
rect 17655 1208 17689 1242
rect 17655 1139 17689 1174
rect 17655 1083 17689 1105
rect 17743 1412 17777 1450
rect 17743 1344 17777 1378
rect 17743 1276 17777 1310
rect 17743 1208 17777 1242
rect 17743 1139 17777 1174
rect 17507 1038 17569 1076
rect 17507 1004 17521 1038
rect 17555 1004 17569 1038
rect 17507 966 17569 1004
rect 17507 932 17521 966
rect 17555 932 17569 966
rect 17507 868 17569 932
rect 17669 1003 17703 1019
rect 16175 330 16237 368
rect 16175 296 16189 330
rect 16223 296 16237 330
rect 16175 258 16237 296
rect 16175 224 16189 258
rect 16223 224 16237 258
rect 16175 186 16237 224
rect 16175 152 16189 186
rect 16223 152 16237 186
rect 16175 114 16237 152
rect 16175 80 16189 114
rect 16223 80 16237 114
rect 16328 361 16362 377
rect 16522 361 16556 377
rect 16362 327 16425 361
rect 16459 327 16522 361
rect 16328 289 16362 327
rect 16328 221 16362 255
rect 16522 289 16556 327
rect 16716 361 16750 377
rect 16328 151 16362 187
rect 16328 101 16362 117
rect 16425 236 16459 252
rect 16175 62 16237 80
rect 16425 62 16459 202
rect 16522 221 16556 255
rect 16619 281 16653 297
rect 16619 245 16653 247
rect 16619 195 16653 211
rect 16716 289 16750 327
rect 16716 221 16750 255
rect 16522 151 16556 187
rect 16716 151 16750 187
rect 16556 117 16619 151
rect 16653 117 16716 151
rect 16522 101 16556 117
rect 16716 101 16750 117
rect 16841 368 16855 402
rect 16889 368 16903 402
rect 16841 330 16903 368
rect 16841 296 16855 330
rect 16889 296 16903 330
rect 16841 258 16903 296
rect 16841 224 16855 258
rect 16889 224 16903 258
rect 16841 186 16903 224
rect 16841 152 16855 186
rect 16889 152 16903 186
rect 16841 114 16903 152
rect 16841 80 16855 114
rect 16889 80 16903 114
rect 16994 361 17028 377
rect 17188 361 17222 377
rect 17373 374 17407 797
rect 17669 831 17703 969
rect 17743 979 17777 1105
rect 17831 1412 17865 1492
rect 17831 1344 17865 1378
rect 17831 1276 17865 1310
rect 17831 1208 17865 1242
rect 17831 1139 17865 1174
rect 17831 1083 17865 1105
rect 17951 1470 18013 1492
rect 17951 1436 17965 1470
rect 17999 1436 18013 1470
rect 17951 1398 18013 1436
rect 17951 1364 17965 1398
rect 17999 1364 18013 1398
rect 17951 1326 18013 1364
rect 17951 1292 17965 1326
rect 17999 1292 18013 1326
rect 17951 1254 18013 1292
rect 17951 1220 17965 1254
rect 17999 1220 18013 1254
rect 17951 1182 18013 1220
rect 17951 1148 17965 1182
rect 17999 1148 18013 1182
rect 17951 1110 18013 1148
rect 17951 1076 17965 1110
rect 17999 1076 18013 1110
rect 17951 1038 18013 1076
rect 17951 1004 17965 1038
rect 17999 1004 18013 1038
rect 17743 945 17851 979
rect 17028 327 17091 361
rect 17125 327 17188 361
rect 16994 289 17028 327
rect 16994 221 17028 255
rect 17188 289 17222 327
rect 16994 151 17028 187
rect 16994 101 17028 117
rect 17091 236 17125 252
rect 16841 62 16903 80
rect 17091 62 17125 202
rect 17188 221 17222 255
rect 17285 340 17407 374
rect 17507 546 17569 572
rect 17507 512 17521 546
rect 17555 512 17569 546
rect 17507 474 17569 512
rect 17507 440 17521 474
rect 17555 440 17569 474
rect 17507 402 17569 440
rect 17669 461 17703 797
rect 17817 831 17851 945
rect 17951 966 18013 1004
rect 17951 932 17965 966
rect 17999 932 18013 966
rect 17951 868 18013 932
rect 17817 461 17851 797
rect 17669 411 17703 427
rect 17743 427 17851 461
rect 17951 546 18013 572
rect 17951 512 17965 546
rect 17999 512 18013 546
rect 17951 474 18013 512
rect 17951 440 17965 474
rect 17999 440 18013 474
rect 17507 368 17521 402
rect 17555 368 17569 402
rect 17285 281 17319 340
rect 17507 330 17569 368
rect 17285 245 17319 247
rect 17285 195 17319 211
rect 17382 289 17416 306
rect 17382 221 17416 255
rect 17188 151 17222 187
rect 17382 151 17416 187
rect 17222 117 17285 151
rect 17319 117 17382 151
rect 17188 101 17222 117
rect 17382 101 17416 117
rect 17507 296 17521 330
rect 17555 296 17569 330
rect 17507 258 17569 296
rect 17507 224 17521 258
rect 17555 224 17569 258
rect 17507 186 17569 224
rect 17507 152 17521 186
rect 17555 152 17569 186
rect 17507 114 17569 152
rect 17507 80 17521 114
rect 17555 80 17569 114
rect 17507 62 17569 80
rect 17647 361 17681 377
rect 17647 289 17681 327
rect 17647 221 17681 255
rect 17743 245 17777 427
rect 17951 402 18013 440
rect 17743 195 17777 211
rect 17841 361 17875 377
rect 17841 289 17875 327
rect 17841 221 17875 255
rect 17647 151 17681 187
rect 17841 151 17875 187
rect 17681 117 17743 151
rect 17777 117 17841 151
rect 17647 62 17681 117
rect 17744 62 17778 117
rect 17841 62 17875 117
rect 17951 368 17965 402
rect 17999 368 18013 402
rect 17951 330 18013 368
rect 17951 296 17965 330
rect 17999 296 18013 330
rect 17951 258 18013 296
rect 17951 224 17965 258
rect 17999 224 18013 258
rect 17951 186 18013 224
rect 17951 152 17965 186
rect 17999 152 18013 186
rect 17951 114 18013 152
rect 17951 80 17965 114
rect 17999 80 18013 114
rect 17951 62 18013 80
rect -31 47 16619 62
rect 16653 47 18013 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 343 47
rect 377 13 415 47
rect 449 13 513 47
rect 547 13 585 47
rect 619 13 657 47
rect 691 13 729 47
rect 763 13 801 47
rect 835 13 873 47
rect 907 13 1017 47
rect 1051 13 1089 47
rect 1123 13 1161 47
rect 1195 13 1233 47
rect 1267 13 1305 47
rect 1339 13 1377 47
rect 1411 13 1475 47
rect 1509 13 1547 47
rect 1581 13 1619 47
rect 1653 13 1691 47
rect 1725 13 1763 47
rect 1797 13 1835 47
rect 1869 13 1979 47
rect 2013 13 2051 47
rect 2085 13 2123 47
rect 2157 13 2195 47
rect 2229 13 2285 47
rect 2319 13 2357 47
rect 2391 13 2429 47
rect 2463 13 2501 47
rect 2535 13 2645 47
rect 2679 13 2717 47
rect 2751 13 2789 47
rect 2823 13 2861 47
rect 2895 13 2933 47
rect 2967 13 3005 47
rect 3039 13 3103 47
rect 3137 13 3175 47
rect 3209 13 3247 47
rect 3281 13 3319 47
rect 3353 13 3391 47
rect 3425 13 3463 47
rect 3497 13 3607 47
rect 3641 13 3679 47
rect 3713 13 3751 47
rect 3785 13 3823 47
rect 3857 13 3895 47
rect 3929 13 3967 47
rect 4001 13 4065 47
rect 4099 13 4137 47
rect 4171 13 4209 47
rect 4243 13 4281 47
rect 4315 13 4353 47
rect 4387 13 4425 47
rect 4459 13 4569 47
rect 4603 13 4641 47
rect 4675 13 4713 47
rect 4747 13 4785 47
rect 4819 13 4875 47
rect 4909 13 4947 47
rect 4981 13 5019 47
rect 5053 13 5091 47
rect 5125 13 5235 47
rect 5269 13 5307 47
rect 5341 13 5379 47
rect 5413 13 5451 47
rect 5485 13 5523 47
rect 5557 13 5595 47
rect 5629 13 5693 47
rect 5727 13 5765 47
rect 5799 13 5837 47
rect 5871 13 5909 47
rect 5943 13 5981 47
rect 6015 13 6053 47
rect 6087 13 6197 47
rect 6231 13 6269 47
rect 6303 13 6341 47
rect 6375 13 6413 47
rect 6447 13 6485 47
rect 6519 13 6557 47
rect 6591 13 6655 47
rect 6689 13 6727 47
rect 6761 13 6799 47
rect 6833 13 6871 47
rect 6905 13 6943 47
rect 6977 13 7015 47
rect 7049 13 7159 47
rect 7193 13 7231 47
rect 7265 13 7303 47
rect 7337 13 7375 47
rect 7409 13 7465 47
rect 7499 13 7537 47
rect 7571 13 7609 47
rect 7643 13 7681 47
rect 7715 13 7825 47
rect 7859 13 7897 47
rect 7931 13 7969 47
rect 8003 13 8041 47
rect 8075 13 8113 47
rect 8147 13 8185 47
rect 8219 13 8283 47
rect 8317 13 8355 47
rect 8389 13 8427 47
rect 8461 13 8499 47
rect 8533 13 8571 47
rect 8605 13 8643 47
rect 8677 13 8787 47
rect 8821 13 8859 47
rect 8893 13 8931 47
rect 8965 13 9003 47
rect 9037 13 9075 47
rect 9109 13 9147 47
rect 9181 13 9245 47
rect 9279 13 9317 47
rect 9351 13 9389 47
rect 9423 13 9461 47
rect 9495 13 9533 47
rect 9567 13 9605 47
rect 9639 13 9749 47
rect 9783 13 9821 47
rect 9855 13 9893 47
rect 9927 13 9965 47
rect 9999 13 10055 47
rect 10089 13 10127 47
rect 10161 13 10199 47
rect 10233 13 10271 47
rect 10305 13 10415 47
rect 10449 13 10487 47
rect 10521 13 10559 47
rect 10593 13 10631 47
rect 10665 13 10703 47
rect 10737 13 10775 47
rect 10809 13 10873 47
rect 10907 13 10945 47
rect 10979 13 11017 47
rect 11051 13 11089 47
rect 11123 13 11161 47
rect 11195 13 11233 47
rect 11267 13 11377 47
rect 11411 13 11449 47
rect 11483 13 11521 47
rect 11555 13 11593 47
rect 11627 13 11665 47
rect 11699 13 11737 47
rect 11771 13 11835 47
rect 11869 13 11907 47
rect 11941 13 11979 47
rect 12013 13 12051 47
rect 12085 13 12123 47
rect 12157 13 12195 47
rect 12229 13 12339 47
rect 12373 13 12411 47
rect 12445 13 12483 47
rect 12517 13 12555 47
rect 12589 13 12645 47
rect 12679 13 12717 47
rect 12751 13 12789 47
rect 12823 13 12861 47
rect 12895 13 13005 47
rect 13039 13 13077 47
rect 13111 13 13149 47
rect 13183 13 13221 47
rect 13255 13 13293 47
rect 13327 13 13365 47
rect 13399 13 13463 47
rect 13497 13 13535 47
rect 13569 13 13607 47
rect 13641 13 13679 47
rect 13713 13 13751 47
rect 13785 13 13823 47
rect 13857 13 13967 47
rect 14001 13 14039 47
rect 14073 13 14111 47
rect 14145 13 14183 47
rect 14217 13 14255 47
rect 14289 13 14327 47
rect 14361 13 14425 47
rect 14459 13 14497 47
rect 14531 13 14569 47
rect 14603 13 14641 47
rect 14675 13 14713 47
rect 14747 13 14785 47
rect 14819 13 14929 47
rect 14963 13 15001 47
rect 15035 13 15073 47
rect 15107 13 15145 47
rect 15179 13 15235 47
rect 15269 13 15307 47
rect 15341 13 15379 47
rect 15413 13 15451 47
rect 15485 13 15595 47
rect 15629 13 15667 47
rect 15701 13 15739 47
rect 15773 13 15811 47
rect 15845 13 15901 47
rect 15935 13 15973 47
rect 16007 13 16045 47
rect 16079 13 16117 47
rect 16151 13 16261 47
rect 16295 13 16333 47
rect 16367 13 16405 47
rect 16439 13 16477 47
rect 16511 13 16567 47
rect 16601 13 16639 47
rect 16673 13 16711 47
rect 16745 13 16783 47
rect 16817 13 16927 47
rect 16961 13 16999 47
rect 17033 13 17071 47
rect 17105 13 17143 47
rect 17177 13 17233 47
rect 17267 13 17305 47
rect 17339 13 17377 47
rect 17411 13 17449 47
rect 17483 13 17593 47
rect 17627 13 17665 47
rect 17699 13 17743 47
rect 17777 13 17821 47
rect 17855 13 17893 47
rect 17927 13 18013 47
rect -31 0 18013 13
<< viali >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 343 1505 377 1539
rect 415 1505 449 1539
rect 513 1505 547 1539
rect 585 1505 619 1539
rect 657 1505 691 1539
rect 729 1505 763 1539
rect 801 1505 835 1539
rect 873 1505 907 1539
rect 1017 1505 1051 1539
rect 1089 1505 1123 1539
rect 1161 1505 1195 1539
rect 1233 1505 1267 1539
rect 1305 1505 1339 1539
rect 1377 1505 1411 1539
rect 1475 1505 1509 1539
rect 1547 1505 1581 1539
rect 1619 1505 1653 1539
rect 1691 1505 1725 1539
rect 1763 1505 1797 1539
rect 1835 1505 1869 1539
rect 1979 1505 2013 1539
rect 2051 1505 2085 1539
rect 2123 1505 2157 1539
rect 2195 1505 2229 1539
rect 2285 1505 2319 1539
rect 2357 1505 2391 1539
rect 2429 1505 2463 1539
rect 2501 1505 2535 1539
rect 2645 1505 2679 1539
rect 2717 1505 2751 1539
rect 2789 1505 2823 1539
rect 2861 1505 2895 1539
rect 2933 1505 2967 1539
rect 3005 1505 3039 1539
rect 3103 1505 3137 1539
rect 3175 1505 3209 1539
rect 3247 1505 3281 1539
rect 3319 1505 3353 1539
rect 3391 1505 3425 1539
rect 3463 1505 3497 1539
rect 3607 1505 3641 1539
rect 3679 1505 3713 1539
rect 3751 1505 3785 1539
rect 3823 1505 3857 1539
rect 3895 1505 3929 1539
rect 3967 1505 4001 1539
rect 4065 1505 4099 1539
rect 4137 1505 4171 1539
rect 4209 1505 4243 1539
rect 4281 1505 4315 1539
rect 4353 1505 4387 1539
rect 4425 1505 4459 1539
rect 4569 1505 4603 1539
rect 4641 1505 4675 1539
rect 4713 1505 4747 1539
rect 4785 1505 4819 1539
rect 4875 1505 4909 1539
rect 4947 1505 4981 1539
rect 5019 1505 5053 1539
rect 5091 1505 5125 1539
rect 5235 1505 5269 1539
rect 5307 1505 5341 1539
rect 5379 1505 5413 1539
rect 5451 1505 5485 1539
rect 5523 1505 5557 1539
rect 5595 1505 5629 1539
rect 5693 1505 5727 1539
rect 5765 1505 5799 1539
rect 5837 1505 5871 1539
rect 5909 1505 5943 1539
rect 5981 1505 6015 1539
rect 6053 1505 6087 1539
rect 6197 1505 6231 1539
rect 6269 1505 6303 1539
rect 6341 1505 6375 1539
rect 6413 1505 6447 1539
rect 6485 1505 6519 1539
rect 6557 1505 6591 1539
rect 6655 1505 6689 1539
rect 6727 1505 6761 1539
rect 6799 1505 6833 1539
rect 6871 1505 6905 1539
rect 6943 1505 6977 1539
rect 7015 1505 7049 1539
rect 7159 1505 7193 1539
rect 7231 1505 7265 1539
rect 7303 1505 7337 1539
rect 7375 1505 7409 1539
rect 7465 1505 7499 1539
rect 7537 1505 7571 1539
rect 7609 1505 7643 1539
rect 7681 1505 7715 1539
rect 7825 1505 7859 1539
rect 7897 1505 7931 1539
rect 7969 1505 8003 1539
rect 8041 1505 8075 1539
rect 8113 1505 8147 1539
rect 8185 1505 8219 1539
rect 8283 1505 8317 1539
rect 8355 1505 8389 1539
rect 8427 1505 8461 1539
rect 8499 1505 8533 1539
rect 8571 1505 8605 1539
rect 8643 1505 8677 1539
rect 8787 1505 8821 1539
rect 8859 1505 8893 1539
rect 8931 1505 8965 1539
rect 9003 1505 9037 1539
rect 9075 1505 9109 1539
rect 9147 1505 9181 1539
rect 9245 1505 9279 1539
rect 9317 1505 9351 1539
rect 9389 1505 9423 1539
rect 9461 1505 9495 1539
rect 9533 1505 9567 1539
rect 9605 1505 9639 1539
rect 9749 1505 9783 1539
rect 9821 1505 9855 1539
rect 9893 1505 9927 1539
rect 9965 1505 9999 1539
rect 10055 1505 10089 1539
rect 10127 1505 10161 1539
rect 10199 1505 10233 1539
rect 10271 1505 10305 1539
rect 10415 1505 10449 1539
rect 10487 1505 10521 1539
rect 10559 1505 10593 1539
rect 10631 1505 10665 1539
rect 10703 1505 10737 1539
rect 10775 1505 10809 1539
rect 10873 1505 10907 1539
rect 10945 1505 10979 1539
rect 11017 1505 11051 1539
rect 11089 1505 11123 1539
rect 11161 1505 11195 1539
rect 11233 1505 11267 1539
rect 11377 1505 11411 1539
rect 11449 1505 11483 1539
rect 11521 1505 11555 1539
rect 11593 1505 11627 1539
rect 11665 1505 11699 1539
rect 11737 1505 11771 1539
rect 11835 1505 11869 1539
rect 11907 1505 11941 1539
rect 11979 1505 12013 1539
rect 12051 1505 12085 1539
rect 12123 1505 12157 1539
rect 12195 1505 12229 1539
rect 12339 1505 12373 1539
rect 12411 1505 12445 1539
rect 12483 1505 12517 1539
rect 12555 1505 12589 1539
rect 12645 1505 12679 1539
rect 12717 1505 12751 1539
rect 12789 1505 12823 1539
rect 12861 1505 12895 1539
rect 13005 1505 13039 1539
rect 13077 1505 13111 1539
rect 13149 1505 13183 1539
rect 13221 1505 13255 1539
rect 13293 1505 13327 1539
rect 13365 1505 13399 1539
rect 13463 1505 13497 1539
rect 13535 1505 13569 1539
rect 13607 1505 13641 1539
rect 13679 1505 13713 1539
rect 13751 1505 13785 1539
rect 13823 1505 13857 1539
rect 13967 1505 14001 1539
rect 14039 1505 14073 1539
rect 14111 1505 14145 1539
rect 14183 1505 14217 1539
rect 14255 1505 14289 1539
rect 14327 1505 14361 1539
rect 14425 1505 14459 1539
rect 14497 1505 14531 1539
rect 14569 1505 14603 1539
rect 14641 1505 14675 1539
rect 14713 1505 14747 1539
rect 14785 1505 14819 1539
rect 14929 1505 14963 1539
rect 15001 1505 15035 1539
rect 15073 1505 15107 1539
rect 15145 1505 15179 1539
rect 15235 1505 15269 1539
rect 15307 1505 15341 1539
rect 15379 1505 15413 1539
rect 15451 1505 15485 1539
rect 15595 1505 15629 1539
rect 15667 1505 15701 1539
rect 15739 1505 15773 1539
rect 15811 1505 15845 1539
rect 15901 1505 15935 1539
rect 15973 1505 16007 1539
rect 16045 1505 16079 1539
rect 16117 1505 16151 1539
rect 16261 1505 16295 1539
rect 16333 1505 16367 1539
rect 16405 1505 16439 1539
rect 16477 1505 16511 1539
rect 16567 1505 16601 1539
rect 16639 1505 16673 1539
rect 16711 1505 16745 1539
rect 16783 1505 16817 1539
rect 16927 1505 16961 1539
rect 16999 1505 17033 1539
rect 17071 1505 17105 1539
rect 17143 1505 17177 1539
rect 17233 1505 17267 1539
rect 17305 1505 17339 1539
rect 17377 1505 17411 1539
rect 17449 1505 17483 1539
rect 17593 1505 17627 1539
rect 17665 1505 17699 1539
rect 17743 1505 17777 1539
rect 17821 1505 17855 1539
rect 17893 1505 17927 1539
rect 205 723 239 757
rect 427 797 461 831
rect 649 575 683 609
rect 797 871 831 905
rect 1167 871 1201 905
rect 1389 427 1423 461
rect 1611 649 1645 683
rect 1759 575 1793 609
rect 2129 575 2163 609
rect 2277 723 2311 757
rect 2425 575 2459 609
rect 2795 575 2829 609
rect 3017 797 3051 831
rect 3239 649 3273 683
rect 3757 871 3791 905
rect 3387 723 3421 757
rect 3979 649 4013 683
rect 4201 969 4235 979
rect 4201 945 4235 969
rect 4349 871 4383 905
rect 4719 871 4753 905
rect 4867 723 4901 757
rect 5015 945 5049 979
rect 5385 723 5419 757
rect 5607 797 5641 831
rect 5829 575 5863 609
rect 5977 871 6011 905
rect 6347 871 6381 905
rect 6569 427 6603 461
rect 6791 649 6825 683
rect 6939 575 6973 609
rect 7309 575 7343 609
rect 7457 723 7491 757
rect 7605 575 7639 609
rect 7975 575 8009 609
rect 8197 797 8231 831
rect 8419 649 8453 683
rect 8937 871 8971 905
rect 8567 723 8601 757
rect 9159 649 9193 683
rect 9381 501 9415 535
rect 9529 871 9563 905
rect 9899 871 9933 905
rect 10047 723 10081 757
rect 10565 723 10599 757
rect 10195 501 10229 535
rect 10787 797 10821 831
rect 11009 575 11043 609
rect 11157 871 11191 905
rect 11527 871 11561 905
rect 11749 427 11783 461
rect 11971 649 12005 683
rect 12119 575 12153 609
rect 12489 575 12523 609
rect 12637 723 12671 757
rect 12785 575 12819 609
rect 13155 575 13189 609
rect 13377 797 13411 831
rect 13599 649 13633 683
rect 14117 871 14151 905
rect 13747 723 13781 757
rect 14339 649 14373 683
rect 14709 871 14743 905
rect 15079 871 15113 905
rect 15227 723 15261 757
rect 15945 1071 15979 1105
rect 16345 1071 16379 1105
rect 16609 1071 16643 1105
rect 15671 871 15705 905
rect 15375 723 15409 757
rect 15671 501 15705 535
rect 15893 970 15901 979
rect 15901 970 15927 979
rect 15893 945 15927 970
rect 17013 1071 17047 1105
rect 16411 871 16445 905
rect 16707 871 16741 905
rect 15893 797 15927 831
rect 17003 871 17037 905
rect 16707 723 16741 757
rect 16411 501 16445 535
rect 17225 797 17259 831
rect 16707 501 16741 535
rect 15953 247 15987 281
rect 17003 501 17037 535
rect 17373 797 17407 831
rect 16619 247 16653 281
rect 17669 797 17703 831
rect 17817 797 17851 831
rect 17285 247 17319 281
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 343 13 377 47
rect 415 13 449 47
rect 513 13 547 47
rect 585 13 619 47
rect 657 13 691 47
rect 729 13 763 47
rect 801 13 835 47
rect 873 13 907 47
rect 1017 13 1051 47
rect 1089 13 1123 47
rect 1161 13 1195 47
rect 1233 13 1267 47
rect 1305 13 1339 47
rect 1377 13 1411 47
rect 1475 13 1509 47
rect 1547 13 1581 47
rect 1619 13 1653 47
rect 1691 13 1725 47
rect 1763 13 1797 47
rect 1835 13 1869 47
rect 1979 13 2013 47
rect 2051 13 2085 47
rect 2123 13 2157 47
rect 2195 13 2229 47
rect 2285 13 2319 47
rect 2357 13 2391 47
rect 2429 13 2463 47
rect 2501 13 2535 47
rect 2645 13 2679 47
rect 2717 13 2751 47
rect 2789 13 2823 47
rect 2861 13 2895 47
rect 2933 13 2967 47
rect 3005 13 3039 47
rect 3103 13 3137 47
rect 3175 13 3209 47
rect 3247 13 3281 47
rect 3319 13 3353 47
rect 3391 13 3425 47
rect 3463 13 3497 47
rect 3607 13 3641 47
rect 3679 13 3713 47
rect 3751 13 3785 47
rect 3823 13 3857 47
rect 3895 13 3929 47
rect 3967 13 4001 47
rect 4065 13 4099 47
rect 4137 13 4171 47
rect 4209 13 4243 47
rect 4281 13 4315 47
rect 4353 13 4387 47
rect 4425 13 4459 47
rect 4569 13 4603 47
rect 4641 13 4675 47
rect 4713 13 4747 47
rect 4785 13 4819 47
rect 4875 13 4909 47
rect 4947 13 4981 47
rect 5019 13 5053 47
rect 5091 13 5125 47
rect 5235 13 5269 47
rect 5307 13 5341 47
rect 5379 13 5413 47
rect 5451 13 5485 47
rect 5523 13 5557 47
rect 5595 13 5629 47
rect 5693 13 5727 47
rect 5765 13 5799 47
rect 5837 13 5871 47
rect 5909 13 5943 47
rect 5981 13 6015 47
rect 6053 13 6087 47
rect 6197 13 6231 47
rect 6269 13 6303 47
rect 6341 13 6375 47
rect 6413 13 6447 47
rect 6485 13 6519 47
rect 6557 13 6591 47
rect 6655 13 6689 47
rect 6727 13 6761 47
rect 6799 13 6833 47
rect 6871 13 6905 47
rect 6943 13 6977 47
rect 7015 13 7049 47
rect 7159 13 7193 47
rect 7231 13 7265 47
rect 7303 13 7337 47
rect 7375 13 7409 47
rect 7465 13 7499 47
rect 7537 13 7571 47
rect 7609 13 7643 47
rect 7681 13 7715 47
rect 7825 13 7859 47
rect 7897 13 7931 47
rect 7969 13 8003 47
rect 8041 13 8075 47
rect 8113 13 8147 47
rect 8185 13 8219 47
rect 8283 13 8317 47
rect 8355 13 8389 47
rect 8427 13 8461 47
rect 8499 13 8533 47
rect 8571 13 8605 47
rect 8643 13 8677 47
rect 8787 13 8821 47
rect 8859 13 8893 47
rect 8931 13 8965 47
rect 9003 13 9037 47
rect 9075 13 9109 47
rect 9147 13 9181 47
rect 9245 13 9279 47
rect 9317 13 9351 47
rect 9389 13 9423 47
rect 9461 13 9495 47
rect 9533 13 9567 47
rect 9605 13 9639 47
rect 9749 13 9783 47
rect 9821 13 9855 47
rect 9893 13 9927 47
rect 9965 13 9999 47
rect 10055 13 10089 47
rect 10127 13 10161 47
rect 10199 13 10233 47
rect 10271 13 10305 47
rect 10415 13 10449 47
rect 10487 13 10521 47
rect 10559 13 10593 47
rect 10631 13 10665 47
rect 10703 13 10737 47
rect 10775 13 10809 47
rect 10873 13 10907 47
rect 10945 13 10979 47
rect 11017 13 11051 47
rect 11089 13 11123 47
rect 11161 13 11195 47
rect 11233 13 11267 47
rect 11377 13 11411 47
rect 11449 13 11483 47
rect 11521 13 11555 47
rect 11593 13 11627 47
rect 11665 13 11699 47
rect 11737 13 11771 47
rect 11835 13 11869 47
rect 11907 13 11941 47
rect 11979 13 12013 47
rect 12051 13 12085 47
rect 12123 13 12157 47
rect 12195 13 12229 47
rect 12339 13 12373 47
rect 12411 13 12445 47
rect 12483 13 12517 47
rect 12555 13 12589 47
rect 12645 13 12679 47
rect 12717 13 12751 47
rect 12789 13 12823 47
rect 12861 13 12895 47
rect 13005 13 13039 47
rect 13077 13 13111 47
rect 13149 13 13183 47
rect 13221 13 13255 47
rect 13293 13 13327 47
rect 13365 13 13399 47
rect 13463 13 13497 47
rect 13535 13 13569 47
rect 13607 13 13641 47
rect 13679 13 13713 47
rect 13751 13 13785 47
rect 13823 13 13857 47
rect 13967 13 14001 47
rect 14039 13 14073 47
rect 14111 13 14145 47
rect 14183 13 14217 47
rect 14255 13 14289 47
rect 14327 13 14361 47
rect 14425 13 14459 47
rect 14497 13 14531 47
rect 14569 13 14603 47
rect 14641 13 14675 47
rect 14713 13 14747 47
rect 14785 13 14819 47
rect 14929 13 14963 47
rect 15001 13 15035 47
rect 15073 13 15107 47
rect 15145 13 15179 47
rect 15235 13 15269 47
rect 15307 13 15341 47
rect 15379 13 15413 47
rect 15451 13 15485 47
rect 15595 13 15629 47
rect 15667 13 15701 47
rect 15739 13 15773 47
rect 15811 13 15845 47
rect 15901 13 15935 47
rect 15973 13 16007 47
rect 16045 13 16079 47
rect 16117 13 16151 47
rect 16261 13 16295 47
rect 16333 13 16367 47
rect 16405 13 16439 47
rect 16477 13 16511 47
rect 16567 13 16601 47
rect 16639 13 16673 47
rect 16711 13 16745 47
rect 16783 13 16817 47
rect 16927 13 16961 47
rect 16999 13 17033 47
rect 17071 13 17105 47
rect 17143 13 17177 47
rect 17233 13 17267 47
rect 17305 13 17339 47
rect 17377 13 17411 47
rect 17449 13 17483 47
rect 17593 13 17627 47
rect 17665 13 17699 47
rect 17743 13 17777 47
rect 17821 13 17855 47
rect 17893 13 17927 47
<< metal1 >>
rect -31 1539 18013 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 343 1539
rect 377 1505 415 1539
rect 449 1505 513 1539
rect 547 1505 585 1539
rect 619 1505 657 1539
rect 691 1505 729 1539
rect 763 1505 801 1539
rect 835 1505 873 1539
rect 907 1505 1017 1539
rect 1051 1505 1089 1539
rect 1123 1505 1161 1539
rect 1195 1505 1233 1539
rect 1267 1505 1305 1539
rect 1339 1505 1377 1539
rect 1411 1505 1475 1539
rect 1509 1505 1547 1539
rect 1581 1505 1619 1539
rect 1653 1505 1691 1539
rect 1725 1505 1763 1539
rect 1797 1505 1835 1539
rect 1869 1505 1979 1539
rect 2013 1505 2051 1539
rect 2085 1505 2123 1539
rect 2157 1505 2195 1539
rect 2229 1505 2285 1539
rect 2319 1505 2357 1539
rect 2391 1505 2429 1539
rect 2463 1505 2501 1539
rect 2535 1505 2645 1539
rect 2679 1505 2717 1539
rect 2751 1505 2789 1539
rect 2823 1505 2861 1539
rect 2895 1505 2933 1539
rect 2967 1505 3005 1539
rect 3039 1505 3103 1539
rect 3137 1505 3175 1539
rect 3209 1505 3247 1539
rect 3281 1505 3319 1539
rect 3353 1505 3391 1539
rect 3425 1505 3463 1539
rect 3497 1505 3607 1539
rect 3641 1505 3679 1539
rect 3713 1505 3751 1539
rect 3785 1505 3823 1539
rect 3857 1505 3895 1539
rect 3929 1505 3967 1539
rect 4001 1505 4065 1539
rect 4099 1505 4137 1539
rect 4171 1505 4209 1539
rect 4243 1505 4281 1539
rect 4315 1505 4353 1539
rect 4387 1505 4425 1539
rect 4459 1505 4569 1539
rect 4603 1505 4641 1539
rect 4675 1505 4713 1539
rect 4747 1505 4785 1539
rect 4819 1505 4875 1539
rect 4909 1505 4947 1539
rect 4981 1505 5019 1539
rect 5053 1505 5091 1539
rect 5125 1505 5235 1539
rect 5269 1505 5307 1539
rect 5341 1505 5379 1539
rect 5413 1505 5451 1539
rect 5485 1505 5523 1539
rect 5557 1505 5595 1539
rect 5629 1505 5693 1539
rect 5727 1505 5765 1539
rect 5799 1505 5837 1539
rect 5871 1505 5909 1539
rect 5943 1505 5981 1539
rect 6015 1505 6053 1539
rect 6087 1505 6197 1539
rect 6231 1505 6269 1539
rect 6303 1505 6341 1539
rect 6375 1505 6413 1539
rect 6447 1505 6485 1539
rect 6519 1505 6557 1539
rect 6591 1505 6655 1539
rect 6689 1505 6727 1539
rect 6761 1505 6799 1539
rect 6833 1505 6871 1539
rect 6905 1505 6943 1539
rect 6977 1505 7015 1539
rect 7049 1505 7159 1539
rect 7193 1505 7231 1539
rect 7265 1505 7303 1539
rect 7337 1505 7375 1539
rect 7409 1505 7465 1539
rect 7499 1505 7537 1539
rect 7571 1505 7609 1539
rect 7643 1505 7681 1539
rect 7715 1505 7825 1539
rect 7859 1505 7897 1539
rect 7931 1505 7969 1539
rect 8003 1505 8041 1539
rect 8075 1505 8113 1539
rect 8147 1505 8185 1539
rect 8219 1505 8283 1539
rect 8317 1505 8355 1539
rect 8389 1505 8427 1539
rect 8461 1505 8499 1539
rect 8533 1505 8571 1539
rect 8605 1505 8643 1539
rect 8677 1505 8787 1539
rect 8821 1505 8859 1539
rect 8893 1505 8931 1539
rect 8965 1505 9003 1539
rect 9037 1505 9075 1539
rect 9109 1505 9147 1539
rect 9181 1505 9245 1539
rect 9279 1505 9317 1539
rect 9351 1505 9389 1539
rect 9423 1505 9461 1539
rect 9495 1505 9533 1539
rect 9567 1505 9605 1539
rect 9639 1505 9749 1539
rect 9783 1505 9821 1539
rect 9855 1505 9893 1539
rect 9927 1505 9965 1539
rect 9999 1505 10055 1539
rect 10089 1505 10127 1539
rect 10161 1505 10199 1539
rect 10233 1505 10271 1539
rect 10305 1505 10415 1539
rect 10449 1505 10487 1539
rect 10521 1505 10559 1539
rect 10593 1505 10631 1539
rect 10665 1505 10703 1539
rect 10737 1505 10775 1539
rect 10809 1505 10873 1539
rect 10907 1505 10945 1539
rect 10979 1505 11017 1539
rect 11051 1505 11089 1539
rect 11123 1505 11161 1539
rect 11195 1505 11233 1539
rect 11267 1505 11377 1539
rect 11411 1505 11449 1539
rect 11483 1505 11521 1539
rect 11555 1505 11593 1539
rect 11627 1505 11665 1539
rect 11699 1505 11737 1539
rect 11771 1505 11835 1539
rect 11869 1505 11907 1539
rect 11941 1505 11979 1539
rect 12013 1505 12051 1539
rect 12085 1505 12123 1539
rect 12157 1505 12195 1539
rect 12229 1505 12339 1539
rect 12373 1505 12411 1539
rect 12445 1505 12483 1539
rect 12517 1505 12555 1539
rect 12589 1505 12645 1539
rect 12679 1505 12717 1539
rect 12751 1505 12789 1539
rect 12823 1505 12861 1539
rect 12895 1505 13005 1539
rect 13039 1505 13077 1539
rect 13111 1505 13149 1539
rect 13183 1505 13221 1539
rect 13255 1505 13293 1539
rect 13327 1505 13365 1539
rect 13399 1505 13463 1539
rect 13497 1505 13535 1539
rect 13569 1505 13607 1539
rect 13641 1505 13679 1539
rect 13713 1505 13751 1539
rect 13785 1505 13823 1539
rect 13857 1505 13967 1539
rect 14001 1505 14039 1539
rect 14073 1505 14111 1539
rect 14145 1505 14183 1539
rect 14217 1505 14255 1539
rect 14289 1505 14327 1539
rect 14361 1505 14425 1539
rect 14459 1505 14497 1539
rect 14531 1505 14569 1539
rect 14603 1505 14641 1539
rect 14675 1505 14713 1539
rect 14747 1505 14785 1539
rect 14819 1505 14929 1539
rect 14963 1505 15001 1539
rect 15035 1505 15073 1539
rect 15107 1505 15145 1539
rect 15179 1505 15235 1539
rect 15269 1505 15307 1539
rect 15341 1505 15379 1539
rect 15413 1505 15451 1539
rect 15485 1505 15595 1539
rect 15629 1505 15667 1539
rect 15701 1505 15739 1539
rect 15773 1505 15811 1539
rect 15845 1505 15901 1539
rect 15935 1505 15973 1539
rect 16007 1505 16045 1539
rect 16079 1505 16117 1539
rect 16151 1505 16261 1539
rect 16295 1505 16333 1539
rect 16367 1505 16405 1539
rect 16439 1505 16477 1539
rect 16511 1505 16567 1539
rect 16601 1505 16639 1539
rect 16673 1505 16711 1539
rect 16745 1505 16783 1539
rect 16817 1505 16927 1539
rect 16961 1505 16999 1539
rect 17033 1505 17071 1539
rect 17105 1505 17143 1539
rect 17177 1505 17233 1539
rect 17267 1505 17305 1539
rect 17339 1505 17377 1539
rect 17411 1505 17449 1539
rect 17483 1505 17593 1539
rect 17627 1505 17665 1539
rect 17699 1505 17743 1539
rect 17777 1505 17821 1539
rect 17855 1505 17893 1539
rect 17927 1505 18013 1539
rect -31 1492 18013 1505
rect 15939 1105 15985 1111
rect 16339 1105 16385 1111
rect 16603 1105 16649 1111
rect 17007 1105 17053 1111
rect 15933 1071 15945 1105
rect 15979 1071 16345 1105
rect 16379 1071 16391 1105
rect 16597 1071 16609 1105
rect 16643 1071 17013 1105
rect 17047 1071 17059 1105
rect 15939 1065 15985 1071
rect 16339 1065 16385 1071
rect 16603 1065 16649 1071
rect 17007 1065 17053 1071
rect 4195 979 4241 985
rect 5009 979 5055 985
rect 15887 979 15933 985
rect 4189 945 4201 979
rect 4235 945 5015 979
rect 5049 945 15893 979
rect 15927 945 15939 979
rect 4195 939 4241 945
rect 5009 939 5055 945
rect 15887 939 15933 945
rect 791 905 837 911
rect 1161 905 1207 911
rect 3751 905 3797 911
rect 4343 905 4389 911
rect 4713 905 4759 911
rect 5971 905 6017 911
rect 6341 905 6387 911
rect 8931 905 8977 911
rect 9523 905 9569 911
rect 9893 905 9939 911
rect 11151 905 11197 911
rect 11521 905 11567 911
rect 14111 905 14157 911
rect 14703 905 14749 911
rect 15073 905 15119 911
rect 15665 905 15711 911
rect 16405 905 16451 911
rect 16701 905 16747 911
rect 16997 905 17043 911
rect 785 871 797 905
rect 831 871 1167 905
rect 1201 871 3757 905
rect 3791 871 3803 905
rect 4337 871 4349 905
rect 4383 871 4719 905
rect 4753 871 4765 905
rect 5965 871 5977 905
rect 6011 871 6347 905
rect 6381 871 8937 905
rect 8971 871 8983 905
rect 9517 871 9529 905
rect 9563 871 9899 905
rect 9933 871 9945 905
rect 11145 871 11157 905
rect 11191 871 11527 905
rect 11561 871 14117 905
rect 14151 871 14163 905
rect 14697 871 14709 905
rect 14743 871 15079 905
rect 15113 871 15125 905
rect 15659 871 15671 905
rect 15705 871 16411 905
rect 16445 871 16457 905
rect 16695 871 16707 905
rect 16741 871 17003 905
rect 17037 871 17049 905
rect 791 865 837 871
rect 1161 865 1207 871
rect 3751 865 3797 871
rect 4343 865 4389 871
rect 4713 865 4759 871
rect 5971 865 6017 871
rect 6341 865 6387 871
rect 8931 865 8977 871
rect 9523 865 9569 871
rect 9893 865 9939 871
rect 11151 865 11197 871
rect 11521 865 11567 871
rect 14111 865 14157 871
rect 14703 865 14749 871
rect 15073 865 15119 871
rect 15665 865 15711 871
rect 16405 865 16451 871
rect 16701 865 16747 871
rect 16997 865 17043 871
rect 421 831 467 837
rect 3011 831 3057 837
rect 5601 831 5647 837
rect 8191 831 8237 837
rect 10781 831 10827 837
rect 13371 831 13417 837
rect 15887 831 15933 837
rect 17219 831 17265 837
rect 17367 831 17413 837
rect 17663 831 17709 837
rect 17811 831 17857 837
rect 415 797 427 831
rect 461 797 3017 831
rect 3051 797 5607 831
rect 5641 797 8197 831
rect 8231 797 10787 831
rect 10821 797 13377 831
rect 13411 797 13423 831
rect 15881 797 15893 831
rect 15927 797 17225 831
rect 17259 797 17271 831
rect 17361 797 17373 831
rect 17407 797 17669 831
rect 17703 797 17715 831
rect 17805 797 17817 831
rect 17851 797 17887 831
rect 421 791 467 797
rect 3011 791 3057 797
rect 5601 791 5647 797
rect 8191 791 8237 797
rect 10781 791 10827 797
rect 13371 791 13417 797
rect 15887 791 15933 797
rect 17219 791 17265 797
rect 17367 791 17413 797
rect 17663 791 17709 797
rect 17811 791 17857 797
rect 199 757 245 763
rect 2271 757 2317 763
rect 3381 757 3427 763
rect 4861 757 4907 763
rect 5379 757 5425 763
rect 7451 757 7497 763
rect 8561 757 8607 763
rect 10041 757 10087 763
rect 10559 757 10605 763
rect 12631 757 12677 763
rect 13741 757 13787 763
rect 15221 757 15267 763
rect 15369 757 15415 763
rect 16701 757 16747 763
rect 193 723 205 757
rect 239 723 2277 757
rect 2311 723 3387 757
rect 3421 723 4867 757
rect 4901 723 4913 757
rect 5373 723 5385 757
rect 5419 723 7457 757
rect 7491 723 8567 757
rect 8601 723 10047 757
rect 10081 723 10093 757
rect 10553 723 10565 757
rect 10599 723 12637 757
rect 12671 723 13747 757
rect 13781 723 15227 757
rect 15261 723 15273 757
rect 15363 723 15375 757
rect 15409 723 16707 757
rect 16741 723 16753 757
rect 199 717 245 723
rect 2271 717 2317 723
rect 3381 717 3427 723
rect 4861 717 4907 723
rect 5379 717 5425 723
rect 7451 717 7497 723
rect 8561 717 8607 723
rect 10041 717 10087 723
rect 10559 717 10605 723
rect 12631 717 12677 723
rect 13741 717 13787 723
rect 15221 717 15267 723
rect 15369 717 15415 723
rect 16701 717 16747 723
rect 1605 683 1651 689
rect 3233 683 3279 689
rect 3973 683 4019 689
rect 6785 683 6831 689
rect 8413 683 8459 689
rect 9153 683 9199 689
rect 11965 683 12011 689
rect 13593 683 13639 689
rect 14333 683 14379 689
rect 1599 649 1611 683
rect 1645 649 3239 683
rect 3273 649 3979 683
rect 4013 649 6791 683
rect 6825 649 8419 683
rect 8453 649 9159 683
rect 9193 649 11971 683
rect 12005 649 13599 683
rect 13633 649 14339 683
rect 14373 649 14385 683
rect 1605 643 1651 649
rect 3233 643 3279 649
rect 3973 643 4019 649
rect 6785 643 6831 649
rect 8413 643 8459 649
rect 9153 643 9199 649
rect 11965 643 12011 649
rect 13593 643 13639 649
rect 14333 643 14379 649
rect 643 609 689 615
rect 1753 609 1799 615
rect 2123 609 2169 615
rect 2419 609 2465 615
rect 2789 609 2835 615
rect 5823 609 5869 615
rect 6933 609 6979 615
rect 7303 609 7349 615
rect 7599 609 7645 615
rect 7969 609 8015 615
rect 11003 609 11049 615
rect 12113 609 12159 615
rect 12483 609 12529 615
rect 12779 609 12825 615
rect 13149 609 13195 615
rect 637 575 649 609
rect 683 575 1759 609
rect 1793 575 2129 609
rect 2163 575 2175 609
rect 2413 575 2425 609
rect 2459 575 2795 609
rect 2829 575 2841 609
rect 5817 575 5829 609
rect 5863 575 6939 609
rect 6973 575 7309 609
rect 7343 575 7355 609
rect 7593 575 7605 609
rect 7639 575 7975 609
rect 8009 575 8021 609
rect 10997 575 11009 609
rect 11043 575 12119 609
rect 12153 575 12489 609
rect 12523 575 12535 609
rect 12773 575 12785 609
rect 12819 575 13155 609
rect 13189 575 13201 609
rect 643 569 689 575
rect 1753 569 1799 575
rect 2123 569 2169 575
rect 2419 569 2465 575
rect 2789 569 2835 575
rect 5823 569 5869 575
rect 6933 569 6979 575
rect 7303 569 7349 575
rect 7599 569 7645 575
rect 7969 569 8015 575
rect 11003 569 11049 575
rect 12113 569 12159 575
rect 12483 569 12529 575
rect 12779 569 12825 575
rect 13149 569 13195 575
rect 9375 535 9421 541
rect 10189 535 10235 541
rect 15665 535 15711 541
rect 16405 535 16451 541
rect 16701 535 16747 541
rect 16997 535 17043 541
rect 9369 501 9381 535
rect 9415 501 10195 535
rect 10229 501 15671 535
rect 15705 501 16411 535
rect 16445 501 16457 535
rect 16695 501 16707 535
rect 16741 501 17003 535
rect 17037 501 17049 535
rect 9375 495 9421 501
rect 10189 495 10235 501
rect 15665 495 15711 501
rect 16405 495 16451 501
rect 16701 495 16747 501
rect 16997 495 17043 501
rect 1383 461 1429 467
rect 6563 461 6609 467
rect 11743 461 11789 467
rect 1353 427 1389 461
rect 1423 427 6569 461
rect 6603 427 11749 461
rect 11783 427 11795 461
rect 1383 421 1429 427
rect 6563 421 6609 427
rect 11743 421 11789 427
rect 15947 281 15993 287
rect 16613 281 16659 287
rect 17279 281 17325 287
rect 15941 247 15953 281
rect 15987 247 16619 281
rect 16653 247 17285 281
rect 17319 247 17331 281
rect 15947 241 15993 247
rect 16613 241 16659 247
rect 17279 241 17325 247
rect -31 47 18013 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 343 47
rect 377 13 415 47
rect 449 13 513 47
rect 547 13 585 47
rect 619 13 657 47
rect 691 13 729 47
rect 763 13 801 47
rect 835 13 873 47
rect 907 13 1017 47
rect 1051 13 1089 47
rect 1123 13 1161 47
rect 1195 13 1233 47
rect 1267 13 1305 47
rect 1339 13 1377 47
rect 1411 13 1475 47
rect 1509 13 1547 47
rect 1581 13 1619 47
rect 1653 13 1691 47
rect 1725 13 1763 47
rect 1797 13 1835 47
rect 1869 13 1979 47
rect 2013 13 2051 47
rect 2085 13 2123 47
rect 2157 13 2195 47
rect 2229 13 2285 47
rect 2319 13 2357 47
rect 2391 13 2429 47
rect 2463 13 2501 47
rect 2535 13 2645 47
rect 2679 13 2717 47
rect 2751 13 2789 47
rect 2823 13 2861 47
rect 2895 13 2933 47
rect 2967 13 3005 47
rect 3039 13 3103 47
rect 3137 13 3175 47
rect 3209 13 3247 47
rect 3281 13 3319 47
rect 3353 13 3391 47
rect 3425 13 3463 47
rect 3497 13 3607 47
rect 3641 13 3679 47
rect 3713 13 3751 47
rect 3785 13 3823 47
rect 3857 13 3895 47
rect 3929 13 3967 47
rect 4001 13 4065 47
rect 4099 13 4137 47
rect 4171 13 4209 47
rect 4243 13 4281 47
rect 4315 13 4353 47
rect 4387 13 4425 47
rect 4459 13 4569 47
rect 4603 13 4641 47
rect 4675 13 4713 47
rect 4747 13 4785 47
rect 4819 13 4875 47
rect 4909 13 4947 47
rect 4981 13 5019 47
rect 5053 13 5091 47
rect 5125 13 5235 47
rect 5269 13 5307 47
rect 5341 13 5379 47
rect 5413 13 5451 47
rect 5485 13 5523 47
rect 5557 13 5595 47
rect 5629 13 5693 47
rect 5727 13 5765 47
rect 5799 13 5837 47
rect 5871 13 5909 47
rect 5943 13 5981 47
rect 6015 13 6053 47
rect 6087 13 6197 47
rect 6231 13 6269 47
rect 6303 13 6341 47
rect 6375 13 6413 47
rect 6447 13 6485 47
rect 6519 13 6557 47
rect 6591 13 6655 47
rect 6689 13 6727 47
rect 6761 13 6799 47
rect 6833 13 6871 47
rect 6905 13 6943 47
rect 6977 13 7015 47
rect 7049 13 7159 47
rect 7193 13 7231 47
rect 7265 13 7303 47
rect 7337 13 7375 47
rect 7409 13 7465 47
rect 7499 13 7537 47
rect 7571 13 7609 47
rect 7643 13 7681 47
rect 7715 13 7825 47
rect 7859 13 7897 47
rect 7931 13 7969 47
rect 8003 13 8041 47
rect 8075 13 8113 47
rect 8147 13 8185 47
rect 8219 13 8283 47
rect 8317 13 8355 47
rect 8389 13 8427 47
rect 8461 13 8499 47
rect 8533 13 8571 47
rect 8605 13 8643 47
rect 8677 13 8787 47
rect 8821 13 8859 47
rect 8893 13 8931 47
rect 8965 13 9003 47
rect 9037 13 9075 47
rect 9109 13 9147 47
rect 9181 13 9245 47
rect 9279 13 9317 47
rect 9351 13 9389 47
rect 9423 13 9461 47
rect 9495 13 9533 47
rect 9567 13 9605 47
rect 9639 13 9749 47
rect 9783 13 9821 47
rect 9855 13 9893 47
rect 9927 13 9965 47
rect 9999 13 10055 47
rect 10089 13 10127 47
rect 10161 13 10199 47
rect 10233 13 10271 47
rect 10305 13 10415 47
rect 10449 13 10487 47
rect 10521 13 10559 47
rect 10593 13 10631 47
rect 10665 13 10703 47
rect 10737 13 10775 47
rect 10809 13 10873 47
rect 10907 13 10945 47
rect 10979 13 11017 47
rect 11051 13 11089 47
rect 11123 13 11161 47
rect 11195 13 11233 47
rect 11267 13 11377 47
rect 11411 13 11449 47
rect 11483 13 11521 47
rect 11555 13 11593 47
rect 11627 13 11665 47
rect 11699 13 11737 47
rect 11771 13 11835 47
rect 11869 13 11907 47
rect 11941 13 11979 47
rect 12013 13 12051 47
rect 12085 13 12123 47
rect 12157 13 12195 47
rect 12229 13 12339 47
rect 12373 13 12411 47
rect 12445 13 12483 47
rect 12517 13 12555 47
rect 12589 13 12645 47
rect 12679 13 12717 47
rect 12751 13 12789 47
rect 12823 13 12861 47
rect 12895 13 13005 47
rect 13039 13 13077 47
rect 13111 13 13149 47
rect 13183 13 13221 47
rect 13255 13 13293 47
rect 13327 13 13365 47
rect 13399 13 13463 47
rect 13497 13 13535 47
rect 13569 13 13607 47
rect 13641 13 13679 47
rect 13713 13 13751 47
rect 13785 13 13823 47
rect 13857 13 13967 47
rect 14001 13 14039 47
rect 14073 13 14111 47
rect 14145 13 14183 47
rect 14217 13 14255 47
rect 14289 13 14327 47
rect 14361 13 14425 47
rect 14459 13 14497 47
rect 14531 13 14569 47
rect 14603 13 14641 47
rect 14675 13 14713 47
rect 14747 13 14785 47
rect 14819 13 14929 47
rect 14963 13 15001 47
rect 15035 13 15073 47
rect 15107 13 15145 47
rect 15179 13 15235 47
rect 15269 13 15307 47
rect 15341 13 15379 47
rect 15413 13 15451 47
rect 15485 13 15595 47
rect 15629 13 15667 47
rect 15701 13 15739 47
rect 15773 13 15811 47
rect 15845 13 15901 47
rect 15935 13 15973 47
rect 16007 13 16045 47
rect 16079 13 16117 47
rect 16151 13 16261 47
rect 16295 13 16333 47
rect 16367 13 16405 47
rect 16439 13 16477 47
rect 16511 13 16567 47
rect 16601 13 16639 47
rect 16673 13 16711 47
rect 16745 13 16783 47
rect 16817 13 16927 47
rect 16961 13 16999 47
rect 17033 13 17071 47
rect 17105 13 17143 47
rect 17177 13 17233 47
rect 17267 13 17305 47
rect 17339 13 17377 47
rect 17411 13 17449 47
rect 17483 13 17593 47
rect 17627 13 17665 47
rect 17699 13 17743 47
rect 17777 13 17821 47
rect 17855 13 17893 47
rect 17927 13 18013 47
rect -31 0 18013 13
<< labels >>
rlabel metal1 17817 797 17851 831 1 Q
port 1 n
rlabel metal1 1389 427 1423 461 1 D
port 2 n
rlabel metal1 427 797 461 831 1 CLK
port 3 n
rlabel metal1 1611 649 1645 683 1 RN
port 4 n
rlabel metal1 72 1522 72 1522 1 VDD
port 5 n
rlabel metal1 72 30 72 30 1 VSS
port 6 n
rlabel metal1 15671 461 15705 988 1 voter3x1_pcell_0/votern3x1_pcell_0/B
rlabel space 15672 501 16411 535 1 voter3x1_pcell_0/votern3x1_pcell_0/B
rlabel space 15893 461 15927 970 1 voter3x1_pcell_0/votern3x1_pcell_0/A
rlabel metal1 16707 461 16741 988 1 voter3x1_pcell_0/votern3x1_pcell_0/C
rlabel metal1 17225 461 17259 1020 1 voter3x1_pcell_0/votern3x1_pcell_0/A
rlabel space 15927 797 17230 831 1 voter3x1_pcell_0/votern3x1_pcell_0/A
rlabel space 16741 871 17003 905 1 voter3x1_pcell_0/votern3x1_pcell_0/C
rlabel space 16741 501 17003 535 1 voter3x1_pcell_0/votern3x1_pcell_0/C
rlabel space 15705 871 16457 905 1 voter3x1_pcell_0/votern3x1_pcell_0/B
<< end >>
