magic
tech sky130A
magscale 1 2
timestamp 1648067205
<< nwell >>
rect -84 833 2082 1576
<< nmos >>
rect 168 317 198 378
tri 198 317 214 333 sw
rect 362 325 392 378
tri 392 325 408 341 sw
rect 168 287 274 317
tri 274 287 304 317 sw
rect 362 295 468 325
tri 468 295 498 325 sw
rect 168 186 198 287
tri 198 271 214 287 nw
tri 258 271 274 287 ne
tri 198 186 214 202 sw
tri 258 186 274 202 se
rect 274 186 304 287
rect 362 194 392 295
tri 392 279 408 295 nw
tri 452 279 468 295 ne
tri 392 194 408 210 sw
tri 452 194 468 210 se
rect 468 194 498 295
tri 168 156 198 186 ne
rect 198 156 274 186
tri 274 156 304 186 nw
tri 362 164 392 194 ne
rect 392 164 468 194
tri 468 164 498 194 nw
rect 834 317 864 378
tri 864 317 880 333 sw
tri 1118 325 1134 341 se
rect 1134 325 1164 378
rect 834 287 940 317
tri 940 287 970 317 sw
tri 1028 295 1058 325 se
rect 1058 295 1164 325
rect 834 186 864 287
tri 864 271 880 287 nw
tri 924 271 940 287 ne
tri 864 186 880 202 sw
tri 924 186 940 202 se
rect 940 186 970 287
rect 1028 194 1058 295
tri 1058 279 1074 295 nw
tri 1118 279 1134 295 ne
tri 1058 194 1074 210 sw
tri 1118 194 1134 210 se
rect 1134 194 1164 295
tri 834 156 864 186 ne
rect 864 156 940 186
tri 940 156 970 186 nw
tri 1028 164 1058 194 ne
rect 1058 164 1134 194
tri 1134 164 1164 194 nw
rect 1500 317 1530 378
tri 1530 317 1546 333 sw
rect 1694 325 1724 378
tri 1724 325 1740 341 sw
rect 1500 287 1606 317
tri 1606 287 1636 317 sw
rect 1694 295 1800 325
tri 1800 295 1830 325 sw
rect 1500 186 1530 287
tri 1530 271 1546 287 nw
tri 1590 271 1606 287 ne
tri 1530 186 1546 202 sw
tri 1590 186 1606 202 se
rect 1606 186 1636 287
rect 1694 280 1725 295
tri 1725 280 1740 295 nw
tri 1784 280 1799 295 ne
rect 1799 280 1830 295
rect 1694 194 1724 280
tri 1724 194 1740 210 sw
tri 1784 194 1800 210 se
rect 1800 194 1830 280
tri 1500 156 1530 186 ne
rect 1530 156 1606 186
tri 1606 156 1636 186 nw
tri 1694 164 1724 194 ne
rect 1724 164 1800 194
tri 1800 164 1830 194 nw
<< pmos >>
rect 187 1052 217 1452
rect 275 1052 305 1452
rect 363 1052 393 1452
rect 451 1052 481 1452
rect 851 1052 881 1452
rect 939 1052 969 1452
rect 1027 1052 1057 1452
rect 1115 1052 1145 1452
rect 1519 1052 1549 1452
rect 1607 1052 1637 1452
rect 1695 1052 1725 1452
rect 1783 1052 1813 1452
<< ndiff >>
rect 112 362 168 378
rect 112 328 122 362
rect 156 328 168 362
rect 112 290 168 328
rect 198 362 362 378
rect 198 333 219 362
tri 198 317 214 333 ne
rect 214 328 219 333
rect 253 328 316 362
rect 350 328 362 362
rect 214 317 362 328
rect 392 362 552 378
rect 392 341 510 362
tri 392 325 408 341 ne
rect 408 328 510 341
rect 544 328 552 362
rect 408 325 552 328
rect 112 256 122 290
rect 156 256 168 290
tri 274 287 304 317 ne
rect 304 290 362 317
tri 468 295 498 325 ne
rect 112 222 168 256
rect 112 188 122 222
rect 156 188 168 222
rect 112 156 168 188
tri 198 271 214 287 se
rect 214 271 258 287
tri 258 271 274 287 sw
rect 198 237 274 271
rect 198 203 219 237
rect 253 203 274 237
rect 198 202 274 203
tri 198 186 214 202 ne
rect 214 186 258 202
tri 258 186 274 202 nw
rect 304 256 316 290
rect 350 256 362 290
rect 304 222 362 256
rect 304 188 316 222
rect 350 188 362 222
tri 392 279 408 295 se
rect 408 279 452 295
tri 452 279 468 295 sw
rect 392 246 468 279
rect 392 212 412 246
rect 446 212 468 246
rect 392 210 468 212
tri 392 194 408 210 ne
rect 408 194 452 210
tri 452 194 468 210 nw
rect 498 290 552 325
rect 498 256 510 290
rect 544 256 552 290
rect 498 222 552 256
tri 168 156 198 186 sw
tri 274 156 304 186 se
rect 304 164 362 188
tri 362 164 392 194 sw
tri 468 164 498 194 se
rect 498 188 510 222
rect 544 188 552 222
rect 498 164 552 188
rect 304 156 552 164
rect 112 152 552 156
rect 112 118 122 152
rect 156 118 316 152
rect 350 118 412 152
rect 446 118 510 152
rect 544 118 552 152
rect 112 102 552 118
rect 778 362 834 378
rect 778 328 788 362
rect 822 328 834 362
rect 778 290 834 328
rect 864 362 1134 378
rect 864 333 885 362
tri 864 317 880 333 ne
rect 880 328 885 333
rect 919 328 982 362
rect 1016 341 1134 362
rect 1016 328 1118 341
rect 880 325 1118 328
tri 1118 325 1134 341 nw
rect 1164 362 1220 378
rect 1164 328 1176 362
rect 1210 328 1220 362
rect 880 317 1028 325
rect 778 256 788 290
rect 822 256 834 290
tri 940 287 970 317 ne
rect 970 290 1028 317
tri 1028 295 1058 325 nw
rect 778 222 834 256
rect 778 188 788 222
rect 822 188 834 222
rect 778 156 834 188
tri 864 271 880 287 se
rect 880 271 924 287
tri 924 271 940 287 sw
rect 864 237 940 271
rect 864 203 885 237
rect 919 203 940 237
rect 864 202 940 203
tri 864 186 880 202 ne
rect 880 186 924 202
tri 924 186 940 202 nw
rect 970 256 982 290
rect 1016 256 1028 290
rect 970 222 1028 256
rect 970 188 982 222
rect 1016 188 1028 222
tri 1058 279 1074 295 se
rect 1074 279 1118 295
tri 1118 279 1134 295 sw
rect 1058 246 1134 279
rect 1058 212 1079 246
rect 1113 212 1134 246
rect 1058 210 1134 212
tri 1058 194 1074 210 ne
rect 1074 194 1118 210
tri 1118 194 1134 210 nw
rect 1164 290 1220 328
rect 1164 256 1176 290
rect 1210 256 1220 290
rect 1164 222 1220 256
tri 834 156 864 186 sw
tri 940 156 970 186 se
rect 970 164 1028 188
tri 1028 164 1058 194 sw
tri 1134 164 1164 194 se
rect 1164 188 1176 222
rect 1210 188 1220 222
rect 1164 164 1220 188
rect 970 156 1220 164
rect 778 152 1220 156
rect 778 118 788 152
rect 822 118 982 152
rect 1016 118 1079 152
rect 1113 118 1176 152
rect 1210 118 1220 152
rect 778 102 1220 118
rect 1444 362 1500 378
rect 1444 328 1454 362
rect 1488 328 1500 362
rect 1444 290 1500 328
rect 1530 362 1694 378
rect 1530 333 1551 362
tri 1530 317 1546 333 ne
rect 1546 328 1551 333
rect 1585 328 1648 362
rect 1682 328 1694 362
rect 1546 317 1694 328
rect 1724 341 1886 378
tri 1724 325 1740 341 ne
rect 1740 325 1886 341
rect 1444 256 1454 290
rect 1488 256 1500 290
tri 1606 287 1636 317 ne
rect 1636 290 1694 317
tri 1800 295 1830 325 ne
rect 1444 222 1500 256
rect 1444 188 1454 222
rect 1488 188 1500 222
rect 1444 156 1500 188
tri 1530 271 1546 287 se
rect 1546 271 1590 287
tri 1590 271 1606 287 sw
rect 1530 237 1606 271
rect 1530 203 1551 237
rect 1585 203 1606 237
rect 1530 202 1606 203
tri 1530 186 1546 202 ne
rect 1546 186 1590 202
tri 1590 186 1606 202 nw
rect 1636 256 1648 290
rect 1682 256 1694 290
tri 1725 280 1740 295 se
rect 1740 280 1784 295
tri 1784 280 1799 295 sw
rect 1830 290 1886 325
rect 1636 222 1694 256
rect 1636 188 1648 222
rect 1682 188 1694 222
rect 1724 246 1800 280
rect 1724 212 1745 246
rect 1779 212 1800 246
rect 1724 210 1800 212
tri 1724 194 1740 210 ne
rect 1740 194 1784 210
tri 1784 194 1800 210 nw
rect 1830 256 1842 290
rect 1876 256 1886 290
rect 1830 222 1886 256
tri 1500 156 1530 186 sw
tri 1606 156 1636 186 se
rect 1636 164 1694 188
tri 1694 164 1724 194 sw
tri 1800 164 1830 194 se
rect 1830 188 1842 222
rect 1876 188 1886 222
rect 1830 164 1886 188
rect 1636 156 1886 164
rect 1444 152 1886 156
rect 1444 118 1454 152
rect 1488 118 1648 152
rect 1682 118 1745 152
rect 1779 118 1842 152
rect 1876 118 1886 152
rect 1444 102 1886 118
<< pdiff >>
rect 131 1412 187 1452
rect 131 1378 141 1412
rect 175 1378 187 1412
rect 131 1344 187 1378
rect 131 1310 141 1344
rect 175 1310 187 1344
rect 131 1276 187 1310
rect 131 1242 141 1276
rect 175 1242 187 1276
rect 131 1208 187 1242
rect 131 1174 141 1208
rect 175 1174 187 1208
rect 131 1140 187 1174
rect 131 1106 141 1140
rect 175 1106 187 1140
rect 131 1052 187 1106
rect 217 1412 275 1452
rect 217 1378 229 1412
rect 263 1378 275 1412
rect 217 1344 275 1378
rect 217 1310 229 1344
rect 263 1310 275 1344
rect 217 1276 275 1310
rect 217 1242 229 1276
rect 263 1242 275 1276
rect 217 1208 275 1242
rect 217 1174 229 1208
rect 263 1174 275 1208
rect 217 1140 275 1174
rect 217 1106 229 1140
rect 263 1106 275 1140
rect 217 1052 275 1106
rect 305 1412 363 1452
rect 305 1378 317 1412
rect 351 1378 363 1412
rect 305 1344 363 1378
rect 305 1310 317 1344
rect 351 1310 363 1344
rect 305 1276 363 1310
rect 305 1242 317 1276
rect 351 1242 363 1276
rect 305 1208 363 1242
rect 305 1174 317 1208
rect 351 1174 363 1208
rect 305 1052 363 1174
rect 393 1412 451 1452
rect 393 1378 405 1412
rect 439 1378 451 1412
rect 393 1344 451 1378
rect 393 1310 405 1344
rect 439 1310 451 1344
rect 393 1276 451 1310
rect 393 1242 405 1276
rect 439 1242 451 1276
rect 393 1208 451 1242
rect 393 1174 405 1208
rect 439 1174 451 1208
rect 393 1052 451 1174
rect 481 1412 535 1452
rect 481 1378 493 1412
rect 527 1378 535 1412
rect 481 1344 535 1378
rect 481 1310 493 1344
rect 527 1310 535 1344
rect 481 1276 535 1310
rect 481 1242 493 1276
rect 527 1242 535 1276
rect 481 1208 535 1242
rect 481 1174 493 1208
rect 527 1174 535 1208
rect 481 1140 535 1174
rect 481 1106 493 1140
rect 527 1106 535 1140
rect 481 1052 535 1106
rect 797 1412 851 1452
rect 797 1378 805 1412
rect 839 1378 851 1412
rect 797 1344 851 1378
rect 797 1310 805 1344
rect 839 1310 851 1344
rect 797 1276 851 1310
rect 797 1242 805 1276
rect 839 1242 851 1276
rect 797 1208 851 1242
rect 797 1174 805 1208
rect 839 1174 851 1208
rect 797 1052 851 1174
rect 881 1344 939 1452
rect 881 1310 893 1344
rect 927 1310 939 1344
rect 881 1276 939 1310
rect 881 1242 893 1276
rect 927 1242 939 1276
rect 881 1208 939 1242
rect 881 1174 893 1208
rect 927 1174 939 1208
rect 881 1140 939 1174
rect 881 1106 893 1140
rect 927 1106 939 1140
rect 881 1052 939 1106
rect 969 1412 1027 1452
rect 969 1378 981 1412
rect 1015 1378 1027 1412
rect 969 1344 1027 1378
rect 969 1310 981 1344
rect 1015 1310 1027 1344
rect 969 1276 1027 1310
rect 969 1242 981 1276
rect 1015 1242 1027 1276
rect 969 1208 1027 1242
rect 969 1174 981 1208
rect 1015 1174 1027 1208
rect 969 1052 1027 1174
rect 1057 1344 1115 1452
rect 1057 1310 1069 1344
rect 1103 1310 1115 1344
rect 1057 1276 1115 1310
rect 1057 1242 1069 1276
rect 1103 1242 1115 1276
rect 1057 1208 1115 1242
rect 1057 1174 1069 1208
rect 1103 1174 1115 1208
rect 1057 1052 1115 1174
rect 1145 1412 1201 1452
rect 1145 1378 1157 1412
rect 1191 1378 1201 1412
rect 1145 1344 1201 1378
rect 1145 1310 1157 1344
rect 1191 1310 1201 1344
rect 1145 1276 1201 1310
rect 1145 1242 1157 1276
rect 1191 1242 1201 1276
rect 1145 1208 1201 1242
rect 1145 1174 1157 1208
rect 1191 1174 1201 1208
rect 1145 1052 1201 1174
rect 1463 1412 1519 1452
rect 1463 1378 1473 1412
rect 1507 1378 1519 1412
rect 1463 1344 1519 1378
rect 1463 1310 1473 1344
rect 1507 1310 1519 1344
rect 1463 1276 1519 1310
rect 1463 1242 1473 1276
rect 1507 1242 1519 1276
rect 1463 1208 1519 1242
rect 1463 1174 1473 1208
rect 1507 1174 1519 1208
rect 1463 1052 1519 1174
rect 1549 1344 1607 1452
rect 1549 1310 1561 1344
rect 1595 1310 1607 1344
rect 1549 1276 1607 1310
rect 1549 1242 1561 1276
rect 1595 1242 1607 1276
rect 1549 1208 1607 1242
rect 1549 1174 1561 1208
rect 1595 1174 1607 1208
rect 1549 1140 1607 1174
rect 1549 1106 1561 1140
rect 1595 1106 1607 1140
rect 1549 1052 1607 1106
rect 1637 1412 1695 1452
rect 1637 1378 1649 1412
rect 1683 1378 1695 1412
rect 1637 1344 1695 1378
rect 1637 1310 1649 1344
rect 1683 1310 1695 1344
rect 1637 1276 1695 1310
rect 1637 1242 1649 1276
rect 1683 1242 1695 1276
rect 1637 1208 1695 1242
rect 1637 1174 1649 1208
rect 1683 1174 1695 1208
rect 1637 1052 1695 1174
rect 1725 1344 1783 1452
rect 1725 1310 1737 1344
rect 1771 1310 1783 1344
rect 1725 1276 1783 1310
rect 1725 1242 1737 1276
rect 1771 1242 1783 1276
rect 1725 1208 1783 1242
rect 1725 1174 1737 1208
rect 1771 1174 1783 1208
rect 1725 1140 1783 1174
rect 1725 1106 1737 1140
rect 1771 1106 1783 1140
rect 1725 1052 1783 1106
rect 1813 1412 1867 1452
rect 1813 1378 1825 1412
rect 1859 1378 1867 1412
rect 1813 1344 1867 1378
rect 1813 1310 1825 1344
rect 1859 1310 1867 1344
rect 1813 1276 1867 1310
rect 1813 1242 1825 1276
rect 1859 1242 1867 1276
rect 1813 1208 1867 1242
rect 1813 1174 1825 1208
rect 1859 1174 1867 1208
rect 1813 1052 1867 1174
<< ndiffc >>
rect 122 328 156 362
rect 219 328 253 362
rect 316 328 350 362
rect 510 328 544 362
rect 122 256 156 290
rect 122 188 156 222
rect 219 203 253 237
rect 316 256 350 290
rect 316 188 350 222
rect 412 212 446 246
rect 510 256 544 290
rect 510 188 544 222
rect 122 118 156 152
rect 316 118 350 152
rect 412 118 446 152
rect 510 118 544 152
rect 788 328 822 362
rect 885 328 919 362
rect 982 328 1016 362
rect 1176 328 1210 362
rect 788 256 822 290
rect 788 188 822 222
rect 885 203 919 237
rect 982 256 1016 290
rect 982 188 1016 222
rect 1079 212 1113 246
rect 1176 256 1210 290
rect 1176 188 1210 222
rect 788 118 822 152
rect 982 118 1016 152
rect 1079 118 1113 152
rect 1176 118 1210 152
rect 1454 328 1488 362
rect 1551 328 1585 362
rect 1648 328 1682 362
rect 1454 256 1488 290
rect 1454 188 1488 222
rect 1551 203 1585 237
rect 1648 256 1682 290
rect 1648 188 1682 222
rect 1745 212 1779 246
rect 1842 256 1876 290
rect 1842 188 1876 222
rect 1454 118 1488 152
rect 1648 118 1682 152
rect 1745 118 1779 152
rect 1842 118 1876 152
<< pdiffc >>
rect 141 1378 175 1412
rect 141 1310 175 1344
rect 141 1242 175 1276
rect 141 1174 175 1208
rect 141 1106 175 1140
rect 229 1378 263 1412
rect 229 1310 263 1344
rect 229 1242 263 1276
rect 229 1174 263 1208
rect 229 1106 263 1140
rect 317 1378 351 1412
rect 317 1310 351 1344
rect 317 1242 351 1276
rect 317 1174 351 1208
rect 405 1378 439 1412
rect 405 1310 439 1344
rect 405 1242 439 1276
rect 405 1174 439 1208
rect 493 1378 527 1412
rect 493 1310 527 1344
rect 493 1242 527 1276
rect 493 1174 527 1208
rect 493 1106 527 1140
rect 805 1378 839 1412
rect 805 1310 839 1344
rect 805 1242 839 1276
rect 805 1174 839 1208
rect 893 1310 927 1344
rect 893 1242 927 1276
rect 893 1174 927 1208
rect 893 1106 927 1140
rect 981 1378 1015 1412
rect 981 1310 1015 1344
rect 981 1242 1015 1276
rect 981 1174 1015 1208
rect 1069 1310 1103 1344
rect 1069 1242 1103 1276
rect 1069 1174 1103 1208
rect 1157 1378 1191 1412
rect 1157 1310 1191 1344
rect 1157 1242 1191 1276
rect 1157 1174 1191 1208
rect 1473 1378 1507 1412
rect 1473 1310 1507 1344
rect 1473 1242 1507 1276
rect 1473 1174 1507 1208
rect 1561 1310 1595 1344
rect 1561 1242 1595 1276
rect 1561 1174 1595 1208
rect 1561 1106 1595 1140
rect 1649 1378 1683 1412
rect 1649 1310 1683 1344
rect 1649 1242 1683 1276
rect 1649 1174 1683 1208
rect 1737 1310 1771 1344
rect 1737 1242 1771 1276
rect 1737 1174 1771 1208
rect 1737 1106 1771 1140
rect 1825 1378 1859 1412
rect 1825 1310 1859 1344
rect 1825 1242 1859 1276
rect 1825 1174 1859 1208
<< psubdiff >>
rect -31 547 2029 573
rect -31 513 -17 547
rect 17 513 649 547
rect 683 513 1315 547
rect 1349 513 1981 547
rect 2015 513 2029 547
rect -31 511 2029 513
rect -31 475 31 511
rect -31 441 -17 475
rect 17 441 31 475
rect -31 403 31 441
rect 635 475 697 511
rect 635 441 649 475
rect 683 441 697 475
rect -31 369 -17 403
rect 17 369 31 403
rect 635 403 697 441
rect -31 331 31 369
rect -31 297 -17 331
rect 17 297 31 331
rect -31 259 31 297
rect -31 225 -17 259
rect 17 225 31 259
rect -31 187 31 225
rect -31 153 -17 187
rect 17 153 31 187
rect -31 115 31 153
rect -31 81 -17 115
rect 17 81 31 115
rect 635 369 649 403
rect 683 369 697 403
rect 1301 475 1363 511
rect 1301 441 1315 475
rect 1349 441 1363 475
rect 1301 403 1363 441
rect 1967 475 2029 511
rect 1967 441 1981 475
rect 2015 441 2029 475
rect 635 331 697 369
rect 635 297 649 331
rect 683 297 697 331
rect 635 259 697 297
rect 635 225 649 259
rect 683 225 697 259
rect 635 187 697 225
rect 635 153 649 187
rect 683 153 697 187
rect 635 115 697 153
rect -31 48 31 81
rect 635 81 649 115
rect 683 81 697 115
rect 1301 369 1315 403
rect 1349 369 1363 403
rect 1967 403 2029 441
rect 1301 331 1363 369
rect 1301 297 1315 331
rect 1349 297 1363 331
rect 1301 259 1363 297
rect 1301 225 1315 259
rect 1349 225 1363 259
rect 1301 187 1363 225
rect 1301 153 1315 187
rect 1349 153 1363 187
rect 1301 115 1363 153
rect 635 48 697 81
rect 1301 81 1315 115
rect 1349 81 1363 115
rect 1967 369 1981 403
rect 2015 369 2029 403
rect 1967 331 2029 369
rect 1967 297 1981 331
rect 2015 297 2029 331
rect 1967 259 2029 297
rect 1967 225 1981 259
rect 2015 225 2029 259
rect 1967 187 2029 225
rect 1967 153 1981 187
rect 2015 153 2029 187
rect 1967 115 2029 153
rect 1301 48 1363 81
rect 1967 81 1981 115
rect 2015 81 2029 115
rect 1967 48 2029 81
rect -31 14 55 48
rect 89 14 127 48
rect 161 14 199 48
rect 233 14 271 48
rect 305 14 361 48
rect 395 14 433 48
rect 467 14 505 48
rect 539 14 577 48
rect 611 14 721 48
rect 755 14 793 48
rect 827 14 865 48
rect 899 14 937 48
rect 971 14 1027 48
rect 1061 14 1099 48
rect 1133 14 1171 48
rect 1205 14 1243 48
rect 1277 14 1387 48
rect 1421 14 1459 48
rect 1493 14 1531 48
rect 1565 14 1603 48
rect 1637 14 1693 48
rect 1727 14 1765 48
rect 1799 14 1837 48
rect 1871 14 1909 48
rect 1943 14 2029 48
rect -31 12 31 14
rect 635 12 697 14
rect 1301 12 1363 14
rect 1967 12 2029 14
<< nsubdiff >>
rect -31 1506 55 1540
rect 89 1506 127 1540
rect 161 1506 199 1540
rect 233 1506 271 1540
rect 305 1506 361 1540
rect 395 1506 433 1540
rect 467 1506 505 1540
rect 539 1506 577 1540
rect 611 1506 721 1540
rect 755 1506 793 1540
rect 827 1506 865 1540
rect 899 1506 937 1540
rect 971 1506 1027 1540
rect 1061 1506 1099 1540
rect 1133 1506 1171 1540
rect 1205 1506 1243 1540
rect 1277 1506 1387 1540
rect 1421 1506 1459 1540
rect 1493 1506 1531 1540
rect 1565 1506 1603 1540
rect 1637 1506 1693 1540
rect 1727 1506 1765 1540
rect 1799 1506 1837 1540
rect 1871 1506 1909 1540
rect 1943 1506 2029 1540
rect -31 1471 31 1506
rect -31 1437 -17 1471
rect 17 1437 31 1471
rect 635 1471 697 1506
rect -31 1399 31 1437
rect -31 1365 -17 1399
rect 17 1365 31 1399
rect -31 1327 31 1365
rect -31 1293 -17 1327
rect 17 1293 31 1327
rect -31 1255 31 1293
rect -31 1221 -17 1255
rect 17 1221 31 1255
rect -31 1183 31 1221
rect -31 1149 -17 1183
rect 17 1149 31 1183
rect -31 1111 31 1149
rect -31 1077 -17 1111
rect 17 1077 31 1111
rect -31 1039 31 1077
rect 635 1437 649 1471
rect 683 1437 697 1471
rect 1301 1471 1363 1506
rect 635 1399 697 1437
rect 635 1365 649 1399
rect 683 1365 697 1399
rect 635 1327 697 1365
rect 635 1293 649 1327
rect 683 1293 697 1327
rect 635 1255 697 1293
rect 635 1221 649 1255
rect 683 1221 697 1255
rect 635 1183 697 1221
rect 635 1149 649 1183
rect 683 1149 697 1183
rect 635 1111 697 1149
rect 635 1077 649 1111
rect 683 1077 697 1111
rect -31 1005 -17 1039
rect 17 1005 31 1039
rect -31 967 31 1005
rect -31 933 -17 967
rect 17 933 31 967
rect 635 1039 697 1077
rect 1301 1437 1315 1471
rect 1349 1437 1363 1471
rect 1967 1471 2029 1506
rect 1301 1399 1363 1437
rect 1301 1365 1315 1399
rect 1349 1365 1363 1399
rect 1301 1327 1363 1365
rect 1301 1293 1315 1327
rect 1349 1293 1363 1327
rect 1301 1255 1363 1293
rect 1301 1221 1315 1255
rect 1349 1221 1363 1255
rect 1301 1183 1363 1221
rect 1301 1149 1315 1183
rect 1349 1149 1363 1183
rect 1301 1111 1363 1149
rect 1301 1077 1315 1111
rect 1349 1077 1363 1111
rect 635 1005 649 1039
rect 683 1005 697 1039
rect 635 967 697 1005
rect -31 931 31 933
rect 635 933 649 967
rect 683 933 697 967
rect 1301 1039 1363 1077
rect 1967 1437 1981 1471
rect 2015 1437 2029 1471
rect 1967 1399 2029 1437
rect 1967 1365 1981 1399
rect 2015 1365 2029 1399
rect 1967 1327 2029 1365
rect 1967 1293 1981 1327
rect 2015 1293 2029 1327
rect 1967 1255 2029 1293
rect 1967 1221 1981 1255
rect 2015 1221 2029 1255
rect 1967 1183 2029 1221
rect 1967 1149 1981 1183
rect 2015 1149 2029 1183
rect 1967 1111 2029 1149
rect 1967 1077 1981 1111
rect 2015 1077 2029 1111
rect 1301 1005 1315 1039
rect 1349 1005 1363 1039
rect 1301 967 1363 1005
rect 635 931 697 933
rect 1301 933 1315 967
rect 1349 933 1363 967
rect 1967 1039 2029 1077
rect 1967 1005 1981 1039
rect 2015 1005 2029 1039
rect 1967 967 2029 1005
rect 1301 931 1363 933
rect 1967 933 1981 967
rect 2015 933 2029 967
rect 1967 931 2029 933
rect -31 869 2029 931
<< psubdiffcont >>
rect -17 513 17 547
rect 649 513 683 547
rect 1315 513 1349 547
rect 1981 513 2015 547
rect -17 441 17 475
rect 649 441 683 475
rect -17 369 17 403
rect -17 297 17 331
rect -17 225 17 259
rect -17 153 17 187
rect -17 81 17 115
rect 649 369 683 403
rect 1315 441 1349 475
rect 1981 441 2015 475
rect 649 297 683 331
rect 649 225 683 259
rect 649 153 683 187
rect 649 81 683 115
rect 1315 369 1349 403
rect 1315 297 1349 331
rect 1315 225 1349 259
rect 1315 153 1349 187
rect 1315 81 1349 115
rect 1981 369 2015 403
rect 1981 297 2015 331
rect 1981 225 2015 259
rect 1981 153 2015 187
rect 1981 81 2015 115
rect 55 14 89 48
rect 127 14 161 48
rect 199 14 233 48
rect 271 14 305 48
rect 361 14 395 48
rect 433 14 467 48
rect 505 14 539 48
rect 577 14 611 48
rect 721 14 755 48
rect 793 14 827 48
rect 865 14 899 48
rect 937 14 971 48
rect 1027 14 1061 48
rect 1099 14 1133 48
rect 1171 14 1205 48
rect 1243 14 1277 48
rect 1387 14 1421 48
rect 1459 14 1493 48
rect 1531 14 1565 48
rect 1603 14 1637 48
rect 1693 14 1727 48
rect 1765 14 1799 48
rect 1837 14 1871 48
rect 1909 14 1943 48
<< nsubdiffcont >>
rect 55 1506 89 1540
rect 127 1506 161 1540
rect 199 1506 233 1540
rect 271 1506 305 1540
rect 361 1506 395 1540
rect 433 1506 467 1540
rect 505 1506 539 1540
rect 577 1506 611 1540
rect 721 1506 755 1540
rect 793 1506 827 1540
rect 865 1506 899 1540
rect 937 1506 971 1540
rect 1027 1506 1061 1540
rect 1099 1506 1133 1540
rect 1171 1506 1205 1540
rect 1243 1506 1277 1540
rect 1387 1506 1421 1540
rect 1459 1506 1493 1540
rect 1531 1506 1565 1540
rect 1603 1506 1637 1540
rect 1693 1506 1727 1540
rect 1765 1506 1799 1540
rect 1837 1506 1871 1540
rect 1909 1506 1943 1540
rect -17 1437 17 1471
rect -17 1365 17 1399
rect -17 1293 17 1327
rect -17 1221 17 1255
rect -17 1149 17 1183
rect -17 1077 17 1111
rect 649 1437 683 1471
rect 649 1365 683 1399
rect 649 1293 683 1327
rect 649 1221 683 1255
rect 649 1149 683 1183
rect 649 1077 683 1111
rect -17 1005 17 1039
rect -17 933 17 967
rect 1315 1437 1349 1471
rect 1315 1365 1349 1399
rect 1315 1293 1349 1327
rect 1315 1221 1349 1255
rect 1315 1149 1349 1183
rect 1315 1077 1349 1111
rect 649 1005 683 1039
rect 649 933 683 967
rect 1981 1437 2015 1471
rect 1981 1365 2015 1399
rect 1981 1293 2015 1327
rect 1981 1221 2015 1255
rect 1981 1149 2015 1183
rect 1981 1077 2015 1111
rect 1315 1005 1349 1039
rect 1315 933 1349 967
rect 1981 1005 2015 1039
rect 1981 933 2015 967
<< poly >>
rect 187 1452 217 1478
rect 275 1452 305 1478
rect 363 1452 393 1478
rect 451 1452 481 1478
rect 851 1452 881 1478
rect 939 1452 969 1478
rect 1027 1452 1057 1478
rect 1115 1452 1145 1478
rect 187 1021 217 1052
rect 275 1021 305 1052
rect 363 1021 393 1052
rect 451 1021 481 1052
rect 121 1005 305 1021
rect 121 971 131 1005
rect 165 991 305 1005
rect 351 1005 481 1021
rect 165 971 175 991
rect 121 955 175 971
rect 351 971 361 1005
rect 395 991 481 1005
rect 1519 1452 1549 1478
rect 1607 1452 1637 1478
rect 1695 1452 1725 1478
rect 1783 1452 1813 1478
rect 395 971 405 991
rect 351 955 405 971
rect 851 1021 881 1052
rect 939 1021 969 1052
rect 851 1005 969 1021
rect 851 991 871 1005
rect 861 971 871 991
rect 905 991 969 1005
rect 1027 1021 1057 1052
rect 1115 1021 1145 1052
rect 1027 1005 1211 1021
rect 1027 991 1167 1005
rect 905 971 915 991
rect 861 955 915 971
rect 1157 971 1167 991
rect 1201 971 1211 1005
rect 1157 955 1211 971
rect 1519 1021 1549 1052
rect 1607 1021 1637 1052
rect 1695 1021 1725 1052
rect 1783 1021 1813 1052
rect 1453 1005 1637 1021
rect 1453 971 1463 1005
rect 1497 991 1637 1005
rect 1679 1005 1813 1021
rect 1497 971 1507 991
rect 1453 955 1507 971
rect 1679 971 1689 1005
rect 1723 991 1813 1005
rect 1723 971 1733 991
rect 1679 955 1733 971
rect 121 462 175 478
rect 121 428 131 462
rect 165 442 175 462
rect 343 462 397 478
rect 165 428 198 442
rect 121 412 198 428
rect 343 428 353 462
rect 387 428 397 462
rect 343 412 397 428
rect 861 462 915 478
rect 861 442 871 462
rect 168 378 198 412
rect 362 378 392 412
rect 834 428 871 442
rect 905 428 915 462
rect 1157 462 1211 478
rect 1157 442 1167 462
rect 834 412 915 428
rect 1134 428 1167 442
rect 1201 428 1211 462
rect 1134 412 1211 428
rect 834 378 864 412
rect 1134 378 1164 412
rect 1453 462 1507 478
rect 1453 428 1463 462
rect 1497 442 1507 462
rect 1675 462 1729 478
rect 1497 428 1530 442
rect 1453 412 1530 428
rect 1675 428 1685 462
rect 1719 428 1729 462
rect 1675 412 1729 428
rect 1500 378 1530 412
rect 1694 378 1724 412
<< polycont >>
rect 131 971 165 1005
rect 361 971 395 1005
rect 871 971 905 1005
rect 1167 971 1201 1005
rect 1463 971 1497 1005
rect 1689 971 1723 1005
rect 131 428 165 462
rect 353 428 387 462
rect 871 428 905 462
rect 1167 428 1201 462
rect 1463 428 1497 462
rect 1685 428 1719 462
<< locali >>
rect -31 1540 2029 1555
rect -31 1506 55 1540
rect 89 1506 127 1540
rect 161 1506 199 1540
rect 233 1506 271 1540
rect 305 1506 361 1540
rect 395 1506 433 1540
rect 467 1506 505 1540
rect 539 1506 577 1540
rect 611 1506 721 1540
rect 755 1506 793 1540
rect 827 1506 865 1540
rect 899 1506 937 1540
rect 971 1506 1027 1540
rect 1061 1506 1099 1540
rect 1133 1506 1171 1540
rect 1205 1506 1243 1540
rect 1277 1506 1387 1540
rect 1421 1506 1459 1540
rect 1493 1506 1531 1540
rect 1565 1506 1603 1540
rect 1637 1506 1693 1540
rect 1727 1506 1765 1540
rect 1799 1506 1837 1540
rect 1871 1506 1909 1540
rect 1943 1506 2029 1540
rect -31 1493 2029 1506
rect -31 1471 31 1493
rect -31 1437 -17 1471
rect 17 1437 31 1471
rect -31 1399 31 1437
rect -31 1365 -17 1399
rect 17 1365 31 1399
rect -31 1327 31 1365
rect -31 1293 -17 1327
rect 17 1293 31 1327
rect -31 1255 31 1293
rect -31 1221 -17 1255
rect 17 1221 31 1255
rect -31 1183 31 1221
rect -31 1149 -17 1183
rect 17 1149 31 1183
rect -31 1111 31 1149
rect -31 1077 -17 1111
rect 17 1077 31 1111
rect -31 1039 31 1077
rect 141 1412 175 1493
rect 141 1344 175 1378
rect 141 1276 175 1310
rect 141 1208 175 1242
rect 141 1140 175 1174
rect 141 1072 175 1106
rect 229 1412 265 1446
rect 317 1412 351 1493
rect 229 1344 263 1378
rect 229 1276 263 1310
rect 229 1208 263 1242
rect 229 1140 263 1174
rect 317 1344 351 1378
rect 317 1276 351 1310
rect 317 1208 351 1242
rect 317 1158 351 1174
rect 405 1412 439 1446
rect 405 1344 439 1378
rect 405 1276 439 1310
rect 405 1208 439 1242
rect 405 1106 439 1174
rect 229 1072 405 1106
rect 493 1412 527 1493
rect 493 1344 527 1378
rect 493 1276 527 1310
rect 493 1208 527 1242
rect 493 1140 527 1174
rect 493 1072 527 1106
rect 635 1471 697 1493
rect 635 1437 649 1471
rect 683 1437 697 1471
rect 1301 1471 1363 1493
rect 635 1399 697 1437
rect 635 1365 649 1399
rect 683 1365 697 1399
rect 635 1327 697 1365
rect 635 1293 649 1327
rect 683 1293 697 1327
rect 635 1255 697 1293
rect 635 1221 649 1255
rect 683 1221 697 1255
rect 635 1183 697 1221
rect 635 1149 649 1183
rect 683 1149 697 1183
rect 635 1111 697 1149
rect 635 1077 649 1111
rect 683 1077 697 1111
rect 405 1056 439 1072
rect -31 1005 -17 1039
rect 17 1005 31 1039
rect 635 1039 697 1077
rect 805 1412 1191 1446
rect 805 1344 839 1378
rect 805 1276 839 1310
rect 805 1208 839 1242
rect 805 1106 839 1174
rect 893 1344 927 1360
rect 893 1276 927 1310
rect 893 1208 927 1242
rect 893 1140 927 1174
rect 981 1344 1015 1378
rect 981 1276 1015 1310
rect 981 1208 1015 1242
rect 981 1158 1015 1174
rect 1069 1344 1103 1360
rect 1069 1276 1103 1310
rect 1069 1208 1103 1242
rect 1069 1106 1103 1174
rect 1157 1344 1191 1378
rect 1157 1276 1191 1310
rect 1157 1208 1191 1242
rect 1157 1122 1191 1174
rect 1301 1437 1315 1471
rect 1349 1437 1363 1471
rect 1967 1471 2029 1493
rect 1301 1399 1363 1437
rect 1301 1365 1315 1399
rect 1349 1365 1363 1399
rect 1301 1327 1363 1365
rect 1301 1293 1315 1327
rect 1349 1293 1363 1327
rect 1301 1255 1363 1293
rect 1301 1221 1315 1255
rect 1349 1221 1363 1255
rect 1301 1183 1363 1221
rect 1301 1149 1315 1183
rect 1349 1149 1363 1183
rect 893 1072 1069 1106
rect 805 1056 839 1072
rect 1069 1056 1103 1072
rect 1301 1111 1363 1149
rect 1301 1077 1315 1111
rect 1349 1077 1363 1111
rect -31 967 31 1005
rect -31 933 -17 967
rect 17 933 31 967
rect -31 869 31 933
rect 131 1005 165 1021
rect 361 1005 395 1021
rect 131 906 165 971
rect -31 547 31 573
rect -31 513 -17 547
rect 17 513 31 547
rect -31 475 31 513
rect -31 441 -17 475
rect 17 441 31 475
rect -31 403 31 441
rect 131 462 165 872
rect 353 971 361 989
rect 353 955 395 971
rect 635 1005 649 1039
rect 683 1005 697 1039
rect 1301 1039 1363 1077
rect 1473 1412 1859 1446
rect 1473 1344 1507 1378
rect 1473 1276 1507 1310
rect 1473 1208 1507 1242
rect 1473 1106 1507 1174
rect 1561 1344 1595 1360
rect 1561 1276 1595 1310
rect 1561 1208 1595 1242
rect 1561 1140 1595 1174
rect 1649 1344 1683 1378
rect 1649 1276 1683 1310
rect 1649 1208 1683 1242
rect 1649 1158 1683 1174
rect 1737 1344 1771 1360
rect 1737 1276 1771 1310
rect 1737 1208 1771 1242
rect 1737 1140 1771 1174
rect 1825 1344 1859 1378
rect 1825 1276 1859 1310
rect 1825 1208 1859 1242
rect 1825 1158 1859 1174
rect 1967 1437 1981 1471
rect 2015 1437 2029 1471
rect 1967 1399 2029 1437
rect 1967 1365 1981 1399
rect 2015 1365 2029 1399
rect 1967 1327 2029 1365
rect 1967 1293 1981 1327
rect 2015 1293 2029 1327
rect 1967 1255 2029 1293
rect 1967 1221 1981 1255
rect 2015 1221 2029 1255
rect 1967 1183 2029 1221
rect 1967 1149 1981 1183
rect 2015 1149 2029 1183
rect 1967 1111 2029 1149
rect 1561 1072 1867 1106
rect 1473 1056 1507 1072
rect 635 967 697 1005
rect 353 832 387 955
rect 635 933 649 967
rect 683 933 697 967
rect 635 869 697 933
rect 871 1005 905 1021
rect 353 782 387 798
rect 871 832 905 971
rect 871 782 905 798
rect 1167 1005 1201 1021
rect 1167 832 1201 971
rect 1301 1005 1315 1039
rect 1349 1005 1363 1039
rect 1301 967 1363 1005
rect 1301 933 1315 967
rect 1349 933 1363 967
rect 1301 869 1363 933
rect 1463 1005 1497 1021
rect 1167 782 1201 798
rect 1463 832 1497 971
rect 1463 782 1497 798
rect 1685 1005 1723 1021
rect 1685 971 1689 1005
rect 1685 955 1723 971
rect 1685 906 1719 955
rect 131 412 165 428
rect 353 536 387 552
rect 353 462 387 502
rect 353 412 387 428
rect 635 547 697 573
rect 635 513 649 547
rect 683 513 697 547
rect 635 475 697 513
rect 635 441 649 475
rect 683 441 697 475
rect -31 369 -17 403
rect 17 369 31 403
rect 635 403 697 441
rect 871 536 905 552
rect 871 462 905 502
rect 871 412 905 428
rect 1167 536 1201 552
rect 1167 462 1201 502
rect 1167 412 1201 428
rect 1301 547 1363 573
rect 1301 513 1315 547
rect 1349 513 1363 547
rect 1301 475 1363 513
rect 1301 441 1315 475
rect 1349 441 1363 475
rect -31 331 31 369
rect -31 297 -17 331
rect 17 297 31 331
rect -31 259 31 297
rect -31 225 -17 259
rect 17 225 31 259
rect -31 187 31 225
rect -31 153 -17 187
rect 17 153 31 187
rect -31 115 31 153
rect -31 81 -17 115
rect 17 81 31 115
rect 122 362 156 378
rect 316 362 350 378
rect 156 328 219 362
rect 253 328 316 362
rect 122 290 156 328
rect 122 222 156 256
rect 316 290 350 328
rect 510 362 544 378
rect 413 282 447 298
rect 122 152 156 188
rect 122 102 156 118
rect 219 237 253 253
rect -31 63 31 81
rect 219 63 253 203
rect 316 222 350 256
rect 412 248 413 263
rect 412 246 447 248
rect 446 232 447 246
rect 510 290 544 328
rect 412 196 446 212
rect 510 222 544 256
rect 316 152 350 188
rect 510 152 544 188
rect 350 118 412 152
rect 446 118 510 152
rect 316 102 350 118
rect 510 102 544 118
rect 635 369 649 403
rect 683 369 697 403
rect 1301 403 1363 441
rect 1463 536 1497 552
rect 1463 462 1497 502
rect 1463 412 1497 428
rect 1685 462 1719 872
rect 1685 412 1719 428
rect 1833 831 1867 1072
rect 1967 1077 1981 1111
rect 2015 1077 2029 1111
rect 1967 1039 2029 1077
rect 1967 1005 1981 1039
rect 2015 1005 2029 1039
rect 1967 967 2029 1005
rect 1967 933 1981 967
rect 2015 933 2029 967
rect 1967 869 2029 933
rect 635 331 697 369
rect 635 297 649 331
rect 683 297 697 331
rect 635 259 697 297
rect 635 225 649 259
rect 683 225 697 259
rect 635 187 697 225
rect 635 153 649 187
rect 683 153 697 187
rect 635 115 697 153
rect 635 81 649 115
rect 683 81 697 115
rect 788 362 822 378
rect 982 362 1016 378
rect 822 328 885 362
rect 919 328 982 362
rect 788 290 822 328
rect 788 222 822 256
rect 982 290 1016 328
rect 1176 362 1210 378
rect 788 152 822 188
rect 788 102 822 118
rect 885 237 919 253
rect 635 63 697 81
rect 885 63 919 203
rect 982 222 1016 256
rect 1079 282 1113 298
rect 1079 246 1113 248
rect 1079 196 1113 212
rect 1176 290 1210 328
rect 1176 222 1210 256
rect 982 152 1016 188
rect 1176 152 1210 188
rect 1016 118 1079 152
rect 1113 118 1176 152
rect 982 102 1016 118
rect 1176 102 1210 118
rect 1301 369 1315 403
rect 1349 369 1363 403
rect 1301 331 1363 369
rect 1301 297 1315 331
rect 1349 297 1363 331
rect 1301 259 1363 297
rect 1301 225 1315 259
rect 1349 225 1363 259
rect 1301 187 1363 225
rect 1301 153 1315 187
rect 1349 153 1363 187
rect 1301 115 1363 153
rect 1301 81 1315 115
rect 1349 81 1363 115
rect 1454 362 1488 378
rect 1648 362 1682 378
rect 1833 375 1867 797
rect 1488 328 1551 362
rect 1585 328 1648 362
rect 1454 290 1488 328
rect 1454 222 1488 256
rect 1648 290 1682 328
rect 1454 152 1488 188
rect 1454 102 1488 118
rect 1551 237 1585 253
rect 1301 63 1363 81
rect 1551 63 1585 203
rect 1648 222 1682 256
rect 1745 341 1867 375
rect 1967 547 2029 573
rect 1967 513 1981 547
rect 2015 513 2029 547
rect 1967 475 2029 513
rect 1967 441 1981 475
rect 2015 441 2029 475
rect 1967 403 2029 441
rect 1967 369 1981 403
rect 2015 369 2029 403
rect 1745 282 1779 341
rect 1967 331 2029 369
rect 1745 246 1779 248
rect 1745 196 1779 212
rect 1842 290 1876 307
rect 1842 222 1876 256
rect 1648 152 1682 188
rect 1842 152 1876 188
rect 1682 118 1745 152
rect 1779 118 1842 152
rect 1648 102 1682 118
rect 1842 102 1876 118
rect 1967 297 1981 331
rect 2015 297 2029 331
rect 1967 259 2029 297
rect 1967 225 1981 259
rect 2015 225 2029 259
rect 1967 187 2029 225
rect 1967 153 1981 187
rect 2015 153 2029 187
rect 1967 115 2029 153
rect 1967 81 1981 115
rect 2015 81 2029 115
rect 1967 63 2029 81
rect -31 48 1079 63
rect 1113 48 2029 63
rect -31 14 55 48
rect 89 14 127 48
rect 161 14 199 48
rect 233 14 271 48
rect 305 14 361 48
rect 395 14 433 48
rect 467 14 505 48
rect 539 14 577 48
rect 611 14 721 48
rect 755 14 793 48
rect 827 14 865 48
rect 899 14 937 48
rect 971 14 1027 48
rect 1061 14 1099 48
rect 1133 14 1171 48
rect 1205 14 1243 48
rect 1277 14 1387 48
rect 1421 14 1459 48
rect 1493 14 1531 48
rect 1565 14 1603 48
rect 1637 14 1693 48
rect 1727 14 1765 48
rect 1799 14 1837 48
rect 1871 14 1909 48
rect 1943 14 2029 48
rect -31 1 2029 14
<< viali >>
rect 55 1506 89 1540
rect 127 1506 161 1540
rect 199 1506 233 1540
rect 271 1506 305 1540
rect 361 1506 395 1540
rect 433 1506 467 1540
rect 505 1506 539 1540
rect 577 1506 611 1540
rect 721 1506 755 1540
rect 793 1506 827 1540
rect 865 1506 899 1540
rect 937 1506 971 1540
rect 1027 1506 1061 1540
rect 1099 1506 1133 1540
rect 1171 1506 1205 1540
rect 1243 1506 1277 1540
rect 1387 1506 1421 1540
rect 1459 1506 1493 1540
rect 1531 1506 1565 1540
rect 1603 1506 1637 1540
rect 1693 1506 1727 1540
rect 1765 1506 1799 1540
rect 1837 1506 1871 1540
rect 1909 1506 1943 1540
rect 405 1072 439 1106
rect 805 1072 839 1106
rect 1069 1072 1103 1106
rect 131 872 165 906
rect 1473 1072 1507 1106
rect 353 798 387 832
rect 871 798 905 832
rect 1167 798 1201 832
rect 1463 798 1497 832
rect 1685 872 1719 906
rect 353 502 387 536
rect 871 502 905 536
rect 1167 502 1201 536
rect 413 248 447 282
rect 1463 502 1497 536
rect 1833 797 1867 831
rect 1079 248 1113 282
rect 1745 248 1779 282
rect 55 14 89 48
rect 127 14 161 48
rect 199 14 233 48
rect 271 14 305 48
rect 361 14 395 48
rect 433 14 467 48
rect 505 14 539 48
rect 577 14 611 48
rect 721 14 755 48
rect 793 14 827 48
rect 865 14 899 48
rect 937 14 971 48
rect 1027 14 1061 48
rect 1099 14 1133 48
rect 1171 14 1205 48
rect 1243 14 1277 48
rect 1387 14 1421 48
rect 1459 14 1493 48
rect 1531 14 1565 48
rect 1603 14 1637 48
rect 1693 14 1727 48
rect 1765 14 1799 48
rect 1837 14 1871 48
rect 1909 14 1943 48
<< metal1 >>
rect -31 1540 2029 1555
rect -31 1506 55 1540
rect 89 1506 127 1540
rect 161 1506 199 1540
rect 233 1506 271 1540
rect 305 1506 361 1540
rect 395 1506 433 1540
rect 467 1506 505 1540
rect 539 1506 577 1540
rect 611 1506 721 1540
rect 755 1506 793 1540
rect 827 1506 865 1540
rect 899 1506 937 1540
rect 971 1506 1027 1540
rect 1061 1506 1099 1540
rect 1133 1506 1171 1540
rect 1205 1506 1243 1540
rect 1277 1506 1387 1540
rect 1421 1506 1459 1540
rect 1493 1506 1531 1540
rect 1565 1506 1603 1540
rect 1637 1506 1693 1540
rect 1727 1506 1765 1540
rect 1799 1506 1837 1540
rect 1871 1506 1909 1540
rect 1943 1506 2029 1540
rect -31 1493 2029 1506
rect 399 1106 445 1112
rect 799 1106 845 1112
rect 1063 1106 1109 1112
rect 1467 1106 1513 1112
rect 393 1072 405 1106
rect 439 1072 805 1106
rect 839 1072 851 1106
rect 1057 1072 1069 1106
rect 1103 1072 1473 1106
rect 1507 1072 1519 1106
rect 399 1066 445 1072
rect 799 1066 845 1072
rect 1063 1066 1109 1072
rect 1467 1066 1513 1072
rect 125 906 171 912
rect 1679 906 1725 912
rect 119 872 131 906
rect 165 872 1685 906
rect 1719 872 1731 906
rect 125 866 171 872
rect 1679 866 1725 872
rect 347 832 393 838
rect 865 832 911 838
rect 1161 832 1207 838
rect 1457 832 1503 838
rect 341 798 353 832
rect 387 798 871 832
rect 905 798 917 832
rect 1155 798 1167 832
rect 1201 798 1463 832
rect 1497 798 1509 832
rect 1827 831 1873 837
rect 347 792 393 798
rect 865 792 911 798
rect 1161 792 1207 798
rect 1457 792 1503 798
rect 1821 797 1833 831
rect 1867 797 1903 831
rect 1827 791 1873 797
rect 347 536 393 542
rect 865 536 911 542
rect 1161 536 1207 542
rect 1457 536 1503 542
rect 341 502 353 536
rect 387 502 871 536
rect 905 502 917 536
rect 1155 502 1167 536
rect 1201 502 1463 536
rect 1497 502 1509 536
rect 347 496 393 502
rect 865 496 911 502
rect 1161 496 1207 502
rect 1457 496 1503 502
rect 407 282 453 288
rect 1073 282 1119 288
rect 1739 282 1785 288
rect 401 248 413 282
rect 447 248 1079 282
rect 1113 248 1745 282
rect 1779 248 1791 282
rect 407 242 453 248
rect 1073 242 1119 248
rect 1739 242 1785 248
rect -31 48 2029 63
rect -31 14 55 48
rect 89 14 127 48
rect 161 14 199 48
rect 233 14 271 48
rect 305 14 361 48
rect 395 14 433 48
rect 467 14 505 48
rect 539 14 577 48
rect 611 14 721 48
rect 755 14 793 48
rect 827 14 865 48
rect 899 14 937 48
rect 971 14 1027 48
rect 1061 14 1099 48
rect 1133 14 1171 48
rect 1205 14 1243 48
rect 1277 14 1387 48
rect 1421 14 1459 48
rect 1493 14 1531 48
rect 1565 14 1603 48
rect 1637 14 1693 48
rect 1727 14 1765 48
rect 1799 14 1837 48
rect 1871 14 1909 48
rect 1943 14 2029 48
rect -31 1 2029 14
<< labels >>
rlabel metal1 1833 797 1867 831 1 YN
port 1 n
rlabel metal1 1167 797 1201 831 1 C
port 2 n
rlabel metal1 353 797 387 831 1 B
port 3 n
rlabel metal1 131 871 165 905 1 A
port 4 n
rlabel metal1 55 13 89 47 1 VSS
port 5 n
rlabel metal1 55 1505 89 1539 1 VDD
port 6 n
<< end >>
