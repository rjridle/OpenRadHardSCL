magic
tech sky130A
magscale 1 2
timestamp 1648232089
<< nwell >>
rect 84 1554 1100 1575
rect 84 1492 1153 1554
rect 84 1487 1100 1492
rect 84 1421 878 1487
rect 84 1408 316 1421
rect 317 1408 878 1421
rect 84 1376 878 1408
rect 84 1358 526 1376
rect 527 1358 878 1376
rect 84 1022 878 1358
rect 1036 1022 1100 1487
rect 84 930 1100 1022
rect 84 903 1154 930
rect 83 868 1154 903
rect 83 832 1100 868
<< pdiffc >>
rect 147 1377 181 1411
rect 235 1377 269 1411
rect 323 1377 357 1411
rect 411 1377 445 1413
rect 499 1377 533 1411
rect 675 1377 709 1411
rect 783 1377 817 1411
rect 959 1377 993 1411
rect 235 1105 269 1139
rect 411 1105 445 1139
<< psubdiff >>
rect 31 510 1153 572
rect 31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 343 47
rect 377 13 415 47
rect 449 13 487 47
rect 521 13 585 47
rect 619 13 663 47
rect 697 13 735 47
rect 769 13 807 47
rect 841 13 879 47
rect 913 13 951 47
rect 985 13 1023 47
rect 1057 13 1095 47
rect 1129 13 1153 47
<< nsubdiff >>
rect 31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 343 1539
rect 377 1505 415 1539
rect 449 1505 487 1539
rect 521 1505 585 1539
rect 619 1505 663 1539
rect 697 1505 735 1539
rect 769 1505 807 1539
rect 841 1505 879 1539
rect 913 1505 951 1539
rect 985 1505 1023 1539
rect 1057 1505 1095 1539
rect 1129 1505 1153 1539
rect 31 868 1154 930
<< psubdiffcont >>
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 343 13 377 47
rect 415 13 449 47
rect 487 13 521 47
rect 585 13 619 47
rect 663 13 697 47
rect 735 13 769 47
rect 807 13 841 47
rect 879 13 913 47
rect 951 13 985 47
rect 1023 13 1057 47
rect 1095 13 1129 47
<< nsubdiffcont >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 343 1505 377 1539
rect 415 1505 449 1539
rect 487 1505 521 1539
rect 585 1505 619 1539
rect 663 1505 697 1539
rect 735 1505 769 1539
rect 807 1505 841 1539
rect 879 1505 913 1539
rect 951 1505 985 1539
rect 1023 1505 1057 1539
rect 1095 1505 1129 1539
<< poly >>
rect 164 411 206 441
rect 164 403 194 411
rect 358 410 388 434
rect 662 410 692 444
rect 856 403 886 444
<< locali >>
rect 31 1539 1153 1554
rect 31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 343 1539
rect 377 1505 415 1539
rect 449 1505 487 1539
rect 521 1505 585 1539
rect 619 1505 663 1539
rect 697 1505 735 1539
rect 769 1505 807 1539
rect 841 1505 879 1539
rect 913 1505 951 1539
rect 985 1505 1023 1539
rect 1057 1505 1095 1539
rect 1129 1505 1153 1539
rect 31 1492 1153 1505
rect 147 1411 181 1492
rect 147 1343 181 1377
rect 235 1411 269 1445
rect 235 1343 269 1377
rect 323 1411 357 1492
rect 323 1343 357 1377
rect 411 1413 445 1429
rect 411 1343 445 1377
rect 499 1411 533 1492
rect 499 1359 533 1377
rect 675 1411 709 1492
rect 675 1343 709 1377
rect 783 1411 993 1445
rect 783 1343 817 1377
rect 959 1343 993 1377
rect 235 1139 269 1158
rect 235 1071 269 1105
rect 411 1139 445 1173
rect 587 1105 621 1163
rect 783 1105 817 1157
rect 411 1071 817 1105
rect 205 461 239 954
rect 353 469 387 988
rect 649 477 683 958
rect 353 461 357 469
rect 409 339 616 373
rect 409 261 443 339
rect 723 213 757 492
rect 871 462 905 970
rect 215 62 249 195
rect 907 62 941 186
rect 31 47 1153 62
rect 31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 343 47
rect 377 13 415 47
rect 449 13 487 47
rect 521 13 585 47
rect 619 13 663 47
rect 697 13 735 47
rect 769 13 807 47
rect 841 13 879 47
rect 913 13 951 47
rect 985 13 1023 47
rect 1057 13 1095 47
rect 1129 13 1153 47
rect 31 0 1153 13
<< viali >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 343 1505 377 1539
rect 415 1505 449 1539
rect 487 1505 521 1539
rect 585 1505 619 1539
rect 663 1505 697 1539
rect 735 1505 769 1539
rect 807 1505 841 1539
rect 879 1505 913 1539
rect 951 1505 985 1539
rect 1023 1505 1057 1539
rect 1095 1505 1129 1539
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 343 13 377 47
rect 415 13 449 47
rect 487 13 521 47
rect 585 13 619 47
rect 663 13 697 47
rect 735 13 769 47
rect 807 13 841 47
rect 879 13 913 47
rect 951 13 985 47
rect 1023 13 1057 47
rect 1095 13 1129 47
<< metal1 >>
rect 31 1539 1153 1554
rect 31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 343 1539
rect 377 1505 415 1539
rect 449 1505 487 1539
rect 521 1505 585 1539
rect 619 1505 663 1539
rect 697 1505 735 1539
rect 769 1505 807 1539
rect 841 1505 879 1539
rect 913 1505 951 1539
rect 985 1505 1023 1539
rect 1057 1505 1095 1539
rect 1129 1505 1153 1539
rect 31 1492 1153 1505
rect 759 501 1284 535
rect 31 47 1153 62
rect 31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 343 47
rect 377 13 415 47
rect 449 13 487 47
rect 521 13 585 47
rect 619 13 663 47
rect 697 13 735 47
rect 769 13 807 47
rect 841 13 879 47
rect 913 13 951 47
rect 985 13 1023 47
rect 1057 13 1095 47
rect 1129 13 1153 47
rect 31 0 1153 13
use diff_ring_side  diff_ring_side_1
timestamp 1648063806
transform 1 0 0 0 1 0
box -84 0 84 1575
use nmos_bottom  nmos_bottom_0
timestamp 1648062456
transform -1 0 356 0 1 101
box 0 0 248 302
use pmos2_1  pmos2_1_0
timestamp 1647326732
transform 1 0 49 0 1 1450
box 52 -460 352 37
use poly_li1_contact  poly_li1_contact_0
timestamp 1648060378
transform 0 1 223 -1 0 988
box -32 -28 34 26
use poly_li1_contact  poly_li1_contact_1
timestamp 1648060378
transform 0 1 223 -1 0 445
box -32 -28 34 26
use pmos2_1  pmos2_1_3
timestamp 1647326732
transform 1 0 401 0 1 1450
box 52 -460 352 37
use nmos_top_trim1  nmos_top_trim1_0
timestamp 1648061897
transform -1 0 550 0 1 101
box 0 0 248 309
use poly_li1_contact  poly_li1_contact_3
timestamp 1648060378
transform 0 1 387 -1 0 988
box -32 -28 34 26
use pmos2_1  pmos2_1_1
timestamp 1647326732
transform 1 0 225 0 1 1450
box 52 -460 352 37
use poly_li1_contact  poly_li1_contact_2
timestamp 1648060378
transform 0 -1 369 1 0 443
box -32 -28 34 26
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform -1 0 740 0 -1 518
box -53 -33 29 33
use poly_li1_contact  poly_li1_contact_6
timestamp 1648060378
transform 0 1 667 -1 0 988
box -32 -28 34 26
use poly_li1_contact  poly_li1_contact_7
timestamp 1648060378
transform 0 -1 665 1 0 443
box -32 -28 34 26
use pmos2_1  pmos2_1_2
timestamp 1647326732
transform 1 0 685 0 1 1450
box 52 -460 352 37
use poly_li1_contact  poly_li1_contact_4
timestamp 1648060378
transform 0 1 889 -1 0 988
box -32 -28 34 26
use poly_li1_contact  poly_li1_contact_5
timestamp 1648060378
transform 0 -1 887 1 0 443
box -32 -28 34 26
use nmos_top_trim1  nmos_top_trim1_1
timestamp 1648061897
transform -1 0 854 0 1 101
box 0 0 248 309
use nmos_bottom  nmos_bottom_1
timestamp 1648062456
transform -1 0 1048 0 1 101
box 0 0 248 302
use li1_M1_contact  li1_M1_contact_2
timestamp 1648061256
transform 1 0 1332 0 1 518
box -53 -33 29 33
use invx1_pcell  invx1_pcell_0
timestamp 1648064504
transform 1 0 1184 0 1 0
box -84 0 528 1575
<< labels >>
rlabel space 205 461 239 970 1 C
port 1 n
rlabel space 353 461 387 988 1 B
port 2 n
rlabel space 871 461 905 970 1 A
port 3 n
rlabel space 649 461 683 970 1 D
port 4 n
rlabel space 1463 427 1497 979 1 Y
port 5 n
<< end >>
