magic
tech sky130
magscale 1 2
timestamp 1651261136
<< nwell >>
rect 55 1505 89 1539
<< pwell >>
rect 55 13 89 47
<< psubdiffcont >>
rect 55 13 89 47
<< nsubdiffcont >>
rect 55 1505 89 1539
<< viali >>
rect 55 1505 89 1539
rect 55 13 89 47
<< metal1 >>
rect -31 1539 17569 1554
rect -31 1505 55 1539
rect 89 1505 17569 1539
rect -31 1492 17569 1505
rect 427 945 461 979
rect 2906 945 13416 979
rect 4386 797 4727 831
rect 9565 797 9877 831
rect 14745 797 15075 831
rect 17373 797 17407 831
rect 14595 723 15884 757
rect 9383 649 15669 683
rect 4207 575 16706 609
rect 1611 501 1645 535
rect 3891 501 14375 535
rect 1389 427 1423 461
rect 1425 427 11807 461
rect -31 47 17569 62
rect -31 13 55 47
rect 89 13 17569 47
rect -31 0 17569 13
use dffrnx1_pcell  dffrnx1_pcell_1 pcells
timestamp 1651259642
transform 1 0 5180 0 1 0
box -84 0 5264 1575
use dffrnx1_pcell  dffrnx1_pcell_0
timestamp 1651259642
transform 1 0 0 0 1 0
box -84 0 5264 1575
use li1_M1_contact  li1_M1_contact_4 pcells
timestamp 1648061256
transform -1 0 1406 0 -1 444
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_8
timestamp 1648061256
transform -1 0 4218 0 -1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_13
timestamp 1648061256
transform 1 0 5032 0 1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform 1 0 4736 0 1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform -1 0 4366 0 -1 814
box -53 -33 29 33
use dffrnx1_pcell  dffrnx1_pcell_2
timestamp 1651259642
transform 1 0 10360 0 1 0
box -84 0 5264 1575
use li1_M1_contact  li1_M1_contact_16
timestamp 1648061256
transform -1 0 6586 0 -1 444
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_7
timestamp 1648061256
transform 1 0 10212 0 1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_6
timestamp 1648061256
transform -1 0 9398 0 -1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_5
timestamp 1648061256
transform -1 0 9546 0 -1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_3
timestamp 1648061256
transform 1 0 9916 0 1 814
box -53 -33 29 33
use votern3x1_pcell  votern3x1_pcell_0 pcells
timestamp 1651259610
transform 1 0 15540 0 1 0
box -84 0 2082 1575
use li1_M1_contact  li1_M1_contact_17
timestamp 1648061256
transform -1 0 11766 0 -1 444
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_14
timestamp 1648061256
transform 1 0 15910 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_12
timestamp 1648061256
transform 1 0 15392 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_11
timestamp 1648061256
transform -1 0 14578 0 -1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_10
timestamp 1648061256
transform -1 0 14726 0 -1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_9
timestamp 1648061256
transform 1 0 15096 0 1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_15
timestamp 1648061256
transform 1 0 15688 0 -1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_18
timestamp 1648061256
transform -1 0 17390 0 -1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_2
timestamp 1648061256
transform 1 0 16724 0 1 592
box -53 -33 29 33
<< labels >>
rlabel metal1 17373 797 17407 831 1 QN
port 1 nsew signal output
rlabel metal1 1389 427 1423 461 1 D
port 2 nsew signal input
rlabel metal1 427 945 461 979 1 CLK
port 3 nsew signal input
rlabel metal1 1611 501 1645 535 1 RN
port 4 nsew signal input
rlabel metal1 -31 1492 17569 1554 1 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 -31 0 17569 62 1 VGND
port 6 nsew ground bidirectional abutment
rlabel nwell 55 1505 89 1539 1 VPB
port 7 nsew power bidirectional
rlabel pwell 55 13 89 47 1 VNB
port 8 nsew ground bidirectional
<< end >>
