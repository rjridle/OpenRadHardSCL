magic
tech sky130
magscale 1 2
timestamp 1645051190
<< nwell >>
rect -36 -287 352 37
<< pmos >>
rect 56 -251 86 1
rect 144 -251 174 1
rect 232 -251 262 1
<< pdiff >>
rect 0 -39 56 1
rect 0 -73 10 -39
rect 44 -73 56 -39
rect 0 -107 56 -73
rect 0 -141 10 -107
rect 44 -141 56 -107
rect 0 -175 56 -141
rect 0 -209 10 -175
rect 44 -209 56 -175
rect 0 -251 56 -209
rect 86 -39 144 1
rect 86 -73 98 -39
rect 132 -73 144 -39
rect 86 -107 144 -73
rect 86 -141 98 -107
rect 132 -141 144 -107
rect 86 -251 144 -141
rect 174 -39 232 1
rect 174 -73 186 -39
rect 220 -73 232 -39
rect 174 -107 232 -73
rect 174 -141 186 -107
rect 220 -141 232 -107
rect 174 -175 232 -141
rect 174 -209 186 -175
rect 220 -209 232 -175
rect 174 -251 232 -209
rect 262 -39 316 1
rect 262 -73 274 -39
rect 308 -73 316 -39
rect 262 -107 316 -73
rect 262 -141 274 -107
rect 308 -141 316 -107
rect 262 -251 316 -141
<< pdiffc >>
rect 10 -73 44 -39
rect 10 -141 44 -107
rect 10 -209 44 -175
rect 98 -73 132 -39
rect 98 -141 132 -107
rect 186 -73 220 -39
rect 186 -141 220 -107
rect 186 -209 220 -175
rect 274 -73 308 -39
rect 274 -141 308 -107
<< poly >>
rect 56 1 86 27
rect 144 1 174 27
rect 232 1 262 27
rect 56 -282 86 -251
rect 144 -282 174 -251
rect 232 -282 262 -251
rect 56 -312 262 -282
<< locali >>
rect 10 -39 44 42
rect 10 -107 44 -73
rect 10 -175 44 -141
rect 10 -227 44 -209
rect 98 -39 132 1
rect 98 -107 132 -73
rect 98 -227 132 -141
rect 186 -39 220 42
rect 186 -107 220 -73
rect 186 -175 220 -141
rect 186 -227 220 -209
rect 274 -39 308 1
rect 274 -107 308 -73
rect 274 -227 308 -141
<< end >>
