* HSPICE file created from tmp.ext - technology: sky130A

.option scale=5000u

.subckt tmp Y A B C VDD VSS
X0 Y C VDD VDD sky130_fd_pr__pfet_01v8 ad=34800 pd=1374 as=45200 ps=1826 w=400 l=30 M=2
X1 VDD A Y VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=400 l=30 M=2
X2 Y C a_372_210 VSS sky130_fd_pr__nfet_01v8 ad=7088 pd=312 as=0 ps=0 w=598 l=30
X3 VDD B Y VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=400 l=30 M=2
X4 a_372_210 B a_91_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=600 l=30
X5 VSS A a_91_103 VSS sky130_fd_pr__nfet_01v8 ad=7088 pd=312 as=0 ps=0 w=598 l=30
C0 VDD Y 2.50fF
.ends

** hspice subcircuit dictionary
