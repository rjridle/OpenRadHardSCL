* SPICE3 file created from OR2X1.ext - technology: sky130A

.subckt OR2X1 Y A B VDD GND
X0 Y.t1 a_198_209.t4 VDD.t7 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X1 a_131_1051.t1 A.t0 VDD.t1  |�0� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X2 a_131_1051.t3 B.t0 a_198_209.t2 �{�0� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X3 VDD.t5 a_198_209.t6 Y.t0  |�0� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X4 VDD.t3 A.t2 a_131_1051.t0 �{�0� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X5 a_198_209.t1 B.t2 a_131_1051.t2  |�0� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X6 Y a_198_209.t5 GND.t1 GND sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=0p ps=0u w=0u l=0u
C0 Y VDD 1.04fF
C1 A B 0.26fF
C2 VDD B 0.32fF
C3 VDD A 0.36fF
R0 a_198_209.n2 a_198_209.t6 512.525
R1 a_198_209.n2 a_198_209.t4 371.139
R2 a_198_209.n4 a_198_209.n1 287.966
R3 a_198_209.n3 a_198_209.t5 282.852
R4 a_198_209.n3 a_198_209.n2 247.347
R5 a_198_209.n9 a_198_209.n8 208.452
R6 a_198_209.n9 a_198_209.n4 142.305
R7 a_198_209.n11 a_198_209.n9 135.417
R8 a_198_209.n12 a_198_209.n0 55.263
R9 a_198_209.n8 a_198_209.n7 30
R10 a_198_209.n11 a_198_209.n10 30
R11 a_198_209.n12 a_198_209.n11 25.263
R12 a_198_209.n6 a_198_209.n5 24.383
R13 a_198_209.n8 a_198_209.n6 23.684
R14 a_198_209.n1 a_198_209.t2 14.282
R15 a_198_209.n1 a_198_209.t1 14.282
R16 a_198_209.n4 a_198_209.n3 10.343
R17 VDD.n66 VDD.n55 144.705
R18 VDD.n35 VDD.t7 135.17
R19 VDD.n24 VDD.t5 135.17
R20 VDD.n97 VDD.n96 129.849
R21 VDD.n51 VDD.n50 92.5
R22 VDD.n49 VDD.n48 92.5
R23 VDD.n47 VDD.n46 92.5
R24 VDD.n45 VDD.n44 92.5
R25 VDD.n53 VDD.n52 92.5
R26 VDD.n80 VDD.n79 92.5
R27 VDD.n78 VDD.n77 92.5
R28 VDD.n76 VDD.n75 92.5
R29 VDD.n74 VDD.n73 92.5
R30 VDD.n82 VDD.n81 92.5
R31 VDD.n14 VDD.n1 92.5
R32 VDD.n5 VDD.n4 92.5
R33 VDD.n7 VDD.n6 92.5
R34 VDD.n9 VDD.n8 92.5
R35 VDD.n11 VDD.n10 92.5
R36 VDD.n13 VDD.n12 92.5
R37 VDD.n21 VDD.n20 92.059
R38 VDD.n65 VDD.n64 92.059
R39 VDD.n88 VDD.n87 92.059
R40 VDD.n20 VDD.n16 67.194
R41 VDD.n20 VDD.n17 67.194
R42 VDD.n20 VDD.n18 67.194
R43 VDD.n20 VDD.n19 67.194
R44 VDD.n72 VDD.n71 44.141
R45 VDD.n5 VDD.n3 44.141
R46 VDD.n71 VDD.n69 44.107
R47 VDD.n3 VDD.n2 44.107
R48 VDD.n25  |�0� 43.472
R49 VDD.n33 VDD.t6 43.472
R50 VDD.n20 VDD.n15 41.052
R51 VDD.n84 VDD.n83 39.742
R52 VDD.n63 VDD.n60 39.742
R53 VDD.n63 VDD.n62 39.742
R54 VDD.n59 VDD.n58 39.742
R55 VDD.n71 VDD.n70 38
R56 VDD.n62 VDD.n61 36.774
R57 VDD.n1 VDD.n0 30.923
R58 VDD.n87 VDD.n85 26.38
R59 VDD.n87 VDD.n84 26.38
R60 VDD.n87 VDD.n86 26.38
R61 VDD.n64 VDD.n63 26.38
R62 VDD.n64 VDD.n59 26.38
R63 VDD.n64 VDD.n57 26.38
R64 VDD.n64 VDD.n56 26.38
R65 VDD.n90 VDD.n82 22.915
R66 VDD.n23 VDD.n14 22.915
R67 VDD.n109 �{�0� 20.457
R68 VDD.n98 �{�0� 17.9
R69 VDD.n82 VDD.n80 14.864
R70 VDD.n80 VDD.n78 14.864
R71 VDD.n78 VDD.n76 14.864
R72 VDD.n76 VDD.n74 14.864
R73 VDD.n74 VDD.n72 14.864
R74 VDD.n53 VDD.n51 14.864
R75 VDD.n51 VDD.n49 14.864
R76 VDD.n49 VDD.n47 14.864
R77 VDD.n47 VDD.n45 14.864
R78 VDD.n45 VDD.n43 14.864
R79 VDD.n43 VDD.n42 14.864
R80 VDD.n14 VDD.n13 14.864
R81 VDD.n13 VDD.n11 14.864
R82 VDD.n11 VDD.n9 14.864
R83 VDD.n9 VDD.n7 14.864
R84 VDD.n7 VDD.n5 14.864
R85 VDD.n67 VDD.n54 14.864
R86 VDD.n96 VDD.t1 14.282
R87 VDD.n96 VDD.t3 14.282
R88 VDD.n23 VDD.n22 8.855
R89 VDD.n22 VDD.n21 8.855
R90 VDD.n27 VDD.n26 8.855
R91 VDD.n26 VDD.n25 8.855
R92 VDD.n31 VDD.n30 8.855
R93 VDD.n30 VDD.n29 8.855
R94 VDD.n36 VDD.n34 8.855
R95 VDD.n34 VDD.n33 8.855
R96 VDD.n40 VDD.n39 8.855
R97 VDD.n39 VDD.n38 8.855
R98 VDD.n67 VDD.n66 8.855
R99 VDD.n66 VDD.n65 8.855
R100 VDD.n115 VDD.n114 8.855
R101 VDD.n114 VDD.n113 8.855
R102 VDD.n111 VDD.n110 8.855
R103 VDD.n110 VDD.n109 8.855
R104 VDD.n107 VDD.n106 8.855
R105 VDD.n106  |�0� 8.855
R106 VDD.n104 VDD.n103 8.855
R107 VDD.n103 VDD.n102 8.855
R108 VDD.n100 VDD.n99 8.855
R109 VDD.n99 VDD.n98 8.855
R110 VDD.n94 VDD.n93 8.855
R111 VDD.n93 VDD.n92 8.855
R112 VDD.n90 VDD.n89 8.855
R113 VDD.n89 VDD.n88 8.855
R114 VDD.n54 VDD.n53 8.051
R115 VDD.n100 VDD.n97 6.193
R116 VDD.n28 VDD.n23 4.795
R117 VDD.n28 VDD.n27 4.65
R118 VDD.n32 VDD.n31 4.65
R119 VDD.n37 VDD.n36 4.65
R120 VDD.n41 VDD.n40 4.65
R121 VDD.n68 VDD.n67 4.65
R122 VDD.n116 VDD.n115 4.65
R123 VDD.n112 VDD.n111 4.65
R124 VDD.n108 VDD.n107 4.65
R125 VDD.n105 VDD.n104 4.65
R126 VDD.n101 VDD.n100 4.65
R127 VDD.n95 VDD.n94 4.65
R128 VDD.n91 VDD.n90 4.65
R129 VDD.n102  |�0� 2.557
R130 VDD.n27 VDD.n24 2.064
R131 VDD.n36 VDD.n35 2.064
R132 VDD.n68 VDD.n41 0.29
R133 VDD.n91 VDD 0.207
R134 VDD.n108 VDD.n105 0.181
R135 VDD.n32 VDD.n28 0.157
R136 VDD.n37 VDD.n32 0.157
R137 VDD.n41 VDD.n37 0.145
R138 VDD.n116 VDD.n112 0.145
R139 VDD.n112 VDD.n108 0.145
R140 VDD.n105 VDD.n101 0.145
R141 VDD.n101 VDD.n95 0.145
R142 VDD.n95 VDD.n91 0.145
R143 VDD VDD.n68 0.078
R144 VDD VDD.n116 0.066
R145 Y.n5 Y.n4 272.451
R146 Y.n5 Y.n0 271.281
R147 Y.n4 Y.n3 30
R148 Y.n2 Y.n1 24.383
R149 Y.n4 Y.n2 23.684
R150 Y.n0 Y.t0 14.282
R151 Y.n0 Y.t1 14.282
R152 Y Y.n5 4.65
R153 GND.n32 GND.n31 237.558
R154 GND.n29 GND.n28 210.82
R155 GND.n56 GND.n55 40.431
R156 GND.n67 GND.n66 40.003
R157 GND.n21 GND.n20 37.582
R158 GND.n41 GND.n40 37.582
R159 GND.t1 GND.n18 32.601
R160 GND.n18 GND.n17 21.734
R161 GND.n4 GND.n3 20.705
R162 GND.n10 GND.n9 20.705
R163 GND.n22 GND.n21 20.705
R164 GND.n46 GND.n45 20.705
R165 GND.n57 GND.n56 20.705
R166 GND.n62 GND.n61 20.705
R167 GND.n68 GND.n67 20.705
R168 GND.n42 GND.n41 20.705
R169 GND.n3 GND.n2 19.952
R170 GND.n30 GND.n29 18.953
R171 GND.n66 GND.n65 17.258
R172 GND.n20 GND.t1 15.644
R173 GND.n40 GND.t2 15.644
R174 GND.n33 GND.n30 14.864
R175 GND.n55 GND.t0 13.654
R176 GND.n20 GND.n19 13.541
R177 GND.n40 GND.n39 13.541
R178 GND.n58 GND.n57 9.29
R179 GND.n43 GND.n38 9.154
R180 GND.n48 GND.n47 9.154
R181 GND.n51 GND.n50 9.154
R182 GND.n58 GND.n53 9.154
R183 GND.n63 GND.n60 9.154
R184 GND.n70 GND.n69 9.154
R185 GND.n33 GND.n32 9.154
R186 GND.n26 GND.n25 9.154
R187 GND.n23 GND.n14 9.154
R188 GND.n12 GND.n11 9.154
R189 GND.n6 GND.n5 9.154
R190 GND.t0 GND.n54 7.04
R191 GND.n7 GND.n1 4.795
R192 GND.n37 GND.n36 4.65
R193 GND.n7 GND.n6 4.65
R194 GND.n13 GND.n12 4.65
R195 GND.n24 GND.n23 4.65
R196 GND.n27 GND.n26 4.65
R197 GND.n34 GND.n33 4.65
R198 GND.n71 GND.n70 4.65
R199 GND.n64 GND.n63 4.65
R200 GND.n59 GND.n58 4.65
R201 GND.n52 GND.n51 4.65
R202 GND.n49 GND.n48 4.65
R203 GND.n44 GND.n43 4.65
R204 GND.n16 GND.n15 4.504
R205 GND.n6 GND.n4 4.129
R206 GND.n63 GND.n62 4.129
R207 GND.n48 GND.n46 4.129
R208 GND.n23 GND.n22 3.716
R209 GND.t1 GND.n16 2.452
R210 GND.n70 GND.n68 1.032
R211 GND.n43 GND.n42 1.032
R212 GND.n1 GND.n0 0.474
R213 GND.n36 GND.n35 0.474
R214 GND.n9 GND.n8 0.376
R215 GND.n34 GND.n27 0.29
R216 GND.n37 GND 0.207
R217 GND.n12 GND.n10 0.206
R218 GND.n59 GND.n52 0.181
R219 GND.n13 GND.n7 0.157
R220 GND.n24 GND.n13 0.157
R221 GND.n27 GND.n24 0.145
R222 GND.n71 GND.n64 0.145
R223 GND.n64 GND.n59 0.145
R224 GND.n52 GND.n49 0.145
R225 GND.n49 GND.n44 0.145
R226 GND.n44 GND.n37 0.145
R227 GND GND.n34 0.078
R228 GND GND.n71 0.066
R229 A.n0 A.t0 486.819
R230 A.n0 A.t2 384.527
R231 A.n1 A.t1 378.637
R232 A.n1 A.n0 151.269
R233 A A.n1 4.65
R234 a_131_1051.n0 a_131_1051.t3 228.369
R235 a_131_1051.n0 a_131_1051.t0 219.778
R236 a_131_1051.n1 a_131_1051.n0 42.29
R237 a_131_1051.n1 a_131_1051.t2 14.282
R238 a_131_1051.t1 a_131_1051.n1 14.282
R239 B.n0 B.t0 470.752
R240 B.n0 B.t2 384.527
R241 B.n1 B.t1 314.896
R242 B.n1 B.n0 182.932
R243 B B.n1 4.65
C4 VDD GND 2.30fF
C5 a_131_1051.n0 GND 0.50fF
C6 a_131_1051.n1 GND 0.21fF
C7 Y.n0 GND 0.65fF
C8 Y.n1 GND 0.04fF
C9 Y.n2 GND 0.05fF
C10 Y.n3 GND 0.03fF
C11 Y.n4 GND 0.19fF
C12 Y.n5 GND 0.63fF
C13 VDD.n1 GND 0.03fF
C14 VDD.n2 GND 0.08fF
C15 VDD.n3 GND 0.02fF
C16 VDD.n4 GND 0.02fF
C17 VDD.n5 GND 0.05fF
C18 VDD.n6 GND 0.02fF
C19 VDD.n7 GND 0.02fF
C20 VDD.n8 GND 0.02fF
C21 VDD.n9 GND 0.02fF
C22 VDD.n10 GND 0.02fF
C23 VDD.n11 GND 0.02fF
C24 VDD.n12 GND 0.02fF
C25 VDD.n13 GND 0.02fF
C26 VDD.n14 GND 0.03fF
C27 VDD.n15 GND 0.01fF
C28 VDD.n20 GND 0.37fF
C29 VDD.n21 GND 0.22fF
C30 VDD.n22 GND 0.02fF
C31 VDD.n23 GND 0.03fF
C32 VDD.n24 GND 0.05fF
C33 VDD.n25 GND 0.16fF
C34 VDD.n26 GND 0.01