* SPICE3 file created from NOR2X2.ext - technology: sky130A

.subckt NOR2X2 VDD VSS A B YN
M1000 a_92_629# A YN VDD pshort w=3u l=0.15u
+  ad=0.87p pd=6.58u as=1.74p ps=13.16u
M1001 a_276_629# B VDD VDD pshort w=3u l=0.15u
+  ad=0.87p pd=6.58u as=0.99p ps=6.66u
M1002 YN A VSS VSS nshort w=3u l=0.15u
+  ad=0.3176p pd=3u as=1.85625p ps=12.67u
M1003 YN B VSS VSS nshort w=3u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 VDD A a_92_629# VDD pshort w=3u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 YN B a_276_629# VDD pshort w=3u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
.ends
