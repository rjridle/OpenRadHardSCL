magic
tech sky130
magscale 1 2
timestamp 1645051291
<< nwell >>
rect 52 -287 352 37
<< pmos >>
rect 144 -251 174 1
rect 232 -251 262 1
<< pdiff >>
rect 88 -39 144 1
rect 88 -73 98 -39
rect 132 -73 144 -39
rect 88 -107 144 -73
rect 88 -141 98 -107
rect 132 -141 144 -107
rect 88 -175 144 -141
rect 88 -209 98 -175
rect 132 -209 144 -175
rect 88 -251 144 -209
rect 174 -39 232 1
rect 174 -73 186 -39
rect 220 -73 232 -39
rect 174 -107 232 -73
rect 174 -141 186 -107
rect 220 -141 232 -107
rect 174 -251 232 -141
rect 262 -39 316 1
rect 262 -73 274 -39
rect 308 -73 316 -39
rect 262 -107 316 -73
rect 262 -141 274 -107
rect 308 -141 316 -107
rect 262 -175 316 -141
rect 262 -209 274 -175
rect 308 -209 316 -175
rect 262 -251 316 -209
<< pdiffc >>
rect 98 -73 132 -39
rect 98 -141 132 -107
rect 98 -209 132 -175
rect 186 -73 220 -39
rect 186 -141 220 -107
rect 274 -73 308 -39
rect 274 -141 308 -107
rect 274 -209 308 -175
<< poly >>
rect 144 1 174 27
rect 232 1 262 27
rect 144 -282 174 -251
rect 232 -282 262 -251
rect 144 -312 262 -282
<< locali >>
rect 98 -39 132 42
rect 98 -107 132 -73
rect 98 -175 132 -141
rect 98 -227 132 -209
rect 186 -39 220 1
rect 186 -107 220 -73
rect 186 -227 220 -141
rect 274 -39 308 42
rect 274 -107 308 -73
rect 274 -175 308 -141
rect 274 -227 308 -209
<< end >>
