* SPICE3 file created from AND2X1.ext - technology: sky130A

.subckt AND2X1 Y A B VDD VSS
X0 VDD A a_217_1050 VDD sky130_fd_pr__pfet_01v8 ad=2.78e+12p pd=2.278e+07u as=0p ps=0u w=2e+06u l=150000u M=2
X1 Y a_217_1050 VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=150000u M=2
X2 Y a_217_1050 VSS VSS sky130_fd_pr__nfet_01v8 ad=1.791e+11p pd=1.57e+06u as=1.3199e+12p ps=9.67e+06u w=3e+06u l=150000u
X3 VDD B a_217_1050 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X4 VSS A a_112_101 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X5 a_217_1050 B a_112_101 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
C0 VDD a_217_1050 2.24fF
.ends
