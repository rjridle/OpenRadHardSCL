magic
tech sky130
magscale 1 2
timestamp 1651259490
<< nwell >>
rect 84 903 582 1575
rect 83 832 582 903
<< pwell >>
rect -31 0 697 572
<< pdiffc >>
rect 141 1377 175 1411
rect 229 1377 263 1411
rect 317 1377 351 1411
rect 493 1377 527 1411
rect 141 1105 175 1139
rect 317 1105 351 1139
rect 405 1105 439 1139
<< psubdiff >>
rect 31 510 635 572
rect 31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 361 47
rect 395 13 433 47
rect 467 13 505 47
rect 539 13 577 47
rect 611 13 635 47
<< nsubdiff >>
rect 31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 361 1539
rect 395 1505 433 1539
rect 467 1505 505 1539
rect 539 1505 577 1539
rect 611 1505 635 1539
rect 31 868 635 930
<< psubdiffcont >>
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 361 13 395 47
rect 433 13 467 47
rect 505 13 539 47
rect 577 13 611 47
<< nsubdiffcont >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 361 1505 395 1539
rect 433 1505 467 1539
rect 505 1505 539 1539
rect 577 1505 611 1539
<< poly >>
rect 168 403 198 441
rect 362 410 392 411
<< locali >>
rect 31 1539 635 1554
rect 31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 361 1539
rect 395 1505 433 1539
rect 467 1505 505 1539
rect 539 1505 577 1539
rect 611 1505 635 1539
rect 31 1492 635 1505
rect 141 1411 175 1451
rect 141 1359 175 1377
rect 229 1411 263 1492
rect 229 1359 263 1377
rect 317 1411 527 1445
rect 317 1359 351 1377
rect 493 1359 527 1377
rect 141 1139 175 1157
rect 317 1139 351 1157
rect 141 1071 351 1105
rect 405 1139 439 1157
rect 405 1071 535 1105
rect 205 461 239 988
rect 353 954 361 988
rect 353 469 387 954
rect 353 461 357 469
rect 501 376 535 1071
rect 219 342 535 376
rect 219 261 253 342
rect 413 261 447 342
rect 122 62 156 101
rect 219 62 253 117
rect 316 62 350 101
rect 413 62 447 117
rect 510 62 544 101
rect 31 47 635 62
rect 31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 361 47
rect 395 13 433 47
rect 467 13 505 47
rect 539 13 577 47
rect 611 13 635 47
rect 31 0 635 13
<< viali >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 361 1505 395 1539
rect 433 1505 467 1539
rect 505 1505 539 1539
rect 577 1505 611 1539
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 361 13 395 47
rect 433 13 467 47
rect 505 13 539 47
rect 577 13 611 47
<< metal1 >>
rect 31 1539 635 1554
rect 31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 361 1539
rect 395 1505 433 1539
rect 467 1505 505 1539
rect 539 1505 577 1539
rect 611 1505 635 1539
rect 31 1492 635 1505
rect 31 47 635 62
rect 31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 361 47
rect 395 13 433 47
rect 467 13 505 47
rect 539 13 577 47
rect 611 13 635 47
rect 31 0 635 13
use diff_ring_side  diff_ring_side_1
timestamp 1651259451
transform 1 0 0 0 1 0
box -84 0 84 1575
use nmos_top_trim1  nmos_top_trim1_1
timestamp 1651256895
transform -1 0 360 0 1 101
box 0 0 248 309
use poly_li1_contact  poly_li1_contact_0
timestamp 1648060378
transform 0 1 192 -1 0 988
box -32 -28 34 26
use poly_li1_contact  poly_li1_contact_1
timestamp 1648060378
transform 0 1 223 -1 0 445
box -32 -28 34 26
use pmos2_1  pmos2_1_0
timestamp 1647326732
transform 1 0 43 0 1 1450
box 52 -460 352 37
use nmos_top_trim2  nmos_top_trim2_0
timestamp 1651256905
transform -1 0 554 0 1 101
box 0 0 248 309
use poly_li1_contact  poly_li1_contact_3
timestamp 1648060378
transform 0 1 378 -1 0 988
box -32 -28 34 26
use poly_li1_contact  poly_li1_contact_2
timestamp 1648060378
transform 0 -1 369 1 0 443
box -32 -28 34 26
use pmos2_1  pmos2_1_1
timestamp 1647326732
transform 1 0 219 0 1 1450
box 52 -460 352 37
use diff_ring_side  diff_ring_side_0
timestamp 1651259451
transform 1 0 666 0 1 0
box -84 0 84 1575
<< end >>
