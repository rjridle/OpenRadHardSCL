* HSPICE file created from tmp.ext - technology: sky130A

.option scale=5000u

.subckt tmp B A Y VDD VSS
X0 a_575_1051 a_184_209 Y VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=23200 ps=916 w=400 l=30 M=2
X1 VDD a_612_186 B VDD sky130_fd_pr__pfet_01v8 ad=67200 pd=2736 as=11600 ps=458 w=400 l=30 M=2
X2 VSS B a_1222_101 VSS sky130_fd_pr__nfet_01v8 ad=106756 pd=3872 as=0 ps=0 w=598 l=30
X3 Y a_184_209 a_1222_101 VSS sky130_fd_pr__nfet_01v8 ad=14176 pd=624 as=0 ps=0 w=598 l=30
X4 a_1241_1051 B VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=400 l=30 M=2
X5 a_184_209 A VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=400 l=30 M=2
X6 VSS a_612_186 a_556_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=598 l=30
X7 B a_612_186 VSS VSS sky130_fd_pr__nfet_01v8 ad=7088 pd=312 as=0 ps=0 w=598 l=30
X8 a_1241_1051 A Y VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=400 l=30 M=2
X9 Y A a_556_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=598 l=30
X10 VDD a_612_186 a_575_1051 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=400 l=30 M=2
X11 a_184_209 A VSS VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=598 l=30
C0 VDD a_184_209 2.56fF
.ends

** hspice subcircuit dictionary
