* SPICE3 file created from FA.ext - technology: sky130A

.subckt FA SUM COUT A B CIN VDD GND
X0 GND A.t1 a_556_101.t0 GND sky130_fd_pr__nfet_01v8 ad=1.09968p pd=7.906u as=0p ps=0u w=0u l=0u
X1 VDD.t16 a_836_209.t6 a_2405_209.t2 VDD.t15 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X2 a_807_990.t1 B.t0 VDD.t66  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X3 VDD.t24 a_4657_1050.t6 a_5291_209.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X4 a_185_209.t1 A.t0 VDD.t55  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X5 a_3027_990.t1 CIN.t1 VDD.t46 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X6 SUM.t0 a_3027_990.t3 a_2795_1051.t3  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X7 COUT.t1 a_6858_209.t4 VDD.t30 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X8 GND a_3027_990.t4 a_3442_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X9 a_3461_1051.t3 a_2405_209.t3 SUM.t4  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X10 VDD.t69 B.t2 a_5767_1050.t4 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X11 VDD.t14 a_836_209.t8 a_4657_1050.t1  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X12 COUT a_6858_209.t5 GND.t19 GND sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=0p ps=0u w=0u l=0u
X13 a_575_1051.t3 a_807_990.t3 a_836_209.t2 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X14 a_2795_1051.t1 a_836_209.t9 VDD.t12  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X15 VDD.t18 CIN.t2 a_3461_1051.t1 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X16 a_4657_1050.t4 CIN.t3 VDD.t20  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X17 a_1241_1051.t3 B.t3 VDD.t34 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X18 VDD.t36 a_5291_209.t4 a_6791_1051.t3  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X19 VDD.t48 a_5767_1050.t6 a_6401_209.t1 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X20 a_6791_1051.t1 a_6401_209.t4 a_6858_209.t2  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X21 a_2405_209.t1 a_836_209.t10 VDD.t10 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X22 a_4657_1050.t0 a_836_209.t11 VDD.t8  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X23 a_836_209.t5 a_807_990.t4 a_575_1051.t2 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X24 a_5291_209.t0 a_4657_1050.t7 VDD.t22  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X25 a_1241_1051.t1 a_185_209.t4 a_836_209.t1 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X26 SUM a_2405_209.t5 a_3442_101.t1 GND sky130_fd_pr__nfet_01v8 ad=3.582p pd=3.14u as=0p ps=0u w=0u l=0u
X27 VDD.t40 A.t4 a_575_1051.t1  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X28 VDD.t28 A.t5 a_185_209.t0 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X29 SUM.t3 a_2405_209.t4 a_3461_1051.t2  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X30 VDD.t53 CIN.t5 a_3027_990.t0 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X31 a_5767_1050.t3 B.t6 VDD.t64  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X32 GND CIN.t6 a_4552_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X33 VDD.t1 A.t6 a_5767_1050.t1 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X34 GND a_836_209.t12 a_2776_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X35 a_2795_1051.t2 a_3027_990.t5 SUM.t1  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X36 VDD.t32 B.t7 a_1241_1051.t2 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X37 a_5767_1050.t0 A.t7 VDD.t4  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X38 VDD.t43 a_6858_209.t6 COUT.t0 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X39 GND a_807_990.t5 a_1222_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X40 a_3461_1051.t0 CIN.t7 VDD.t59  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X41 a_6401_209.t0 a_5767_1050.t7 VDD.t50 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X42 a_6858_209.t1 a_6401_209.t5 a_6791_1051.t0  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X43 SUM CIN.t0 a_2776_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X44 VDD.t71 CIN.t8 a_4657_1050.t3 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X45 GND B.t1 a_5662_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X46 a_575_1051.t0 A.t8 VDD.t38  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X47 a_836_209.t0 a_185_209.t5 a_1241_1051.t0 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X48 VDD.t26 B.t8 a_807_990.t0  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X49 a_6791_1051.t2 a_5291_209.t5 VDD.t57 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X50 VDD.t6 a_836_209.t14 a_2795_1051.t0  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
C0 COUT VDD 1.04fF
C1 SUM A 0.26fF
C2 VDD A 1.59fF
C3 SUM B 0.24fF
C4 VDD B 3.94fF
C5 CIN A 0.54fF
C6 CIN B 1.51fF
C7 SUM VDD 1.04fF
C8 SUM CIN 0.62fF
C9 A B 0.85fF
C10 CIN VDD 2.13fF
R0 a_836_209.n1 a_836_209.t6 512.525
R1 a_836_209.n2 a_836_209.t9 480.392
R2 a_836_209.n5 a_836_209.t8 472.359
R3 a_836_209.n3 a_836_209.t12 412.921
R4 a_836_209.n2 a_836_209.t14 403.272
R5 a_836_209.n5 a_836_209.t11 384.527
R6 a_836_209.n1 a_836_209.t10 371.139
R7 a_836_209.n11 a_836_209.n10 327.32
R8 a_836_209.n15 a_836_209.n13 312.103
R9 a_836_209.n6 a_836_209.n5 294.249
R10 a_836_209.n11 a_836_209.n9 260.107
R11 a_836_209.n13 a_836_209.n0 260.107
R12 a_836_209.n4 a_836_209.n1 163.771
R13 a_836_209.n6 a_836_209.t7 136.225
R14 a_836_209.n7 a_836_209.t13 132.04
R15 a_836_209.n3 a_836_209.n2 115.947
R16 a_836_209.n8 a_836_209.n7 111.435
R17 a_836_209.n8 a_836_209.n4 55.717
R18 a_836_209.n7 a_836_209.n6 18.232
R19 a_836_209.n15 a_836_209.n14 15.218
R20 a_836_209.n9 a_836_209.t1 14.282
R21 a_836_209.n9 a_836_209.t0 14.282
R22 a_836_209.n0 a_836_209.t2 14.282
R23 a_836_209.n0 a_836_209.t5 14.282
R24 a_836_209.n16 a_836_209.n15 12.014
R25 a_836_209.n4 a_836_209.n3 11.159
R26 a_836_209.n12 a_836_209.n8 7.325
R27 a_836_209.n13 a_836_209.n12 7.053
R28 a_836_209.n12 a_836_209.n11 4.65
R29 a_2405_209.n2 a_2405_209.t4 477.179
R30 a_2405_209.n2 a_2405_209.t3 406.485
R31 a_2405_209.n3 a_2405_209.t5 341.566
R32 a_2405_209.n6 a_2405_209.n4 272.451
R33 a_2405_209.n4 a_2405_209.n1 271.281
R34 a_2405_209.n3 a_2405_209.n2 199.524
R35 a_2405_209.n6 a_2405_209.n5 30
R36 a_2405_209.n7 a_2405_209.n0 24.383
R37 a_2405_209.n7 a_2405_209.n6 23.684
R38 a_2405_209.n1 a_2405_209.t2 14.282
R39 a_2405_209.n1 a_2405_209.t1 14.282
R40 a_2405_209.n4 a_2405_209.n3 13.879
R41 VDD.n443 VDD.n442 173.148
R42 VDD.n498 VDD.n497 173.148
R43 VDD.n641 VDD.n640 173.148
R44 VDD.n696 VDD.n695 173.148
R45 VDD.n422 VDD.n411 144.705
R46 VDD.n474 VDD.n467 144.705
R47 VDD.n529 VDD.n522 144.705
R48 VDD.n589 VDD.n582 144.705
R49 VDD.n617 VDD.n610 144.705
R50 VDD.n367 VDD.n360 144.705
R51 VDD.n672 VDD.n665 144.705
R52 VDD.n323 VDD.n316 144.705
R53 VDD.n266 VDD.n259 144.705
R54 VDD.n222 VDD.n215 144.705
R55 VDD.n165 VDD.n158 144.705
R56 VDD.n121 VDD.n114 144.705
R57 VDD.n66 VDD.n55 144.705
R58 VDD.n269 VDD.t14 143.754
R59 VDD.n170 VDD.t1 143.754
R60 VDD.n395 VDD.t55 135.17
R61 VDD.n402 VDD.t28 135.17
R62 VDD.n548 VDD.t66 135.17
R63 VDD.n557 VDD.t26 135.17
R64 VDD.n594 VDD.t10 135.17
R65 VDD.n601 VDD.t16 135.17
R66 VDD.n335 VDD.t46 135.17
R67 VDD.n326 VDD.t53 135.17
R68 VDD.n291 VDD.t20 135.17
R69 VDD.n236 VDD.t22 135.17
R70 VDD.n225 VDD.t24 135.17
R71 VDD.n190 VDD.t64 135.17
R72 VDD.n133 VDD.t50 135.17
R73 VDD.n124 VDD.t48 135.17
R74 VDD.n35 VDD.t30 135.17
R75 VDD.n24 VDD.t43 135.17
R76 VDD.n85 VDD.n84 129.849
R77 VDD.n279 VDD.n278 129.472
R78 VDD.n179 VDD.n178 129.472
R79 VDD.n51 VDD.n50 92.5
R80 VDD.n49 VDD.n48 92.5
R81 VDD.n47 VDD.n46 92.5
R82 VDD.n45 VDD.n44 92.5
R83 VDD.n53 VDD.n52 92.5
R84 VDD.n110 VDD.n109 92.5
R85 VDD.n108 VDD.n107 92.5
R86 VDD.n106 VDD.n105 92.5
R87 VDD.n104 VDD.n103 92.5
R88 VDD.n112 VDD.n111 92.5
R89 VDD.n154 VDD.n153 92.5
R90 VDD.n152 VDD.n151 92.5
R91 VDD.n150 VDD.n149 92.5
R92 VDD.n148 VDD.n147 92.5
R93 VDD.n156 VDD.n155 92.5
R94 VDD.n211 VDD.n210 92.5
R95 VDD.n209 VDD.n208 92.5
R96 VDD.n207 VDD.n206 92.5
R97 VDD.n205 VDD.n204 92.5
R98 VDD.n213 VDD.n212 92.5
R99 VDD.n255 VDD.n254 92.5
R100 VDD.n253 VDD.n252 92.5
R101 VDD.n251 VDD.n250 92.5
R102 VDD.n249 VDD.n248 92.5
R103 VDD.n257 VDD.n256 92.5
R104 VDD.n312 VDD.n311 92.5
R105 VDD.n310 VDD.n309 92.5
R106 VDD.n308 VDD.n307 92.5
R107 VDD.n306 VDD.n305 92.5
R108 VDD.n314 VDD.n313 92.5
R109 VDD.n356 VDD.n355 92.5
R110 VDD.n354 VDD.n353 92.5
R111 VDD.n352 VDD.n351 92.5
R112 VDD.n350 VDD.n349 92.5
R113 VDD.n358 VDD.n357 92.5
R114 VDD.n685 VDD.n684 92.5
R115 VDD.n683 VDD.n682 92.5
R116 VDD.n681 VDD.n680 92.5
R117 VDD.n679 VDD.n678 92.5
R118 VDD.n687 VDD.n686 92.5
R119 VDD.n630 VDD.n629 92.5
R120 VDD.n628 VDD.n627 92.5
R121 VDD.n626 VDD.n625 92.5
R122 VDD.n624 VDD.n623 92.5
R123 VDD.n632 VDD.n631 92.5
R124 VDD.n578 VDD.n577 92.5
R125 VDD.n576 VDD.n575 92.5
R126 VDD.n574 VDD.n573 92.5
R127 VDD.n572 VDD.n571 92.5
R128 VDD.n580 VDD.n579 92.5
R129 VDD.n542 VDD.n541 92.5
R130 VDD.n540 VDD.n539 92.5
R131 VDD.n538 VDD.n537 92.5
R132 VDD.n536 VDD.n535 92.5
R133 VDD.n544 VDD.n543 92.5
R134 VDD.n487 VDD.n486 92.5
R135 VDD.n485 VDD.n484 92.5
R136 VDD.n483 VDD.n482 92.5
R137 VDD.n481 VDD.n480 92.5
R138 VDD.n489 VDD.n488 92.5
R139 VDD.n432 VDD.n431 92.5
R140 VDD.n430 VDD.n429 92.5
R141 VDD.n428 VDD.n427 92.5
R142 VDD.n426 VDD.n425 92.5
R143 VDD.n434 VDD.n433 92.5
R144 VDD.n381 VDD.n380 92.5
R145 VDD.n379 VDD.n378 92.5
R146 VDD.n377 VDD.n376 92.5
R147 VDD.n375 VDD.n374 92.5
R148 VDD.n383 VDD.n382 92.5
R149 VDD.n14 VDD.n1 92.5
R150 VDD.n5 VDD.n4 92.5
R151 VDD.n7 VDD.n6 92.5
R152 VDD.n9 VDD.n8 92.5
R153 VDD.n11 VDD.n10 92.5
R154 VDD.n13 VDD.n12 92.5
R155 VDD.n21 VDD.n20 92.059
R156 VDD.n65 VDD.n64 92.059
R157 VDD.n120 VDD.n119 92.059
R158 VDD.n164 VDD.n163 92.059
R159 VDD.n221 VDD.n220 92.059
R160 VDD.n265 VDD.n264 92.059
R161 VDD.n322 VDD.n321 92.059
R162 VDD.n366 VDD.n365 92.059
R163 VDD.n671 VDD.n670 92.059
R164 VDD.n616 VDD.n615 92.059
R165 VDD.n588 VDD.n587 92.059
R166 VDD.n528 VDD.n527 92.059
R167 VDD.n473 VDD.n472 92.059
R168 VDD.n421 VDD.n420 92.059
R169 VDD.n389 VDD.n388 92.059
R170 VDD.n20 VDD.n16 67.194
R171 VDD.n20 VDD.n17 67.194
R172 VDD.n20 VDD.n18 67.194
R173 VDD.n20 VDD.n19 67.194
R174 VDD.n373 VDD.n372 44.141
R175 VDD.n479 VDD.n478 44.141
R176 VDD.n534 VDD.n533 44.141
R177 VDD.n570 VDD.n569 44.141
R178 VDD.n622 VDD.n621 44.141
R179 VDD.n677 VDD.n676 44.141
R180 VDD.n348 VDD.n347 44.141
R181 VDD.n304 VDD.n303 44.141
R182 VDD.n247 VDD.n246 44.141
R183 VDD.n203 VDD.n202 44.141
R184 VDD.n146 VDD.n145 44.141
R185 VDD.n102 VDD.n101 44.141
R186 VDD.n5 VDD.n3 44.141
R187 VDD.n478 VDD.n476 44.107
R188 VDD.n533 VDD.n531 44.107
R189 VDD.n569 VDD.n567 44.107
R190 VDD.n621 VDD.n619 44.107
R191 VDD.n676 VDD.n674 44.107
R192 VDD.n347 VDD.n345 44.107
R193 VDD.n303 VDD.n301 44.107
R194 VDD.n246 VDD.n244 44.107
R195 VDD.n202 VDD.n200 44.107
R196 VDD.n145 VDD.n143 44.107
R197 VDD.n101 VDD.n99 44.107
R198 VDD.n372 VDD.n370 44.107
R199 VDD.n3 VDD.n2 44.107
R200 VDD.n25 �{�� 43.472
R201 VDD.n33 �{�� 43.472
R202 VDD.n125 �{�� 43.472
R203 VDD.n134 �{�� 43.472
R204 VDD.n226  43.472
R205 VDD.n234  |�� 43.472
R206 VDD.n327 �{�� 43.472
R207 VDD.n336 �{�� 43.472
R208 VDD.n602 VDD.t15 43.472
R209 VDD.n592 �{�� 43.472
R210 VDD.n558  |�� 43.472
R211 VDD.n549  43.472
R212 VDD.n403 �{�� 43.472
R213 VDD.n393  |�� 43.472
R214 VDD.n20 VDD.n15 41.052
R215 VDD.n59 VDD.n57 39.742
R216 VDD.n59 VDD.n58 39.742
R217 VDD.n61 VDD.n60 39.742
R218 VDD.n116 VDD.n115 39.742
R219 VDD.n160 VDD.n159 39.742
R220 VDD.n217 VDD.n216 39.742
R221 VDD.n261 VDD.n260 39.742
R222 VDD.n318 VDD.n317 39.742
R223 VDD.n362 VDD.n361 39.742
R224 VDD.n667 VDD.n666 39.742
R225 VDD.n612 VDD.n611 39.742
R226 VDD.n584 VDD.n583 39.742
R227 VDD.n524 VDD.n523 39.742
R228 VDD.n469 VDD.n468 39.742
R229 VDD.n385 VDD.n384 39.742
R230 VDD.n419 VDD.n416 39.742
R231 VDD.n419 VDD.n418 39.742
R232 VDD.n415 VDD.n414 39.742
R233 VDD.n101 VDD.n100 38
R234 VDD.n145 VDD.n144 38
R235 VDD.n202 VDD.n201 38
R236 VDD.n246 VDD.n245 38
R237 VDD.n303 VDD.n302 38
R238 VDD.n347 VDD.n346 38
R239 VDD.n676 VDD.n675 38
R240 VDD.n621 VDD.n620 38
R241 VDD.n569 VDD.n568 38
R242 VDD.n533 VDD.n532 38
R243 VDD.n478 VDD.n477 38
R244 VDD.n372 VDD.n371 38
R245 VDD.n476 VDD.n475 36.774
R246 VDD.n531 VDD.n530 36.774
R247 VDD.n567 VDD.n566 36.774
R248 VDD.n619 VDD.n618 36.774
R249 VDD.n674 VDD.n673 36.774
R250 VDD.n345 VDD.n344 36.774
R251 VDD.n301 VDD.n300 36.774
R252 VDD.n244 VDD.n243 36.774
R253 VDD.n200 VDD.n199 36.774
R254 VDD.n143 VDD.n142 36.774
R255 VDD.n99 VDD.n98 36.774
R256 VDD.n57 VDD.n56 36.774
R257 VDD.n418 VDD.n417 36.774
R258 VDD.n1 VDD.n0 30.923
R259 VDD.n64 VDD.n62 26.38
R260 VDD.n64 VDD.n61 26.38
R261 VDD.n64 VDD.n59 26.38
R262 VDD.n64 VDD.n63 26.38
R263 VDD.n119 VDD.n117 26.38
R264 VDD.n119 VDD.n116 26.38
R265 VDD.n119 VDD.n118 26.38
R266 VDD.n163 VDD.n161 26.38
R267 VDD.n163 VDD.n160 26.38
R268 VDD.n163 VDD.n162 26.38
R269 VDD.n220 VDD.n218 26.38
R270 VDD.n220 VDD.n217 26.38
R271 VDD.n220 VDD.n219 26.38
R272 VDD.n264 VDD.n262 26.38
R273 VDD.n264 VDD.n261 26.38
R274 VDD.n264 VDD.n263 26.38
R275 VDD.n321 VDD.n319 26.38
R276 VDD.n321 VDD.n318 26.38
R277 VDD.n321 VDD.n320 26.38
R278 VDD.n365 VDD.n363 26.38
R279 VDD.n365 VDD.n362 26.38
R280 VDD.n365 VDD.n364 26.38
R281 VDD.n670 VDD.n668 26.38
R282 VDD.n670 VDD.n667 26.38
R283 VDD.n670 VDD.n669 26.38
R284 VDD.n615 VDD.n613 26.38
R285 VDD.n615 VDD.n612 26.38
R286 VDD.n615 VDD.n614 26.38
R287 VDD.n587 VDD.n585 26.38
R288 VDD.n587 VDD.n584 26.38
R289 VDD.n587 VDD.n586 26.38
R290 VDD.n527 VDD.n525 26.38
R291 VDD.n527 VDD.n524 26.38
R292 VDD.n527 VDD.n526 26.38
R293 VDD.n472 VDD.n470 26.38
R294 VDD.n472 VDD.n469 26.38
R295 VDD.n472 VDD.n471 26.38
R296 VDD.n388 VDD.n386 26.38
R297 VDD.n388 VDD.n385 26.38
R298 VDD.n388 VDD.n387 26.38
R299 VDD.n420 VDD.n419 26.38
R300 VDD.n420 VDD.n415 26.38
R301 VDD.n420 VDD.n413 26.38
R302 VDD.n420 VDD.n412 26.38
R303 VDD.n391 VDD.n383 22.915
R304 VDD.n23 VDD.n14 22.915
R305 VDD.n73  |�� 20.457
R306 VDD.n173 �{�� 20.457
R307 VDD.n274  |�� 20.457
R308 VDD.n708  |�� 20.457
R309 VDD.n653  |�� 20.457
R310 VDD.n510 �{�� 20.457
R311 VDD.n455 �{�� 20.457
R312 VDD.n86  |�� 17.9
R313 VDD.n186  |�� 17.9
R314 VDD.n287  |�� 17.9
R315 VDD.n697 �{�� 17.9
R316 VDD.n642  |�� 17.9
R317 VDD.n499 �{�� 17.9
R318 VDD.n444  |�� 17.9
R319 VDD.n383 VDD.n381 14.864
R320 VDD.n381 VDD.n379 14.864
R321 VDD.n379 VDD.n377 14.864
R322 VDD.n377 VDD.n375 14.864
R323 VDD.n375 VDD.n373 14.864
R324 VDD.n489 VDD.n487 14.864
R325 VDD.n487 VDD.n485 14.864
R326 VDD.n485 VDD.n483 14.864
R327 VDD.n483 VDD.n481 14.864
R328 VDD.n481 VDD.n479 14.864
R329 VDD.n544 VDD.n542 14.864
R330 VDD.n542 VDD.n540 14.864
R331 VDD.n540 VDD.n538 14.864
R332 VDD.n538 VDD.n536 14.864
R333 VDD.n536 VDD.n534 14.864
R334 VDD.n580 VDD.n578 14.864
R335 VDD.n578 VDD.n576 14.864
R336 VDD.n576 VDD.n574 14.864
R337 VDD.n574 VDD.n572 14.864
R338 VDD.n572 VDD.n570 14.864
R339 VDD.n632 VDD.n630 14.864
R340 VDD.n630 VDD.n628 14.864
R341 VDD.n628 VDD.n626 14.864
R342 VDD.n626 VDD.n624 14.864
R343 VDD.n624 VDD.n622 14.864
R344 VDD.n687 VDD.n685 14.864
R345 VDD.n685 VDD.n683 14.864
R346 VDD.n683 VDD.n681 14.864
R347 VDD.n681 VDD.n679 14.864
R348 VDD.n679 VDD.n677 14.864
R349 VDD.n358 VDD.n356 14.864
R350 VDD.n356 VDD.n354 14.864
R351 VDD.n354 VDD.n352 14.864
R352 VDD.n352 VDD.n350 14.864
R353 VDD.n350 VDD.n348 14.864
R354 VDD.n314 VDD.n312 14.864
R355 VDD.n312 VDD.n310 14.864
R356 VDD.n310 VDD.n308 14.864
R357 VDD.n308 VDD.n306 14.864
R358 VDD.n306 VDD.n304 14.864
R359 VDD.n257 VDD.n255 14.864
R360 VDD.n255 VDD.n253 14.864
R361 VDD.n253 VDD.n251 14.864
R362 VDD.n251 VDD.n249 14.864
R363 VDD.n249 VDD.n247 14.864
R364 VDD.n213 VDD.n211 14.864
R365 VDD.n211 VDD.n209 14.864
R366 VDD.n209 VDD.n207 14.864
R367 VDD.n207 VDD.n205 14.864
R368 VDD.n205 VDD.n203 14.864
R369 VDD.n156 VDD.n154 14.864
R370 VDD.n154 VDD.n152 14.864
R371 VDD.n152 VDD.n150 14.864
R372 VDD.n150 VDD.n148 14.864
R373 VDD.n148 VDD.n146 14.864
R374 VDD.n112 VDD.n110 14.864
R375 VDD.n110 VDD.n108 14.864
R376 VDD.n108 VDD.n106 14.864
R377 VDD.n106 VDD.n104 14.864
R378 VDD.n104 VDD.n102 14.864
R379 VDD.n53 VDD.n51 14.864
R380 VDD.n51 VDD.n49 14.864
R381 VDD.n49 VDD.n47 14.864
R382 VDD.n47 VDD.n45 14.864
R383 VDD.n45 VDD.n43 14.864
R384 VDD.n43 VDD.n42 14.864
R385 VDD.n434 VDD.n432 14.864
R386 VDD.n432 VDD.n430 14.864
R387 VDD.n430 VDD.n428 14.864
R388 VDD.n428 VDD.n426 14.864
R389 VDD.n426 VDD.n424 14.864
R390 VDD.n424 VDD.n423 14.864
R391 VDD.n14 VDD.n13 14.864
R392 VDD.n13 VDD.n11 14.864
R393 VDD.n11 VDD.n9 14.864
R394 VDD.n9 VDD.n7 14.864
R395 VDD.n7 VDD.n5 14.864
R396 VDD.n67 VDD.n54 14.864
R397 VDD.n122 VDD.n113 14.864
R398 VDD.n166 VDD.n157 14.864
R399 VDD.n223 VDD.n214 14.864
R400 VDD.n267 VDD.n258 14.864
R401 VDD.n324 VDD.n315 14.864
R402 VDD.n368 VDD.n359 14.864
R403 VDD.n689 VDD.n688 14.864
R404 VDD.n634 VDD.n633 14.864
R405 VDD.n590 VDD.n581 14.864
R406 VDD.n546 VDD.n545 14.864
R407 VDD.n491 VDD.n490 14.864
R408 VDD.n436 VDD.n435 14.864
R409 VDD.n442 VDD.t38 14.282
R410 VDD.n442 VDD.t40 14.282
R411 VDD.n497 VDD.t34 14.282
R412 VDD.n497 VDD.t32 14.282
R413 VDD.n640 VDD.t12 14.282
R414 VDD.n640 VDD.t6 14.282
R415 VDD.n695 VDD.t59 14.282
R416 VDD.n695 VDD.t18 14.282
R417 VDD.n278 VDD.t8 14.282
R418 VDD.n278 VDD.t71 14.282
R419 VDD.n178 VDD.t4 14.282
R420 VDD.n178 VDD.t69 14.282
R421 VDD.n84 VDD.t57 14.282
R422 VDD.n84 VDD.t36 14.282
R423 VDD.n180 VDD.n179 9.083
R424 VDD.n281 VDD.n279 9.083
R425 VDD.n23 VDD.n22 8.855
R426 VDD.n22 VDD.n21 8.855
R427 VDD.n27 VDD.n26 8.855
R428 VDD.n26 VDD.n25 8.855
R429 VDD.n31 VDD.n30 8.855
R430 VDD.n30 VDD.n29 8.855
R431 VDD.n36 VDD.n34 8.855
R432 VDD.n34 VDD.n33 8.855
R433 VDD.n40 VDD.n39 8.855
R434 VDD.n39 VDD.n38 8.855
R435 VDD.n67 VDD.n66 8.855
R436 VDD.n66 VDD.n65 8.855
R437 VDD.n71 VDD.n70 8.855
R438 VDD.n70 VDD.n69 8.855
R439 VDD.n75 VDD.n74 8.855
R440 VDD.n74 VDD.n73 8.855
R441 VDD.n78 VDD.n77 8.855
R442 VDD.n77  |�� 8.855
R443 VDD.n82 VDD.n81 8.855
R444 VDD.n81 VDD.n80 8.855
R445 VDD.n88 VDD.n87 8.855
R446 VDD.n87 VDD.n86 8.855
R447 VDD.n92 VDD.n91 8.855
R448 VDD.n91 VDD.n90 8.855
R449 VDD.n96 VDD.n95 8.855
R450 VDD.n95 VDD.n94 8.855
R451 VDD.n122 VDD.n121 8.855
R452 VDD.n121 VDD.n120 8.855
R453 VDD.n127 VDD.n126 8.855
R454 VDD.n126 VDD.n125 8.855
R455 VDD.n131 VDD.n130 8.855
R456 VDD.n130 VDD.n129 8.855
R457 VDD.n136 VDD.n135 8.855
R458 VDD.n135 VDD.n134 8.855
R459 VDD.n140 VDD.n139 8.855
R460 VDD.n139 VDD.n138 8.855
R461 VDD.n166 VDD.n165 8.855
R462 VDD.n165 VDD.n164 8.855
R463 VDD.n171 VDD.n169 8.855
R464 VDD.n169 VDD.n168 8.855
R465 VDD.n175 VDD.n174 8.855
R466 VDD.n174 VDD.n173 8.855
R467 VDD.n180 VDD.n177 8.855
R468 VDD.n177  |�� 8.855
R469 VDD.n184 VDD.n183 8.855
R470 VDD.n183 VDD.n182 8.855
R471 VDD.n188 VDD.n187 8.855
R472 VDD.n187 VDD.n186 8.855
R473 VDD.n193 VDD.n192 8.855
R474 VDD.n192 VDD.n191 8.855
R475 VDD.n197 VDD.n196 8.855
R476 VDD.n196 VDD.n195 8.855
R477 VDD.n223 VDD.n222 8.855
R478 VDD.n222 VDD.n221 8.855
R479 VDD.n228 VDD.n227 8.855
R480 VDD.n227 VDD.n226 8.855
R481 VDD.n232 VDD.n231 8.855
R482 VDD.n231 VDD.n230 8.855
R483 VDD.n237 VDD.n235 8.855
R484 VDD.n235 VDD.n234 8.855
R485 VDD.n241 VDD.n240 8.855
R486 VDD.n240 VDD.n239 8.855
R487 VDD.n267 VDD.n266 8.855
R488 VDD.n266 VDD.n265 8.855
R489 VDD.n272 VDD.n271 8.855
R490 VDD.n271 VDD.n270 8.855
R491 VDD.n276 VDD.n275 8.855
R492 VDD.n275 VDD.n274 8.855
R493 VDD.n281 VDD.n280 8.855
R494 VDD.n280  |�� 8.855
R495 VDD.n285 VDD.n284 8.855
R496 VDD.n284 VDD.n283 8.855
R497 VDD.n289 VDD.n288 8.855
R498 VDD.n288 VDD.n287 8.855
R499 VDD.n294 VDD.n293 8.855
R500 VDD.n293 VDD.n292 8.855
R501 VDD.n298 VDD.n297 8.855
R502 VDD.n297 VDD.n296 8.855
R503 VDD.n324 VDD.n323 8.855
R504 VDD.n323 VDD.n322 8.855
R505 VDD.n329 VDD.n328 8.855
R506 VDD.n328 VDD.n327 8.855
R507 VDD.n333 VDD.n332 8.855
R508 VDD.n332 VDD.n331 8.855
R509 VDD.n338 VDD.n337 8.855
R510 VDD.n337 VDD.n336 8.855
R511 VDD.n342 VDD.n341 8.855
R512 VDD.n341 VDD.n340 8.855
R513 VDD.n368 VDD.n367 8.855
R514 VDD.n367 VDD.n366 8.855
R515 VDD.n714 VDD.n713 8.855
R516 VDD.n713 VDD.n712 8.855
R517 VDD.n710 VDD.n709 8.855
R518 VDD.n709 VDD.n708 8.855
R519 VDD.n706 VDD.n705 8.855
R520 VDD.n705  |�� 8.855
R521 VDD.n703 VDD.n702 8.855
R522 VDD.n702 VDD.n701 8.855
R523 VDD.n699 VDD.n698 8.855
R524 VDD.n698 VDD.n697 8.855
R525 VDD.n693 VDD.n692 8.855
R526 VDD.n692 VDD.n691 8.855
R527 VDD.n689 VDD.n672 8.855
R528 VDD.n672 VDD.n671 8.855
R529 VDD.n663 VDD.n662 8.855
R530 VDD.n662 VDD.n661 8.855
R531 VDD.n659 VDD.n658 8.855
R532 VDD.n658 VDD.n657 8.855
R533 VDD.n655 VDD.n654 8.855
R534 VDD.n654 VDD.n653 8.855
R535 VDD.n651 VDD.n650 8.855
R536 VDD.n650  |�� 8.855
R537 VDD.n648 VDD.n647 8.855
R538 VDD.n647 VDD.n646 8.855
R539 VDD.n644 VDD.n643 8.855
R540 VDD.n643 VDD.n642 8.855
R541 VDD.n638 VDD.n637 8.855
R542 VDD.n637 VDD.n636 8.855
R543 VDD.n634 VDD.n617 8.855
R544 VDD.n617 VDD.n616 8.855
R545 VDD.n608 VDD.n607 8.855
R546 VDD.n607 VDD.n606 8.855
R547 VDD.n604 VDD.n603 8.855
R548 VDD.n603 VDD.n602 8.855
R549 VDD.n599 VDD.n598 8.855
R550 VDD.n598 VDD.n597 8.855
R551 VDD.n595 VDD.n593 8.855
R552 VDD.n593 VDD.n592 8.855
R553 VDD.n590 VDD.n589 8.855
R554 VDD.n589 VDD.n588 8.855
R555 VDD.n564 VDD.n563 8.855
R556 VDD.n563 VDD.n562 8.855
R557 VDD.n560 VDD.n559 8.855
R558 VDD.n559 VDD.n558 8.855
R559 VDD.n555 VDD.n554 8.855
R560 VDD.n554 VDD.n553 8.855
R561 VDD.n551 VDD.n550 8.855
R562 VDD.n550 VDD.n549 8.855
R563 VDD.n546 VDD.n529 8.855
R564 VDD.n529 VDD.n528 8.855
R565 VDD.n520 VDD.n519 8.855
R566 VDD.n519 VDD.n518 8.855
R567 VDD.n516 VDD.n515 8.855
R568 VDD.n515 VDD.n514 8.855
R569 VDD.n512 VDD.n511 8.855
R570 VDD.n511 VDD.n510 8.855
R571 VDD.n508 VDD.n507 8.855
R572 VDD.n507 �{�� 8.855
R573 VDD.n505 VDD.n504 8.855
R574 VDD.n504 VDD.n503 8.855
R575 VDD.n501 VDD.n500 8.855
R576 VDD.n500 VDD.n499 8.855
R577 VDD.n495 VDD.n494 8.855
R578 VDD.n494 VDD.n493 8.855
R579 VDD.n491 VDD.n474 8.855
R580 VDD.n474 VDD.n473 8.855
R581 VDD.n465 VDD.n464 8.855
R582 VDD.n464 VDD.n463 8.855
R583 VDD.n461 VDD.n460 8.855
R584 VDD.n460 VDD.n459 8.855
R585 VDD.n457 VDD.n456 8.855
R586 VDD.n456 VDD.n455 8.855
R587 VDD.n453 VDD.n452 8.855
R588 VDD.n452 �{�� 8.855
R589 VDD.n450 VDD.n449 8.855
R590 VDD.n449 VDD.n448 8.855
R591 VDD.n446 VDD.n445 8.855
R592 VDD.n445 VDD.n444 8.855
R593 VDD.n440 VDD.n439 8.855
R594 VDD.n439 VDD.n438 8.855
R595 VDD.n436 VDD.n422 8.855
R596 VDD.n422 VDD.n421 8.855
R597 VDD.n409 VDD.n408 8.855
R598 VDD.n408 VDD.n407 8.855
R599 VDD.n405 VDD.n404 8.855
R600 VDD.n404 VDD.n403 8.855
R601 VDD.n400 VDD.n399 8.855
R602 VDD.n399 VDD.n398 8.855
R603 VDD.n396 VDD.n394 8.855
R604 VDD.n394 VDD.n393 8.855
R605 VDD.n391 VDD.n390 8.855
R606 VDD.n390 VDD.n389 8.855
R607 VDD.n490 VDD.n489 8.051
R608 VDD.n545 VDD.n544 8.051
R609 VDD.n581 VDD.n580 8.051
R610 VDD.n633 VDD.n632 8.051
R611 VDD.n688 VDD.n687 8.051
R612 VDD.n359 VDD.n358 8.051
R613 VDD.n315 VDD.n314 8.051
R614 VDD.n258 VDD.n257 8.051
R615 VDD.n214 VDD.n213 8.051
R616 VDD.n157 VDD.n156 8.051
R617 VDD.n113 VDD.n112 8.051
R618 VDD.n54 VDD.n53 8.051
R619 VDD.n435 VDD.n434 8.051
R620 VDD.n88 VDD.n85 6.193
R621 VDD.n699 VDD.n696 6.193
R622 VDD.n644 VDD.n641 6.193
R623 VDD.n501 VDD.n498 6.193
R624 VDD.n446 VDD.n443 6.193
R625 VDD.n28 VDD.n23 4.795
R626 VDD.n28 VDD.n27 4.65
R627 VDD.n32 VDD.n31 4.65
R628 VDD.n37 VDD.n36 4.65
R629 VDD.n41 VDD.n40 4.65
R630 VDD.n68 VDD.n67 4.65
R631 VDD.n72 VDD.n71 4.65
R632 VDD.n76 VDD.n75 4.65
R633 VDD.n79 VDD.n78 4.65
R634 VDD.n83 VDD.n82 4.65
R635 VDD.n89 VDD.n88 4.65
R636 VDD.n93 VDD.n92 4.65
R637 VDD.n97 VDD.n96 4.65
R638 VDD.n123 VDD.n122 4.65
R639 VDD.n128 VDD.n127 4.65
R640 VDD.n132 VDD.n131 4.65
R641 VDD.n137 VDD.n136 4.65
R642 VDD.n141 VDD.n140 4.65
R643 VDD.n167 VDD.n166 4.65
R644 VDD.n172 VDD.n171 4.65
R645 VDD.n176 VDD.n175 4.65
R646 VDD.n181 VDD.n180 4.65
R647 VDD.n185 VDD.n184 4.65
R648 VDD.n189 VDD.n188 4.65
R649 VDD.n194 VDD.n193 4.65
R650 VDD.n198 VDD.n197 4.65
R651 VDD.n224 VDD.n223 4.65
R652 VDD.n229 VDD.n228 4.65
R653 VDD.n233 VDD.n232 4.65
R654 VDD.n238 VDD.n237 4.65
R655 VDD.n242 VDD.n241 4.65
R656 VDD.n268 VDD.n267 4.65
R657 VDD.n273 VDD.n272 4.65
R658 VDD.n277 VDD.n276 4.65
R659 VDD.n282 VDD.n281 4.65
R660 VDD.n286 VDD.n285 4.65
R661 VDD.n290 VDD.n289 4.65
R662 VDD.n295 VDD.n294 4.65
R663 VDD.n299 VDD.n298 4.65
R664 VDD.n325 VDD.n324 4.65
R665 VDD.n330 VDD.n329 4.65
R666 VDD.n334 VDD.n333 4.65
R667 VDD.n339 VDD.n338 4.65
R668 VDD.n343 VDD.n342 4.65
R669 VDD.n369 VDD.n368 4.65
R670 VDD.n715 VDD.n714 4.65
R671 VDD.n711 VDD.n710 4.65
R672 VDD.n707 VDD.n706 4.65
R673 VDD.n704 VDD.n703 4.65
R674 VDD.n700 VDD.n699 4.65
R675 VDD.n694 VDD.n693 4.65
R676 VDD.n690 VDD.n689 4.65
R677 VDD.n664 VDD.n663 4.65
R678 VDD.n660 VDD.n659 4.65
R679 VDD.n656 VDD.n655 4.65
R680 VDD.n652 VDD.n651 4.65
R681 VDD.n649 VDD.n648 4.65
R682 VDD.n645 VDD.n644 4.65
R683 VDD.n639 VDD.n638 4.65
R684 VDD.n635 VDD.n634 4.65
R685 VDD.n609 VDD.n608 4.65
R686 VDD.n605 VDD.n604 4.65
R687 VDD.n600 VDD.n599 4.65
R688 VDD.n596 VDD.n595 4.65
R689 VDD.n591 VDD.n590 4.65
R690 VDD.n565 VDD.n564 4.65
R691 VDD.n561 VDD.n560 4.65
R692 VDD.n556 VDD.n555 4.65
R693 VDD.n552 VDD.n551 4.65
R694 VDD.n547 VDD.n546 4.65
R695 VDD.n521 VDD.n520 4.65
R696 VDD.n517 VDD.n516 4.65
R697 VDD.n513 VDD.n512 4.65
R698 VDD.n509 VDD.n508 4.65
R699 VDD.n506 VDD.n505 4.65
R700 VDD.n502 VDD.n501 4.65
R701 VDD.n496 VDD.n495 4.65
R702 VDD.n492 VDD.n491 4.65
R703 VDD.n466 VDD.n465 4.65
R704 VDD.n462 VDD.n461 4.65
R705 VDD.n458 VDD.n457 4.65
R706 VDD.n454 VDD.n453 4.65
R707 VDD.n451 VDD.n450 4.65
R708 VDD.n447 VDD.n446 4.65
R709 VDD.n441 VDD.n440 4.65
R710 VDD.n437 VDD.n436 4.65
R711 VDD.n410 VDD.n409 4.65
R712 VDD.n406 VDD.n405 4.65
R713 VDD.n401 VDD.n400 4.65
R714 VDD.n397 VDD.n396 4.65
R715 VDD.n392 VDD.n391 4.65
R716 VDD.n193 VDD.n190 2.89
R717 VDD.n294 VDD.n291 2.89
R718 VDD.n80 �{�� 2.557
R719 VDD.n182 �{�� 2.557
R720 VDD.n283 �{�� 2.557
R721 VDD.n701  |�� 2.557
R722 VDD.n646  |�� 2.557
R723 VDD.n503 �{�� 2.557
R724 VDD.n448  |�� 2.557
R725 VDD.n171 VDD.n170 2.477
R726 VDD.n272 VDD.n269 2.477
R727 VDD.n27 VDD.n24 2.064
R728 VDD.n36 VDD.n35 2.064
R729 VDD.n127 VDD.n124 2.064
R730 VDD.n136 VDD.n133 2.064
R731 VDD.n228 VDD.n225 2.064
R732 VDD.n237 VDD.n236 2.064
R733 VDD.n329 VDD.n326 2.064
R734 VDD.n338 VDD.n335 2.064
R735 VDD.n604 VDD.n601 2.064
R736 VDD.n595 VDD.n594 2.064
R737 VDD.n560 VDD.n557 2.064
R738 VDD.n551 VDD.n548 2.064
R739 VDD.n405 VDD.n402 2.064
R740 VDD.n396 VDD.n395 2.064
R741 VDD.n68 VDD.n41 0.29
R742 VDD.n123 VDD.n97 0.29
R743 VDD.n167 VDD.n141 0.29
R744 VDD.n224 VDD.n198 0.29
R745 VDD.n268 VDD.n242 0.29
R746 VDD.n325 VDD.n299 0.29
R747 VDD.n369 VDD.n343 0.29
R748 VDD.n690 VDD.n664 0.29
R749 VDD.n635 VDD.n609 0.29
R750 VDD.n591 VDD.n565 0.29
R751 VDD.n547 VDD.n521 0.29
R752 VDD.n492 VDD.n466 0.29
R753 VDD.n437 VDD.n410 0.29
R754 VDD.n392 VDD 0.207
R755 VDD.n83 VDD.n79 0.181
R756 VDD.n185 VDD.n181 0.181
R757 VDD.n286 VDD.n282 0.181
R758 VDD.n707 VDD.n704 0.181
R759 VDD.n652 VDD.n649 0.181
R760 VDD.n509 VDD.n506 0.181
R761 VDD.n454 VDD.n451 0.181
R762 VDD.n32 VDD.n28 0.157
R763 VDD.n37 VDD.n32 0.157
R764 VDD.n132 VDD.n128 0.157
R765 VDD.n137 VDD.n132 0.157
R766 VDD.n233 VDD.n229 0.157
R767 VDD.n238 VDD.n233 0.157
R768 VDD.n334 VDD.n330 0.157
R769 VDD.n339 VDD.n334 0.157
R770 VDD.n605 VDD.n600 0.157
R771 VDD.n600 VDD.n596 0.157
R772 VDD.n561 VDD.n556 0.157
R773 VDD.n556 VDD.n552 0.157
R774 VDD.n406 VDD.n401 0.157
R775 VDD.n401 VDD.n397 0.157
R776 VDD.n41 VDD.n37 0.145
R777 VDD.n72 VDD.n68 0.145
R778 VDD.n76 VDD.n72 0.145
R779 VDD.n79 VDD.n76 0.145
R780 VDD.n89 VDD.n83 0.145
R781 VDD.n93 VDD.n89 0.145
R782 VDD.n97 VDD.n93 0.145
R783 VDD.n128 VDD.n123 0.145
R784 VDD.n141 VDD.n137 0.145
R785 VDD.n172 VDD.n167 0.145
R786 VDD.n176 VDD.n172 0.145
R787 VDD.n181 VDD.n176 0.145
R788 VDD.n189 VDD.n185 0.145
R789 VDD.n194 VDD.n189 0.145
R790 VDD.n198 VDD.n194 0.145
R791 VDD.n229 VDD.n224 0.145
R792 VDD.n242 VDD.n238 0.145
R793 VDD.n273 VDD.n268 0.145
R794 VDD.n277 VDD.n273 0.145
R795 VDD.n282 VDD.n277 0.145
R796 VDD.n290 VDD.n286 0.145
R797 VDD.n295 VDD.n290 0.145
R798 VDD.n299 VDD.n295 0.145
R799 VDD.n330 VDD.n325 0.145
R800 VDD.n343 VDD.n339 0.145
R801 VDD.n715 VDD.n711 0.145
R802 VDD.n711 VDD.n707 0.145
R803 VDD.n704 VDD.n700 0.145
R804 VDD.n700 VDD.n694 0.145
R805 VDD.n694 VDD.n690 0.145
R806 VDD.n664 VDD.n660 0.145
R807 VDD.n660 VDD.n656 0.145
R808 VDD.n656 VDD.n652 0.145
R809 VDD.n649 VDD.n645 0.145
R810 VDD.n645 VDD.n639 0.145
R811 VDD.n639 VDD.n635 0.145
R812 VDD.n609 VDD.n605 0.145
R813 VDD.n596 VDD.n591 0.145
R814 VDD.n565 VDD.n561 0.145
R815 VDD.n552 VDD.n547 0.145
R816 VDD.n521 VDD.n517 0.145
R817 VDD.n517 VDD.n513 0.145
R818 VDD.n513 VDD.n509 0.145
R819 VDD.n506 VDD.n502 0.145
R820 VDD.n502 VDD.n496 0.145
R821 VDD.n496 VDD.n492 0.145
R822 VDD.n466 VDD.n462 0.145
R823 VDD.n462 VDD.n458 0.145
R824 VDD.n458 VDD.n454 0.145
R825 VDD.n451 VDD.n447 0.145
R826 VDD.n447 VDD.n441 0.145
R827 VDD.n441 VDD.n437 0.145
R828 VDD.n410 VDD.n406 0.145
R829 VDD.n397 VDD.n392 0.145
R830 VDD VDD.n369 0.078
R831 VDD VDD.n715 0.066
R832 CIN.n2 CIN.t1 512.525
R833 CIN.n0 CIN.t8 480.392
R834 CIN.n5 CIN.t7 480.392
R835 CIN.n1 CIN.t6 412.921
R836 CIN.n0 CIN.t3 403.272
R837 CIN.n5 CIN.t2 403.272
R838 CIN.n2 CIN.t5 371.139
R839 CIN.n3 CIN.t0 299.455
R840 CIN.n3 CIN.t4 227.134
R841 CIN.n4 CIN.n2 163.771
R842 CIN.n4 CIN.n3 139.294
R843 CIN.n6 CIN.n5 123.272
R844 CIN.n1 CIN.n0 115.571
R845 CIN.n6 CIN.n4 4.65
R846 CIN.n7 CIN.n1 4.65
R847 CIN CIN.n6 1.269
R848 CIN.n7 CIN 0.046
R849 a_2776_101.t0 a_2776_101.n6 93.333
R850 a_2776_101.n5 a_2776_101.n4 51.907
R851 a_2776_101.n5 a_2776_101.n3 51.594
R852 a_2776_101.n2 a_2776_101.n0 41.528
R853 a_2776_101.t0 a_2776_101.n5 38.864
R854 a_2776_101.t0 a_2776_101.n7 8.137
R855 a_2776_101.n2 a_2776_101.n1 3.644
R856 a_2776_101.t0 a_2776_101.n2 1.093
R857 SUM.n8 SUM.n7 327.32
R858 SUM.n5 SUM.n4 305.581
R859 SUM.n5 SUM.n0 260.107
R860 SUM.n8 SUM.n6 260.107
R861 SUM.n4 SUM.n3 30
R862 SUM.n2 SUM.n1 24.383
R863 SUM.n4 SUM.n2 23.684
R864 SUM.n0 SUM.t4 14.282
R865 SUM.n0 SUM.t3 14.282
R866 SUM.n6 SUM.t1 14.282
R867 SUM.n6 SUM.t0 14.282
R868 SUM SUM.n8 7.007
R869 SUM.n9 SUM.n5 4.65
R870 SUM.n9 SUM 0.046
R871 GND.n271 GND.n270 237.558
R872 GND.n301 GND.n300 237.558
R873 GND.n331 GND.n330 237.558
R874 GND.n361 GND.n360 237.558
R875 GND.n394 GND.n393 237.558
R876 GND.n238 GND.n237 237.558
R877 GND.n424 GND.n423 237.558
R878 GND.n206 GND.n205 237.558
R879 GND.n173 GND.n172 237.558
R880 GND.n140 GND.n139 237.558
R881 GND.n110 GND.n109 237.558
R882 GND.n77 GND.n76 237.558
R883 GND.n32 GND.n31 237.558
R884 GND.n29 GND.n28 210.82
R885 GND.n273 GND.n272 210.82
R886 GND.n303 GND.n302 210.82
R887 GND.n333 GND.n332 210.82
R888 GND.n363 GND.n362 210.82
R889 GND.n396 GND.n395 210.82
R890 GND.n426 GND.n425 210.82
R891 GND.n235 GND.n234 210.82
R892 GND.n203 GND.n202 210.82
R893 GND.n170 GND.n169 210.82
R894 GND.n137 GND.n136 210.82
R895 GND.n107 GND.n106 210.82
R896 GND.n74 GND.n73 210.82
R897 GND.n126 GND.n125 172.612
R898 GND.n434 GND.n433 172.612
R899 GND.n404 GND.n403 172.612
R900 GND.n311 GND.n310 172.612
R901 GND.n281 GND.n280 172.612
R902 GND.n192 GND.n191 151.605
R903 GND.n44 GND.n43 92.5
R904 GND.n219 GND.n218 92.5
R905 GND.n210 GND.t14 45.414
R906 GND.n53 GND.n52 40.431
R907 GND.n226 GND.n225 40.414
R908 GND.n210 GND.n209 39.307
R909 GND.n340 GND.n339 38.384
R910 GND.n21 GND.n20 37.582
R911 GND.n66 GND.n65 37.582
R912 GND.n99 GND.n98 37.582
R913 GND.n162 GND.n161 37.582
R914 GND.n374 GND.n373 37.582
R915 GND.n251 GND.n250 37.582
R916 GND.n36 GND.n35 35.865
R917 GND.n352 GND.n351 34.159
R918 GND.t19 GND.n18 32.601
R919 GND.t9 GND.n96 32.601
R920 GND.t20 GND.n159 32.601
R921 GND.t2 GND.n371 32.601
R922 GND.t8 GND.n248 32.601
R923 GND.n37 GND.n36 28.503
R924 GND.n191 GND.n190 28.421
R925 GND.n191 GND.n189 25.263
R926 GND.n189 GND.n188 24.383
R927 GND.n227 GND.n226 23.961
R928 GND.n211 GND.n210 23.77
R929 GND.n18 GND.n17 21.734
R930 GND.n96 GND.n95 21.734
R931 GND.n159 GND.n158 21.734
R932 GND.n371 GND.n370 21.734
R933 GND.n248 GND.n247 21.734
R934 GND.n4 GND.n3 20.705
R935 GND.n10 GND.n9 20.705
R936 GND.n22 GND.n21 20.705
R937 GND.n59 GND.n58 20.705
R938 GND.n54 GND.n53 20.705
R939 GND.n45 GND.n44 20.705
R940 GND.n38 GND.n37 20.705
R941 GND.n67 GND.n66 20.705
R942 GND.n82 GND.n81 20.705
R943 GND.n88 GND.n87 20.705
R944 GND.n100 GND.n99 20.705
R945 GND.n145 GND.n144 20.705
R946 GND.n151 GND.n150 20.705
R947 GND.n163 GND.n162 20.705
R948 GND.n212 GND.n211 20.705
R949 GND.n221 GND.n220 20.705
R950 GND.n228 GND.n227 20.705
R951 GND.n386 GND.n385 20.705
R952 GND.n380 GND.n379 20.705
R953 GND.n375 GND.n374 20.705
R954 GND.n353 GND.n352 20.705
R955 GND.n347 GND.n346 20.705
R956 GND.n341 GND.n340 20.705
R957 GND.n263 GND.n262 20.705
R958 GND.n257 GND.n256 20.705
R959 GND.n252 GND.n251 20.705
R960 GND.n3 GND.n2 19.952
R961 GND.n81 GND.n80 19.952
R962 GND.n144 GND.n143 19.952
R963 GND.n385 GND.n384 19.952
R964 GND.n262 GND.n261 19.952
R965 GND.n351 GND.n350 19.926
R966 GND.n30 GND.n29 18.953
R967 GND.n274 GND.n273 18.953
R968 GND.n304 GND.n303 18.953
R969 GND.n334 GND.n333 18.953
R970 GND.n364 GND.n363 18.953
R971 GND.n397 GND.n396 18.953
R972 GND.n427 GND.n426 18.953
R973 GND.n236 GND.n235 18.953
R974 GND.n204 GND.n203 18.953
R975 GND.n171 GND.n170 18.953
R976 GND.n138 GND.n137 18.953
R977 GND.n108 GND.n107 18.953
R978 GND.n75 GND.n74 18.953
R979 GND.n339 GND.t5 15.889
R980 GND.n20 GND.t19 15.644
R981 GND.n65 GND.t17 15.644
R982 GND.n98 GND.t9 15.644
R983 GND.n161 GND.t20 15.644
R984 GND.n373 GND.t2 15.644
R985 GND.n250 GND.t8 15.644
R986 GND.n33 GND.n30 14.864
R987 GND.n78 GND.n75 14.864
R988 GND.n111 GND.n108 14.864
R989 GND.n141 GND.n138 14.864
R990 GND.n174 GND.n171 14.864
R991 GND.n207 GND.n204 14.864
R992 GND.n239 GND.n236 14.864
R993 GND.n428 GND.n427 14.864
R994 GND.n398 GND.n397 14.864
R995 GND.n365 GND.n364 14.864
R996 GND.n335 GND.n334 14.864
R997 GND.n305 GND.n304 14.864
R998 GND.n275 GND.n274 14.864
R999 GND.n52 GND.t18 13.654
R1000 GND.n339 GND.n338 13.624
R1001 GND.n20 GND.n19 13.541
R1002 GND.n65 GND.n64 13.541
R1003 GND.n98 GND.n97 13.541
R1004 GND.n161 GND.n160 13.541
R1005 GND.n373 GND.n372 13.541
R1006 GND.n250 GND.n249 13.541
R1007 GND.n56 GND.n54 9.29
R1008 GND.n253 GND.n244 9.154
R1009 GND.n259 GND.n258 9.154
R1010 GND.n265 GND.n264 9.154
R1011 GND.n268 GND.n267 9.154
R1012 GND.n275 GND.n271 9.154
R1013 GND.n278 GND.n277 9.154
R1014 GND.n283 GND.n282 9.154
R1015 GND.n286 GND.n285 9.154
R1016 GND.n289 GND.n288 9.154
R1017 GND.n292 GND.n291 9.154
R1018 GND.n295 GND.n294 9.154
R1019 GND.n298 GND.n297 9.154
R1020 GND.n305 GND.n301 9.154
R1021 GND.n308 GND.n307 9.154
R1022 GND.n313 GND.n312 9.154
R1023 GND.n316 GND.n315 9.154
R1024 GND.n319 GND.n318 9.154
R1025 GND.n322 GND.n321 9.154
R1026 GND.n325 GND.n324 9.154
R1027 GND.n328 GND.n327 9.154
R1028 GND.n335 GND.n331 9.154
R1029 GND.n342 GND.n337 9.154
R1030 GND.n348 GND.n344 9.154
R1031 GND.n355 GND.n354 9.154
R1032 GND.n358 GND.n357 9.154
R1033 GND.n365 GND.n361 9.154
R1034 GND.n376 GND.n367 9.154
R1035 GND.n382 GND.n381 9.154
R1036 GND.n388 GND.n387 9.154
R1037 GND.n391 GND.n390 9.154
R1038 GND.n398 GND.n394 9.154
R1039 GND.n401 GND.n400 9.154
R1040 GND.n406 GND.n405 9.154
R1041 GND.n409 GND.n408 9.154
R1042 GND.n412 GND.n411 9.154
R1043 GND.n415 GND.n414 9.154
R1044 GND.n418 GND.n417 9.154
R1045 GND.n421 GND.n420 9.154
R1046 GND.n428 GND.n424 9.154
R1047 GND.n431 GND.n430 9.154
R1048 GND.n436 GND.n435 9.154
R1049 GND.n439 GND.n438 9.154
R1050 GND.n442 GND.n441 9.154
R1051 GND.n445 GND.n444 9.154
R1052 GND.n448 GND.n447 9.154
R1053 GND.n239 GND.n238 9.154
R1054 GND.n232 GND.n231 9.154
R1055 GND.n229 GND.n224 9.154
R1056 GND.n222 GND.n216 9.154
R1057 GND.n214 GND.n213 9.154
R1058 GND.n207 GND.n206 9.154
R1059 GND.n200 GND.n199 9.154
R1060 GND.n197 GND.n196 9.154
R1061 GND.n194 GND.n193 9.154
R1062 GND.n186 GND.n185 9.154
R1063 GND.n183 GND.n182 9.154
R1064 GND.n180 GND.n179 9.154
R1065 GND.n177 GND.n176 9.154
R1066 GND.n174 GND.n173 9.154
R1067 GND.n167 GND.n166 9.154
R1068 GND.n164 GND.n155 9.154
R1069 GND.n153 GND.n152 9.154
R1070 GND.n147 GND.n146 9.154
R1071 GND.n141 GND.n140 9.154
R1072 GND.n134 GND.n133 9.154
R1073 GND.n131 GND.n130 9.154
R1074 GND.n128 GND.n127 9.154
R1075 GND.n123 GND.n122 9.154
R1076 GND.n120 GND.n119 9.154
R1077 GND.n117 GND.n116 9.154
R1078 GND.n114 GND.n113 9.154
R1079 GND.n111 GND.n110 9.154
R1080 GND.n104 GND.n103 9.154
R1081 GND.n101 GND.n92 9.154
R1082 GND.n90 GND.n89 9.154
R1083 GND.n84 GND.n83 9.154
R1084 GND.n78 GND.n77 9.154
R1085 GND.n71 GND.n70 9.154
R1086 GND.n68 GND.n63 9.154
R1087 GND.n61 GND.n60 9.154
R1088 GND.n56 GND.n55 9.154
R1089 GND.n49 GND.n48 9.154
R1090 GND.n46 GND.n42 9.154
R1091 GND.n40 GND.n39 9.154
R1092 GND.n33 GND.n32 9.154
R1093 GND.n26 GND.n25 9.154
R1094 GND.n23 GND.n14 9.154
R1095 GND.n12 GND.n11 9.154
R1096 GND.n6 GND.n5 9.154
R1097 GND.t18 GND.n51 7.04
R1098 GND.n7 GND.n1 4.795
R1099 GND.n243 GND.n242 4.65
R1100 GND.n7 GND.n6 4.65
R1101 GND.n13 GND.n12 4.65
R1102 GND.n24 GND.n23 4.65
R1103 GND.n27 GND.n26 4.65
R1104 GND.n34 GND.n33 4.65
R1105 GND.n41 GND.n40 4.65
R1106 GND.n47 GND.n46 4.65
R1107 GND.n50 GND.n49 4.65
R1108 GND.n57 GND.n56 4.65
R1109 GND.n62 GND.n61 4.65
R1110 GND.n69 GND.n68 4.65
R1111 GND.n72 GND.n71 4.65
R1112 GND.n79 GND.n78 4.65
R1113 GND.n85 GND.n84 4.65
R1114 GND.n91 GND.n90 4.65
R1115 GND.n102 GND.n101 4.65
R1116 GND.n105 GND.n104 4.65
R1117 GND.n112 GND.n111 4.65
R1118 GND.n115 GND.n114 4.65
R1119 GND.n118 GND.n117 4.65
R1120 GND.n121 GND.n120 4.65
R1121 GND.n124 GND.n123 4.65
R1122 GND.n129 GND.n128 4.65
R1123 GND.n132 GND.n131 4.65
R1124 GND.n135 GND.n134 4.65
R1125 GND.n142 GND.n141 4.65
R1126 GND.n148 GND.n147 4.65
R1127 GND.n154 GND.n153 4.65
R1128 GND.n165 GND.n164 4.65
R1129 GND.n168 GND.n167 4.65
R1130 GND.n175 GND.n174 4.65
R1131 GND.n178 GND.n177 4.65
R1132 GND.n181 GND.n180 4.65
R1133 GND.n184 GND.n183 4.65
R1134 GND.n187 GND.n186 4.65
R1135 GND.n195 GND.n194 4.65
R1136 GND.n198 GND.n197 4.65
R1137 GND.n201 GND.n200 4.65
R1138 GND.n208 GND.n207 4.65
R1139 GND.n215 GND.n214 4.65
R1140 GND.n223 GND.n222 4.65
R1141 GND.n230 GND.n229 4.65
R1142 GND.n233 GND.n232 4.65
R1143 GND.n240 GND.n239 4.65
R1144 GND.n449 GND.n448 4.65
R1145 GND.n446 GND.n445 4.65
R1146 GND.n443 GND.n442 4.65
R1147 GND.n440 GND.n439 4.65
R1148 GND.n437 GND.n436 4.65
R1149 GND.n432 GND.n431 4.65
R1150 GND.n429 GND.n428 4.65
R1151 GND.n422 GND.n421 4.65
R1152 GND.n419 GND.n418 4.65
R1153 GND.n416 GND.n415 4.65
R1154 GND.n413 GND.n412 4.65
R1155 GND.n410 GND.n409 4.65
R1156 GND.n407 GND.n406 4.65
R1157 GND.n402 GND.n401 4.65
R1158 GND.n399 GND.n398 4.65
R1159 GND.n392 GND.n391 4.65
R1160 GND.n389 GND.n388 4.65
R1161 GND.n383 GND.n382 4.65
R1162 GND.n377 GND.n376 4.65
R1163 GND.n366 GND.n365 4.65
R1164 GND.n359 GND.n358 4.65
R1165 GND.n356 GND.n355 4.65
R1166 GND.n349 GND.n348 4.65
R1167 GND.n343 GND.n342 4.65
R1168 GND.n336 GND.n335 4.65
R1169 GND.n329 GND.n328 4.65
R1170 GND.n326 GND.n325 4.65
R1171 GND.n323 GND.n322 4.65
R1172 GND.n320 GND.n319 4.65
R1173 GND.n317 GND.n316 4.65
R1174 GND.n314 GND.n313 4.65
R1175 GND.n309 GND.n308 4.65
R1176 GND.n306 GND.n305 4.65
R1177 GND.n299 GND.n298 4.65
R1178 GND.n296 GND.n295 4.65
R1179 GND.n293 GND.n292 4.65
R1180 GND.n290 GND.n289 4.65
R1181 GND.n287 GND.n286 4.65
R1182 GND.n284 GND.n283 4.65
R1183 GND.n279 GND.n278 4.65
R1184 GND.n276 GND.n275 4.65
R1185 GND.n269 GND.n268 4.65
R1186 GND.n266 GND.n265 4.65
R1187 GND.n260 GND.n259 4.65
R1188 GND.n254 GND.n253 4.65
R1189 GND.n16 GND.n15 4.504
R1190 GND.n94 GND.n93 4.504
R1191 GND.n157 GND.n156 4.504
R1192 GND.n369 GND.n368 4.504
R1193 GND.n246 GND.n245 4.504
R1194 GND.n6 GND.n4 4.129
R1195 GND.n46 GND.n45 4.129
R1196 GND.n61 GND.n59 4.129
R1197 GND.n84 GND.n82 4.129
R1198 GND.n128 GND.n126 4.129
R1199 GND.n147 GND.n145 4.129
R1200 GND.n194 GND.n192 4.129
R1201 GND.n229 GND.n228 4.129
R1202 GND.n436 GND.n434 4.129
R1203 GND.n406 GND.n404 4.129
R1204 GND.n388 GND.n386 4.129
R1205 GND.n342 GND.n341 4.129
R1206 GND.n313 GND.n311 4.129
R1207 GND.n283 GND.n281 4.129
R1208 GND.n265 GND.n263 4.129
R1209 GND.n23 GND.n22 3.716
R1210 GND.n101 GND.n100 3.716
R1211 GND.n164 GND.n163 3.716
R1212 GND.n214 GND.n212 3.716
R1213 GND.n376 GND.n375 3.716
R1214 GND.n355 GND.n353 3.716
R1215 GND.n253 GND.n252 3.716
R1216 GND.t19 GND.n16 2.452
R1217 GND.t9 GND.n94 2.452
R1218 GND.t20 GND.n157 2.452
R1219 GND.t2 GND.n369 2.452
R1220 GND.t8 GND.n246 2.452
R1221 GND.n218 GND.n217 1.935
R1222 GND.n40 GND.n38 1.032
R1223 GND.n68 GND.n67 1.032
R1224 GND.n1 GND.n0 0.474
R1225 GND.n242 GND.n241 0.474
R1226 GND.n9 GND.n8 0.376
R1227 GND.n87 GND.n86 0.376
R1228 GND.n150 GND.n149 0.376
R1229 GND.n220 GND.n219 0.376
R1230 GND.n379 GND.n378 0.376
R1231 GND.n346 GND.n345 0.376
R1232 GND.n256 GND.n255 0.376
R1233 GND.n34 GND.n27 0.29
R1234 GND.n79 GND.n72 0.29
R1235 GND.n112 GND.n105 0.29
R1236 GND.n142 GND.n135 0.29
R1237 GND.n175 GND.n168 0.29
R1238 GND.n208 GND.n201 0.29
R1239 GND.n240 GND.n233 0.29
R1240 GND.n429 GND.n422 0.29
R1241 GND.n399 GND.n392 0.29
R1242 GND.n366 GND.n359 0.29
R1243 GND.n336 GND.n329 0.29
R1244 GND.n306 GND.n299 0.29
R1245 GND.n276 GND.n269 0.29
R1246 GND.n243 GND 0.207
R1247 GND.n12 GND.n10 0.206
R1248 GND.n90 GND.n88 0.206
R1249 GND.n153 GND.n151 0.206
R1250 GND.n222 GND.n221 0.206
R1251 GND.n382 GND.n380 0.206
R1252 GND.n348 GND.n347 0.206
R1253 GND.n259 GND.n257 0.206
R1254 GND.n57 GND.n50 0.181
R1255 GND.n124 GND.n121 0.181
R1256 GND.n187 GND.n184 0.181
R1257 GND.n443 GND.n440 0.181
R1258 GND.n413 GND.n410 0.181
R1259 GND.n320 GND.n317 0.181
R1260 GND.n290 GND.n287 0.181
R1261 GND.n13 GND.n7 0.157
R1262 GND.n24 GND.n13 0.157
R1263 GND.n91 GND.n85 0.157
R1264 GND.n102 GND.n91 0.157
R1265 GND.n154 GND.n148 0.157
R1266 GND.n165 GND.n154 0.157
R1267 GND.n223 GND.n215 0.157
R1268 GND.n230 GND.n223 0.157
R1269 GND.n389 GND.n383 0.157
R1270 GND.n383 GND.n377 0.157
R1271 GND.n356 GND.n349 0.157
R1272 GND.n349 GND.n343 0.157
R1273 GND.n266 GND.n260 0.157
R1274 GND.n260 GND.n254 0.157
R1275 GND.n27 GND.n24 0.145
R1276 GND.n41 GND.n34 0.145
R1277 GND.n47 GND.n41 0.145
R1278 GND.n50 GND.n47 0.145
R1279 GND.n62 GND.n57 0.145
R1280 GND.n69 GND.n62 0.145
R1281 GND.n72 GND.n69 0.145
R1282 GND.n85 GND.n79 0.145
R1283 GND.n105 GND.n102 0.145
R1284 GND.n115 GND.n112 0.145
R1285 GND.n118 GND.n115 0.145
R1286 GND.n121 GND.n118 0.145
R1287 GND.n129 GND.n124 0.145
R1288 GND.n132 GND.n129 0.145
R1289 GND.n135 GND.n132 0.145
R1290 GND.n148 GND.n142 0.145
R1291 GND.n168 GND.n165 0.145
R1292 GND.n178 GND.n175 0.145
R1293 GND.n181 GND.n178 0.145
R1294 GND.n184 GND.n181 0.145
R1295 GND.n195 GND.n187 0.145
R1296 GND.n198 GND.n195 0.145
R1297 GND.n201 GND.n198 0.145
R1298 GND.n215 GND.n208 0.145
R1299 GND.n233 GND.n230 0.145
R1300 GND.n449 GND.n446 0.145
R1301 GND.n446 GND.n443 0.145
R1302 GND.n440 GND.n437 0.145
R1303 GND.n437 GND.n432 0.145
R1304 GND.n432 GND.n429 0.145
R1305 GND.n422 GND.n419 0.145
R1306 GND.n419 GND.n416 0.145
R1307 GND.n416 GND.n413 0.145
R1308 GND.n410 GND.n407 0.145
R1309 GND.n407 GND.n402 0.145
R1310 GND.n402 GND.n399 0.145
R1311 GND.n392 GND.n389 0.145
R1312 GND.n377 GND.n366 0.145
R1313 GND.n359 GND.n356 0.145
R1314 GND.n343 GND.n336 0.145
R1315 GND.n329 GND.n326 0.145
R1316 GND.n326 GND.n323 0.145
R1317 GND.n323 GND.n320 0.145
R1318 GND.n317 GND.n314 0.145
R1319 GND.n314 GND.n309 0.145
R1320 GND.n309 GND.n306 0.145
R1321 GND.n299 GND.n296 0.145
R1322 GND.n296 GND.n293 0.145
R1323 GND.n293 GND.n290 0.145
R1324 GND.n287 GND.n284 0.145
R1325 GND.n284 GND.n279 0.145
R1326 GND.n279 GND.n276 0.145
R1327 GND.n269 GND.n266 0.145
R1328 GND.n254 GND.n243 0.145
R1329 GND GND.n240 0.078
R1330 GND GND.n449 0.066
R1331 a_4657_1050.n0 a_4657_1050.t6 512.525
R1332 a_4657_1050.n0 a_4657_1050.t7 371.139
R1333 a_4657_1050.n1 a_4657_1050.t5 282.852
R1334 a_4657_1050.n6 a_4657_1050.n5 277.722
R1335 a_4657_1050.n1 a_4657_1050.n0 247.347
R1336 a_4657_1050.n8 a_4657_1050.n6 187.858
R1337 a_4657_1050.n8 a_4657_1050.n7 157.964
R1338 a_4657_1050.n9 a_4657_1050.n8 91.705
R1339 a_4657_1050.n5 a_4657_1050.n4 30
R1340 a_4657_1050.n3 a_4657_1050.n2 24.383
R1341 a_4657_1050.n5 a_4657_1050.n3 23.684
R1342 a_4657_1050.n7 a_4657_1050.t3 14.282
R1343 a_4657_1050.n7 a_4657_1050.t4 14.282
R1344 a_4657_1050.t1 a_4657_1050.n9 14.282
R1345 a_4657_1050.n9 a_4657_1050.t0 14.282
R1346 a_4657_1050.n6 a_4657_1050.n1 10.343
R1347 a_5291_209.n0 a_5291_209.t5 486.819
R1348 a_5291_209.n0 a_5291_209.t4 384.527
R1349 a_5291_209.n4 a_5291_209.n3 299.14
R1350 a_5291_209.n1 a_5291_209.t3 295.06
R1351 a_5291_209.n3 a_5291_209.n2 266.331
R1352 a_5291_209.n1 a_5291_209.n0 234.846
R1353 a_5291_209.n3 a_5291_209.n1 14.696
R1354 a_5291_209.t1 a_5291_209.n4 14.282
R1355 a_5291_209.n4 a_5291_209.t0 14.282
R1356 B.n2 B.t0 512.525
R1357 B.n6 B.t3 480.392
R1358 B.n0 B.t2 480.392
R1359 B.n1 B.t1 440.954
R1360 B.n6 B.t7 403.272
R1361 B.n0 B.t6 403.272
R1362 B.n2 B.t8 371.139
R1363 B.n4 B.t5 299.455
R1364 B.n4 B.t4 227.134
R1365 B.n5 B.n4 139.294
R1366 B.n7 B.n6 120.597
R1367 B.n3 B.n2 69.036
R1368 B.n5 B.n3 28.032
R1369 B.n1 B.n0 20.835
R1370 B.n3 B.n1 17.715
R1371 B.n7 B.n5 7.325
R1372 B.n7 B 0.046
R1373 a_807_990.n0 a_807_990.t4 477.179
R1374 a_807_990.n0 a_807_990.t3 406.485
R1375 a_807_990.n4 a_807_990.t5 312.917
R1376 a_807_990.n4 a_807_990.n3 260.115
R1377 a_807_990.n6 a_807_990.n5 215.563
R1378 a_807_990.n5 a_807_990.n0 156.869
R1379 a_807_990.n5 a_807_990.n4 83.576
R1380 a_807_990.n3 a_807_990.n2 22.578
R1381 a_807_990.n6 a_807_990.t0 14.282
R1382 a_807_990.t1 a_807_990.n6 14.282
R1383 a_807_990.n3 a_807_990.n1 8.58
R1384 a_5662_101.n11 a_5662_101.n10 68.43
R1385 a_5662_101.n3 a_5662_101.n2 62.817
R1386 a_5662_101.n7 a_5662_101.n6 38.626
R1387 a_5662_101.n6 a_5662_101.n5 35.955
R1388 a_5662_101.n3 a_5662_101.n1 26.202
R1389 a_5662_101.t0 a_5662_101.n3 19.737
R1390 a_5662_101.t1 a_5662_101.n8 8.137
R1391 a_5662_101.t0 a_5662_101.n4 7.273
R1392 a_5662_101.t0 a_5662_101.n0 6.109
R1393 a_5662_101.t1 a_5662_101.n7 4.864
R1394 a_5662_101.t0 a_5662_101.n12 2.074
R1395 a_5662_101.n12 a_5662_101.t1 0.937
R1396 a_5662_101.t1 a_5662_101.n11 0.763
R1397 a_5662_101.n11 a_5662_101.n9 0.185
R1398 A.n5 A.t5 512.525
R1399 A.n0 A.t8 480.392
R1400 A.n1 A.t6 472.359
R1401 A.n0 A.t4 403.272
R1402 A.n1 A.t7 384.527
R1403 A.n5 A.t0 371.139
R1404 A.n6 A.t2 366.428
R1405 A.n2 A.n1 291.145
R1406 A.n3 A.t1 178.533
R1407 A.n4 A.n3 164.048
R1408 A.n6 A.n5 163.771
R1409 A.n2 A.t3 136.225
R1410 A.n4 A.n0 115.947
R1411 A.n3 A.n2 28.99
R1412 A.n7 A.n4 6.509
R1413 A.n7 A.n6 4.65
R1414 A.n7 A 0.046
R1415 a_185_209.n0 a_185_209.t5 477.179
R1416 a_185_209.n0 a_185_209.t4 406.485
R1417 a_185_209.n1 a_185_209.t3 341.566
R1418 a_185_209.n3 a_185_209.n2 294.19
R1419 a_185_209.n4 a_185_209.n3 271.281
R1420 a_185_209.n1 a_185_209.n0 199.524
R1421 a_185_209.n4 a_185_209.t0 14.282
R1422 a_185_209.t1 a_185_209.n4 14.282
R1423 a_185_209.n3 a_185_209.n1 13.879
R1424 a_3027_990.n0 a_3027_990.t3 477.179
R1425 a_3027_990.n0 a_3027_990.t5 406.485
R1426 a_3027_990.n4 a_3027_990.t4 312.917
R1427 a_3027_990.n4 a_3027_990.n3 260.115
R1428 a_3027_990.n6 a_3027_990.n5 215.563
R1429 a_3027_990.n5 a_3027_990.n0 156.869
R1430 a_3027_990.n5 a_3027_990.n4 83.576
R1431 a_3027_990.n3 a_3027_990.n2 22.578
R1432 a_3027_990.n6 a_3027_990.t0 14.282
R1433 a_3027_990.t1 a_3027_990.n6 14.282
R1434 a_3027_990.n3 a_3027_990.n1 8.58
R1435 a_556_101.n11 a_556_101.n10 68.43
R1436 a_556_101.n3 a_556_101.n2 62.817
R1437 a_556_101.n7 a_556_101.n6 38.626
R1438 a_556_101.n6 a_556_101.n5 35.955
R1439 a_556_101.n3 a_556_101.n1 26.202
R1440 a_556_101.t0 a_556_101.n3 19.737
R1441 a_556_101.t1 a_556_101.n8 8.137
R1442 a_556_101.t0 a_556_101.n4 7.273
R1443 a_556_101.t0 a_556_101.n0 6.109
R1444 a_556_101.t1 a_556_101.n7 4.864
R1445 a_556_101.t0 a_556_101.n12 2.074
R1446 a_556_101.n12 a_556_101.t1 0.937
R1447 a_556_101.t1 a_556_101.n11 0.763
R1448 a_556_101.n11 a_556_101.n9 0.185
R1449 a_4552_101.n3 a_4552_101.n1 42.788
R1450 a_4552_101.t0 a_4552_101.n0 8.137
R1451 a_4552_101.n3 a_4552_101.n2 4.665
R1452 a_4552_101.t0 a_4552_101.n3 0.06
R1453 a_2795_1051.n0 a_2795_1051.t2 228.369
R1454 a_2795_1051.n0 a_2795_1051.t0 219.778
R1455 a_2795_1051.n1 a_2795_1051.n0 42.29
R1456 a_2795_1051.n1 a_2795_1051.t3 14.282
R1457 a_2795_1051.t1 a_2795_1051.n1 14.282
R1458 a_6858_209.n1 a_6858_209.t6 512.525
R1459 a_6858_209.n1 a_6858_209.t4 371.139
R1460 a_6858_209.n3 a_6858_209.n0 287.966
R1461 a_6858_209.n2 a_6858_209.t5 282.852
R1462 a_6858_209.n2 a_6858_209.n1 247.347
R1463 a_6858_209.n7 a_6858_209.n6 223.975
R1464 a_6858_209.n7 a_6858_209.n3 142.305
R1465 a_6858_209.n9 a_6858_209.n7 142.275
R1466 a_6858_209.n6 a_6858_209.n5 22.578
R1467 a_6858_209.n9 a_6858_209.n8 15.001
R1468 a_6858_209.n0 a_6858_209.t2 14.282
R1469 a_6858_209.n0 a_6858_209.t1 14.282
R1470 a_6858_209.n10 a_6858_209.n9 12.632
R1471 a_6858_209.n3 a_6858_209.n2 10.343
R1472 a_6858_209.n6 a_6858_209.n4 8.58
R1473 COUT.n2 COUT.n1 294.19
R1474 COUT.n2 COUT.n0 271.281
R1475 COUT.n0 COUT.t0 14.282
R1476 COUT.n0 COUT.t1 14.282
R1477 COUT.n3 COUT.n2 4.65
R1478 COUT.n3 COUT 0.046
R1479 a_3461_1051.n1 a_3461_1051.t3 228.368
R1480 a_3461_1051.t1 a_3461_1051.n1 219.777
R1481 a_3461_1051.n1 a_3461_1051.n0 42.29
R1482 a_3461_1051.n0 a_3461_1051.t2 14.282
R1483 a_3461_1051.n0 a_3461_1051.t0 14.282
R1484 a_5767_1050.n0 a_5767_1050.t6 512.525
R1485 a_5767_1050.n0 a_5767_1050.t7 371.139
R1486 a_5767_1050.n3 a_5767_1050.n2 299.461
R1487 a_5767_1050.n1 a_5767_1050.t5 282.852
R1488 a_5767_1050.n1 a_5767_1050.n0 247.347
R1489 a_5767_1050.n5 a_5767_1050.n3 187.858
R1490 a_5767_1050.n5 a_5767_1050.n4 157.964
R1491 a_5767_1050.n6 a_5767_1050.n5 91.705
R1492 a_5767_1050.n4 a_5767_1050.t4 14.282
R1493 a_5767_1050.n4 a_5767_1050.t3 14.282
R1494 a_5767_1050.t1 a_5767_1050.n6 14.282
R1495 a_5767_1050.n6 a_5767_1050.t0 14.282
R1496 a_5767_1050.n3 a_5767_1050.n1 10.343
R1497 a_6401_209.n0 a_6401_209.t4 470.752
R1498 a_6401_209.n0 a_6401_209.t5 384.527
R1499 a_6401_209.n3 a_6401_209.n2 294.19
R1500 a_6401_209.n1 a_6401_209.t3 287.037
R1501 a_6401_209.n4 a_6401_209.n3 271.281
R1502 a_6401_209.n1 a_6401_209.n0 210.791
R1503 a_6401_209.t1 a_6401_209.n4 14.282
R1504 a_6401_209.n4 a_6401_209.t0 14.282
R1505 a_6401_209.n3 a_6401_209.n1 11.159
R1506 a_575_1051.n1 a_575_1051.t3 228.368
R1507 a_575_1051.t1 a_575_1051.n1 219.777
R1508 a_575_1051.n1 a_575_1051.n0 42.29
R1509 a_575_1051.n0 a_575_1051.t2 14.282
R1510 a_575_1051.n0 a_575_1051.t0 14.282
R1511 a_1222_101.n3 a_1222_101.n1 42.788
R1512 a_1222_101.t0 a_1222_101.n0 8.137
R1513 a_1222_101.n3 a_1222_101.n2 4.665
R1514 a_1222_101.t0 a_1222_101.n3 0.06
R1515 a_1241_1051.t1 a_1241_1051.n1 228.371
R1516 a_1241_1051.n1 a_1241_1051.t2 219.777
R1517 a_1241_1051.n1 a_1241_1051.n0 42.29
R1518 a_1241_1051.n0 a_1241_1051.t0 14.282
R1519 a_1241_1051.n0 a_1241_1051.t3 14.282
R1520 a_6791_1051.t1 a_6791_1051.n1 228.371
R1521 a_6791_1051.n1 a_6791_1051.t3 219.777
R1522 a_6791_1051.n1 a_6791_1051.n0 42.29
R1523 a_6791_1051.n0 a_6791_1051.t0 14.282
R1524 a_6791_1051.n0 a_6791_1051.t2 14.282
R1525 a_3442_101.n11 a_3442_101.n10 68.43
R1526 a_3442_101.n3 a_3442_101.n2 62.817
R1527 a_3442_101.n7 a_3442_101.n6 38.626
R1528 a_3442_101.n6 a_3442_101.n5 35.955
R1529 a_3442_101.n3 a_3442_101.n1 26.202
R1530 a_3442_101.t0 a_3442_101.n3 19.737
R1531 a_3442_101.t1 a_3442_101.n8 8.137
R1532 a_3442_101.t0 a_3442_101.n4 7.273
R1533 a_3442_101.t0 a_3442_101.n0 6.109
R1534 a_3442_101.t1 a_3442_101.n7 4.864
R1535 a_3442_101.t0 a_3442_101.n12 2.074
R1536 a_3442_101.n12 a_3442_101.t1 0.937
R1537 a_3442_101.t1 a_3442_101.n11 0.763
R1538 a_3442_101.n11 a_3442_101.n9 0.185
C11 VDD GND 13.24fF
C12 a_3442_101.n0 GND 0.03fF
C13 a_3442_101.n1 GND 0.11fF
C14 a_3442_101.n2 GND 0.09fF
C15 a_3442_101.n3 GND 0.04fF
C16 a_3442_101.n4 GND 0.02fF
C17 a_3442_101.n5 GND 0.04fF
C18 a_3442_101.n6 GND 0.05fF
C19 a_3442_101.n7 GND 0.02fF
C20 a_3442_101.n8 GND 0.06fF
C21 a_3442_101.n9 GND 0.18fF
C22 a_3442_101.n10 GND 0.10fF
C23 a_3442_101.n11 GND 0.10fF
C24 a_3442_101.n12 GND 0.01fF
C25 a_6791_1051.n0 GND 0.22fF
C26 a_6791_1051.n1 GND 0.52fF
C27 a_1241_1051.n0 GND 0.22fF
C28 a_1241_1051.n1 GND 0.50fF
C29 a_1222_101.n0 GND 0.06fF
C30 a_1222_101.n1 GND 0.14fF
C31 a_1222_101.n2 GND 0.05fF
C32 a_1222_101.n3 GND 0.20fF
C33 a_575_1051.n0 GND 0.22fF
C34 a_575_1051.n1 GND 0.50fF
C35 a_6401_209.n0 GND 0.33fF
C36 a_6401_209.t3 GND 0.50fF
C37 a_6401_209.n1 GND 0.63fF
C38 a_6401_209.n2 GND 0.29fF
C39 a_6401_209.n3 GND 0.86fF
C40 a_6401_209.n4 GND 0.63fF
C41 a_5767_1050.n0 GND 0.30fF
C42 a_5767_1050.t5 GND 0.44fF
C43 a_5767_1050.n1 GND 0.50fF
C44 a_5767_1050.n2 GND 0.26fF
C45 a_5767_1050.n3 GND 0.56fF
C46 a_5767_1050.n4 GND 0.42fF
C47 a_5767_1050.n5 GND 0.52fF
C48 a_5767_1050.n6 GND 0.33fF
C49 a_3461_1051.n0 GND 0.22fF
C50 a_3461_1051.n1 GND 0.50fF
C51 a_6858_209.n0 GND 0.46fF
C52 a_6858_209.n1 GND 0.28fF
C53 a_6858_209.n2 GND 0.46fF
C54 a_6858_209.n3 GND 0.50fF
C55 a_6858_209.n4 GND 0.03fF
C56 a_6858_209.n5 GND 0.04fF
C57 a_6858_209.n6 GND 0.11fF
C58 a_6858_209.n7 GND 0.37fF
C59 a_6858_209.n8 GND 0.06fF
C60 a_6858_209.n9 GND 0.04fF
C61 a_6858_209.n10 GND 0.04fF
C62 a_2795_1051.n0 GND 0.50fF
C63 a_2795_1051.n1 GND 0.22fF
C64 a_4552_101.n0 GND 0.06fF
C65 a_4552_101.n1 GND 0.14fF
C66 a_4552_101.n2 GND 0.05fF
C67 a_4552_101.n3 GND 0.20fF
C68 a_556_101.n0 GND 0.03fF
C69 a_556_101.n1 GND 0.11fF
C70 a_556_101.n2 GND 0.09fF
C71 a_556_101.n3 GND 0.04fF
C72 a_556_101.n4 GND 0.02fF
C73 a_556_101.n5 GND 0.04fF
C74 a_556_101.n6 GND 0.05fF
C75 a_556_101.n7 GND 0.02fF
C76 a_556_101.n8 GND 0.06fF
C77 a_556_101.n9 GND 0.18fF
C78 a_556_101.n10 GND 0.10fF
C79 a_556_101.n11 GND 0.10fF
C80 a_556_101.t1 GND 0.27fF
C81 a_556_101.n12 GND 0.01fF
C82 a_3027_990.n0 GND 0.64fF
C83 a_3027_990.n1 GND 0.08fF
C84 a_3027_990.n2 GND 0.10fF
C85 a_3027_990.n3 GND 0.32fF
C86 a_3027_990.n4 GND 1.97fF
C87 a_3027_990.n5 GND 2.47fF
C88 a_3027_990.n6 GND 1.03fF
C89 a_185_209.n0 GND 0.47fF
C90 a_185_209.t3 GND 0.69fF
C91 a_185_209.n1 GND 1.28fF
C92 a_185_209.n2 GND 0.39fF
C93 a_185_209.n3 GND 1.55fF
C94 a_185_209.n4 GND 0.84fF
C95 a_5662_101.n0 GND 0.03fF
C96 a_5662_101.n1 GND 0.11fF
C97 a_5662_101.n2 GND 0.09fF
C98 a_5662_101.n3 GND 0.04fF
C99 a_5662_101.n4 GND 0.02fF
C100 a_5662_101.n5 GND 0.04fF
C101 a_5662_101.n6 GND 0.05fF
C102 a_5662_101.n7 GND 0.02fF
C103 a_5662_101.n8 GND 0.06fF
C104 a_5662_101.n9 GND 0.18fF
C105 a_5662_101.n10 GND 0.10fF
C106 a_5662_101.n11 GND 0.10fF
C107 a_5662_101.t1 GND 0.27fF
C108 a_5662_101.n12 GND 0.01fF
C109 a_807_990.n0 GND 0.59fF
C110 a_807_990.n1 GND 0.07fF
C111 a_807_990.n2 GND 0.09fF
C112 a_807_990.n3 GND 0.30fF
C113 a_807_990.n4 GND 1.82fF
C114 a_807_990.n5 GND 2.29fF
C115 a_807_990.n6 GND 0.95fF
C116 a_5291_209.n0 GND 0.40fF
C117 a_5291_209.t3 GND 0.52fF
C118 a_5291_209.n1 GND 1.09fF
C119 a_5291_209.n2 GND 0.28fF
C120 a_5291_209.n3 GND 1.32fF
C121 a_5291_209.n4 GND 0.71fF
C122 a_4657_1050.n0 GND 0.29fF
C123 a_4657_1050.t5 GND 0.42fF
C124 a_4657_1050.n1 GND 0.48fF
C125 a_4657_1050.n2 GND 0.03fF
C126 a_4657_1050.n3 GND 0.04fF
C127 a_4657_1050.n4 GND 0.03fF
C128 a_4657_1050.n5 GND 0.16fF
C129 a_4657_1050.n6 GND 0.52fF
C130 a_4657_1050.n7 GND 0.40fF
C131 a_4657_1050.n8 GND 0.49fF
C132 a_4657_1050.n9 GND 0.31fF
C133 SUM.n0 GND 0.97fF
C134 SUM.n1 GND 0.07fF
C135 SUM.n2 GND 0.09fF
C136 SUM.n3 GND 0.06fF
C137 SUM.n4 GND 0.39fF
C138 SUM.n5 GND 1.11fF
C139 SUM.n6 GND 0.97fF
C140 SUM.n7 GND 0.59fF
C141 SUM.n8 GND 1.32fF
C142 SUM.n9 GND 0.05fF
C143 a_2776_101.n0 GND 0.10fF
C144 a_2776_101.n1 GND 0.03fF
C145 a_2776_101.n2 GND 0.02fF
C146 a_2776_101.n3 GND 0.11fF
C147 a_2776_101.n4 GND 0.09fF
C148 a_2776_101.n5 GND 0.05fF
C149 a_2776_101.n6 GND 0.03fF
C150 a_2776_101.n7 GND 0.06fF
C151 VDD.n1 GND 0.03fF
C152 VDD.n2 GND 0.09fF
C153 VDD.n3 GND 0.03fF
C154 VDD.n4 GND 0.02fF
C155 VDD.n5 GND 0.06fF
C156 VDD.n6 GND 0.02fF
C157 VDD.n7 GND 0.02fF
C158 VDD.n8 GND 0.02fF
C159 VDD.n9 GND 0.02fF
C160 VDD.n10 GND 0.02fF
C161 VDD.n11 GND 0.02fF
C162 VDD.n12 GND 0.02fF
C163 VDD.n13 GND 0.02fF
C164 VDD.n14 GND 0.03fF
C165 VDD.n15 GND 0.01fF
C166 VDD.n20 GND 0.43fF
C167 VDD.n21 GND 0.26fF
C168 VDD.n22 GND 0.02fF
C169 VDD.n23 GND 0.03fF
C170 VDD.n24 GND 0.06fF
C171 VDD.n25 GND 0.19fF
C172 VDD.n26 GND 0.01fF
C173 VDD.n27 GND 0.01fF
C174 VDD.n28 GND 0.06fF
C175 VDD.n29 GND 0.16fF
C176 VDD.n30 GND 0.01fF
C177 VDD.n31 GND 0.02fF
C178 VDD.n32 GND 0.02fF
C179 VDD.n33 GND 0.19fF
C180 VDD.n34 GND 0.01fF
C181 VDD.n35 GND 0.06fF
C182 VDD.n36 GND 0.01fF
C183 VDD.n37 GND 0.02fF
C184 VDD.n38 GND 0.26fF
C185 VDD.n39 GND 0.01fF
C186 VDD.n40 GND 0.02fF
C187 VDD.n41 GND 0.03fF
C188 VDD.n42 GND 0.05fF
C189 VDD.n43 GND 0.02fF
C190 VDD.n44 GND 0.02fF
C191 VDD.n45 GND 0.02fF
C192 VDD.n46 GND 0.02fF
C193 VDD.n47 GND 0.02fF
C194 VDD.n48 GND 0.02fF
C195 VDD.n49 GND 0.02fF
C196 VDD.n50 GND 0.02fF
C197 VDD.n51 GND 0.02fF
C198 VDD.n52 GND 0.02fF
C199 VDD.n53 GND 0.02fF
C200 VDD.n54 GND 0.03fF
C201 VDD.n55 GND 0.02fF
C202 VDD.n56 GND 0.17fF
C203 VDD.n57 GND 0.02fF
C204 VDD.n58 GND 0.02fF
C205 VDD.n60 GND 0.02fF
C206 VDD.n64 GND 0.26fF
C207 VDD.n65 GND 0.26fF
C208 VDD.n66 GND 0.01fF
C209 VDD.n67 GND 0.02fF
C210 VDD.n68 GND 0.03fF
C211 VDD.n69 GND 0.23fF
C212 VDD.n70 GND 0.01fF
C213 VDD.n71 GND 0.02fF
C214 VDD.n72 GND 0.02fF
C215 VDD.n73 GND 0.16fF
C216 VDD.n74 GND 0.01fF
C217 VDD.n75 GND 0.02fF
C218 VDD.n76 GND 0.02fF
C219 VDD.n77 GND 0.01fF
C220 VDD.n78 GND 0.02fF
C221 VDD.n79 GND 0.02fF
C222 VDD.n80 GND 0.13fF
C223 VDD.n81 GND 0.01fF
C224 VDD.n82 GND 0.02fF
C225 VDD.n83 GND 0.02fF
C226 VDD.n84 GND 0.08fF
C227 VDD.n85 GND 0.05fF
C228 VDD.n86 GND 0.16fF
C229 VDD.n87 GND 0.01fF
C230 VDD.n88 GND 0.02fF
C231 VDD.n89 GND 0.02fF
C232 VDD.n90 GND 0.24fF
C233 VDD.n91 GND 0.01fF
C234 VDD.n92 GND 0.02fF
C235 VDD.n93 GND 0.02fF
C236 VDD.n94 GND 0.26fF
C237 VDD.n95 GND 0.01fF
C238 VDD.n96 GND 0.02fF
C239 VDD.n97 GND 0.03fF
C240 VDD.n98 GND 0.17fF
C241 VDD.n99 GND 0.02fF
C242 VDD.n100 GND 0.02fF
C243 VDD.n101 GND 0.02fF
C244 VDD.n102 GND 0.06fF
C245 VDD.n103 GND 0.02fF
C246 VDD.n104 GND 0.02fF
C247 VDD.n105 GND 0.02fF
C248 VDD.n106 GND 0.02fF
C249 VDD.n107 GND 0.02fF
C250 VDD.n108 GND 0.02fF
C251 VDD.n109 GND 0.02fF
C252 VDD.n110 GND 0.02fF
C253 VDD.n111 GND 0.02fF
C254 VDD.n112 GND 0.02fF
C255 VDD.n113 GND 0.03fF
C256 VDD.n114 GND 0.02fF
C257 VDD.n115 GND 0.02fF
C258 VDD.n119 GND 0.26fF
C259 VDD.n120 GND 0.26fF
C260 VDD.n121 GND 0.01fF
C261 VDD.n122 GND 0.02fF
C262 VDD.n123 GND 0.03fF
C263 VDD.n124 GND 0.06fF
C264 VDD.n125 GND 0.19fF
C265 VDD.n126 GND 0.01fF
C266 VDD.n127 GND 0.01fF
C267 VDD.n128 GND 0.02fF
C268 VDD.n129 GND 0.16fF
C269 VDD.n130 GND 0.01fF
C270 VDD.n131 GND 0.02fF
C271 VDD.n132 GND 0.02fF
C272 VDD.n133 GND 0.06fF
C273 VDD.n134 GND 0.19fF
C274 VDD.n135 GND 0.01fF
C275 VDD.n136 GND 0.01fF
C276 VDD.n137 GND 0.02fF
C277 VDD.n138 GND 0.26fF
C278 VDD.n139 GND 0.01fF
C279 VDD.n140 GND 0.02fF
C280 VDD.n141 GND 0.03fF
C281 VDD.n142 GND 0.17fF
C282 VDD.n143 GND 0.02fF
C283 VDD.n144 GND 0.02fF
C284 VDD.n145 GND 0.02fF
C285 VDD.n146 GND 0.06fF
C286 VDD.n147 GND 0.02fF
C287 VDD.n148 GND 0.02fF
C288 VDD.n149 GND 0.02fF
C289 VDD.n150 GND 0.02fF
C290 VDD.n151 GND 0.02fF
C291 VDD.n152 GND 0.02fF
C292 VDD.n153 GND 0.02fF
C293 VDD.n154 GND 0.02fF
C294 VDD.n155 GND 0.02fF
C295 VDD.n156 GND 0.02fF
C296 VDD.n157 GND 0.03fF
C297 VDD.n158 GND 0.02fF
C298 VDD.n159 GND 0.02fF
C299 VDD.n163 GND 0.26fF
C300 VDD.n164 GND 0.26fF
C301 VDD.n165 GND 0.01fF
C302 VDD.n166 GND 0.02fF
C303 VDD.n167 GND 0.03fF
C304 VDD.n168 GND 0.23fF
C305 VDD.n169 GND 0.01fF
C306 VDD.n170 GND 0.06fF
C307 VDD.n171 GND 0.01fF
C308 VDD.n172 GND 0.02fF
C309 VDD.n173 GND 0.16fF
C310 VDD.n174 GND 0.01fF
C311 VDD.n175 GND 0.02fF
C312 VDD.n176 GND 0.02fF
C313 VDD.n177 GND 0.01fF
C314 VDD.n178 GND 0.08fF
C315 VDD.n179 GND 0.05fF
C316 VDD.n180 GND 0.02fF
C317 VDD.n181 GND 0.02fF
C318 VDD.n182 GND 0.13fF
C319 VDD.n183 GND 0.01fF
C320 VDD.n184 GND 0.02fF
C321 VDD.n185 GND 0.02fF
C322 VDD.n186 GND 0.16fF
C323 VDD.n187 GND 0.01fF
C324 VDD.n188 GND 0.02fF
C325 VDD.n189 GND 0.02fF
C326 VDD.n190 GND 0.06fF
C327 VDD.n191 GND 0.24fF
C328 VDD.n192 GND 0.01fF
C329 VDD.n193 GND 0.01fF
C330 VDD.n194 GND 0.02fF
C331 VDD.n195 GND 0.26fF
C332 VDD.n196 GND 0.01fF
C333 VDD.n197 GND 0.02fF
C334 VDD.n198 GND 0.03fF
C335 VDD.n199 GND 0.17fF
C336 VDD.n200 GND 0.02fF
C337 VDD.n201 GND 0.02fF
C338 VDD.n202 GND 0.02fF
C339 VDD.n203 GND 0.06fF
C340 VDD.n204 GND 0.02fF
C341 VDD.n205 GND 0.02fF
C342 VDD.n206 GND 0.02fF
C343 VDD.n207 GND 0.02fF
C344 VDD.n208 GND 0.02fF
C345 VDD.n209 GND 0.02fF
C346 VDD.n210 GND 0.02fF
C347 VDD.n211 GND 0.02fF
C348 VDD.n212 GND 0.02fF
C349 VDD.n213 GND 0.02fF
C350 VDD.n214 GND 0.03fF
C351 VDD.n215 GND 0.02fF
C352 VDD.n216 GND 0.02fF
C353 VDD.n220 GND 0.26fF
C354 VDD.n221 GND 0.26fF
C355 VDD.n222 GND 0.01fF
C356 VDD.n223 GND 0.02fF
C357 VDD.n224 GND 0.03fF
C358 VDD.n225 GND 0.06fF
C359 VDD.n226 GND 0.19fF
C360 VDD.n227 GND 0.01fF
C361 VDD.n228 GND 0.01fF
C362 VDD.n229 GND 0.02fF
C363 VDD.n230 GND 0.16fF
C364 VDD.n231 GND 0.01fF
C365 VDD.n232 GND 0.02fF
C366 VDD.n233 GND 0.02fF
C367 VDD.n234 GND 0.19fF
C368 VDD.n235 GND 0.01fF
C369 VDD.n236 GND 0.06fF
C370 VDD.n237 GND 0.01fF
C371 VDD.n238 GND 0.02fF
C372 VDD.n239 GND 0.26fF
C373 VDD.n240 GND 0.01fF
C374 VDD.n241 GND 0.02fF
C375 VDD.n242 GND 0.03fF
C376 VDD.n243 GND 0.17fF
C377 VDD.n244 GND 0.02fF
C378 VDD.n245 GND 0.02fF
C379 VDD.n246 GND 0.02fF
C380 VDD.n247 GND 0.06fF
C381 VDD.n248 GND 0.02fF
C382 VDD.n249 GND 0.02fF
C383 VDD.n250 GND 0.02fF
C384 VDD.n251 GND 0.02fF
C385 VDD.n252 GND 0.02fF
C386 VDD.n253 GND 0.02fF
C387 VDD.n254 GND 0.02fF
C388 VDD.n255 GND 0.02fF
C389 VDD.n256 GND 0.02fF
C390 VDD.n257 GND 0.02fF
C391 VDD.n258 GND 0.03fF
C392 VDD.n259 GND 0.02fF
C393 VDD.n260 GND 0.02fF
C394 VDD.n264 GND 0.26fF
C395 VDD.n265 GND 0.26fF
C396 VDD.n266 GND 0.01fF
C397 VDD.n267 GND 0.02fF
C398 VDD.n268 GND 0.03fF
C399 VDD.n269 GND 0.06fF
C400 VDD.n270 GND 0.23fF
C401 VDD.n271 GND 0.01fF
C402 VDD.n272 GND 0.01fF
C403 VDD.n273 GND 0.02fF
C404 VDD.n274 GND 0.16fF
C405 VDD.n275 GND 0.01fF
C406 VDD.n276 GND 0.02fF
C407 VDD.n277 GND 0.02fF
C408 VDD.n278 GND 0.08fF
C409 VDD.n279 GND 0.05fF
C410 VDD.n280 GND 0.01fF
C411 VDD.n281 GND 0.02fF
C412 VDD.n282 GND 0.02fF
C413 VDD.n283 GND 0.13fF
C414 VDD.n284 GND 0.01fF
C415 VDD.n285 GND 0.02fF
C416 VDD.n286 GND 0.02fF
C417 VDD.n287 GND 0.16fF
C418 VDD.n288 GND 0.01fF
C419 VDD.n289 GND 0.02fF
C420 VDD.n290 GND 0.02fF
C421 VDD.n291 GND 0.06fF
C422 VDD.n292 GND 0.24fF
C423 VDD.n293 GND 0.01fF
C424 VDD.n294 GND 0.01fF
C425 VDD.n295 GND 0.02fF
C426 VDD.n296 GND 0.26fF
C427 VDD.n297 GND 0.01fF
C428 VDD.n298 GND 0.02fF
C429 VDD.n299 GND 0.03fF
C430 VDD.n300 GND 0.17fF
C431 VDD.n301 GND 0.02fF
C432 VDD.n302 GND 0.02fF
C433 VDD.n303 GND 0.02fF
C434 VDD.n304 GND 0.06fF
C435 VDD.n305 GND 0.02fF
C436 VDD.n306 GND 0.02fF
C437 VDD.n307 GND 0.02fF
C438 VDD.n308 GND 0.02fF
C439 VDD.n309 GND 0.02fF
C440 VDD.n310 GND 0.02fF
C441 VDD.n311 GND 0.02fF
C442 VDD.n312 GND 0.02fF
C443 VDD.n313 GND 0.02fF
C444 VDD.n314 GND 0.02fF
C445 VDD.n315 GND 0.03fF
C446 VDD.n316 GND 0.02fF
C447 VDD.n317 GND 0.02fF
C448 VDD.n321 GND 0.26fF
C449 VDD.n322 GND 0.26fF
C450 VDD.n323 GND 0.01fF
C451 VDD.n324 GND 0.02fF
C452 VDD.n325 GND 0.03fF
C453 VDD.n326 GND 0.06fF
C454 VDD.n327 GND 0.19fF
C455 VDD.n328 GND 0.01fF
C456 VDD.n329 GND 0.01fF
C457 VDD.n330 GND 0.02fF
C458 VDD.n331 GND 0.16fF
C459 VDD.n332 GND 0.01fF
C460 VDD.n333 GND 0.02fF
C461 VDD.n334 GND 0.02fF
C462 VDD.n335 GND 0.06fF
C463 VDD.n336 GND 0.19fF
C464 VDD.n337 GND 0.01fF
C465 VDD.n338 GND 0.01fF
C466 VDD.n339 GND 0.02fF
C467 VDD.n340 GND 0.26fF
C468 VDD.n341 GND 0.01fF
C469 VDD.n342 GND 0.02fF
C470 VDD.n343 GND 0.03fF
C471 VDD.n344 GND 0.17fF
C472 VDD.n345 GND 0.02fF
C473 VDD.n346 GND 0.02fF
C474 VDD.n347 GND 0.02fF
C475 VDD.n348 GND 0.06fF
C476 VDD.n349 GND 0.02fF
C477 VDD.n350 GND 0.02fF
C478 VDD.n351 GND 0.02fF
C479 VDD.n352 GND 0.02fF
C480 VDD.n353 GND 0.02fF
C481 VDD.n354 GND 0.02fF
C482 VDD.n355 GND 0.02fF
C483 VDD.n356 GND 0.02fF
C484 VDD.n357 GND 0.02fF
C485 VDD.n358 GND 0.02fF
C486 VDD.n359 GND 0.03fF
C487 VDD.n360 GND 0.02fF
C488 VDD.n361 GND 0.02fF
C489 VDD.n365 GND 0.26fF
C490 VDD.n366 GND 0.26fF
C491 VDD.n367 GND 0.01fF
C492 VDD.n368 GND 0.02fF
C493 VDD.n369 GND 0.03fF
C494 VDD.n370 GND 0.09fF
C495 VDD.n371 GND 0.02fF
C496 VDD.n372 GND 0.02fF
C497 VDD.n373 GND 0.06fF
C498 VDD.n374 GND 0.02fF
C499 VDD.n375 GND 0.02fF
C500 VDD.n376 GND 0.02fF
C501 VDD.n377 GND 0.02fF
C502 VDD.n378 GND 0.02fF
C503 VDD.n379 GND 0.02fF
C504 VDD.n380 GND 0.02fF
C505 VDD.n381 GND 0.02fF
C506 VDD.n382 GND 0.03fF
C507 VDD.n383 GND 0.03fF
C508 VDD.n384 GND 0.02fF
C509 VDD.n388 GND 0.43fF
C510 VDD.n389 GND 0.26fF
C511 VDD.n390 GND 0.02fF
C512 VDD.n391 GND 0.03fF
C513 VDD.n392 GND 0.03fF
C514 VDD.n393 GND 0.19fF
C515 VDD.n394 GND 0.01fF
C516 VDD.n395 GND 0.06fF
C517 VDD.n396 GND 0.01fF
C518 VDD.n397 GND 0.02fF
C519 VDD.n398 GND 0.16fF
C520 VDD.n399 GND 0.01fF
C521 VDD.n400 GND 0.02fF
C522 VDD.n401 GND 0.02fF
C523 VDD.n402 GND 0.06fF
C524 VDD.n403 GND 0.19fF
C525 VDD.n404 GND 0.01fF
C526 VDD.n405 GND 0.01fF
C527 VDD.n406 GND 0.02fF
C528 VDD.n407 GND 0.26fF
C529 VDD.n408 GND 0.01fF
C530 VDD.n409 GND 0.02fF
C531 VDD.n410 GND 0.03fF
C532 VDD.n411 GND 0.02fF
C533 VDD.n414 GND 0.02fF
C534 VDD.n416 GND 0.02fF
C535 VDD.n417 GND 0.17fF
C536 VDD.n418 GND 0.02fF
C537 VDD.n420 GND 0.26fF
C538 VDD.n421 GND 0.26fF
C539 VDD.n422 GND 0.01fF
C540 VDD.n423 GND 0.05fF
C541 VDD.n424 GND 0.02fF
C542 VDD.n425 GND 0.02fF
C543 VDD.n426 GND 0.02fF
C544 VDD.n427 GND 0.02fF
C545 VDD.n428 GND 0.02fF
C546 VDD.n429 GND 0.02fF
C547 VDD.n430 GND 0.02fF
C548 VDD.n431 GND 0.02fF
C549 VDD.n432 GND 0.02fF
C550 VDD.n433 GND 0.02fF
C551 VDD.n434 GND 0.02fF
C552 VDD.n435 GND 0.03fF
C553 VDD.n436 GND 0.02fF
C554 VDD.n437 GND 0.03fF
C555 VDD.n438 GND 0.24fF
C556 VDD.n439 GND 0.01fF
C557 VDD.n440 GND 0.02fF
C558 VDD.n441 GND 0.02fF
C559 VDD.n442 GND 0.07fF
C560 VDD.n443 GND 0.05fF
C561 VDD.n444 GND 0.16fF
C562 VDD.n445 GND 0.01fF
C563 VDD.n446 GND 0.02fF
C564 VDD.n447 GND 0.02fF
C565 VDD.n448 GND 0.13fF
C566 VDD.n449 GND 0.01fF
C567 VDD.n450 GND 0.02fF
C568 VDD.n451 GND 0.02fF
C569 VDD.n452 GND 0.01fF
C570 VDD.n453 GND 0.02fF
C571 VDD.n454 GND 0.02fF
C572 VDD.n455 GND 0.16fF
C573 VDD.n456 GND 0.01fF
C574 VDD.n457 GND 0.02fF
C575 VDD.n458 GND 0.02fF
C576 VDD.n459 GND 0.23fF
C577 VDD.n460 GND 0.01fF
C578 VDD.n461 GND 0.02fF
C579 VDD.n462 GND 0.02fF
C580 VDD.n463 GND 0.26fF
C581 VDD.n464 GND 0.01fF
C582 VDD.n465 GND 0.02fF
C583 VDD.n466 GND 0.03fF
C584 VDD.n467 GND 0.02fF
C585 VDD.n468 GND 0.02fF
C586 VDD.n472 GND 0.26fF
C587 VDD.n473 GND 0.26fF
C588 VDD.n474 GND 0.01fF
C589 VDD.n475 GND 0.20fF
C590 VDD.n476 GND 0.02fF
C591 VDD.n477 GND 0.02fF
C592 VDD.n478 GND 0.02fF
C593 VDD.n479 GND 0.06fF
C594 VDD.n480 GND 0.02fF
C595 VDD.n481 GND 0.02fF
C596 VDD.n482 GND 0.02fF
C597 VDD.n483 GND 0.02fF
C598 VDD.n484 GND 0.02fF
C599 VDD.n485 GND 0.02fF
C600 VDD.n486 GND 0.02fF
C601 VDD.n487 GND 0.02fF
C602 VDD.n488 GND 0.02fF
C603 VDD.n489 GND 0.02fF
C604 VDD.n490 GND 0.03fF
C605 VDD.n491 GND 0.02fF
C606 VDD.n492 GND 0.03fF
C607 VDD.n493 GND 0.24fF
C608 VDD.n494 GND 0.01fF
C609 VDD.n495 GND 0.02fF
C610 VDD.n496 GND 0.02fF
C611 VDD.n497 GND 0.07fF
C612 VDD.n498 GND 0.05fF
C613 VDD.n499 GND 0.16fF
C614 VDD.n500 GND 0.01fF
C615 VDD.n501 GND 0.02fF
C616 VDD.n502 GND 0.02fF
C617 VDD.n503 GND 0.13fF
C618 VDD.n504 GND 0.01fF
C619 VDD.n505 GND 0.02fF
C620 VDD.n506 GND 0.02fF
C621 VDD.n507 GND 0.01fF
C622 VDD.n508 GND 0.02fF
C623 VDD.n509 GND 0.02fF
C624 VDD.n510 GND 0.16fF
C625 VDD.n511 GND 0.01fF
C626 VDD.n512 GND 0.02fF
C627 VDD.n513 GND 0.02fF
C628 VDD.n514 GND 0.23fF
C629 VDD.n515 GND 0.01fF
C630 VDD.n516 GND 0.02fF
C631 VDD.n517 GND 0.02fF
C632 VDD.n518 GND 0.26fF
C633 VDD.n519 GND 0.01fF
C634 VDD.n520 GND 0.02fF
C635 VDD.n521 GND 0.03fF
C636 VDD.n522 GND 0.02fF
C637 VDD.n523 GND 0.02fF
C638 VDD.n527 GND 0.26fF
C639 VDD.n528 GND 0.26fF
C640 VDD.n529 GND 0.01fF
C641 VDD.n530 GND 0.17fF
C642 VDD.n531 GND 0.02fF
C643 VDD.n532 GND 0.02fF
C644 VDD.n533 GND 0.02fF
C645 VDD.n534 GND 0.06fF
C646 VDD.n535 GND 0.02fF
C647 VDD.n536 GND 0.02fF
C648 VDD.n537 GND 0.02fF
C649 VDD.n538 GND 0.02fF
C650 VDD.n539 GND 0.02fF
C651 VDD.n540 GND 0.02fF
C652 VDD.n541 GND 0.02fF
C653 VDD.n542 GND 0.02fF
C654 VDD.n543 GND 0.02fF
C655 VDD.n544 GND 0.02fF
C656 VDD.n545 GND 0.03fF
C657 VDD.n546 GND 0.02fF
C658 VDD.n547 GND 0.03fF
C659 VDD.n548 GND 0.06fF
C660 VDD.n549 GND 0.19fF
C661 VDD.n550 GND 0.01fF
C662 VDD.n551 GND 0.01fF
C663 VDD.n552 GND 0.02fF
C664 VDD.n553 GND 0.16fF
C665 VDD.n554 GND 0.01fF
C666 VDD.n555 GND 0.02fF
C667 VDD.n556 GND 0.02fF
C668 VDD.n557 GND 0.06fF
C669 VDD.n558 GND 0.19fF
C670 VDD.n559 GND 0.01fF
C671 VDD.n560 GND 0.01fF
C672 VDD.n561 GND 0.02fF
C673 VDD.n562 GND 0.26fF
C674 VDD.n563 GND 0.01fF
C675 VDD.n564 GND 0.02fF
C676 VDD.n565 GND 0.03fF
C677 VDD.n566 GND 0.14fF
C678 VDD.n567 GND 0.02fF
C679 VDD.n568 GND 0.02fF
C680 VDD.n569 GND 0.02fF
C681 VDD.n570 GND 0.06fF
C682 VDD.n571 GND 0.02fF
C683 VDD.n572 GND 0.02fF
C684 VDD.n573 GND 0.02fF
C685 VDD.n574 GND 0.02fF
C686 VDD.n575 GND 0.02fF
C687 VDD.n576 GND 0.02fF
C688 VDD.n577 GND 0.02fF
C689 VDD.n578 GND 0.02fF
C690 VDD.n579 GND 0.02fF
C691 VDD.n580 GND 0.02fF
C692 VDD.n581 GND 0.03fF
C693 VDD.n582 GND 0.02fF
C694 VDD.n583 GND 0.02fF
C695 VDD.n587 GND 0.26fF
C696 VDD.n588 GND 0.26fF
C697 VDD.n589 GND 0.01fF
C698 VDD.n590 GND 0.02fF
C699 VDD.n591 GND 0.03fF
C700 VDD.n592 GND 0.19fF
C701 VDD.n593 GND 0.01fF
C702 VDD.n594 GND 0.06fF
C703 VDD.n595 GND 0.01fF
C704 VDD.n596 GND 0.02fF
C705 VDD.n597 GND 0.16fF
C706 VDD.n598 GND 0.01fF
C707 VDD.n599 GND 0.02fF
C708 VDD.n600 GND 0.02fF
C709 VDD.n601 GND 0.06fF
C710 VDD.n602 GND 0.19fF
C711 VDD.n603 GND 0.01fF
C712 VDD.n604 GND 0.01fF
C713 VDD.n605 GND 0.02fF
C714 VDD.n606 GND 0.26fF
C715 VDD.n607 GND 0.01fF
C716 VDD.n608 GND 0.02fF
C717 VDD.n609 GND 0.03fF
C718 VDD.n610 GND 0.02fF
C719 VDD.n611 GND 0.02fF
C720 VDD.n615 GND 0.26fF
C721 VDD.n616 GND 0.26fF
C722 VDD.n617 GND 0.01fF
C723 VDD.n618 GND 0.17fF
C724 VDD.n619 GND 0.02fF
C725 VDD.n620 GND 0.02fF
C726 VDD.n621 GND 0.02fF
C727 VDD.n622 GND 0.06fF
C728 VDD.n623 GND 0.02fF
C729 VDD.n624 GND 0.02fF
C730 VDD.n625 GND 0.02fF
C731 VDD.n626 GND 0.02fF
C732 VDD.n627 GND 0.02fF
C733 VDD.n628 GND 0.02fF
C734 VDD.n629 GND 0.02fF
C735 VDD.n630 GND 0.02fF
C736 VDD.n631 GND 0.02fF
C737 VDD.n632 GND 0.02fF
C738 VDD.n633 GND 0.03fF
C739 VDD.n634 GND 0.02fF
C740 VDD.n635 GND 0.03fF
C741 VDD.n636 GND 0.24fF
C742 VDD.n637 GND 0.01fF
C743 VDD.n638 GND 0.02fF
C744 VDD.n639 GND 0.02fF
C745 VDD.n640 GND 0.07fF
C746 VDD.n641 GND 0.05fF
C747 VDD.n642 GND 0.16fF
C748 VDD.n643 GND 0.01fF
C749 VDD.n644 GND 0.02fF
C750 VDD.n645 GND 0.02fF
C751 VDD.n646 GND 0.13fF
C752 VDD.n647 GND 0.01fF
C753 VDD.n648 GND 0.02fF
C754 VDD.n649 GND 0.02fF
C755 VDD.n650 GND 0.01fF
C756 VDD.n651 GND 0.02fF
C757 VDD.n652 GND 0.02fF
C758 VDD.n653 GND 0.16fF
C759 VDD.n654 GND 0.01fF
C760 VDD.n655 GND 0.02fF
C761 VDD.n656 GND 0.02fF
C762 VDD.n657 GND 0.23fF
C763 VDD.n658 GND 0.01fF
C764 VDD.n659 GND 0.02fF
C765 VDD.n660 GND 0.02fF
C766 VDD.n661 GND 0.26fF
C767 VDD.n662 GND 0.01fF
C768 VDD.n663 GND 0.02fF
C769 VDD.n664 GND 0.03fF
C770 VDD.n665 GND 0.02fF
C771 VDD.n666 GND 0.02fF
C772 VDD.n670 GND 0.26fF
C773 VDD.n671 GND 0.26fF
C774 VDD.n672 GND 0.01fF
C775 VDD.n673 GND 0.20fF
C776 VDD.n674 GND 0.02fF
C777 VDD.n675 GND 0.02fF
C778 VDD.n676 GND 0.02fF
C779 VDD.n677 GND 0.06fF
C780 VDD.n678 GND 0.02fF
C781 VDD.n679 GND 0.02fF
C782 VDD.n680 GND 0.02fF
C783 VDD.n681 GND 0.02fF
C784 VDD.n682 GND 0.02fF
C785 VDD.n683 GND 0.02fF
C786 VDD.n684 GND 0.02fF
C787 VDD.n685 GND 0.02fF
C788 VDD.n686 GND 0.02fF
C789 VDD.n687 GND 0.02fF
C790 VDD.n688 GND 0.03fF
C791 VDD.n689 GND 0.02fF
C792 VDD.n690 GND 0.03fF
C793 VDD.n691 GND 0.24fF
C794 VDD.n692 GND 0.01fF
C795 VDD.n693 GND 0.02fF
C796 VDD.n694 GND 0.02fF
C797 VDD.n695 GND 0.07fF
C798 VDD.n696 GND 0.05fF
C799 VDD.n697 GND 0.16fF
C800 VDD.n698 GND 0.01fF
C801 VDD.n699 GND 0.02fF
C802 VDD.n700 GND 0.02fF
C803 VDD.n701 GND 0.13fF
C804 VDD.n702 GND 0.01fF
C805 VDD.n703 GND 0.02fF
C806 VDD.n704 GND 0.02fF
C807 VDD.n705 GND 0.01fF
C808 VDD.n706 GND 0.02fF
C809 VDD.n707 GND 0.02fF
C810 VDD.n708 GND 0.16fF
C811 VDD.n709 GND 0.01fF
C812 VDD.n710 GND 0.02fF
C813 VDD.n711 GND 0.02fF
C814 VDD.n712 GND 0.23fF
C815 VDD.n713 GND 0.01fF
C816 VDD.n714 GND 0.02fF
C817 VDD.n715 GND 0.02fF
C818 a_2405_209.n0 GND 0.06fF
C819 a_2405_209.n1 GND 0.97fF
C820 a_2405_209.n2 GND 0.54fF
C821 a_2405_209.n3 GND 1.47fF
C822 a_2405_209.n4 GND 1.75fF
C823 a_2405_209.n5 GND 0.05fF
C824 a_2405_209.n6 GND 0.28fF
C825 a_2405_209.n7 GND 0.08fF
C826 a_836_209.n0 GND 0.86fF
C827 a_836_209.n1 GND 0.44fF
C828 a_836_209.n2 GND 0.44fF
C829 a_836_209.n3 GND 1.05fF
C830 a_836_209.n4 GND 0.64fF
C831 a_836_209.n5 GND 0.65fF
C832 a_836_209.t7 GND 0.67fF
C833 a_836_209.n6 GND 2.22fF
C834 a_836_209.t13 GND 0.67fF
C835 a_836_209.n7 GND 1.97fF
C836 a_836_209.n8 GND 0.47fF
C837 a_836_209.n9 GND 0.86fF
C838 a_836_209.n10 GND 0.52fF
C839 a_836_209.n11 GND 1.01fF
C840 a_836_209.n12 GND 1.54fF
C841 a_836_209.n13 GND 1.15f