magic
tech sky130A
magscale 1 2
timestamp 1645051401
<< nwell >>
rect 52 -287 264 37
<< pmos >>
rect 144 -251 174 1
<< pdiff >>
rect 88 -39 144 1
rect 88 -73 98 -39
rect 132 -73 144 -39
rect 88 -107 144 -73
rect 88 -141 98 -107
rect 132 -141 144 -107
rect 88 -175 144 -141
rect 88 -209 98 -175
rect 132 -209 144 -175
rect 88 -251 144 -209
rect 174 -39 228 1
rect 174 -73 186 -39
rect 220 -73 228 -39
rect 174 -107 228 -73
rect 174 -141 186 -107
rect 220 -141 228 -107
rect 174 -251 228 -141
<< pdiffc >>
rect 98 -73 132 -39
rect 98 -141 132 -107
rect 98 -209 132 -175
rect 186 -73 220 -39
rect 186 -141 220 -107
<< poly >>
rect 144 1 174 27
rect 144 -277 174 -251
<< locali >>
rect 98 -39 132 42
rect 98 -107 132 -73
rect 98 -175 132 -141
rect 98 -227 132 -209
rect 186 -39 220 1
rect 186 -107 220 -73
rect 186 -227 220 -141
<< end >>
