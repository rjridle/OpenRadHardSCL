* SPICE3 file created from AO3X1.ext - technology: sky130A

.subckt AO3X1 A B C Y VDD GND
X0 VDD.t15 A.t0 a_217_1050.t4  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X1 VDD.t11 a_217_1050.t5 a_797_1051.t3 VDD.t10 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X2 VDD.t17 a_864_209.t4 Y.t1  U�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X3 VDD.t2 B.t0 a_217_1050.t1 �U�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X4 GND A.t1 a_112_101.t0 GND sky130_fd_pr__nfet_01v8 ad=3.2565p pd=2.261u as=0p ps=0u w=0u l=0u
X5 a_797_1051.t0 C.t0 a_864_209.t0  U�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X6 a_217_1050.t3 A.t2 VDD.t13 �U�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X7 Y.t0 a_864_209.t5 VDD.t7  U�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X8 a_797_1051.t2 a_217_1050.t7 VDD.t9 �U�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X9 a_217_1050.t2 B.t1 VDD.t5  U�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X10 Y a_864_209.t6 GND.t0 GND sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=0p ps=0u w=0u l=0u
X11 a_864_209.t2 C.t1 a_797_1051.t1 �U�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
C0 A VDD 0.32fF
C1 Y VDD 1.05fF
C2 C VDD 0.32fF
C3 B A 0.27fF
C4 B VDD 0.32fF
R0 A.n0 A.t0 480.392
R1 A.n0 A.t2 403.272
R2 A.n1 A.t1 301.486
R3 A.n1 A.n0 227.006
R4 A.n2 A.n1 4.65
R5 A.n2 A 0.046
R6 a_217_1050.n3 a_217_1050.t7 486.819
R7 a_217_1050.n3 a_217_1050.t5 384.527
R8 a_217_1050.n4 a_217_1050.t6 267.201
R9 a_217_1050.n4 a_217_1050.n3 262.705
R10 a_217_1050.n5 a_217_1050.n2 243.576
R11 a_217_1050.n7 a_217_1050.n5 228.526
R12 a_217_1050.n2 a_217_1050.n1 157.964
R13 a_217_1050.n2 a_217_1050.n0 91.706
R14 a_217_1050.n7 a_217_1050.n6 15.218
R15 a_217_1050.n0 a_217_1050.t1 14.282
R16 a_217_1050.n0 a_217_1050.t2 14.282
R17 a_217_1050.n1 a_217_1050.t4 14.282
R18 a_217_1050.n1 a_217_1050.t3 14.282
R19 a_217_1050.n8 a_217_1050.n7 12.014
R20 a_217_1050.n5 a_217_1050.n4 10.615
R21 VDD.n66 VDD.n55 144.705
R22 VDD.n162 VDD.n151 144.705
R23 VDD.n129 VDD.t2 143.754
R24 VDD.n107 VDD.t13 135.17
R25 VDD.n35 VDD.t7 135.17
R26 VDD.n24 VDD.t17 135.17
R27 VDD.n170 VDD.n169 129.849
R28 VDD.n121 VDD.n120 129.472
R29 VDD.n51 VDD.n50 92.5
R30 VDD.n49 VDD.n48 92.5
R31 VDD.n47 VDD.n46 92.5
R32 VDD.n45 VDD.n44 92.5
R33 VDD.n53 VDD.n52 92.5
R34 VDD.n147 VDD.n146 92.5
R35 VDD.n145 VDD.n144 92.5
R36 VDD.n143 VDD.n142 92.5
R37 VDD.n141 VDD.n140 92.5
R38 VDD.n149 VDD.n148 92.5
R39 VDD.n95 VDD.n94 92.5
R40 VDD.n93 VDD.n92 92.5
R41 VDD.n91 VDD.n90 92.5
R42 VDD.n89 VDD.n88 92.5
R43 VDD.n97 VDD.n96 92.5
R44 VDD.n14 VDD.n1 92.5
R45 VDD.n5 VDD.n4 92.5
R46 VDD.n7 VDD.n6 92.5
R47 VDD.n9 VDD.n8 92.5
R48 VDD.n11 VDD.n10 92.5
R49 VDD.n13 VDD.n12 92.5
R50 VDD.n21 VDD.n20 92.059
R51 VDD.n65 VDD.n64 92.059
R52 VDD.n161 VDD.n160 92.059
R53 VDD.n103 VDD.n102 92.059
R54 VDD.n20 VDD.n16 67.194
R55 VDD.n20 VDD.n17 67.194
R56 VDD.n20 VDD.n18 67.194
R57 VDD.n20 VDD.n19 67.194
R58 VDD.n87 VDD.n86 44.141
R59 VDD.n5 VDD.n3 44.141
R60 VDD.n86 VDD.n84 44.107
R61 VDD.n3 VDD.n2 44.107
R62 VDD.n25  U�� 43.472
R63 VDD.n33  U�� 43.472
R64 VDD.n20 VDD.n15 41.052
R65 VDD.n59 VDD.n57 39.742
R66 VDD.n59 VDD.n58 39.742
R67 VDD.n61 VDD.n60 39.742
R68 VDD.n99 VDD.n98 39.742
R69 VDD.n159 VDD.n156 39.742
R70 VDD.n159 VDD.n158 39.742
R71 VDD.n155 VDD.n154 39.742
R72 VDD.n86 VDD.n85 38
R73 VDD.n57 VDD.n56 36.774
R74 VDD.n158 VDD.n157 36.774
R75 VDD.n1 VDD.n0 30.923
R76 VDD.n64 VDD.n62 26.38
R77 VDD.n64 VDD.n61 26.38
R78 VDD.n64 VDD.n59 26.38
R79 VDD.n64 VDD.n63 26.38
R80 VDD.n102 VDD.n100 26.38
R81 VDD.n102 VDD.n99 26.38
R82 VDD.n102 VDD.n101 26.38
R83 VDD.n160 VDD.n159 26.38
R84 VDD.n160 VDD.n155 26.38
R85 VDD.n160 VDD.n153 26.38
R86 VDD.n160 VDD.n152 26.38
R87 VDD.n105 VDD.n97 22.915
R88 VDD.n23 VDD.n14 22.915
R89 VDD.n73  U�� 20.457
R90 VDD.n125 �U�� 20.457
R91 VDD.n171 VDD.t10 17.9
R92 VDD.n112 �U�� 17.9
R93 VDD.n97 VDD.n95 14.864
R94 VDD.n95 VDD.n93 14.864
R95 VDD.n93 VDD.n91 14.864
R96 VDD.n91 VDD.n89 14.864
R97 VDD.n89 VDD.n87 14.864
R98 VDD.n53 VDD.n51 14.864
R99 VDD.n51 VDD.n49 14.864
R100 VDD.n49 VDD.n47 14.864
R101 VDD.n47 VDD.n45 14.864
R102 VDD.n45 VDD.n43 14.864
R103 VDD.n43 VDD.n42 14.864
R104 VDD.n149 VDD.n147 14.864
R105 VDD.n147 VDD.n145 14.864
R106 VDD.n145 VDD.n143 14.864
R107 VDD.n143 VDD.n141 14.864
R108 VDD.n141 VDD.n139 14.864
R109 VDD.n139 VDD.n138 14.864
R110 VDD.n14 VDD.n13 14.864
R111 VDD.n13 VDD.n11 14.864
R112 VDD.n11 VDD.n9 14.864
R113 VDD.n9 VDD.n7 14.864
R114 VDD.n7 VDD.n5 14.864
R115 VDD.n67 VDD.n54 14.864
R116 VDD.n163 VDD.n150 14.864
R117 VDD.n120 VDD.t5 14.282
R118 VDD.n120 VDD.t15 14.282
R119 VDD.n169 VDD.t9 14.282
R120 VDD.n169 VDD.t11 14.282
R121 VDD.n123 VDD.n121 9.083
R122 VDD.n23 VDD.n22 8.855
R123 VDD.n22 VDD.n21 8.855
R124 VDD.n27 VDD.n26 8.855
R125 VDD.n26 VDD.n25 8.855
R126 VDD.n31 VDD.n30 8.855
R127 VDD.n30 VDD.n29 8.855
R128 VDD.n36 VDD.n34 8.855
R129 VDD.n34 VDD.n33 8.855
R130 VDD.n40 VDD.n39 8.855
R131 VDD.n39 VDD.n38 8.855
R132 VDD.n67 VDD.n66 8.855
R133 VDD.n66 VDD.n65 8.855
R134 VDD.n71 VDD.n70 8.855
R135 VDD.n70 VDD.n69 8.855
R136 VDD.n75 VDD.n74 8.855
R137 VDD.n74 VDD.n73 8.855
R138 VDD.n78 VDD.n77 8.855
R139 VDD.n77 �U�� 8.855
R140 VDD.n82 VDD.n81 8.855
R141 VDD.n81 VDD.n80 8.855
R142 VDD.n173 VDD.n172 8.855
R143 VDD.n172 VDD.n171 8.855
R144 VDD.n167 VDD.n166 8.855
R145 VDD.n166 VDD.n165 8.855
R146 VDD.n163 VDD.n162 8.855
R147 VDD.n162 VDD.n161 8.855
R148 VDD.n136 VDD.n135 8.855
R149 VDD.n135 VDD.n134 8.855
R150 VDD.n132 VDD.n131 8.855
R151 VDD.n131 VDD.n130 8.855
R152 VDD.n127 VDD.n126 8.855
R153 VDD.n126 VDD.n125 8.855
R154 VDD.n123 VDD.n122 8.855
R155 VDD.n122  U�� 8.855
R156 VDD.n118 VDD.n117 8.855
R157 VDD.n117 VDD.n116 8.855
R158 VDD.n114 VDD.n113 8.855
R159 VDD.n113 VDD.n112 8.855
R160 VDD.n110 VDD.n109 8.855
R161 VDD.n109 VDD.n108 8.855
R162 VDD.n105 VDD.n104 8.855
R163 VDD.n104 VDD.n103 8.855
R164 VDD.n54 VDD.n53 8.051
R165 VDD.n150 VDD.n149 8.051
R166 VDD.n173 VDD.n170 6.193
R167 VDD.n28 VDD.n23 4.795
R168 VDD.n28 VDD.n27 4.65
R169 VDD.n32 VDD.n31 4.65
R170 VDD.n37 VDD.n36 4.65
R171 VDD.n41 VDD.n40 4.65
R172 VDD.n68 VDD.n67 4.65
R173 VDD.n72 VDD.n71 4.65
R174 VDD.n76 VDD.n75 4.65
R175 VDD.n79 VDD.n78 4.65
R176 VDD.n83 VDD.n82 4.65
R177 VDD.n174 VDD.n173 4.65
R178 VDD.n168 VDD.n167 4.65
R179 VDD.n164 VDD.n163 4.65
R180 VDD.n137 VDD.n136 4.65
R181 VDD.n133 VDD.n132 4.65
R182 VDD.n128 VDD.n127 4.65
R183 VDD.n124 VDD.n123 4.65
R184 VDD.n119 VDD.n118 4.65
R185 VDD.n115 VDD.n114 4.65
R186 VDD.n111 VDD.n110 4.65
R187 VDD.n106 VDD.n105 4.65
R188 VDD.n110 VDD.n107 2.89
R189 VDD.n80 �U�� 2.557
R190 VDD.n116 @i�]!V 2.557
R191 VDD.n132 VDD.n129 2.477
R192 VDD.n27 VDD.n24 2.064
R193 VDD.n36 VDD.n35 2.064
R194 VDD.n68 VDD.n41 0.29
R195 VDD.n164 VDD.n137 0.29
R196 VDD.n106 VDD 0.207
R197 VDD.n83 VDD.n79 0.181
R198 VDD.n124 VDD.n119 0.181
R199 VDD.n32 VDD.n28 0.157
R200 VDD.n37 VDD.n32 0.157
R201 VDD.n41 VDD.n37 0.145
R202 VDD.n72 VDD.n68 0.145
R203 VDD.n76 VDD.n72 0.145
R204 VDD.n79 VDD.n76 0.145
R205 VDD.n174 VDD.n168 0.145
R206 VDD.n168 VDD.n164 0.145
R207 VDD.n137 VDD.n133 0.145
R208 VDD.n133 VDD.n128 0.145
R209 VDD.n128 VDD.n124 0.145
R210 VDD.n119 VDD.n115 0.145
R211 VDD.n115 VDD.n111 0.145
R212 VDD.n111 VDD.n106 0.145
R213 VDD VDD.n83 0.133
R214 VDD VDD.n174 0.012
R215 a_797_1051.n0 a_797_1051.t0 228.369
R216 a_797_1051.n0 a_797_1051.t3 219.778
R217 a_797_1051.n1 a_797_1051.n0 42.29
R218 a_797_1051.n1 a_797_1051.t1 14.282
R219 a_797_1051.t2 a_797_1051.n1 14.282
R220 a_864_209.n1 a_864_209.t4 512.525
R221 a_864_209.n1 a_864_209.t5 371.139
R222 a_864_209.n3 a_864_209.n0 343.684
R223 a_864_209.n2 a_864_209.n1 303.065
R224 a_864_209.n2 a_864_209.t6 227.134
R225 a_864_209.n8 a_864_209.n7 208.452
R226 a_864_209.n10 a_864_209.n8 142.275
R227 a_864_209.n8 a_864_209.n3 86.587
R228 a_864_209.n7 a_864_209.n6 30
R229 a_864_209.n5 a_864_209.n4 24.383
R230 a_864_209.n7 a_864_209.n5 23.684
R231 a_864_209.n10 a_864_209.n9 15.001
R232 a_864_209.n0 a_864_209.t0 14.282
R233 a_864_209.n0 a_864_209.t2 14.282
R234 a_864_209.n11 a_864_209.n10 12.632
R235 a_864_209.n3 a_864_209.n2 10.343
R236 Y.n5 Y.n4 328.169
R237 Y.n5 Y.n0 215.564
R238 Y.n4 Y.n3 30
R239 Y.n2 Y.n1 24.383
R240 Y.n4 Y.n2 23.684
R241 Y.n0 Y.t1 14.282
R242 Y.n0 Y.t0 14.282
R243 Y.n6 Y.n5 4.65
R244 Y.n6 Y 0.046
R245 B.n0 B.t0 472.359
R246 B.n0 B.t1 384.527
R247 B.n1 B.t2 287.037
R248 B.n1 B.n0 210.673
R249 B.n2 B.n1 4.65
R250 B.n2 B 0.046
R251 C.n0 C.t0 470.752
R252 C.n0 C.t1 384.527
R253 C.n1 C.t2 314.896
R254 C.n1 C.n0 182.932
R255 C.n2 C.n1 4.65
R256 C.n2 C 0.046
R257 a_112_101.n10 a_112_101.n9 93.333
R258 a_112_101.n12 a_112_101.n11 68.43
R259 a_112_101.n3 a_112_101.n2 51.907
R260 a_112_101.n3 a_112_101.n1 51.594
R261 a_112_101.t0 a_112_101.n3 38.864
R262 a_112_101.n7 a_112_101.n6 38.626
R263 a_112_101.n6 a_112_101.n5 35.955
R264 a_112_101.t1 a_112_101.n8 8.137
R265 a_112_101.t0 a_112_101.n0 6.109
R266 a_112_101.t1 a_112_101.n7 4.864
R267 a_112_101.t0 a_112_101.n4 3.871
R268 a_112_101.t0 a_112_101.n13 2.535
R269 a_112_101.n13 a_112_101.t1 1.145
R270 a_112_101.t1 a_112_101.n12 0.763
R271 a_112_101.n12 a_112_101.n10 0.185
R272 GND.n32 GND.n31 237.558
R273 GND.n84 GND.n83 237.558
R274 GND.n29 GND.n28 210.82
R275 GND.n86 GND.n85 210.82
R276 GND.n64 GND.n63 172.612
R277 GND.n52 GND.n51 40.431
R278 GND.n37 GND.n36 40.003
R279 GND.n21 GND.n20 37.582
R280 GND.n93 GND.n92 37.582
R281 GND.t0 GND.n18 32.601
R282 GND.n18 GND.n17 21.734
R283 GND.n4 GND.n3 20.705
R284 GND.n10 GND.n9 20.705
R285 GND.n22 GND.n21 20.705
R286 GND.n98 GND.n97 20.705
R287 GND.n53 GND.n52 20.705
R288 GND.n44 GND.n43 20.705
R289 GND.n38 GND.n37 20.705
R290 GND.n94 GND.n93 20.705
R291 GND.n3 GND.n2 19.952
R292 GND.n30 GND.n29 18.953
R293 GND.n87 GND.n86 18.953
R294 GND.n36 GND.n35 17.258
R295 GND.n20 GND.t0 15.644
R296 GND.n92 GND.t1 15.644
R297 GND.n33 GND.n30 14.864
R298 GND.n88 GND.n87 14.864
R299 GND.n51 GND.t4 13.654
R300 GND.n20 GND.n19 13.541
R301 GND.n92 GND.n91 13.541
R302 GND.n55 GND.n53 9.29
R303 GND.n61 GND.n60 9.154
R304 GND.n66 GND.n65 9.154
R305 GND.n69 GND.n68 9.154
R306 GND.n72 GND.n71 9.154
R307 GND.n75 GND.n74 9.154
R308 GND.n78 GND.n77 9.154
R309 GND.n81 GND.n80 9.154
R310 GND.n88 GND.n84 9.154
R311 GND.n95 GND.n90 9.154
R312 GND.n100 GND.n99 9.154
R313 GND.n55 GND.n54 9.154
R314 GND.n48 GND.n47 9.154
R315 GND.n45 GND.n42 9.154
R316 GND.n40 GND.n39 9.154
R317 GND.n33 GND.n32 9.154
R318 GND.n26 GND.n25 9.154
R319 GND.n23 GND.n14 9.154
R320 GND.n12 GND.n11 9.154
R321 GND.n6 GND.n5 9.154
R322 GND.t4 GND.n50 7.04
R323 GND.n7 GND.n1 4.795
R324 GND.n59 GND.n58 4.65
R325 GND.n7 GND.n6 4.65
R326 GND.n13 GND.n12 4.65
R327 GND.n24 GND.n23 4.65
R328 GND.n27 GND.n26 4.65
R329 GND.n34 GND.n33 4.65
R330 GND.n41 GND.n40 4.65
R331 GND.n46 GND.n45 4.65
R332 GND.n49 GND.n48 4.65
R333 GND.n56 GND.n55 4.65
R334 GND.n101 GND.n100 4.65
R335 GND.n96 GND.n95 4.65
R336 GND.n89 GND.n88 4.65
R337 GND.n82 GND.n81 4.65
R338 GND.n79 GND.n78 4.65
R339 GND.n76 GND.n75 4.65
R340 GND.n73 GND.n72 4.65
R341 GND.n70 GND.n69 4.65
R342 GND.n67 GND.n66 4.65
R343 GND.n62 GND.n61 4.65
R344 GND.n16 GND.n15 4.504
R345 GND.n6 GND.n4 4.129
R346 GND.n45 GND.n44 4.129
R347 GND.n100 GND.n98 4.129
R348 GND.n66 GND.n64 4.129
R349 GND.n23 GND.n22 3.716
R350 GND.t0 GND.n16 2.452
R351 GND.n40 GND.n38 1.032
R352 GND.n95 GND.n94 1.032
R353 GND.n1 GND.n0 0.474
R354 GND.n58 GND.n57 0.474
R355 GND.n9 GND.n8 0.376
R356 GND.n34 GND.n27 0.29
R357 GND.n89 GND.n82 0.29
R358 GND.n59 GND 0.207
R359 GND.n12 GND.n10 0.206
R360 GND.n56 GND.n49 0.181
R361 GND.n73 GND.n70 0.181
R362 GND.n13 GND.n7 0.157
R363 GND.n24 GND.n13 0.157
R364 GND.n27 GND.n24 0.145
R365 GND.n41 GND.n34 0.145
R366 GND.n46 GND.n41 0.145
R367 GND.n49 GND.n46 0.145
R368 GND.n101 GND.n96 0.145
R369 GND.n96 GND.n89 0.145
R370 GND.n82 GND.n79 0.145
R371 GND.n79 GND.n76 0.145
R372 GND.n76 GND.n73 0.145
R373 GND.n70 GND.n67 0.145
R374 GND.n67 GND.n62 0.145
R375 GND.n62 GND.n59 0.145
R376 GND GND.n56 0.133
R377 GND GND.n101 0.012
C5 VDD GND 3.31fF
C6 a_112_101.n0 GND 0.02fF
C7 a_112_101.n1 GND 0.09fF
C8 a_112_101.n2 GND 0.07fF
C9 a_112_101.n3 GND 0.04fF
C10 a_112_101.n4 GND 0.01fF
C11 a_112_101.n5 GND 0.04fF
C12 a_112_101.n6 GND 0.04fF
C13 a_112_101.n7 GND 0.02fF
C14 a_112_101.n8 GND 0.05fF
C15 a_112_101.n9 GND 0.02fF
C16 a_112_101.n10 GND 0.14fF
C17 a_112_101.n11 GND 0.08fF
C18 a_112_101.n12 GND 0.08fF
C19 a_112_101.t1 GND 0.22fF
C20 a_112_101.n13 GND 0.01fF
C21 Y.n0 GND 0.57fF
C22 Y.n1 GND 0.04fF
C23 Y.n2 GND 0.05fF
C24 Y.n3 GND 0.03fF
C25 Y.n4 GND 0.25fF
C26 Y.n5 GND 0.63fF
C27 Y.n6 GND 0.01fF
C28 a_864_209.n0 GND 0.50fF
C29 a_864_209.n1 GND 0.32fF
C30 a_864_209.n2 GND 0.45fF
C31 a_864_209.n3 GND 0.50fF
C32 a_864_209.n4 GND 0.03fF
C33 a_864_209.n5 GND 0.04fF
C34 a_864_209.n6 GND 0.03fF
C35 a_864_209.n7 GND 0.09fF
C36 a_864_209.n8 GND 0.31fF
C37 a_864_209.n9 GND 0.06fF
C38 a_864_209.n10 GND 0.04fF
C39 a_864_209.n11 GND 0.04fF
C40 a_797_1051.n0 GND 0.52fF
C41 a_797_1051.n1 GND 0.22fF
C42 VDD.n1 GND 0.03fF
C43 VDD.n2 GND 0.08fF
C44 VDD.n3 GND 0.02fF
C45 VDD.n4 GND 0.02fF
C46 VDD.n5 GND 0.05fF
C47 VDD.n6 GND 0.02fF
C48 VDD.n7 GND 0.02fF
C49 VDD.n8 GND 0.02fF
C50 VDD.n9 GND 0.02fF
C51 VDD.n10 GND 0.02fF
C52 VDD.n11 GND 0.02fF
C53 VDD.n12 GND 0.02fF
C54 VDD.n13 GND 0.02fF
C55 VDD.n14 GND 0.03fF
C56 VDD.n15 GND 0.01fF
C57 VDD.n20 GND 0.37fF
C58 VDD.n21 GND 0.22fF
C59 VDD.n22 GND 0.02fF
C60 VDD.n23 GND 0.03fF
C61 VDD.n24 GND 0.05fF
C62 VDD.n25 GND 0.17fF
C63 VDD.n26 GND 0.01fF
C64 VDD.n27 GND 0.01fF
C65 VDD.n28 GND 0.05fF
C66 VDD.n29 GND 0.14fF
C67 VDD.n30 GND 0.01fF
C68 VDD.n31 GND 0.02fF
C69 VDD.n32 GND 0.02fF
C70 VDD.n33 GND 0.17fF
C71 VDD.n34 GND 0.01fF
C72 VDD.n35 GND 0.05fF
C73 VDD.n36 GND 0.01fF
C74 VDD.n37 GND 0.02fF
C75 VDD.n38 GND 0.22fF
C76 VDD.n39 GND 0.01fF
C77 VDD.n40 GND 0.02fF
C78 VDD.n41 GND 0.03fF
C79 VDD.n42 GND 0.05fF
C80 VDD.n43 GND 0.02fF
C81 VDD.n44 GND 0.02fF
C82 VDD.n45 GND 0.02fF
C83 VDD.n46 GND 0.02fF
C84 VDD.n47 GND 0.02fF
C85 VDD.n48 GND 0.02fF
C86 VDD.n49 GND 0.02fF
C87 VDD.n50 GND 0.02fF
C88 VDD.n51 GND 0.02fF
C89 VDD.n52 GND 0.02fF
C90 VDD.n53 GND 0.01fF
C91 VDD.n54 GND 0.02fF
C92 VDD.n55 GND 0.02fF
C93 VDD.n56 GND 0.15fF
C94 VDD.n57 GND 0.02fF
C95 VDD.n58 GND 0.02fF
C96 VDD.n60 GND 0.02fF
C97 VDD.n64 GND 0.22fF
C98 VDD.n65 GND 0.22fF
C99 VDD.n66 GND 0.01fF
C100 VDD.n67 GND 0.02fF
C101 VDD.n68 GND 0.03fF
C102 VDD.n69 GND 0.20fF
C103 VDD.n70 GND 0.01fF
C104 VDD.n71 GND 0.02fF
C105 VDD.n72 GND 0.02fF
C106 VDD.n73 GND 0.14fF
C107 VDD.n74 GND 0.01fF
C108 VDD.n75 GND 0.02fF
C109 VDD.n76 GND 0.02fF
C110 VDD.n77 GND 0.01fF
C111 VDD.n78 GND 0.02fF
C112 VDD.n79 GND 0.02fF
C113 VDD.n80 GND 0.12fF
C114 VDD.n81 GND 0.01fF
C115 VDD.n82 GND 0.02fF
C116 VDD.n83 GND 0.02fF
C117 VDD.n84 GND 0.11fF
C118 VDD.n85 GND 0.02fF
C119 VDD.n86 GND 0.02fF
C120 VDD.n87 GND 0.05fF
C121 VDD.n88 GND 0.02fF
C122 VDD.n89 GND 0.02fF
C123 VDD.n90 GND 0.02fF
C124 VDD.n91 GND 0.02fF
C125 VDD.n92 GND 0.02fF
C126 VDD.n93 GND 0.02fF
C127 VDD.n94 GND 0.02fF
C128 VDD.n95 GND 0.02fF
C129 VDD.n96 GND 0.03fF
C130 VDD.n97 GND 0.03fF
C131 VDD.n98 GND 0.02fF
C132 VDD.n102 GND 0.37fF
C133 VDD.n103 GND 0.22fF
C134 VDD.n104 GND 0.02fF
C135 VDD.n105 GND 0.03fF
C136 VDD.n106 GND 0.02fF
C137 VDD.n107 GND 0.05fF
C138 VDD.n108 GND 0.20fF
C139 VDD.n109 GND 0.01fF
C140 VDD.n110 GND 0.01fF
C141 VDD.n111 GND 0.02fF
C142 VDD.n112 GND 0.13fF
C143 VDD.n113 GND 0.01fF
C144 VDD.n114 GND 0.02fF
C145 VDD.n115 GND 0.02fF
C146 VDD.n116 GND 0.12fF
C147 VDD.n117 GND 0.01fF
C148 VDD.n118 GND 0.02fF
C149 VDD.n119 GND 0.02fF
C150 VDD.n120 GND 0.07fF
C151 VDD.n121 GND 0.04fF
C152 VDD.n122 GND 0.01fF
C153 VDD.n123 GND 0.02fF
C154 VDD.n124 GND 0.02fF
C155 VDD.n125 GND 0.14fF
C156 VDD.n126 GND 0.01fF
C157 VDD.n127 GND 0.02fF
C158 VDD.n128 GND 0.02fF
C159 VDD.n129 GND 0.05fF
C160 VDD.n130 GND 0.20fF
C161 VDD.n131 GND 0.01fF
C162 VDD.n132 GND 0.01fF
C163 VDD.n133 GND 0.02fF
C164 VDD.n134 GND 0.22fF
C165 VDD.n135 GND 0.01fF
C166 VDD.n136 GND 0.02fF
C167 VDD.n137 GND 0.03fF
C168 VDD.n138 GND 0.05fF
C169 VDD.n139 GND 0.02fF
C170 VDD.n140 GND 0.02fF
C171 VDD.n141 GND 0.02fF
C172 VDD.n142 GND 0.02fF
C173 VDD.n143 GND 0.02fF
C174 VDD.n144 GND 0.02fF
C175 VDD.n145 GND 0.02fF
C176 VDD.n146 GND 0.02fF
C177 VDD.n147 GND 0.02fF
C178 VDD.n148 GND 0.02fF
C179 VDD.n149 GND 0.01fF
C1