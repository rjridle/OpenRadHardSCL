magic
tech sky130A
magscale 1 2
timestamp 1647814309
<< metal1 >>
rect 55 1505 89 1539
rect 131 871 165 905
rect 353 797 387 831
rect 1167 797 1201 831
rect 1833 797 1867 831
rect 55 13 89 47
use votern3x1_pcell  votern3x1_pcell_0 pcells
timestamp 1647814117
transform 1 0 0 0 1 1
box -84 0 2082 1575
use li1_M1_contact  li1_M1_contact_3 pcells
timestamp 1646004885
transform -1 0 1850 0 -1 814
box -53 -33 29 33
<< labels >>
rlabel metal1 1833 797 1867 831 1 YN
rlabel metal1 1167 797 1201 831 1 C
rlabel metal1 353 797 387 831 1 B
rlabel metal1 131 871 165 905 1 A
rlabel metal1 55 13 89 47 1 VSS
rlabel metal1 55 1505 89 1539 1 VDD
<< end >>
