* SPICE3 file created from TMRDFFRNQX1.ext - technology: sky130A

.subckt TMRDFFRNQX1 Q D CLK RN VDD GND
X0 VDD.t171 RN.t0 a_10507_187.t4 VDD.t170 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X1 GND a_10507_187.t7 a_10451_103.t0 GND sky130_fd_pr__nfet_01v8 ad=4.9019p pd=4.107u as=0p ps=0u w=0u l=0u
X2 a_14189_1050.t2 a_10637_1050.t7 VDD.t127 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X3 a_10959_989.t1 a_10637_1050.t8 VDD.t95  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X4 a_599_989.t2 D.t0 VDD.t1 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X5 a_16421_1051.t5 a_14511_989.t5 a_15932_209.t4  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X6 a_5327_187.t3 CLK.t0 VDD.t52 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X7 VDD.t5 a_599_989.t7 a_2141_1050.t4  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X8 a_9331_989.t4 a_9009_1050.t7 VDD.t60 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X9 VDD.t131 CLK.t1 a_277_1050.t6  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X10 VDD.t44 a_5457_1050.t7 a_5779_989.t6 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X11 VDD.t42 a_5457_1050.t8 a_9009_1050.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X12 VDD.t109 a_277_1050.t7 a_3829_1050.t3 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X13 VDD.t169 RN.t2 a_5779_989.t3  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X14 VDD.t191 a_9331_989.t5 a_9009_1050.t5 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X15 VDD.t101 CLK.t2 a_10637_1050.t3  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X16 VDD.t79 CLK.t3 a_10507_187.t2 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X17 a_9331_989.t2 a_5327_187.t7 VDD.t29  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X18 a_14189_1050.t4 RN.t3 VDD.t167 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X19 a_10959_989.t5 D.t2 VDD.t173  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X20 GND a_9331_989.t7 a_16318_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X21 a_599_989.t5 RN.t4 VDD.t165 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X22 a_3829_1050.t6 a_4151_989.t5 VDD.t3  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X23 VDD.t177 a_14511_989.t6 a_15757_1051.t3 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X24 a_10637_1050.t5 a_10507_187.t8 VDD.t123  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X25 a_147_187.t6 CLK.t4 VDD.t193 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X26 a_4151_989.t1 a_3829_1050.t7 VDD.t25  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X27 GND a_5457_1050.t10 a_8823_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X28 a_9009_1050.t1 a_5457_1050.t9 VDD.t54 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X29 a_15757_1051.t5 a_9331_989.t6 VDD.t27  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X30 VDD.t72 a_14189_1050.t7 a_14511_989.t1 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X31 VDD.t15 a_10959_989.t8 a_12501_1050.t4  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X32 GND a_5457_1050.t11 a_6233_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X33 VDD.t81 a_147_187.t9 a_2141_1050.t1 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X34 VDD.t66 a_599_989.t8 a_277_1050.t2  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X35 VDD.t87 D.t4 a_5779_989.t1 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X36 VDD.t163 RN.t6 a_9009_1050.t3  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X37 VDD.t211 a_2141_1050.t5 a_147_187.t4 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X38 VDD.t19 a_5327_187.t8 a_5457_1050.t4  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X39 VDD.t31 a_7321_1050.t5 a_5327_187.t0 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X40 GND a_9009_1050.t9 a_9806_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X41 a_14189_1050.t5 a_14511_989.t8 VDD.t175  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X42 a_10959_989.t4 RN.t8 VDD.t161 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X43 a_147_187.t2 RN.t9 VDD.t159  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X44 GND a_5779_989.t8 a_7216_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X45 GND a_147_187.t12 a_91_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X46 GND a_7321_1050.t6 a_7861_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X47 a_4151_989.t3 a_147_187.t10 VDD.t203 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X48 a_7321_1050.t3 a_5327_187.t9 VDD.t97  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X49 a_15932_209.t2 a_4151_989.t6 a_16421_1051.t3 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X50 Q a_15932_209.t8 GND.t4 GND sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=0p ps=0u w=0u l=0u
X51 VDD.t58 a_10959_989.t9 a_10637_1050.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X52 GND a_5327_187.t10 a_5271_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X53 a_15757_1051.t2 a_14511_989.t9 VDD.t17 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X54 VDD.t121 a_10507_187.t10 a_14511_989.t4  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X55 VDD.t119 a_10507_187.t11 a_12501_1050.t1 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X56 VDD.t83 a_15932_209.t7 Q.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X57 a_277_1050.t4 a_147_187.t11 VDD.t68 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X58 a_16421_1051.t7 a_4151_989.t7 a_15757_1051.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X59 VDD.t195 a_9009_1050.t8 a_9331_989.t3 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X60 a_10507_187.t0 a_12501_1050.t5 VDD.t56  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X61 a_10637_1050.t6 a_10959_989.t10 VDD.t199 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X62 a_10507_187.t5 RN.t11 VDD.t157  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X63 a_7321_1050.t1 a_5779_989.t9 VDD.t189 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X64 VDD.t205 a_277_1050.t8 a_599_989.t6  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X65 a_15932_209.t3 a_14511_989.t11 a_16421_1051.t4 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X66 VDD.t155 RN.t12 a_599_989.t4  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X67 VDD.t38 a_4151_989.t8 a_3829_1050.t5 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X68 GND a_12501_1050.t6 a_13041_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X69 GND a_277_1050.t11 a_3643_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X70 VDD.t33 a_5779_989.t10 a_5457_1050.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X71 VDD.t153 RN.t14 a_5327_187.t5 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X72 a_16421_1051.t0 a_9331_989.t8 a_15757_1051.t7  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X73 a_2141_1050.t3 a_599_989.t10 VDD.t85 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X74 a_277_1050.t5 CLK.t7 VDD.t70  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X75 a_3829_1050.t2 a_277_1050.t9 VDD.t9 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X76 a_5779_989.t5 a_5457_1050.t12 VDD.t13  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X77 a_10637_1050.t2 CLK.t8 VDD.t74 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X78 a_10507_187.t6 CLK.t9 VDD.t183  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X79 VDD.t50 a_10637_1050.t10 a_14189_1050.t1 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X80 VDD.t129 a_10637_1050.t11 a_10959_989.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X81 GND a_3829_1050.t8 a_4626_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X82 VDD.t151 RN.t15 a_3829_1050.t1 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X83 VDD.t179 D.t6 a_599_989.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X84 GND a_599_989.t12 a_2036_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X85 GND a_10637_1050.t12 a_14003_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X86 GND a_2141_1050.t7 a_2681_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X87 a_599_989.t0 a_277_1050.t10 VDD.t11 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X88 VDD.t21 CLK.t11 a_5457_1050.t6  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X89 VDD.t40 CLK.t12 a_5327_187.t1 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X90 a_2141_1050.t0 a_147_187.t13 VDD.t76  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X91 a_277_1050.t1 a_599_989.t11 VDD.t93 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X92 a_3829_1050.t0 RN.t16 VDD.t149  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X93 a_5779_989.t0 D.t7 VDD.t7 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X94 a_9009_1050.t2 RN.t17 VDD.t147  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X95 a_5327_187.t2 a_7321_1050.t7 VDD.t48 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X96 VDD.t207 a_5327_187.t12 a_9331_989.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X97 GND a_9331_989.t11 a_15652_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X98 GND a_14189_1050.t8 a_14986_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X99 a_147_187.t3 a_2141_1050.t6 VDD.t125 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X100 a_5457_1050.t3 a_5327_187.t13 VDD.t89  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X101 VDD.t145 RN.t18 a_14189_1050.t3 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X102 VDD.t181 D.t8 a_10959_989.t6  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X103 VDD.t91 CLK.t14 a_147_187.t5 0�3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X104 VDD.t135 a_5779_989.t11 a_7321_1050.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X105 VDD.t23 a_3829_1050.t9 a_4151_989.t0 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X106 VDD.t62 a_9331_989.t9 a_15757_1051.t4 VDD.t61 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X107 GND a_277_1050.t12 a_1053_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X108 a_14511_989.t3 a_10507_187.t13 VDD.t117 �3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X109 a_12501_1050.t0 a_10507_187.t14 VDD.t115 �3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X110 a_9009_1050.t6 a_9331_989.t10 VDD.t197 �3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X111 a_5779_989.t2 RN.t21 VDD.t143 �3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X112 Q.t0 a_15932_209.t9 VDD.t111 �3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X113 a_5457_1050.t5 CLK.t16 VDD.t99 �3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X114 a_15757_1051.t6 a_9331_989.t12 a_16421_1051.t6 �3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X115 VDD.t201 a_14511_989.t13 a_14189_1050.t6 �3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X116 GND a_4151_989.t13 a_16984_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X117 VDD.t141 RN.t23 a_147_187.t1 �3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X118 VDD.t187 a_147_187.t14 a_4151_989.t2 VDD.t186 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X119 VDD.t105 a_5327_187.t15 a_7321_1050.t2 �3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X120 a_16421_1051.t2 a_4151_989.t11 a_15932_209.t1 VDD.t106 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X121 GND a_10637_1050.t9 a_11413_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X122 a_14511_989.t0 a_14189_1050.t9 VDD.t35 �3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X123 a_12501_1050.t3 a_10959_989.t12 VDD.t185  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X124 VDD.t139 RN.t25 a_10959_989.t3 VDD.t138 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X125 a_5457_1050.t2 a_5779_989.t12 VDD.t133 �3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X126 a_5327_187.t4 RN.t26 VDD.t137  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X127 VDD.t103 a_147_187.t15 a_277_1050.t3 VDD.t102 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X128 a_15757_1051.t0 a_4151_989.t12 a_16421_1051.t1 �3� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X129 GND a_10959_989.t7 a_12396_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X130 VDD.t113 a_10507_187.t15 a_10637_1050.t4  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X131 VDD.t64 a_12501_1050.t7 a_10507_187.t1 VDD.t63 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
C0 CLK D 0.45fF
C1 CLK RN 1.13fF
C2 CLK VDD 8.54fF
C3 D RN 12.60fF
C4 D VDD 0.88fF
C5 RN VDD 2.66fF
C6 Q VDD 1.05fF
R0 RN.n17 RN.t15 479.223
R1 RN.n8 RN.t6 479.223
R2 RN.n0 RN.t18 479.223
R3 RN.n23 RN.t4 454.685
R4 RN.n20 RN.t9 454.685
R5 RN.n14 RN.t21 454.685
R6 RN.n11 RN.t26 454.685
R7 RN.n5 RN.t8 454.685
R8 RN.n2 RN.t11 454.685
R9 RN.n23 RN.t12 428.979
R10 RN.n20 RN.t23 428.979
R11 RN.n14 RN.t2 428.979
R12 RN.n11 RN.t14 428.979
R13 RN.n5 RN.t25 428.979
R14 RN.n2 RN.t0 428.979
R15 RN.n17 RN.t16 375.52
R16 RN.n8 RN.t17 375.52
R17 RN.n0 RN.t3 375.52
R18 RN.n24 RN.n23 254.865
R19 RN.n21 RN.n20 254.865
R20 RN.n15 RN.n14 254.865
R21 RN.n12 RN.n11 254.865
R22 RN.n6 RN.n5 254.865
R23 RN.n3 RN.n2 254.865
R24 RN.n18 RN.n17 252.188
R25 RN.n9 RN.n8 252.188
R26 RN.n1 RN.n0 252.188
R27 RN.n18 RN.t20 231.854
R28 RN.n9 RN.t7 231.854
R29 RN.n1 RN.t24 231.854
R30 RN.n24 RN.t19 228.106
R31 RN.n21 RN.t10 228.106
R32 RN.n15 RN.t5 228.106
R33 RN.n12 RN.t1 228.106
R34 RN.n6 RN.t22 228.106
R35 RN.n3 RN.t13 228.106
R36 RN.n10 RN.n7 10.293
R37 RN.n19 RN.n16 10.293
R38 RN.n4 RN.n1 7.325
R39 RN.n7 RN.n4 5.94
R40 RN.n16 RN.n13 5.94
R41 RN.n25 RN.n22 5.94
R42 RN.n4 RN.n3 4.65
R43 RN.n7 RN.n6 4.65
R44 RN.n10 RN.n9 4.65
R45 RN.n13 RN.n12 4.65
R46 RN.n16 RN.n15 4.65
R47 RN.n19 RN.n18 4.65
R48 RN.n22 RN.n21 4.65
R49 RN.n25 RN.n24 4.65
R50 RN.n13 RN.n10 2.675
R51 RN.n22 RN.n19 2.675
R52 RN.n25 RN 0.046
R53 a_10507_187.n10 a_10507_187.t15 512.525
R54 a_10507_187.n8 a_10507_187.t11 472.359
R55 a_10507_187.n6 a_10507_187.t10 472.359
R56 a_10507_187.n11 a_10507_187.t7 417.109
R57 a_10507_187.n8 a_10507_187.t14 384.527
R58 a_10507_187.n6 a_10507_187.t13 384.527
R59 a_10507_187.n10 a_10507_187.t8 371.139
R60 a_10507_187.n9 a_10507_187.t12 370.613
R61 a_10507_187.n7 a_10507_187.t9 370.613
R62 a_10507_187.n16 a_10507_187.n14 363.934
R63 a_10507_187.n11 a_10507_187.n10 179.837
R64 a_10507_187.n4 a_10507_187.n3 161.352
R65 a_10507_187.n9 a_10507_187.n8 127.096
R66 a_10507_187.n7 a_10507_187.n6 127.096
R67 a_10507_187.n14 a_10507_187.n5 123.481
R68 a_10507_187.n5 a_10507_187.n1 95.095
R69 a_10507_187.n4 a_10507_187.n2 95.095
R70 a_10507_187.n5 a_10507_187.n4 66.258
R71 a_10507_187.n16 a_10507_187.n15 30
R72 a_10507_187.n17 a_10507_187.n0 24.383
R73 a_10507_187.n17 a_10507_187.n16 23.684
R74 a_10507_187.n1 a_10507_187.t4 14.282
R75 a_10507_187.n1 a_10507_187.t5 14.282
R76 a_10507_187.n2 a_10507_187.t2 14.282
R77 a_10507_187.n2 a_10507_187.t6 14.282
R78 a_10507_187.n3 a_10507_187.t1 14.282
R79 a_10507_187.n3 a_10507_187.t0 14.282
R80 a_10507_187.n12 a_10507_187.n11 12.222
R81 a_10507_187.n13 a_10507_187.n7 10.046
R82 a_10507_187.n12 a_10507_187.n9 4.65
R83 a_10507_187.n14 a_10507_187.n13 4.65
R84 a_10507_187.n13 a_10507_187.n12 4.035
R85 VDD.n835 VDD.n824 144.705
R86 VDD.n910 VDD.n903 144.705
R87 VDD.n967 VDD.n960 144.705
R88 VDD.n1042 VDD.n1035 144.705
R89 VDD.n1117 VDD.n1110 144.705
R90 VDD.n1174 VDD.n1167 144.705
R91 VDD.n1249 VDD.n1242 144.705
R92 VDD.n1324 VDD.n1317 144.705
R93 VDD.n1381 VDD.n1374 144.705
R94 VDD.n700 VDD.n693 144.705
R95 VDD.n1456 VDD.n1449 144.705
R96 VDD.n643 VDD.n636 144.705
R97 VDD.n568 VDD.n561 144.705
R98 VDD.n493 VDD.n486 144.705
R99 VDD.n436 VDD.n429 144.705
R100 VDD.n361 VDD.n354 144.705
R101 VDD.n286 VDD.n279 144.705
R102 VDD.n229 VDD.n222 144.705
R103 VDD.n172 VDD.n165 144.705
R104 VDD.n119 VDD.n112 144.705
R105 VDD.n66 VDD.n55 144.705
R106 VDD.n801 VDD.t66 143.754
R107 VDD.n877 VDD.t155 143.754
R108 VDD.n1009 VDD.t141 143.754
R109 VDD.n1084 VDD.t38 143.754
R110 VDD.n1216 VDD.t33 143.754
R111 VDD.n1291 VDD.t169 143.754
R112 VDD.n1423 VDD.t153 143.754
R113 VDD.n709 VDD.t191 143.754
R114 VDD.n577 VDD.t58 143.754
R115 VDD.n502 VDD.t139 143.754
R116 VDD.n370 VDD.t171 143.754
R117 VDD.n295 VDD.t201 143.754
R118 VDD.n935 VDD.t81 143.754
R119 VDD.n1142 VDD.t187 143.754
R120 VDD.n1349 VDD.t105 143.754
R121 VDD.n646 VDD.t207 143.754
R122 VDD.n439 VDD.t119 143.754
R123 VDD.n232 VDD.t121 143.754
R124 VDD.n197 VDD.t27 135.539
R125 VDD.n175 VDD.t177 135.539
R126 VDD.n766 VDD.t68 135.17
R127 VDD.n842 VDD.t11 135.17
R128 VDD.n913 VDD.t85 135.17
R129 VDD.n974 VDD.t125 135.17
R130 VDD.n1049 VDD.t9 135.17
R131 VDD.n1120 VDD.t25 135.17
R132 VDD.n1181 VDD.t89 135.17
R133 VDD.n1256 VDD.t13 135.17
R134 VDD.n1327 VDD.t189 135.17
R135 VDD.n1388 VDD.t48 135.17
R136 VDD.n1463 VDD.t54 135.17
R137 VDD.n668 VDD.t60 135.17
R138 VDD.n607 VDD.t123 135.17
R139 VDD.n532 VDD.t95 135.17
R140 VDD.n461 VDD.t185 135.17
R141 VDD.n400 VDD.t56 135.17
R142 VDD.n325 VDD.t127 135.17
R143 VDD.n254 VDD.t35 135.17
R144 VDD.n35 VDD.t111 135.17
R145 VDD.n24 VDD.t83 135.17
R146 VDD.n185 VDD.n184 129.849
R147 VDD.n776 VDD.n775 129.472
R148 VDD.n792 VDD.n791 129.472
R149 VDD.n852 VDD.n851 129.472
R150 VDD.n868 VDD.n867 129.472
R151 VDD.n927 VDD.n926 129.472
R152 VDD.n984 VDD.n983 129.472
R153 VDD.n1000 VDD.n999 129.472
R154 VDD.n1059 VDD.n1058 129.472
R155 VDD.n1075 VDD.n1074 129.472
R156 VDD.n1134 VDD.n1133 129.472
R157 VDD.n1191 VDD.n1190 129.472
R158 VDD.n1207 VDD.n1206 129.472
R159 VDD.n1266 VDD.n1265 129.472
R160 VDD.n1282 VDD.n1281 129.472
R161 VDD.n1341 VDD.n1340 129.472
R162 VDD.n1398 VDD.n1397 129.472
R163 VDD.n1414 VDD.n1413 129.472
R164 VDD.n730 VDD.n729 129.472
R165 VDD.n718 VDD.n717 129.472
R166 VDD.n656 VDD.n655 129.472
R167 VDD.n598 VDD.n597 129.472
R168 VDD.n586 VDD.n585 129.472
R169 VDD.n523 VDD.n522 129.472
R170 VDD.n511 VDD.n510 129.472
R171 VDD.n449 VDD.n448 129.472
R172 VDD.n391 VDD.n390 129.472
R173 VDD.n379 VDD.n378 129.472
R174 VDD.n316 VDD.n315 129.472
R175 VDD.n304 VDD.n303 129.472
R176 VDD.n242 VDD.n241 129.472
R177 VDD.n51 VDD.n50 92.5
R178 VDD.n49 VDD.n48 92.5
R179 VDD.n47 VDD.n46 92.5
R180 VDD.n45 VDD.n44 92.5
R181 VDD.n53 VDD.n52 92.5
R182 VDD.n108 VDD.n107 92.5
R183 VDD.n106 VDD.n105 92.5
R184 VDD.n104 VDD.n103 92.5
R185 VDD.n102 VDD.n101 92.5
R186 VDD.n110 VDD.n109 92.5
R187 VDD.n161 VDD.n160 92.5
R188 VDD.n159 VDD.n158 92.5
R189 VDD.n157 VDD.n156 92.5
R190 VDD.n155 VDD.n154 92.5
R191 VDD.n163 VDD.n162 92.5
R192 VDD.n218 VDD.n217 92.5
R193 VDD.n216 VDD.n215 92.5
R194 VDD.n214 VDD.n213 92.5
R195 VDD.n212 VDD.n211 92.5
R196 VDD.n220 VDD.n219 92.5
R197 VDD.n275 VDD.n274 92.5
R198 VDD.n273 VDD.n272 92.5
R199 VDD.n271 VDD.n270 92.5
R200 VDD.n269 VDD.n268 92.5
R201 VDD.n277 VDD.n276 92.5
R202 VDD.n350 VDD.n349 92.5
R203 VDD.n348 VDD.n347 92.5
R204 VDD.n346 VDD.n345 92.5
R205 VDD.n344 VDD.n343 92.5
R206 VDD.n352 VDD.n351 92.5
R207 VDD.n425 VDD.n424 92.5
R208 VDD.n423 VDD.n422 92.5
R209 VDD.n421 VDD.n420 92.5
R210 VDD.n419 VDD.n418 92.5
R211 VDD.n427 VDD.n426 92.5
R212 VDD.n482 VDD.n481 92.5
R213 VDD.n480 VDD.n479 92.5
R214 VDD.n478 VDD.n477 92.5
R215 VDD.n476 VDD.n475 92.5
R216 VDD.n484 VDD.n483 92.5
R217 VDD.n557 VDD.n556 92.5
R218 VDD.n555 VDD.n554 92.5
R219 VDD.n553 VDD.n552 92.5
R220 VDD.n551 VDD.n550 92.5
R221 VDD.n559 VDD.n558 92.5
R222 VDD.n632 VDD.n631 92.5
R223 VDD.n630 VDD.n629 92.5
R224 VDD.n628 VDD.n627 92.5
R225 VDD.n626 VDD.n625 92.5
R226 VDD.n634 VDD.n633 92.5
R227 VDD.n689 VDD.n688 92.5
R228 VDD.n687 VDD.n686 92.5
R229 VDD.n685 VDD.n684 92.5
R230 VDD.n683 VDD.n682 92.5
R231 VDD.n691 VDD.n690 92.5
R232 VDD.n1445 VDD.n1444 92.5
R233 VDD.n1443 VDD.n1442 92.5
R234 VDD.n1441 VDD.n1440 92.5
R235 VDD.n1439 VDD.n1438 92.5
R236 VDD.n1447 VDD.n1446 92.5
R237 VDD.n1370 VDD.n1369 92.5
R238 VDD.n1368 VDD.n1367 92.5
R239 VDD.n1366 VDD.n1365 92.5
R240 VDD.n1364 VDD.n1363 92.5
R241 VDD.n1372 VDD.n1371 92.5
R242 VDD.n1313 VDD.n1312 92.5
R243 VDD.n1311 VDD.n1310 92.5
R244 VDD.n1309 VDD.n1308 92.5
R245 VDD.n1307 VDD.n1306 92.5
R246 VDD.n1315 VDD.n1314 92.5
R247 VDD.n1238 VDD.n1237 92.5
R248 VDD.n1236 VDD.n1235 92.5
R249 VDD.n1234 VDD.n1233 92.5
R250 VDD.n1232 VDD.n1231 92.5
R251 VDD.n1240 VDD.n1239 92.5
R252 VDD.n1163 VDD.n1162 92.5
R253 VDD.n1161 VDD.n1160 92.5
R254 VDD.n1159 VDD.n1158 92.5
R255 VDD.n1157 VDD.n1156 92.5
R256 VDD.n1165 VDD.n1164 92.5
R257 VDD.n1106 VDD.n1105 92.5
R258 VDD.n1104 VDD.n1103 92.5
R259 VDD.n1102 VDD.n1101 92.5
R260 VDD.n1100 VDD.n1099 92.5
R261 VDD.n1108 VDD.n1107 92.5
R262 VDD.n1031 VDD.n1030 92.5
R263 VDD.n1029 VDD.n1028 92.5
R264 VDD.n1027 VDD.n1026 92.5
R265 VDD.n1025 VDD.n1024 92.5
R266 VDD.n1033 VDD.n1032 92.5
R267 VDD.n956 VDD.n955 92.5
R268 VDD.n954 VDD.n953 92.5
R269 VDD.n952 VDD.n951 92.5
R270 VDD.n950 VDD.n949 92.5
R271 VDD.n958 VDD.n957 92.5
R272 VDD.n899 VDD.n898 92.5
R273 VDD.n897 VDD.n896 92.5
R274 VDD.n895 VDD.n894 92.5
R275 VDD.n893 VDD.n892 92.5
R276 VDD.n901 VDD.n900 92.5
R277 VDD.n820 VDD.n819 92.5
R278 VDD.n818 VDD.n817 92.5
R279 VDD.n816 VDD.n815 92.5
R280 VDD.n814 VDD.n813 92.5
R281 VDD.n822 VDD.n821 92.5
R282 VDD.n750 VDD.n749 92.5
R283 VDD.n748 VDD.n747 92.5
R284 VDD.n746 VDD.n745 92.5
R285 VDD.n744 VDD.n743 92.5
R286 VDD.n752 VDD.n751 92.5
R287 VDD.n14 VDD.n1 92.5
R288 VDD.n5 VDD.n4 92.5
R289 VDD.n7 VDD.n6 92.5
R290 VDD.n9 VDD.n8 92.5
R291 VDD.n11 VDD.n10 92.5
R292 VDD.n13 VDD.n12 92.5
R293 VDD.n21 VDD.n20 92.059
R294 VDD.n65 VDD.n64 92.059
R295 VDD.n118 VDD.n117 92.059
R296 VDD.n171 VDD.n170 92.059
R297 VDD.n228 VDD.n227 92.059
R298 VDD.n285 VDD.n284 92.059
R299 VDD.n360 VDD.n359 92.059
R300 VDD.n435 VDD.n434 92.059
R301 VDD.n492 VDD.n491 92.059
R302 VDD.n567 VDD.n566 92.059
R303 VDD.n642 VDD.n641 92.059
R304 VDD.n699 VDD.n698 92.059
R305 VDD.n1455 VDD.n1454 92.059
R306 VDD.n1380 VDD.n1379 92.059
R307 VDD.n1323 VDD.n1322 92.059
R308 VDD.n1248 VDD.n1247 92.059
R309 VDD.n1173 VDD.n1172 92.059
R310 VDD.n1116 VDD.n1115 92.059
R311 VDD.n1041 VDD.n1040 92.059
R312 VDD.n966 VDD.n965 92.059
R313 VDD.n909 VDD.n908 92.059
R314 VDD.n834 VDD.n833 92.059
R315 VDD.n758 VDD.n757 92.059
R316 VDD.n20 VDD.n16 67.194
R317 VDD.n20 VDD.n17 67.194
R318 VDD.n20 VDD.n18 67.194
R319 VDD.n20 VDD.n19 67.194
R320 VDD.n742 VDD.n741 44.141
R321 VDD.n891 VDD.n890 44.141
R322 VDD.n948 VDD.n947 44.141
R323 VDD.n1023 VDD.n1022 44.141
R324 VDD.n1098 VDD.n1097 44.141
R325 VDD.n1155 VDD.n1154 44.141
R326 VDD.n1230 VDD.n1229 44.141
R327 VDD.n1305 VDD.n1304 44.141
R328 VDD.n1362 VDD.n1361 44.141
R329 VDD.n1437 VDD.n1436 44.141
R330 VDD.n681 VDD.n680 44.141
R331 VDD.n624 VDD.n623 44.141
R332 VDD.n549 VDD.n548 44.141
R333 VDD.n474 VDD.n473 44.141
R334 VDD.n417 VDD.n416 44.141
R335 VDD.n342 VDD.n341 44.141
R336 VDD.n267 VDD.n266 44.141
R337 VDD.n210 VDD.n209 44.141
R338 VDD.n153 VDD.n152 44.141
R339 VDD.n100 VDD.n99 44.141
R340 VDD.n5 VDD.n3 44.141
R341 VDD.n890 VDD.n888 44.107
R342 VDD.n947 VDD.n945 44.107
R343 VDD.n1022 VDD.n1020 44.107
R344 VDD.n1097 VDD.n1095 44.107
R345 VDD.n1154 VDD.n1152 44.107
R346 VDD.n1229 VDD.n1227 44.107
R347 VDD.n1304 VDD.n1302 44.107
R348 VDD.n1361 VDD.n1359 44.107
R349 VDD.n1436 VDD.n1434 44.107
R350 VDD.n680 VDD.n678 44.107
R351 VDD.n623 VDD.n621 44.107
R352 VDD.n548 VDD.n546 44.107
R353 VDD.n473 VDD.n471 44.107
R354 VDD.n416 VDD.n414 44.107
R355 VDD.n341 VDD.n339 44.107
R356 VDD.n266 VDD.n264 44.107
R357 VDD.n209 VDD.n207 44.107
R358 VDD.n152 VDD.n150 44.107
R359 VDD.n99 VDD.n97 44.107
R360 VDD.n741 VDD.n739 44.107
R361 VDD.n3 VDD.n2 44.107
R362 VDD.n25  43.472
R363 VDD.n33 �3� 43.472
R364 VDD.n20 VDD.n15 41.052
R365 VDD.n59 VDD.n57 39.742
R366 VDD.n59 VDD.n58 39.742
R367 VDD.n61 VDD.n60 39.742
R368 VDD.n114 VDD.n113 39.742
R369 VDD.n167 VDD.n166 39.742
R370 VDD.n224 VDD.n223 39.742
R371 VDD.n281 VDD.n280 39.742
R372 VDD.n356 VDD.n355 39.742
R373 VDD.n431 VDD.n430 39.742
R374 VDD.n488 VDD.n487 39.742
R375 VDD.n563 VDD.n562 39.742
R376 VDD.n638 VDD.n637 39.742
R377 VDD.n695 VDD.n694 39.742
R378 VDD.n1451 VDD.n1450 39.742
R379 VDD.n1376 VDD.n1375 39.742
R380 VDD.n1319 VDD.n1318 39.742
R381 VDD.n1244 VDD.n1243 39.742
R382 VDD.n1169 VDD.n1168 39.742
R383 VDD.n1112 VDD.n1111 39.742
R384 VDD.n1037 VDD.n1036 39.742
R385 VDD.n962 VDD.n961 39.742
R386 VDD.n905 VDD.n904 39.742
R387 VDD.n754 VDD.n753 39.742
R388 VDD.n832 VDD.n829 39.742
R389 VDD.n832 VDD.n831 39.742
R390 VDD.n828 VDD.n827 39.742
R391 VDD.n99 VDD.n98 38
R392 VDD.n152 VDD.n151 38
R393 VDD.n209 VDD.n208 38
R394 VDD.n266 VDD.n265 38
R395 VDD.n341 VDD.n340 38
R396 VDD.n416 VDD.n415 38
R397 VDD.n473 VDD.n472 38
R398 VDD.n548 VDD.n547 38
R399 VDD.n623 VDD.n622 38
R400 VDD.n680 VDD.n679 38
R401 VDD.n1436 VDD.n1435 38
R402 VDD.n1361 VDD.n1360 38
R403 VDD.n1304 VDD.n1303 38
R404 VDD.n1229 VDD.n1228 38
R405 VDD.n1154 VDD.n1153 38
R406 VDD.n1097 VDD.n1096 38
R407 VDD.n1022 VDD.n1021 38
R408 VDD.n947 VDD.n946 38
R409 VDD.n890 VDD.n889 38
R410 VDD.n741 VDD.n740 38
R411 VDD.n888 VDD.n887 36.774
R412 VDD.n945 VDD.n944 36.774
R413 VDD.n1020 VDD.n1019 36.774
R414 VDD.n1095 VDD.n1094 36.774
R415 VDD.n1152 VDD.n1151 36.774
R416 VDD.n1227 VDD.n1226 36.774
R417 VDD.n1302 VDD.n1301 36.774
R418 VDD.n1359 VDD.n1358 36.774
R419 VDD.n1434 VDD.n1433 36.774
R420 VDD.n678 VDD.n677 36.774
R421 VDD.n621 VDD.n620 36.774
R422 VDD.n546 VDD.n545 36.774
R423 VDD.n471 VDD.n470 36.774
R424 VDD.n414 VDD.n413 36.774
R425 VDD.n339 VDD.n338 36.774
R426 VDD.n264 VDD.n263 36.774
R427 VDD.n207 VDD.n206 36.774
R428 VDD.n150 VDD.n149 36.774
R429 VDD.n97 VDD.n96 36.774
R430 VDD.n57 VDD.n56 36.774
R431 VDD.n831 VDD.n830 36.774
R432 VDD.n297 �3� 35.8
R433 VDD.n372 VDD.t170 35.8
R434 VDD.n504 VDD.t138 35.8
R435 VDD.n579  35.8
R436 VDD.n711 0�3� 35.8
R437 VDD.n1417 0�3� 35.8
R438 VDD.n1285  35.8
R439 VDD.n1210  35.8
R440 VDD.n1078 0�3� 35.8
R441 VDD.n1003 �3� 35.8
R442 VDD.n871  35.8
R443 VDD.n795  35.8
R444 VDD.n321 0�3� 33.243
R445 VDD.n396  33.243
R446 VDD.n528  33.243
R447 VDD.n603  33.243
R448 VDD.n735 0�3� 33.243
R449 VDD.n1393 0�3� 33.243
R450 VDD.n1261  33.243
R451 VDD.n1186  33.243
R452 VDD.n1054 0�3� 33.243
R453 VDD.n979 0�3� 33.243
R454 VDD.n847 0�3� 33.243
R455 VDD.n771 0�3� 33.243
R456 VDD.n1 VDD.n0 30.923
R457 VDD.n64 VDD.n62 26.38
R458 VDD.n64 VDD.n61 26.38
R459 VDD.n64 VDD.n59 26.38
R460 VDD.n64 VDD.n63 26.38
R461 VDD.n117 VDD.n115 26.38
R462 VDD.n117 VDD.n114 26.38
R463 VDD.n117 VDD.n116 26.38
R464 VDD.n170 VDD.n168 26.38
R465 VDD.n170 VDD.n167 26.38
R466 VDD.n170 VDD.n169 26.38
R467 VDD.n227 VDD.n225 26.38
R468 VDD.n227 VDD.n224 26.38
R469 VDD.n227 VDD.n226 26.38
R470 VDD.n284 VDD.n282 26.38
R471 VDD.n284 VDD.n281 26.38
R472 VDD.n284 VDD.n283 26.38
R473 VDD.n359 VDD.n357 26.38
R474 VDD.n359 VDD.n356 26.38
R475 VDD.n359 VDD.n358 26.38
R476 VDD.n434 VDD.n432 26.38
R477 VDD.n434 VDD.n431 26.38
R478 VDD.n434 VDD.n433 26.38
R479 VDD.n491 VDD.n489 26.38
R480 VDD.n491 VDD.n488 26.38
R481 VDD.n491 VDD.n490 26.38
R482 VDD.n566 VDD.n564 26.38
R483 VDD.n566 VDD.n563 26.38
R484 VDD.n566 VDD.n565 26.38
R485 VDD.n641 VDD.n639 26.38
R486 VDD.n641 VDD.n638 26.38
R487 VDD.n641 VDD.n640 26.38
R488 VDD.n698 VDD.n696 26.38
R489 VDD.n698 VDD.n695 26.38
R490 VDD.n698 VDD.n697 26.38
R491 VDD.n1454 VDD.n1452 26.38
R492 VDD.n1454 VDD.n1451 26.38
R493 VDD.n1454 VDD.n1453 26.38
R494 VDD.n1379 VDD.n1377 26.38
R495 VDD.n1379 VDD.n1376 26.38
R496 VDD.n1379 VDD.n1378 26.38
R497 VDD.n1322 VDD.n1320 26.38
R498 VDD.n1322 VDD.n1319 26.38
R499 VDD.n1322 VDD.n1321 26.38
R500 VDD.n1247 VDD.n1245 26.38
R501 VDD.n1247 VDD.n1244 26.38
R502 VDD.n1247 VDD.n1246 26.38
R503 VDD.n1172 VDD.n1170 26.38
R504 VDD.n1172 VDD.n1169 26.38
R505 VDD.n1172 VDD.n1171 26.38
R506 VDD.n1115 VDD.n1113 26.38
R507 VDD.n1115 VDD.n1112 26.38
R508 VDD.n1115 VDD.n1114 26.38
R509 VDD.n1040 VDD.n1038 26.38
R510 VDD.n1040 VDD.n1037 26.38
R511 VDD.n1040 VDD.n1039 26.38
R512 VDD.n965 VDD.n963 26.38
R513 VDD.n965 VDD.n962 26.38
R514 VDD.n965 VDD.n964 26.38
R515 VDD.n908 VDD.n906 26.38
R516 VDD.n908 VDD.n905 26.38
R517 VDD.n908 VDD.n907 26.38
R518 VDD.n757 VDD.n755 26.38
R519 VDD.n757 VDD.n754 26.38
R520 VDD.n757 VDD.n756 26.38
R521 VDD.n833 VDD.n832 26.38
R522 VDD.n833 VDD.n828 26.38
R523 VDD.n833 VDD.n826 26.38
R524 VDD.n833 VDD.n825 26.38
R525 VDD.n760 VDD.n752 22.915
R526 VDD.n23 VDD.n14 22.915
R527 VDD.n73  20.457
R528 VDD.n137  20.457
R529 VDD.n180 0�3� 20.457
R530 VDD.n237  20.457
R531 VDD.n444 0�3� 20.457
R532 VDD.n651  20.457
R533 VDD.n1345 �3� 20.457
R534 VDD.n1138 VDD.t186 20.457
R535 VDD.n931 0�3� 20.457
R536 VDD.n84 0�3� 17.9
R537 VDD.n126 �3� 17.9
R538 VDD.n193  17.9
R539 VDD.n250 �3� 17.9
R540 VDD.n457 �Ԅ)�U 17.9
R541 VDD.n664 0�3� 17.9
R542 VDD.n1332 0�3� 17.9
R543 VDD.n1125  17.9
R544 VDD.n918 0�3� 17.9
R545 VDD.n301  15.343
R546 VDD.n376  15.343
R547 VDD.n508 0�3� 15.343
R548 VDD.n583 0�3� 15.343
R549 VDD.n715 �3� 15.343
R550 VDD.n1411 ���)�U 15.343
R551 VDD.n1279 �3� 15.343
R552 VDD.n1204 �3� 15.343
R553 VDD.n1072  15.343
R554 VDD.n997  15.343
R555 VDD.n865 0�3� 15.343
R556 VDD.n789 0�3� 15.343
R557 VDD.n752 VDD.n750 14.864
R558 VDD.n750 VDD.n748 14.864
R559 VDD.n748 VDD.n746 14.864
R560 VDD.n746 VDD.n744 14.864
R561 VDD.n744 VDD.n742 14.864
R562 VDD.n901 VDD.n899 14.864
R563 VDD.n899 VDD.n897 14.864
R564 VDD.n897 VDD.n895 14.864
R565 VDD.n895 VDD.n893 14.864
R566 VDD.n893 VDD.n891 14.864
R567 VDD.n958 VDD.n956 14.864
R568 VDD.n956 VDD.n954 14.864
R569 VDD.n954 VDD.n952 14.864
R570 VDD.n952 VDD.n950 14.864
R571 VDD.n950 VDD.n948 14.864
R572 VDD.n1033 VDD.n1031 14.864
R573 VDD.n1031 VDD.n1029 14.864
R574 VDD.n1029 VDD.n1027 14.864
R575 VDD.n1027 VDD.n1025 14.864
R576 VDD.n1025 VDD.n1023 14.864
R577 VDD.n1108 VDD.n1106 14.864
R578 VDD.n1106 VDD.n1104 14.864
R579 VDD.n1104 VDD.n1102 14.864
R580 VDD.n1102 VDD.n1100 14.864
R581 VDD.n1100 VDD.n1098 14.864
R582 VDD.n1165 VDD.n1163 14.864
R583 VDD.n1163 VDD.n1161 14.864
R584 VDD.n1161 VDD.n1159 14.864
R585 VDD.n1159 VDD.n1157 14.864
R586 VDD.n1157 VDD.n1155 14.864
R587 VDD.n1240 VDD.n1238 14.864
R588 VDD.n1238 VDD.n1236 14.864
R589 VDD.n1236 VDD.n1234 14.864
R590 VDD.n1234 VDD.n1232 14.864
R591 VDD.n1232 VDD.n1230 14.864
R592 VDD.n1315 VDD.n1313 14.864
R593 VDD.n1313 VDD.n1311 14.864
R594 VDD.n1311 VDD.n1309 14.864
R595 VDD.n1309 VDD.n1307 14.864
R596 VDD.n1307 VDD.n1305 14.864
R597 VDD.n1372 VDD.n1370 14.864
R598 VDD.n1370 VDD.n1368 14.864
R599 VDD.n1368 VDD.n1366 14.864
R600 VDD.n1366 VDD.n1364 14.864
R601 VDD.n1364 VDD.n1362 14.864
R602 VDD.n1447 VDD.n1445 14.864
R603 VDD.n1445 VDD.n1443 14.864
R604 VDD.n1443 VDD.n1441 14.864
R605 VDD.n1441 VDD.n1439 14.864
R606 VDD.n1439 VDD.n1437 14.864
R607 VDD.n691 VDD.n689 14.864
R608 VDD.n689 VDD.n687 14.864
R609 VDD.n687 VDD.n685 14.864
R610 VDD.n685 VDD.n683 14.864
R611 VDD.n683 VDD.n681 14.864
R612 VDD.n634 VDD.n632 14.864
R613 VDD.n632 VDD.n630 14.864
R614 VDD.n630 VDD.n628 14.864
R615 VDD.n628 VDD.n626 14.864
R616 VDD.n626 VDD.n624 14.864
R617 VDD.n559 VDD.n557 14.864
R618 VDD.n557 VDD.n555 14.864
R619 VDD.n555 VDD.n553 14.864
R620 VDD.n553 VDD.n551 14.864
R621 VDD.n551 VDD.n549 14.864
R622 VDD.n484 VDD.n482 14.864
R623 VDD.n482 VDD.n480 14.864
R624 VDD.n480 VDD.n478 14.864
R625 VDD.n478 VDD.n476 14.864
R626 VDD.n476 VDD.n474 14.864
R627 VDD.n427 VDD.n425 14.864
R628 VDD.n425 VDD.n423 14.864
R629 VDD.n423 VDD.n421 14.864
R630 VDD.n421 VDD.n419 14.864
R631 VDD.n419 VDD.n417 14.864
R632 VDD.n352 VDD.n350 14.864
R633 VDD.n350 VDD.n348 14.864
R634 VDD.n348 VDD.n346 14.864
R635 VDD.n346 VDD.n344 14.864
R636 VDD.n344 VDD.n342 14.864
R637 VDD.n277 VDD.n275 14.864
R638 VDD.n275 VDD.n273 14.864
R639 VDD.n273 VDD.n271 14.864
R640 VDD.n271 VDD.n269 14.864
R641 VDD.n269 VDD.n267 14.864
R642 VDD.n220 VDD.n218 14.864
R643 VDD.n218 VDD.n216 14.864
R644 VDD.n216 VDD.n214 14.864
R645 VDD.n214 VDD.n212 14.864
R646 VDD.n212 VDD.n210 14.864
R647 VDD.n163 VDD.n161 14.864
R648 VDD.n161 VDD.n159 14.864
R649 VDD.n159 VDD.n157 14.864
R650 VDD.n157 VDD.n155 14.864
R651 VDD.n155 VDD.n153 14.864
R652 VDD.n110 VDD.n108 14.864
R653 VDD.n108 VDD.n106 14.864
R654 VDD.n106 VDD.n104 14.864
R655 VDD.n104 VDD.n102 14.864
R656 VDD.n102 VDD.n100 14.864
R657 VDD.n53 VDD.n51 14.864
R658 VDD.n51 VDD.n49 14.864
R659 VDD.n49 VDD.n47 14.864
R660 VDD.n47 VDD.n45 14.864
R661 VDD.n45 VDD.n43 14.864
R662 VDD.n43 VDD.n42 14.864
R663 VDD.n822 VDD.n820 14.864
R664 VDD.n820 VDD.n818 14.864
R665 VDD.n818 VDD.n816 14.864
R666 VDD.n816 VDD.n814 14.864
R667 VDD.n814 VDD.n812 14.864
R668 VDD.n812 VDD.n811 14.864
R669 VDD.n14 VDD.n13 14.864
R670 VDD.n13 VDD.n11 14.864
R671 VDD.n11 VDD.n9 14.864
R672 VDD.n9 VDD.n7 14.864
R673 VDD.n7 VDD.n5 14.864
R674 VDD.n67 VDD.n54 14.864
R675 VDD.n120 VDD.n111 14.864
R676 VDD.n173 VDD.n164 14.864
R677 VDD.n230 VDD.n221 14.864
R678 VDD.n287 VDD.n278 14.864
R679 VDD.n362 VDD.n353 14.864
R680 VDD.n437 VDD.n428 14.864
R681 VDD.n494 VDD.n485 14.864
R682 VDD.n569 VDD.n560 14.864
R683 VDD.n644 VDD.n635 14.864
R684 VDD.n701 VDD.n692 14.864
R685 VDD.n1457 VDD.n1448 14.864
R686 VDD.n1382 VDD.n1373 14.864
R687 VDD.n1325 VDD.n1316 14.864
R688 VDD.n1250 VDD.n1241 14.864
R689 VDD.n1175 VDD.n1166 14.864
R690 VDD.n1118 VDD.n1109 14.864
R691 VDD.n1043 VDD.n1034 14.864
R692 VDD.n968 VDD.n959 14.864
R693 VDD.n911 VDD.n902 14.864
R694 VDD.n836 VDD.n823 14.864
R695 VDD.n775 VDD.t70 14.282
R696 VDD.n775 VDD.t103 14.282
R697 VDD.n791 VDD.t93 14.282
R698 VDD.n791 VDD.t131 14.282
R699 VDD.n851 VDD.t1 14.282
R700 VDD.n851 VDD.t205 14.282
R701 VDD.n867 VDD.t165 14.282
R702 VDD.n867 VDD.t179 14.282
R703 VDD.n926 VDD.t76 14.282
R704 VDD.n926 VDD.t5 14.282
R705 VDD.n983 VDD.t193 14.282
R706 VDD.n983 VDD.t211 14.282
R707 VDD.n999 VDD.t159 14.282
R708 VDD.n999 VDD.t91 14.282
R709 VDD.n1058 VDD.t149 14.282
R710 VDD.n1058 VDD.t109 14.282
R711 VDD.n1074 VDD.t3 14.282
R712 VDD.n1074 VDD.t151 14.282
R713 VDD.n1133 VDD.t203 14.282
R714 VDD.n1133 VDD.t23 14.282
R715 VDD.n1190 VDD.t99 14.282
R716 VDD.n1190 VDD.t19 14.282
R717 VDD.n1206 VDD.t133 14.282
R718 VDD.n1206 VDD.t21 14.282
R719 VDD.n1265 VDD.t7 14.282
R720 VDD.n1265 VDD.t44 14.282
R721 VDD.n1281 VDD.t143 14.282
R722 VDD.n1281 VDD.t87 14.282
R723 VDD.n1340 VDD.t97 14.282
R724 VDD.n1340 VDD.t135 14.282
R725 VDD.n1397 VDD.t52 14.282
R726 VDD.n1397 VDD.t31 14.282
R727 VDD.n1413 VDD.t137 14.282
R728 VDD.n1413 VDD.t40 14.282
R729 VDD.n729 VDD.t147 14.282
R730 VDD.n729 VDD.t42 14.282
R731 VDD.n717 VDD.t197 14.282
R732 VDD.n717 VDD.t163 14.282
R733 VDD.n655 VDD.t29 14.282
R734 VDD.n655 VDD.t195 14.282
R735 VDD.n597 VDD.t74 14.282
R736 VDD.n597 VDD.t113 14.282
R737 VDD.n585 VDD.t199 14.282
R738 VDD.n585 VDD.t101 14.282
R739 VDD.n522 VDD.t173 14.282
R740 VDD.n522 VDD.t129 14.282
R741 VDD.n510 VDD.t161 14.282
R742 VDD.n510 VDD.t181 14.282
R743 VDD.n448 VDD.t115 14.282
R744 VDD.n448 VDD.t15 14.282
R745 VDD.n390 VDD.t183 14.282
R746 VDD.n390 VDD.t64 14.282
R747 VDD.n378 VDD.t157 14.282
R748 VDD.n378 VDD.t79 14.282
R749 VDD.n315 VDD.t167 14.282
R750 VDD.n315 VDD.t50 14.282
R751 VDD.n303 VDD.t175 14.282
R752 VDD.n303 VDD.t145 14.282
R753 VDD.n241 VDD.t117 14.282
R754 VDD.n241 VDD.t72 14.282
R755 VDD.n184 VDD.t17 14.282
R756 VDD.n184 VDD.t62 14.282
R757 VDD.n317 0�3� 12.786
R758 VDD.n392 VDD.t63 12.786
R759 VDD.n524  12.786
R760 VDD.n599 P��(�U 12.786
R761 VDD.n731  12.786
R762 VDD.n1399 0�3� 12.786
R763 VDD.n1267 0�3� 12.786
R764 VDD.n1192  12.786
R765 VDD.n1060 0�3� 12.786
R766 VDD.n985 0�3� 12.786
R767 VDD.n853  12.786
R768 VDD.n777 VDD.t102 12.786
R769 VDD.n187 VDD.n185 9.083
R770 VDD.n244 VDD.n242 9.083
R771 VDD.n451 VDD.n449 9.083
R772 VDD.n658 VDD.n656 9.083
R773 VDD.n1343 VDD.n1341 9.083
R774 VDD.n1136 VDD.n1134 9.083
R775 VDD.n929 VDD.n927 9.083
R776 VDD.n23 VDD.n22 8.855
R777 VDD.n22 VDD.n21 8.855
R778 VDD.n27 VDD.n26 8.855
R779 VDD.n26 VDD.n25 8.855
R780 VDD.n31 VDD.n30 8.855
R781 VDD.n30 VDD.n29 8.855
R782 VDD.n36 VDD.n34 8.855
R783 VDD.n34 VDD.n33 8.855
R784 VDD.n40 VDD.n39 8.855
R785 VDD.n39 VDD.n38 8.855
R786 VDD.n67 VDD.n66 8.855
R787 VDD.n66 VDD.n65 8.855
R788 VDD.n71 VDD.n70 8.855
R789 VDD.n70 VDD.n69 8.855
R790 VDD.n75 VDD.n74 8.855
R791 VDD.n74 VDD.n73 8.855
R792 VDD.n78 VDD.n77 8.855
R793 VDD.n77 0�3� 8.855
R794 VDD.n82 VDD.n81 8.855
R795 VDD.n81 VDD.n80 8.855
R796 VDD.n86 VDD.n85 8.855
R797 VDD.n85 VDD.n84 8.855
R798 VDD.n90 VDD.n89 8.855
R799 VDD.n89 VDD.n88 8.855
R800 VDD.n94 VDD.n93 8.855
R801 VDD.n93 VDD.n92 8.855
R802 VDD.n120 VDD.n119 8.855
R803 VDD.n119 VDD.n118 8.855
R804 VDD.n124 VDD.n123 8.855
R805 VDD.n123 VDD.n122 8.855
R806 VDD.n128 VDD.n127 8.855
R807 VDD.n127 VDD.n126 8.855
R808 VDD.n132 VDD.n131 8.855
R809 VDD.n131 VDD.n130 8.855
R810 VDD.n135 VDD.n134 8.855
R811 VDD.n134 �3� 8.855
R812 VDD.n139 VDD.n138 8.855
R813 VDD.n138 VDD.n137 8.855
R814 VDD.n143 VDD.n142 8.855
R815 VDD.n142 VDD.n141 8.855
R816 VDD.n147 VDD.n146 8.855
R817 VDD.n146 VDD.n145 8.855
R818 VDD.n173 VDD.n172 8.855
R819 VDD.n172 VDD.n171 8.855
R820 VDD.n178 VDD.n177 8.855
R821 VDD.n177 VDD.n176 8.855
R822 VDD.n182 VDD.n181 8.855
R823 VDD.n181 VDD.n180 8.855
R824 VDD.n187 VDD.n186 8.855
R825 VDD.n186 0�3� 8.855
R826 VDD.n191 VDD.n190 8.855
R827 VDD.n190 VDD.n189 8.855
R828 VDD.n195 VDD.n194 8.855
R829 VDD.n194 VDD.n193 8.855
R830 VDD.n200 VDD.n199 8.855
R831 VDD.n199 VDD.n198 8.855
R832 VDD.n204 VDD.n203 8.855
R833 VDD.n203 VDD.n202 8.855
R834 VDD.n230 VDD.n229 8.855
R835 VDD.n229 VDD.n228 8.855
R836 VDD.n235 VDD.n234 8.855
R837 VDD.n234 VDD.n233 8.855
R838 VDD.n239 VDD.n238 8.855
R839 VDD.n238 VDD.n237 8.855
R840 VDD.n244 VDD.n243 8.855
R841 VDD.n243 �3� 8.855
R842 VDD.n248 VDD.n247 8.855
R843 VDD.n247 VDD.n246 8.855
R844 VDD.n252 VDD.n251 8.855
R845 VDD.n251 VDD.n250 8.855
R846 VDD.n257 VDD.n256 8.855
R847 VDD.n256 VDD.n255 8.855
R848 VDD.n261 VDD.n260 8.855
R849 VDD.n260 VDD.n259 8.855
R850 VDD.n287 VDD.n286 8.855
R851 VDD.n286 VDD.n285 8.855
R852 VDD.n291 VDD.n290 8.855
R853 VDD.n290 VDD.n289 8.855
R854 VDD.n295 VDD.n294 8.855
R855 VDD.n294 VDD.n293 8.855
R856 VDD.n299 VDD.n298 8.855
R857 VDD.n298 VDD.n297 8.855
R858 VDD.n305 VDD.n302 8.855
R859 VDD.n302 VDD.n301 8.855
R860 VDD.n309 VDD.n308 8.855
R861 VDD.n308 VDD.n307 8.855
R862 VDD.n313 VDD.n312 8.855
R863 VDD.n312 VDD.n311 8.855
R864 VDD.n319 VDD.n318 8.855
R865 VDD.n318 VDD.n317 8.855
R866 VDD.n323 VDD.n322 8.855
R867 VDD.n322 VDD.n321 8.855
R868 VDD.n328 VDD.n327 8.855
R869 VDD.n327 VDD.n326 8.855
R870 VDD.n332 VDD.n331 8.855
R871 VDD.n331 VDD.n330 8.855
R872 VDD.n336 VDD.n335 8.855
R873 VDD.n335 VDD.n334 8.855
R874 VDD.n362 VDD.n361 8.855
R875 VDD.n361 VDD.n360 8.855
R876 VDD.n366 VDD.n365 8.855
R877 VDD.n365 VDD.n364 8.855
R878 VDD.n370 VDD.n369 8.855
R879 VDD.n369 VDD.n368 8.855
R880 VDD.n374 VDD.n373 8.855
R881 VDD.n373 VDD.n372 8.855
R882 VDD.n380 VDD.n377 8.855
R883 VDD.n377 VDD.n376 8.855
R884 VDD.n384 VDD.n383 8.855
R885 VDD.n383 VDD.n382 8.855
R886 VDD.n388 VDD.n387 8.855
R887 VDD.n387 VDD.n386 8.855
R888 VDD.n394 VDD.n393 8.855
R889 VDD.n393 VDD.n392 8.855
R890 VDD.n398 VDD.n397 8.855
R891 VDD.n397 VDD.n396 8.855
R892 VDD.n403 VDD.n402 8.855
R893 VDD.n402 VDD.n401 8.855
R894 VDD.n407 VDD.n406 8.855
R895 VDD.n406 VDD.n405 8.855
R896 VDD.n411 VDD.n410 8.855
R897 VDD.n410 VDD.n409 8.855
R898 VDD.n437 VDD.n436 8.855
R899 VDD.n436 VDD.n435 8.855
R900 VDD.n442 VDD.n441 8.855
R901 VDD.n441 VDD.n440 8.855
R902 VDD.n446 VDD.n445 8.855
R903 VDD.n445 VDD.n444 8.855
R904 VDD.n451 VDD.n450 8.855
R905 VDD.n450 �3� 8.855
R906 VDD.n455 VDD.n454 8.855
R907 VDD.n454 VDD.n453 8.855
R908 VDD.n459 VDD.n458 8.855
R909 VDD.n458 VDD.n457 8.855
R910 VDD.n464 VDD.n463 8.855
R911 VDD.n463 VDD.n462 8.855
R912 VDD.n468 VDD.n467 8.855
R913 VDD.n467 VDD.n466 8.855
R914 VDD.n494 VDD.n493 8.855
R915 VDD.n493 VDD.n492 8.855
R916 VDD.n498 VDD.n497 8.855
R917 VDD.n497 VDD.n496 8.855
R918 VDD.n502 VDD.n501 8.855
R919 VDD.n501 VDD.n500 8.855
R920 VDD.n506 VDD.n505 8.855
R921 VDD.n505 VDD.n504 8.855
R922 VDD.n512 VDD.n509 8.855
R923 VDD.n509 VDD.n508 8.855
R924 VDD.n516 VDD.n515 8.855
R925 VDD.n515 VDD.n514 8.855
R926 VDD.n520 VDD.n519 8.855
R927 VDD.n519 VDD.n518 8.855
R928 VDD.n526 VDD.n525 8.855
R929 VDD.n525 VDD.n524 8.855
R930 VDD.n530 VDD.n529 8.855
R931 VDD.n529 VDD.n528 8.855
R932 VDD.n535 VDD.n534 8.855
R933 VDD.n534 VDD.n533 8.855
R934 VDD.n539 VDD.n538 8.855
R935 VDD.n538 VDD.n537 8.855
R936 VDD.n543 VDD.n542 8.855
R937 VDD.n542 VDD.n541 8.855
R938 VDD.n569 VDD.n568 8.855
R939 VDD.n568 VDD.n567 8.855
R940 VDD.n573 VDD.n572 8.855
R941 VDD.n572 VDD.n571 8.855
R942 VDD.n577 VDD.n576 8.855
R943 VDD.n576 VDD.n575 8.855
R944 VDD.n581 VDD.n580 8.855
R945 VDD.n580 VDD.n579 8.855
R946 VDD.n587 VDD.n584 8.855
R947 VDD.n584 VDD.n583 8.855
R948 VDD.n591 VDD.n590 8.855
R949 VDD.n590 VDD.n589 8.855
R950 VDD.n595 VDD.n594 8.855
R951 VDD.n594 VDD.n593 8.855
R952 VDD.n601 VDD.n600 8.855
R953 VDD.n600 VDD.n599 8.855
R954 VDD.n605 VDD.n604 8.855
R955 VDD.n604 VDD.n603 8.855
R956 VDD.n610 VDD.n609 8.855
R957 VDD.n609 VDD.n608 8.855
R958 VDD.n614 VDD.n613 8.855
R959 VDD.n613 VDD.n612 8.855
R960 VDD.n618 VDD.n617 8.855
R961 VDD.n617 VDD.n616 8.855
R962 VDD.n644 VDD.n643 8.855
R963 VDD.n643 VDD.n642 8.855
R964 VDD.n649 VDD.n648 8.855
R965 VDD.n648 VDD.n647 8.855
R966 VDD.n653 VDD.n652 8.855
R967 VDD.n652 VDD.n651 8.855
R968 VDD.n658 VDD.n657 8.855
R969 VDD.n657  8.855
R970 VDD.n662 VDD.n661 8.855
R971 VDD.n661 VDD.n660 8.855
R972 VDD.n666 VDD.n665 8.855
R973 VDD.n665 VDD.n664 8.855
R974 VDD.n671 VDD.n670 8.855
R975 VDD.n670 VDD.n669 8.855
R976 VDD.n675 VDD.n674 8.855
R977 VDD.n674 VDD.n673 8.855
R978 VDD.n701 VDD.n700 8.855
R979 VDD.n700 VDD.n699 8.855
R980 VDD.n705 VDD.n704 8.855
R981 VDD.n704 VDD.n703 8.855
R982 VDD.n709 VDD.n708 8.855
R983 VDD.n708 VDD.n707 8.855
R984 VDD.n713 VDD.n712 8.855
R985 VDD.n712 VDD.n711 8.855
R986 VDD.n719 VDD.n716 8.855
R987 VDD.n716 VDD.n715 8.855
R988 VDD.n723 VDD.n722 8.855
R989 VDD.n722 VDD.n721 8.855
R990 VDD.n727 VDD.n726 8.855
R991 VDD.n726 VDD.n725 8.855
R992 VDD.n733 VDD.n732 8.855
R993 VDD.n732 VDD.n731 8.855
R994 VDD.n737 VDD.n736 8.855
R995 VDD.n736 VDD.n735 8.855
R996 VDD.n1466 VDD.n1465 8.855
R997 VDD.n1465 VDD.n1464 8.855
R998 VDD.n1461 VDD.n1460 8.855
R999 VDD.n1460 VDD.n1459 8.855
R1000 VDD.n1457 VDD.n1456 8.855
R1001 VDD.n1456 VDD.n1455 8.855
R1002 VDD.n1431 VDD.n1430 8.855
R1003 VDD.n1430 VDD.n1429 8.855
R1004 VDD.n1427 VDD.n1426 8.855
R1005 VDD.n1426 VDD.n1425 8.855
R1006 VDD.n1423 VDD.n1422 8.855
R1007 VDD.n1422 VDD.n1421 8.855
R1008 VDD.n1419 VDD.n1418 8.855
R1009 VDD.n1418 VDD.n1417 8.855
R1010 VDD.n1415 VDD.n1412 8.855
R1011 VDD.n1412 VDD.n1411 8.855
R1012 VDD.n1409 VDD.n1408 8.855
R1013 VDD.n1408 VDD.n1407 8.855
R1014 VDD.n1405 VDD.n1404 8.855
R1015 VDD.n1404 VDD.n1403 8.855
R1016 VDD.n1401 VDD.n1400 8.855
R1017 VDD.n1400 VDD.n1399 8.855
R1018 VDD.n1395 VDD.n1394 8.855
R1019 VDD.n1394 VDD.n1393 8.855
R1020 VDD.n1391 VDD.n1390 8.855
R1021 VDD.n1390 VDD.n1389 8.855
R1022 VDD.n1386 VDD.n1385 8.855
R1023 VDD.n1385 VDD.n1384 8.855
R1024 VDD.n1382 VDD.n1381 8.855
R1025 VDD.n1381 VDD.n1380 8.855
R1026 VDD.n1356 VDD.n1355 8.855
R1027 VDD.n1355 VDD.n1354 8.855
R1028 VDD.n1352 VDD.n1351 8.855
R1029 VDD.n1351 VDD.n1350 8.855
R1030 VDD.n1347 VDD.n1346 8.855
R1031 VDD.n1346 VDD.n1345 8.855
R1032 VDD.n1343 VDD.n1342 8.855
R1033 VDD.n1342  8.855
R1034 VDD.n1338 VDD.n1337 8.855
R1035 VDD.n1337 VDD.n1336 8.855
R1036 VDD.n1334 VDD.n1333 8.855
R1037 VDD.n1333 VDD.n1332 8.855
R1038 VDD.n1330 VDD.n1329 8.855
R1039 VDD.n1329 VDD.n1328 8.855
R1040 VDD.n1325 VDD.n1324 8.855
R1041 VDD.n1324 VDD.n1323 8.855
R1042 VDD.n1299 VDD.n1298 8.855
R1043 VDD.n1298 VDD.n1297 8.855
R1044 VDD.n1295 VDD.n1294 8.855
R1045 VDD.n1294 VDD.n1293 8.855
R1046 VDD.n1291 VDD.n1290 8.855
R1047 VDD.n1290 VDD.n1289 8.855
R1048 VDD.n1287 VDD.n1286 8.855
R1049 VDD.n1286 VDD.n1285 8.855
R1050 VDD.n1283 VDD.n1280 8.855
R1051 VDD.n1280 VDD.n1279 8.855
R1052 VDD.n1277 VDD.n1276 8.855
R1053 VDD.n1276 VDD.n1275 8.855
R1054 VDD.n1273 VDD.n1272 8.855
R1055 VDD.n1272 VDD.n1271 8.855
R1056 VDD.n1269 VDD.n1268 8.855
R1057 VDD.n1268 VDD.n1267 8.855
R1058 VDD.n1263 VDD.n1262 8.855
R1059 VDD.n1262 VDD.n1261 8.855
R1060 VDD.n1259 VDD.n1258 8.855
R1061 VDD.n1258 VDD.n1257 8.855
R1062 VDD.n1254 VDD.n1253 8.855
R1063 VDD.n1253 VDD.n1252 8.855
R1064 VDD.n1250 VDD.n1249 8.855
R1065 VDD.n1249 VDD.n1248 8.855
R1066 VDD.n1224 VDD.n1223 8.855
R1067 VDD.n1223 VDD.n1222 8.855
R1068 VDD.n1220 VDD.n1219 8.855
R1069 VDD.n1219 VDD.n1218 8.855
R1070 VDD.n1216 VDD.n1215 8.855
R1071 VDD.n1215 VDD.n1214 8.855
R1072 VDD.n1212 VDD.n1211 8.855
R1073 VDD.n1211 VDD.n1210 8.855
R1074 VDD.n1208 VDD.n1205 8.855
R1075 VDD.n1205 VDD.n1204 8.855
R1076 VDD.n1202 VDD.n1201 8.855
R1077 VDD.n1201 VDD.n1200 8.855
R1078 VDD.n1198 VDD.n1197 8.855
R1079 VDD.n1197 VDD.n1196 8.855
R1080 VDD.n1194 VDD.n1193 8.855
R1081 VDD.n1193 VDD.n1192 8.855
R1082 VDD.n1188 VDD.n1187 8.855
R1083 VDD.n1187 VDD.n1186 8.855
R1084 VDD.n1184 VDD.n1183 8.855
R1085 VDD.n1183 VDD.n1182 8.855
R1086 VDD.n1179 VDD.n1178 8.855
R1087 VDD.n1178 VDD.n1177 8.855
R1088 VDD.n1175 VDD.n1174 8.855
R1089 VDD.n1174 VDD.n1173 8.855
R1090 VDD.n1149 VDD.n1148 8.855
R1091 VDD.n1148 VDD.n1147 8.855
R1092 VDD.n1145 VDD.n1144 8.855
R1093 VDD.n1144 VDD.n1143 8.855
R1094 VDD.n1140 VDD.n1139 8.855
R1095 VDD.n1139 VDD.n1138 8.855
R1096 VDD.n1136 VDD.n1135 8.855
R1097 VDD.n1135 0�3� 8.855
R1098 VDD.n1131 VDD.n1130 8.855
R1099 VDD.n1130 VDD.n1129 8.855
R1100 VDD.n1127 VDD.n1126 8.855
R1101 VDD.n1126 VDD.n1125 8.855
R1102 VDD.n1123 VDD.n1122 8.855
R1103 VDD.n1122 VDD.n1121 8.855
R1104 VDD.n1118 VDD.n1117 8.855
R1105 VDD.n1117 VDD.n1116 8.855
R1106 VDD.n1092 VDD.n1091 8.855
R1107 VDD.n1091 VDD.n1090 8.855
R1108 VDD.n1088 VDD.n1087 8.855
R1109 VDD.n1087 VDD.n1086 8.855
R1110 VDD.n1084 VDD.n1083 8.855
R1111 VDD.n1083 VDD.n1082 8.855
R1112 VDD.n1080 VDD.n1079 8.855
R1113 VDD.n1079 VDD.n1078 8.855
R1114 VDD.n1076 VDD.n1073 8.855
R1115 VDD.n1073 VDD.n1072 8.855
R1116 VDD.n1070 VDD.n1069 8.855
R1117 VDD.n1069 VDD.n1068 8.855
R1118 VDD.n1066 VDD.n1065 8.855
R1119 VDD.n1065 VDD.n1064 8.855
R1120 VDD.n1062 VDD.n1061 8.855
R1121 VDD.n1061 VDD.n1060 8.855
R1122 VDD.n1056 VDD.n1055 8.855
R1123 VDD.n1055 VDD.n1054 8.855
R1124 VDD.n1052 VDD.n1051 8.855
R1125 VDD.n1051 VDD.n1050 8.855
R1126 VDD.n1047 VDD.n1046 8.855
R1127 VDD.n1046 VDD.n1045 8.855
R1128 VDD.n1043 VDD.n1042 8.855
R1129 VDD.n1042 VDD.n1041 8.855
R1130 VDD.n1017 VDD.n1016 8.855
R1131 VDD.n1016 VDD.n1015 8.855
R1132 VDD.n1013 VDD.n1012 8.855
R1133 VDD.n1012 VDD.n1011 8.855
R1134 VDD.n1009 VDD.n1008 8.855
R1135 VDD.n1008 VDD.n1007 8.855
R1136 VDD.n1005 VDD.n1004 8.855
R1137 VDD.n1004 VDD.n1003 8.855
R1138 VDD.n1001 VDD.n998 8.855
R1139 VDD.n998 VDD.n997 8.855
R1140 VDD.n995 VDD.n994 8.855
R1141 VDD.n994 VDD.n993 8.855
R1142 VDD.n991 VDD.n990 8.855
R1143 VDD.n990 VDD.n989 8.855
R1144 VDD.n987 VDD.n986 8.855
R1145 VDD.n986 VDD.n985 8.855
R1146 VDD.n981 VDD.n980 8.855
R1147 VDD.n980 VDD.n979 8.855
R1148 VDD.n977 VDD.n976 8.855
R1149 VDD.n976 VDD.n975 8.855
R1150 VDD.n972 VDD.n971 8.855
R1151 VDD.n971 VDD.n970 8.855
R1152 VDD.n968 VDD.n967 8.855
R1153 VDD.n967 VDD.n966 8.855
R1154 VDD.n942 VDD.n941 8.855
R1155 VDD.n941 VDD.n940 8.855
R1156 VDD.n938 VDD.n937 8.855
R1157 VDD.n937 VDD.n936 8.855
R1158 VDD.n933 VDD.n932 8.855
R1159 VDD.n932 VDD.n931 8.855
R1160 VDD.n929 VDD.n928 8.855
R1161 VDD.n928  8.855
R1162 VDD.n924 VDD.n923 8.855
R1163 VDD.n923 VDD.n922 8.855
R1164 VDD.n920 VDD.n919 8.855
R1165 VDD.n919 VDD.n918 8.855
R1166 VDD.n916 VDD.n915 8.855
R1167 VDD.n915 VDD.n914 8.855
R1168 VDD.n911 VDD.n910 8.855
R1169 VDD.n910 VDD.n909 8.855
R1170 VDD.n885 VDD.n884 8.855
R1171 VDD.n884 VDD.n883 8.855
R1172 VDD.n881 VDD.n880 8.855
R1173 VDD.n880 VDD.n879 8.855
R1174 VDD.n877 VDD.n876 8.855
R1175 VDD.n876 VDD.n875 8.855
R1176 VDD.n873 VDD.n872 8.855
R1177 VDD.n872 VDD.n871 8.855
R1178 VDD.n869 VDD.n866 8.855
R1179 VDD.n866 VDD.n865 8.855
R1180 VDD.n863 VDD.n862 8.855
R1181 VDD.n862 VDD.n861 8.855
R1182 VDD.n859 VDD.n858 8.855
R1183 VDD.n858 VDD.n857 8.855
R1184 VDD.n855 VDD.n854 8.855
R1185 VDD.n854 VDD.n853 8.855
R1186 VDD.n849 VDD.n848 8.855
R1187 VDD.n848 VDD.n847 8.855
R1188 VDD.n845 VDD.n844 8.855
R1189 VDD.n844 VDD.n843 8.855
R1190 VDD.n840 VDD.n839 8.855
R1191 VDD.n839 VDD.n838 8.855
R1192 VDD.n836 VDD.n835 8.855
R1193 VDD.n835 VDD.n834 8.855
R1194 VDD.n809 VDD.n808 8.855
R1195 VDD.n808 VDD.n807 8.855
R1196 VDD.n805 VDD.n804 8.855
R1197 VDD.n804 VDD.n803 8.855
R1198 VDD.n801 VDD.n800 8.855
R1199 VDD.n800 VDD.n799 8.855
R1200 VDD.n797 VDD.n796 8.855
R1201 VDD.n796 VDD.n795 8.855
R1202 VDD.n793 VDD.n790 8.855
R1203 VDD.n790 VDD.n789 8.855
R1204 VDD.n787 VDD.n786 8.855
R1205 VDD.n786 VDD.n785 8.855
R1206 VDD.n783 VDD.n782 8.855
R1207 VDD.n782 VDD.n781 8.855
R1208 VDD.n779 VDD.n778 8.855
R1209 VDD.n778 VDD.n777 8.855
R1210 VDD.n773 VDD.n772 8.855
R1211 VDD.n772 VDD.n771 8.855
R1212 VDD.n769 VDD.n768 8.855
R1213 VDD.n768 VDD.n767 8.855
R1214 VDD.n764 VDD.n763 8.855
R1215 VDD.n763 VDD.n762 8.855
R1216 VDD.n760 VDD.n759 8.855
R1217 VDD.n759 VDD.n758 8.855
R1218 VDD.n902 VDD.n901 8.051
R1219 VDD.n959 VDD.n958 8.051
R1220 VDD.n1034 VDD.n1033 8.051
R1221 VDD.n1109 VDD.n1108 8.051
R1222 VDD.n1166 VDD.n1165 8.051
R1223 VDD.n1241 VDD.n1240 8.051
R1224 VDD.n1316 VDD.n1315 8.051
R1225 VDD.n1373 VDD.n1372 8.051
R1226 VDD.n1448 VDD.n1447 8.051
R1227 VDD.n692 VDD.n691 8.051
R1228 VDD.n635 VDD.n634 8.051
R1229 VDD.n560 VDD.n559 8.051
R1230 VDD.n485 VDD.n484 8.051
R1231 VDD.n428 VDD.n427 8.051
R1232 VDD.n353 VDD.n352 8.051
R1233 VDD.n278 VDD.n277 8.051
R1234 VDD.n221 VDD.n220 8.051
R1235 VDD.n164 VDD.n163 8.051
R1236 VDD.n111 VDD.n110 8.051
R1237 VDD.n54 VDD.n53 8.051
R1238 VDD.n823 VDD.n822 8.051
R1239 VDD.n311 0�3� 7.671
R1240 VDD.n386  7.671
R1241 VDD.n518  7.671
R1242 VDD.n593 0�3� 7.671
R1243 VDD.n725  7.671
R1244 VDD.n1403 0�3� 7.671
R1245 VDD.n1271 0�3� 7.671
R1246 VDD.n1196 �3� 7.671
R1247 VDD.n1064  7.671
R1248 VDD.n989 0�3� 7.671
R1249 VDD.n857 0�3� 7.671
R1250 VDD.n781  7.671
R1251 VDD.n319 VDD.n316 7.019
R1252 VDD.n394 VDD.n391 7.019
R1253 VDD.n526 VDD.n523 7.019
R1254 VDD.n601 VDD.n598 7.019
R1255 VDD.n733 VDD.n730 7.019
R1256 VDD.n1401 VDD.n1398 7.019
R1257 VDD.n1269 VDD.n1266 7.019
R1258 VDD.n1194 VDD.n1191 7.019
R1259 VDD.n1062 VDD.n1059 7.019
R1260 VDD.n987 VDD.n984 7.019
R1261 VDD.n855 VDD.n852 7.019
R1262 VDD.n779 VDD.n776 7.019
R1263 VDD.n305 VDD.n304 6.606
R1264 VDD.n380 VDD.n379 6.606
R1265 VDD.n512 VDD.n511 6.606
R1266 VDD.n587 VDD.n586 6.606
R1267 VDD.n719 VDD.n718 6.606
R1268 VDD.n1415 VDD.n1414 6.606
R1269 VDD.n1283 VDD.n1282 6.606
R1270 VDD.n1208 VDD.n1207 6.606
R1271 VDD.n1076 VDD.n1075 6.606
R1272 VDD.n1001 VDD.n1000 6.606
R1273 VDD.n869 VDD.n868 6.606
R1274 VDD.n793 VDD.n792 6.606
R1275 VDD.n307 0�3� 5.114
R1276 VDD.n382 0�3� 5.114
R1277 VDD.n514  5.114
R1278 VDD.n589  5.114
R1279 VDD.n721  5.114
R1280 VDD.n1407 0�3� 5.114
R1281 VDD.n1275 0�3� 5.114
R1282 VDD.n1200  5.114
R1283 VDD.n1068 0�3� 5.114
R1284 VDD.n993 0�3� 5.114
R1285 VDD.n861  5.114
R1286 VDD.n785  5.114
R1287 VDD.n28 VDD.n23 4.795
R1288 VDD.n28 VDD.n27 4.65
R1289 VDD.n32 VDD.n31 4.65
R1290 VDD.n37 VDD.n36 4.65
R1291 VDD.n41 VDD.n40 4.65
R1292 VDD.n68 VDD.n67 4.65
R1293 VDD.n72 VDD.n71 4.65
R1294 VDD.n76 VDD.n75 4.65
R1295 VDD.n79 VDD.n78 4.65
R1296 VDD.n83 VDD.n82 4.65
R1297 VDD.n87 VDD.n86 4.65
R1298 VDD.n91 VDD.n90 4.65
R1299 VDD.n95 VDD.n94 4.65
R1300 VDD.n121 VDD.n120 4.65
R1301 VDD.n125 VDD.n124 4.65
R1302 VDD.n129 VDD.n128 4.65
R1303 VDD.n133 VDD.n132 4.65
R1304 VDD.n136 VDD.n135 4.65
R1305 VDD.n140 VDD.n139 4.65
R1306 VDD.n144 VDD.n143 4.65
R1307 VDD.n148 VDD.n147 4.65
R1308 VDD.n174 VDD.n173 4.65
R1309 VDD.n179 VDD.n178 4.65
R1310 VDD.n183 VDD.n182 4.65
R1311 VDD.n188 VDD.n187 4.65
R1312 VDD.n192 VDD.n191 4.65
R1313 VDD.n196 VDD.n195 4.65
R1314 VDD.n201 VDD.n200 4.65
R1315 VDD.n205 VDD.n204 4.65
R1316 VDD.n231 VDD.n230 4.65
R1317 VDD.n236 VDD.n235 4.65
R1318 VDD.n240 VDD.n239 4.65
R1319 VDD.n245 VDD.n244 4.65
R1320 VDD.n249 VDD.n248 4.65
R1321 VDD.n253 VDD.n252 4.65
R1322 VDD.n258 VDD.n257 4.65
R1323 VDD.n262 VDD.n261 4.65
R1324 VDD.n288 VDD.n287 4.65
R1325 VDD.n292 VDD.n291 4.65
R1326 VDD.n296 VDD.n295 4.65
R1327 VDD.n300 VDD.n299 4.65
R1328 VDD.n306 VDD.n305 4.65
R1329 VDD.n310 VDD.n309 4.65
R1330 VDD.n314 VDD.n313 4.65
R1331 VDD.n320 VDD.n319 4.65
R1332 VDD.n324 VDD.n323 4.65
R1333 VDD.n329 VDD.n328 4.65
R1334 VDD.n333 VDD.n332 4.65
R1335 VDD.n337 VDD.n336 4.65
R1336 VDD.n363 VDD.n362 4.65
R1337 VDD.n367 VDD.n366 4.65
R1338 VDD.n371 VDD.n370 4.65
R1339 VDD.n375 VDD.n374 4.65
R1340 VDD.n381 VDD.n380 4.65
R1341 VDD.n385 VDD.n384 4.65
R1342 VDD.n389 VDD.n388 4.65
R1343 VDD.n395 VDD.n394 4.65
R1344 VDD.n399 VDD.n398 4.65
R1345 VDD.n404 VDD.n403 4.65
R1346 VDD.n408 VDD.n407 4.65
R1347 VDD.n412 VDD.n411 4.65
R1348 VDD.n438 VDD.n437 4.65
R1349 VDD.n443 VDD.n442 4.65
R1350 VDD.n447 VDD.n446 4.65
R1351 VDD.n452 VDD.n451 4.65
R1352 VDD.n456 VDD.n455 4.65
R1353 VDD.n460 VDD.n459 4.65
R1354 VDD.n465 VDD.n464 4.65
R1355 VDD.n469 VDD.n468 4.65
R1356 VDD.n495 VDD.n494 4.65
R1357 VDD.n499 VDD.n498 4.65
R1358 VDD.n503 VDD.n502 4.65
R1359 VDD.n507 VDD.n506 4.65
R1360 VDD.n513 VDD.n512 4.65
R1361 VDD.n517 VDD.n516 4.65
R1362 VDD.n521 VDD.n520 4.65
R1363 VDD.n527 VDD.n526 4.65
R1364 VDD.n531 VDD.n530 4.65
R1365 VDD.n536 VDD.n535 4.65
R1366 VDD.n540 VDD.n539 4.65
R1367 VDD.n544 VDD.n543 4.65
R1368 VDD.n570 VDD.n569 4.65
R1369 VDD.n574 VDD.n573 4.65
R1370 VDD.n578 VDD.n577 4.65
R1371 VDD.n582 VDD.n581 4.65
R1372 VDD.n588 VDD.n587 4.65
R1373 VDD.n592 VDD.n591 4.65
R1374 VDD.n596 VDD.n595 4.65
R1375 VDD.n602 VDD.n601 4.65
R1376 VDD.n606 VDD.n605 4.65
R1377 VDD.n611 VDD.n610 4.65
R1378 VDD.n615 VDD.n614 4.65
R1379 VDD.n619 VDD.n618 4.65
R1380 VDD.n645 VDD.n644 4.65
R1381 VDD.n650 VDD.n649 4.65
R1382 VDD.n654 VDD.n653 4.65
R1383 VDD.n659 VDD.n658 4.65
R1384 VDD.n663 VDD.n662 4.65
R1385 VDD.n667 VDD.n666 4.65
R1386 VDD.n672 VDD.n671 4.65
R1387 VDD.n676 VDD.n675 4.65
R1388 VDD.n702 VDD.n701 4.65
R1389 VDD.n706 VDD.n705 4.65
R1390 VDD.n710 VDD.n709 4.65
R1391 VDD.n714 VDD.n713 4.65
R1392 VDD.n720 VDD.n719 4.65
R1393 VDD.n724 VDD.n723 4.65
R1394 VDD.n728 VDD.n727 4.65
R1395 VDD.n734 VDD.n733 4.65
R1396 VDD.n738 VDD.n737 4.65
R1397 VDD.n1467 VDD.n1466 4.65
R1398 VDD.n1462 VDD.n1461 4.65
R1399 VDD.n1458 VDD.n1457 4.65
R1400 VDD.n1432 VDD.n1431 4.65
R1401 VDD.n1428 VDD.n1427 4.65
R1402 VDD.n1424 VDD.n1423 4.65
R1403 VDD.n1420 VDD.n1419 4.65
R1404 VDD.n1416 VDD.n1415 4.65
R1405 VDD.n1410 VDD.n1409 4.65
R1406 VDD.n1406 VDD.n1405 4.65
R1407 VDD.n1402 VDD.n1401 4.65
R1408 VDD.n1396 VDD.n1395 4.65
R1409 VDD.n1392 VDD.n1391 4.65
R1410 VDD.n1387 VDD.n1386 4.65
R1411 VDD.n1383 VDD.n1382 4.65
R1412 VDD.n1357 VDD.n1356 4.65
R1413 VDD.n1353 VDD.n1352 4.65
R1414 VDD.n1348 VDD.n1347 4.65
R1415 VDD.n1344 VDD.n1343 4.65
R1416 VDD.n1339 VDD.n1338 4.65
R1417 VDD.n1335 VDD.n1334 4.65
R1418 VDD.n1331 VDD.n1330 4.65
R1419 VDD.n1326 VDD.n1325 4.65
R1420 VDD.n1300 VDD.n1299 4.65
R1421 VDD.n1296 VDD.n1295 4.65
R1422 VDD.n1292 VDD.n1291 4.65
R1423 VDD.n1288 VDD.n1287 4.65
R1424 VDD.n1284 VDD.n1283 4.65
R1425 VDD.n1278 VDD.n1277 4.65
R1426 VDD.n1274 VDD.n1273 4.65
R1427 VDD.n1270 VDD.n1269 4.65
R1428 VDD.n1264 VDD.n1263 4.65
R1429 VDD.n1260 VDD.n1259 4.65
R1430 VDD.n1255 VDD.n1254 4.65
R1431 VDD.n1251 VDD.n1250 4.65
R1432 VDD.n1225 VDD.n1224 4.65
R1433 VDD.n1221 VDD.n1220 4.65
R1434 VDD.n1217 VDD.n1216 4.65
R1435 VDD.n1213 VDD.n1212 4.65
R1436 VDD.n1209 VDD.n1208 4.65
R1437 VDD.n1203 VDD.n1202 4.65
R1438 VDD.n1199 VDD.n1198 4.65
R1439 VDD.n1195 VDD.n1194 4.65
R1440 VDD.n1189 VDD.n1188 4.65
R1441 VDD.n1185 VDD.n1184 4.65
R1442 VDD.n1180 VDD.n1179 4.65
R1443 VDD.n1176 VDD.n1175 4.65
R1444 VDD.n1150 VDD.n1149 4.65
R1445 VDD.n1146 VDD.n1145 4.65
R1446 VDD.n1141 VDD.n1140 4.65
R1447 VDD.n1137 VDD.n1136 4.65
R1448 VDD.n1132 VDD.n1131 4.65
R1449 VDD.n1128 VDD.n1127 4.65
R1450 VDD.n1124 VDD.n1123 4.65
R1451 VDD.n1119 VDD.n1118 4.65
R1452 VDD.n1093 VDD.n1092 4.65
R1453 VDD.n1089 VDD.n1088 4.65
R1454 VDD.n1085 VDD.n1084 4.65
R1455 VDD.n1081 VDD.n1080 4.65
R1456 VDD.n1077 VDD.n1076 4.65
R1457 VDD.n1071 VDD.n1070 4.65
R1458 VDD.n1067 VDD.n1066 4.65
R1459 VDD.n1063 VDD.n1062 4.65
R1460 VDD.n1057 VDD.n1056 4.65
R1461 VDD.n1053 VDD.n1052 4.65
R1462 VDD.n1048 VDD.n1047 4.65
R1463 VDD.n1044 VDD.n1043 4.65
R1464 VDD.n1018 VDD.n1017 4.65
R1465 VDD.n1014 VDD.n1013 4.65
R1466 VDD.n1010 VDD.n1009 4.65
R1467 VDD.n1006 VDD.n1005 4.65
R1468 VDD.n1002 VDD.n1001 4.65
R1469 VDD.n996 VDD.n995 4.65
R1470 VDD.n992 VDD.n991 4.65
R1471 VDD.n988 VDD.n987 4.65
R1472 VDD.n982 VDD.n981 4.65
R1473 VDD.n978 VDD.n977 4.65
R1474 VDD.n973 VDD.n972 4.65
R1475 VDD.n969 VDD.n968 4.65
R1476 VDD.n943 VDD.n942 4.65
R1477 VDD.n939 VDD.n938 4.65
R1478 VDD.n934 VDD.n933 4.65
R1479 VDD.n930 VDD.n929 4.65
R1480 VDD.n925 VDD.n924 4.65
R1481 VDD.n921 VDD.n920 4.65
R1482 VDD.n917 VDD.n916 4.65
R1483 VDD.n912 VDD.n911 4.65
R1484 VDD.n886 VDD.n885 4.65
R1485 VDD.n882 VDD.n881 4.65
R1486 VDD.n878 VDD.n877 4.65
R1487 VDD.n874 VDD.n873 4.65
R1488 VDD.n870 VDD.n869 4.65
R1489 VDD.n864 VDD.n863 4.65
R1490 VDD.n860 VDD.n859 4.65
R1491 VDD.n856 VDD.n855 4.65
R1492 VDD.n850 VDD.n849 4.65
R1493 VDD.n846 VDD.n845 4.65
R1494 VDD.n841 VDD.n840 4.65
R1495 VDD.n837 VDD.n836 4.65
R1496 VDD.n810 VDD.n809 4.65
R1497 VDD.n806 VDD.n805 4.65
R1498 VDD.n802 VDD.n801 4.65
R1499 VDD.n798 VDD.n797 4.65
R1500 VDD.n794 VDD.n793 4.65
R1501 VDD.n788 VDD.n787 4.65
R1502 VDD.n784 VDD.n783 4.65
R1503 VDD.n780 VDD.n779 4.65
R1504 VDD.n774 VDD.n773 4.65
R1505 VDD.n770 VDD.n769 4.65
R1506 VDD.n765 VDD.n764 4.65
R1507 VDD.n761 VDD.n760 4.65
R1508 VDD.n200 VDD.n197 2.89
R1509 VDD.n257 VDD.n254 2.89
R1510 VDD.n464 VDD.n461 2.89
R1511 VDD.n671 VDD.n668 2.89
R1512 VDD.n1330 VDD.n1327 2.89
R1513 VDD.n1123 VDD.n1120 2.89
R1514 VDD.n916 VDD.n913 2.89
R1515 VDD.n80 VDD.t106 2.557
R1516 VDD.n130  2.557
R1517 VDD.n189 VDD.t61 2.557
R1518 VDD.n246 0�3� 2.557
R1519 VDD.n453  2.557
R1520 VDD.n660 0�3� 2.557
R1521 VDD.n1336  2.557
R1522 VDD.n1129 VDD.t22 2.557
R1523 VDD.n922  2.557
R1524 VDD.n178 VDD.n175 2.477
R1525 VDD.n235 VDD.n232 2.477
R1526 VDD.n442 VDD.n439 2.477
R1527 VDD.n649 VDD.n646 2.477
R1528 VDD.n1352 VDD.n1349 2.477
R1529 VDD.n1145 VDD.n1142 2.477
R1530 VDD.n938 VDD.n935 2.477
R1531 VDD.n27 VDD.n24 2.064
R1532 VDD.n36 VDD.n35 2.064
R1533 VDD.n328 VDD.n325 0.412
R1534 VDD.n403 VDD.n400 0.412
R1535 VDD.n535 VDD.n532 0.412
R1536 VDD.n610 VDD.n607 0.412
R1537 VDD.n1466 VDD.n1463 0.412
R1538 VDD.n1391 VDD.n1388 0.412
R1539 VDD.n1259 VDD.n1256 0.412
R1540 VDD.n1184 VDD.n1181 0.412
R1541 VDD.n1052 VDD.n1049 0.412
R1542 VDD.n977 VDD.n974 0.412
R1543 VDD.n845 VDD.n842 0.412
R1544 VDD.n769 VDD.n766 0.412
R1545 VDD.n68 VDD.n41 0.29
R1546 VDD.n121 VDD.n95 0.29
R1547 VDD.n174 VDD.n148 0.29
R1548 VDD.n231 VDD.n205 0.29
R1549 VDD.n288 VDD.n262 0.29
R1550 VDD.n363 VDD.n337 0.29
R1551 VDD.n438 VDD.n412 0.29
R1552 VDD.n495 VDD.n469 0.29
R1553 VDD.n570 VDD.n544 0.29
R1554 VDD.n645 VDD.n619 0.29
R1555 VDD.n702 VDD.n676 0.29
R1556 VDD.n1458 VDD.n1432 0.29
R1557 VDD.n1383 VDD.n1357 0.29
R1558 VDD.n1326 VDD.n1300 0.29
R1559 VDD.n1251 VDD.n1225 0.29
R1560 VDD.n1176 VDD.n1150 0.29
R1561 VDD.n1119 VDD.n1093 0.29
R1562 VDD.n1044 VDD.n1018 0.29
R1563 VDD.n969 VDD.n943 0.29
R1564 VDD.n912 VDD.n886 0.29
R1565 VDD.n837 VDD.n810 0.29
R1566 VDD.n761 VDD 0.207
R1567 VDD.n314 VDD.n310 0.197
R1568 VDD.n389 VDD.n385 0.197
R1569 VDD.n521 VDD.n517 0.197
R1570 VDD.n596 VDD.n592 0.197
R1571 VDD.n728 VDD.n724 0.197
R1572 VDD.n1410 VDD.n1406 0.197
R1573 VDD.n1278 VDD.n1274 0.197
R1574 VDD.n1203 VDD.n1199 0.197
R1575 VDD.n1071 VDD.n1067 0.197
R1576 VDD.n996 VDD.n992 0.197
R1577 VDD.n864 VDD.n860 0.197
R1578 VDD.n788 VDD.n784 0.197
R1579 VDD.n83 VDD.n79 0.181
R1580 VDD.n136 VDD.n133 0.181
R1581 VDD.n192 VDD.n188 0.181
R1582 VDD.n249 VDD.n245 0.181
R1583 VDD.n456 VDD.n452 0.181
R1584 VDD.n663 VDD.n659 0.181
R1585 VDD.n1344 VDD.n1339 0.181
R1586 VDD.n1137 VDD.n1132 0.181
R1587 VDD.n930 VDD.n925 0.181
R1588 VDD.n32 VDD.n28 0.157
R1589 VDD.n37 VDD.n32 0.157
R1590 VDD.n41 VDD.n37 0.145
R1591 VDD.n72 VDD.n68 0.145
R1592 VDD.n76 VDD.n72 0.145
R1593 VDD.n79 VDD.n76 0.145
R1594 VDD.n87 VDD.n83 0.145
R1595 VDD.n91 VDD.n87 0.145
R1596 VDD.n95 VDD.n91 0.145
R1597 VDD.n125 VDD.n121 0.145
R1598 VDD.n129 VDD.n125 0.145
R1599 VDD.n133 VDD.n129 0.145
R1600 VDD.n140 VDD.n136 0.145
R1601 VDD.n144 VDD.n140 0.145
R1602 VDD.n148 VDD.n144 0.145
R1603 VDD.n179 VDD.n174 0.145
R1604 VDD.n183 VDD.n179 0.145
R1605 VDD.n188 VDD.n183 0.145
R1606 VDD.n196 VDD.n192 0.145
R1607 VDD.n201 VDD.n196 0.145
R1608 VDD.n205 VDD.n201 0.145
R1609 VDD.n236 VDD.n231 0.145
R1610 VDD.n240 VDD.n236 0.145
R1611 VDD.n245 VDD.n240 0.145
R1612 VDD.n253 VDD.n249 0.145
R1613 VDD.n258 VDD.n253 0.145
R1614 VDD.n262 VDD.n258 0.145
R1615 VDD.n292 VDD.n288 0.145
R1616 VDD.n296 VDD.n292 0.145
R1617 VDD.n300 VDD.n296 0.145
R1618 VDD.n306 VDD.n300 0.145
R1619 VDD.n310 VDD.n306 0.145
R1620 VDD.n320 VDD.n314 0.145
R1621 VDD.n324 VDD.n320 0.145
R1622 VDD.n329 VDD.n324 0.145
R1623 VDD.n333 VDD.n329 0.145
R1624 VDD.n337 VDD.n333 0.145
R1625 VDD.n367 VDD.n363 0.145
R1626 VDD.n371 VDD.n367 0.145
R1627 VDD.n375 VDD.n371 0.145
R1628 VDD.n381 VDD.n375 0.145
R1629 VDD.n385 VDD.n381 0.145
R1630 VDD.n395 VDD.n389 0.145
R1631 VDD.n399 VDD.n395 0.145
R1632 VDD.n404 VDD.n399 0.145
R1633 VDD.n408 VDD.n404 0.145
R1634 VDD.n412 VDD.n408 0.145
R1635 VDD.n443 VDD.n438 0.145
R1636 VDD.n447 VDD.n443 0.145
R1637 VDD.n452 VDD.n447 0.145
R1638 VDD.n460 VDD.n456 0.145
R1639 VDD.n465 VDD.n460 0.145
R1640 VDD.n469 VDD.n465 0.145
R1641 VDD.n499 VDD.n495 0.145
R1642 VDD.n503 VDD.n499 0.145
R1643 VDD.n507 VDD.n503 0.145
R1644 VDD.n513 VDD.n507 0.145
R1645 VDD.n517 VDD.n513 0.145
R1646 VDD.n527 VDD.n521 0.145
R1647 VDD.n531 VDD.n527 0.145
R1648 VDD.n536 VDD.n531 0.145
R1649 VDD.n540 VDD.n536 0.145
R1650 VDD.n544 VDD.n540 0.145
R1651 VDD.n574 VDD.n570 0.145
R1652 VDD.n578 VDD.n574 0.145
R1653 VDD.n582 VDD.n578 0.145
R1654 VDD.n588 VDD.n582 0.145
R1655 VDD.n592 VDD.n588 0.145
R1656 VDD.n602 VDD.n596 0.145
R1657 VDD.n606 VDD.n602 0.145
R1658 VDD.n611 VDD.n606 0.145
R1659 VDD.n615 VDD.n611 0.145
R1660 VDD.n619 VDD.n615 0.145
R1661 VDD.n650 VDD.n645 0.145
R1662 VDD.n654 VDD.n650 0.145
R1663 VDD.n659 VDD.n654 0.145
R1664 VDD.n667 VDD.n663 0.145
R1665 VDD.n672 VDD.n667 0.145
R1666 VDD.n676 VDD.n672 0.145
R1667 VDD.n706 VDD.n702 0.145
R1668 VDD.n710 VDD.n706 0.145
R1669 VDD.n714 VDD.n710 0.145
R1670 VDD.n720 VDD.n714 0.145
R1671 VDD.n724 VDD.n720 0.145
R1672 VDD.n734 VDD.n728 0.145
R1673 VDD.n738 VDD.n734 0.145
R1674 VDD.n1467 VDD.n1462 0.145
R1675 VDD.n1462 VDD.n1458 0.145
R1676 VDD.n1432 VDD.n1428 0.145
R1677 VDD.n1428 VDD.n1424 0.145
R1678 VDD.n1424 VDD.n1420 0.145
R1679 VDD.n1420 VDD.n1416 0.145
R1680 VDD.n1416 VDD.n1410 0.145
R1681 VDD.n1406 VDD.n1402 0.145
R1682 VDD.n1402 VDD.n1396 0.145
R1683 VDD.n1396 VDD.n1392 0.145
R1684 VDD.n1392 VDD.n1387 0.145
R1685 VDD.n1387 VDD.n1383 0.145
R1686 VDD.n1357 VDD.n1353 0.145
R1687 VDD.n1353 VDD.n1348 0.145
R1688 VDD.n1348 VDD.n1344 0.145
R1689 VDD.n1339 VDD.n1335 0.145
R1690 VDD.n1335 VDD.n1331 0.145
R1691 VDD.n1331 VDD.n1326 0.145
R1692 VDD.n1300 VDD.n1296 0.145
R1693 VDD.n1296 VDD.n1292 0.145
R1694 VDD.n1292 VDD.n1288 0.145
R1695 VDD.n1288 VDD.n1284 0.145
R1696 VDD.n1284 VDD.n1278 0.145
R1697 VDD.n1274 VDD.n1270 0.145
R1698 VDD.n1270 VDD.n1264 0.145
R1699 VDD.n1264 VDD.n1260 0.145
R1700 VDD.n1260 VDD.n1255 0.145
R1701 VDD.n1255 VDD.n1251 0.145
R1702 VDD.n1225 VDD.n1221 0.145
R1703 VDD.n1221 VDD.n1217 0.145
R1704 VDD.n1217 VDD.n1213 0.145
R1705 VDD.n1213 VDD.n1209 0.145
R1706 VDD.n1209 VDD.n1203 0.145
R1707 VDD.n1199 VDD.n1195 0.145
R1708 VDD.n1195 VDD.n1189 0.145
R1709 VDD.n1189 VDD.n1185 0.145
R1710 VDD.n1185 VDD.n1180 0.145
R1711 VDD.n1180 VDD.n1176 0.145
R1712 VDD.n1150 VDD.n1146 0.145
R1713 VDD.n1146 VDD.n1141 0.145
R1714 VDD.n1141 VDD.n1137 0.145
R1715 VDD.n1132 VDD.n1128 0.145
R1716 VDD.n1128 VDD.n1124 0.145
R1717 VDD.n1124 VDD.n1119 0.145
R1718 VDD.n1093 VDD.n1089 0.145
R1719 VDD.n1089 VDD.n1085 0.145
R1720 VDD.n1085 VDD.n1081 0.145
R1721 VDD.n1081 VDD.n1077 0.145
R1722 VDD.n1077 VDD.n1071 0.145
R1723 VDD.n1067 VDD.n1063 0.145
R1724 VDD.n1063 VDD.n1057 0.145
R1725 VDD.n1057 VDD.n1053 0.145
R1726 VDD.n1053 VDD.n1048 0.145
R1727 VDD.n1048 VDD.n1044 0.145
R1728 VDD.n1018 VDD.n1014 0.145
R1729 VDD.n1014 VDD.n1010 0.145
R1730 VDD.n1010 VDD.n1006 0.145
R1731 VDD.n1006 VDD.n1002 0.145
R1732 VDD.n1002 VDD.n996 0.145
R1733 VDD.n992 VDD.n988 0.145
R1734 VDD.n988 VDD.n982 0.145
R1735 VDD.n982 VDD.n978 0.145
R1736 VDD.n978 VDD.n973 0.145
R1737 VDD.n973 VDD.n969 0.145
R1738 VDD.n943 VDD.n939 0.145
R1739 VDD.n939 VDD.n934 0.145
R1740 VDD.n934 VDD.n930 0.145
R1741 VDD.n925 VDD.n921 0.145
R1742 VDD.n921 VDD.n917 0.145
R1743 VDD.n917 VDD.n912 0.145
R1744 VDD.n886 VDD.n882 0.145
R1745 VDD.n882 VDD.n878 0.145
R1746 VDD.n878 VDD.n874 0.145
R1747 VDD.n874 VDD.n870 0.145
R1748 VDD.n870 VDD.n864 0.145
R1749 VDD.n860 VDD.n856 0.145
R1750 VDD.n856 VDD.n850 0.145
R1751 VDD.n850 VDD.n846 0.145
R1752 VDD.n846 VDD.n841 0.145
R1753 VDD.n841 VDD.n837 0.145
R1754 VDD.n810 VDD.n806 0.145
R1755 VDD.n806 VDD.n802 0.145
R1756 VDD.n802 VDD.n798 0.145
R1757 VDD.n798 VDD.n794 0.145
R1758 VDD.n794 VDD.n788 0.145
R1759 VDD.n784 VDD.n780 0.145
R1760 VDD.n780 VDD.n774 0.145
R1761 VDD.n774 VDD.n770 0.145
R1762 VDD.n770 VDD.n765 0.145
R1763 VDD.n765 VDD.n761 0.145
R1764 VDD VDD.n1467 0.086
R1765 VDD VDD.n738 0.058
R1766 a_10637_1050.n4 a_10637_1050.t11 512.525
R1767 a_10637_1050.n2 a_10637_1050.t10 512.525
R1768 a_10637_1050.n5 a_10637_1050.t9 389.251
R1769 a_10637_1050.n3 a_10637_1050.t12 389.251
R1770 a_10637_1050.n4 a_10637_1050.t8 371.139
R1771 a_10637_1050.n2 a_10637_1050.t7 371.139
R1772 a_10637_1050.n8 a_10637_1050.n7 357.814
R1773 a_10637_1050.n5 a_10637_1050.n4 207.695
R1774 a_10637_1050.n3 a_10637_1050.n2 207.695
R1775 a_10637_1050.n11 a_10637_1050.n10 161.352
R1776 a_10637_1050.n9 a_10637_1050.n8 151.34
R1777 a_10637_1050.n9 a_10637_1050.n1 95.095
R1778 a_10637_1050.n10 a_10637_1050.n0 95.095
R1779 a_10637_1050.n10 a_10637_1050.n9 66.258
R1780 a_10637_1050.n1 a_10637_1050.t0 14.282
R1781 a_10637_1050.n1 a_10637_1050.t6 14.282
R1782 a_10637_1050.n0 a_10637_1050.t3 14.282
R1783 a_10637_1050.n0 a_10637_1050.t2 14.282
R1784 a_10637_1050.n11 a_10637_1050.t4 14.282
R1785 a_10637_1050.t5 a_10637_1050.n11 14.282
R1786 a_10637_1050.n6 a_10637_1050.n3 14.126
R1787 a_10637_1050.n8 a_10637_1050.n6 5.965
R1788 a_10637_1050.n6 a_10637_1050.n5 4.65
R1789 a_14189_1050.n2 a_14189_1050.t7 480.392
R1790 a_14189_1050.n2 a_14189_1050.t9 403.272
R1791 a_14189_1050.n3 a_14189_1050.t8 385.063
R1792 a_14189_1050.n5 a_14189_1050.n4 357.814
R1793 a_14189_1050.n8 a_14189_1050.n7 161.352
R1794 a_14189_1050.n6 a_14189_1050.n5 151.34
R1795 a_14189_1050.n3 a_14189_1050.n2 143.429
R1796 a_14189_1050.n6 a_14189_1050.n1 95.095
R1797 a_14189_1050.n7 a_14189_1050.n0 95.095
R1798 a_14189_1050.n7 a_14189_1050.n6 66.258
R1799 a_14189_1050.n1 a_14189_1050.t6 14.282
R1800 a_14189_1050.n1 a_14189_1050.t5 14.282
R1801 a_14189_1050.n0 a_14189_1050.t3 14.282
R1802 a_14189_1050.n0 a_14189_1050.t4 14.282
R1803 a_14189_1050.n8 a_14189_1050.t1 14.282
R1804 a_14189_1050.t2 a_14189_1050.n8 14.282
R1805 a_14189_1050.n5 a_14189_1050.n3 10.615
R1806 a_10959_989.n2 a_10959_989.t8 480.392
R1807 a_10959_989.n4 a_10959_989.t10 454.685
R1808 a_10959_989.n4 a_10959_989.t9 428.979
R1809 a_10959_989.n2 a_10959_989.t12 403.272
R1810 a_10959_989.n3 a_10959_989.t7 357.204
R1811 a_10959_989.n5 a_10959_989.t11 311.683
R1812 a_10959_989.n11 a_10959_989.n10 308.216
R1813 a_10959_989.n12 a_10959_989.n11 179.199
R1814 a_10959_989.n5 a_10959_989.n4 171.288
R1815 a_10959_989.n3 a_10959_989.n2 171.288
R1816 a_10959_989.n14 a_10959_989.n13 161.352
R1817 a_10959_989.n12 a_10959_989.n1 95.095
R1818 a_10959_989.n13 a_10959_989.n0 95.095
R1819 a_10959_989.n13 a_10959_989.n12 66.258
R1820 a_10959_989.n10 a_10959_989.n9 30
R1821 a_10959_989.n8 a_10959_989.n7 24.383
R1822 a_10959_989.n10 a_10959_989.n8 23.684
R1823 a_10959_989.n1 a_10959_989.t3 14.282
R1824 a_10959_989.n1 a_10959_989.t4 14.282
R1825 a_10959_989.n0 a_10959_989.t6 14.282
R1826 a_10959_989.n0 a_10959_989.t5 14.282
R1827 a_10959_989.n14 a_10959_989.t0 14.282
R1828 a_10959_989.t1 a_10959_989.n14 14.282
R1829 a_10959_989.n6 a_10959_989.n5 8.685
R1830 a_10959_989.n6 a_10959_989.n3 5.965
R1831 a_10959_989.n11 a_10959_989.n6 4.65
R1832 D.n5 D.t6 479.223
R1833 D.n2 D.t4 479.223
R1834 D.n0 D.t8 479.223
R1835 D.n5 D.t0 375.52
R1836 D.n2 D.t7 375.52
R1837 D.n0 D.t2 375.52
R1838 D.n6 D.n5 280.047
R1839 D.n3 D.n2 280.047
R1840 D.n1 D.n0 280.047
R1841 D.n6 D.t1 136.76
R1842 D.n3 D.t5 136.76
R1843 D.n1 D.t3 136.76
R1844 D.n4 D.n1 23.649
R1845 D.n7 D.n4 18.999
R1846 D.n4 D.n3 4.65
R1847 D.n7 D.n6 4.65
R1848 D.n7 D 0.046
R1849 a_599_989.n1 a_599_989.t7 480.392
R1850 a_599_989.n3 a_599_989.t11 454.685
R1851 a_599_989.n3 a_599_989.t8 428.979
R1852 a_599_989.n1 a_599_989.t10 403.272
R1853 a_599_989.n2 a_599_989.t12 357.204
R1854 a_599_989.n4 a_599_989.t9 311.683
R1855 a_599_989.n10 a_599_989.n9 308.216
R1856 a_599_989.n11 a_599_989.n10 179.199
R1857 a_599_989.n4 a_599_989.n3 171.288
R1858 a_599_989.n2 a_599_989.n1 171.288
R1859 a_599_989.n13 a_599_989.n12 161.352
R1860 a_599_989.n11 a_599_989.n0 95.095
R1861 a_599_989.n14 a_599_989.n13 95.094
R1862 a_599_989.n13 a_599_989.n11 66.258
R1863 a_599_989.n9 a_599_989.n8 30
R1864 a_599_989.n7 a_599_989.n6 24.383
R1865 a_599_989.n9 a_599_989.n7 23.684
R1866 a_599_989.n0 a_599_989.t4 14.282
R1867 a_599_989.n0 a_599_989.t5 14.282
R1868 a_599_989.n12 a_599_989.t6 14.282
R1869 a_599_989.n12 a_599_989.t0 14.282
R1870 a_599_989.n14 a_599_989.t1 14.282
R1871 a_599_989.t2 a_599_989.n14 14.282
R1872 a_599_989.n5 a_599_989.n4 8.685
R1873 a_599_989.n5 a_599_989.n2 5.965
R1874 a_599_989.n10 a_599_989.n5 4.65
R1875 a_11413_103.t0 a_11413_103.n0 117.777
R1876 a_11413_103.n2 a_11413_103.n1 66.629
R1877 a_11413_103.t0 a_11413_103.n8 59.616
R1878 a_11413_103.n5 a_11413_103.n3 54.496
R1879 a_11413_103.n5 a_11413_103.n4 54.496
R1880 a_11413_103.t0 a_11413_103.n2 20.262
R1881 a_11413_103.n7 a_11413_103.n5 7.859
R1882 a_11413_103.t0 a_11413_103.n7 3.034
R1883 a_11413_103.n7 a_11413_103.n6 0.443
R1884 GND.n32 GND.n31 237.558
R1885 GND.n64 GND.n63 237.558
R1886 GND.n470 GND.n469 237.558
R1887 GND.n515 GND.n514 237.558
R1888 GND.n548 GND.n547 237.558
R1889 GND.n590 GND.n589 237.558
R1890 GND.n632 GND.n631 237.558
R1891 GND.n665 GND.n664 237.558
R1892 GND.n707 GND.n706 237.558
R1893 GND.n749 GND.n748 237.558
R1894 GND.n781 GND.n780 237.558
R1895 GND.n402 GND.n401 237.558
R1896 GND.n825 GND.n824 237.558
R1897 GND.n370 GND.n369 237.558
R1898 GND.n325 GND.n324 237.558
R1899 GND.n281 GND.n280 237.558
R1900 GND.n248 GND.n247 237.558
R1901 GND.n206 GND.n205 237.558
R1902 GND.n161 GND.n160 237.558
R1903 GND.n128 GND.n127 237.558
R1904 GND.n96 GND.n95 237.558
R1905 GND.n29 GND.n28 210.82
R1906 GND.n61 GND.n60 210.82
R1907 GND.n93 GND.n92 210.82
R1908 GND.n472 GND.n471 210.82
R1909 GND.n517 GND.n516 210.82
R1910 GND.n550 GND.n549 210.82
R1911 GND.n592 GND.n591 210.82
R1912 GND.n634 GND.n633 210.82
R1913 GND.n667 GND.n666 210.82
R1914 GND.n709 GND.n708 210.82
R1915 GND.n751 GND.n750 210.82
R1916 GND.n783 GND.n782 210.82
R1917 GND.n827 GND.n826 210.82
R1918 GND.n399 GND.n398 210.82
R1919 GND.n367 GND.n366 210.82
R1920 GND.n322 GND.n321 210.82
R1921 GND.n278 GND.n277 210.82
R1922 GND.n245 GND.n244 210.82
R1923 GND.n203 GND.n202 210.82
R1924 GND.n158 GND.n157 210.82
R1925 GND.n125 GND.n124 210.82
R1926 GND.n235 GND.n234 173.365
R1927 GND.n836 GND.n835 173.365
R1928 GND.n718 GND.n717 173.365
R1929 GND.n676 GND.n675 173.365
R1930 GND.n601 GND.n600 173.365
R1931 GND.n559 GND.n558 173.365
R1932 GND.n312 GND.n311 167.358
R1933 GND.n794 GND.n793 167.358
R1934 GND.n439 GND.n438 167.358
R1935 GND.n82 GND.n81 166.605
R1936 GND.n114 GND.n113 166.605
R1937 GND.n388 GND.n387 166.605
R1938 GND.n761 GND.n760 166.605
R1939 GND.n50 GND.n49 166.605
R1940 GND.n193 GND.n192 152.358
R1941 GND.n357 GND.n356 152.358
R1942 GND.n484 GND.n483 152.358
R1943 GND.n147 GND.n146 151.605
R1944 GND.n267 GND.n266 151.605
R1945 GND.n645 GND.n644 151.605
R1946 GND.n528 GND.n527 151.605
R1947 GND.n20 GND.n19 37.582
R1948 GND.t4 GND.n17 32.601
R1949 GND.n146 GND.n145 28.421
R1950 GND.n192 GND.n191 28.421
R1951 GND.n266 GND.n265 28.421
R1952 GND.n356 GND.n355 28.421
R1953 GND.n644 GND.n643 28.421
R1954 GND.n527 GND.n526 28.421
R1955 GND.n483 GND.n482 28.421
R1956 GND.n146 GND.n144 25.263
R1957 GND.n192 GND.n190 25.263
R1958 GND.n266 GND.n264 25.263
R1959 GND.n356 GND.n354 25.263
R1960 GND.n644 GND.n642 25.263
R1961 GND.n527 GND.n525 25.263
R1962 GND.n483 GND.n481 25.263
R1963 GND.n144 GND.n143 24.383
R1964 GND.n190 GND.n189 24.383
R1965 GND.n264 GND.n263 24.383
R1966 GND.n354 GND.n353 24.383
R1967 GND.n642 GND.n641 24.383
R1968 GND.n525 GND.n524 24.383
R1969 GND.n481 GND.n480 24.383
R1970 GND.n81 GND.n79 23.03
R1971 GND.n113 GND.n111 23.03
R1972 GND.n311 GND.n309 23.03
R1973 GND.n387 GND.n385 23.03
R1974 GND.n793 GND.n791 23.03
R1975 GND.n760 GND.n758 23.03
R1976 GND.n438 GND.n436 23.03
R1977 GND.n49 GND.n47 23.03
R1978 GND.n17 GND.n16 21.734
R1979 GND.n4 GND.n3 20.705
R1980 GND.n10 GND.n9 20.705
R1981 GND.n21 GND.n20 20.705
R1982 GND.n3 GND.n2 19.952
R1983 GND.n30 GND.n29 18.953
R1984 GND.n62 GND.n61 18.953
R1985 GND.n94 GND.n93 18.953
R1986 GND.n473 GND.n472 18.953
R1987 GND.n518 GND.n517 18.953
R1988 GND.n551 GND.n550 18.953
R1989 GND.n593 GND.n592 18.953
R1990 GND.n635 GND.n634 18.953
R1991 GND.n668 GND.n667 18.953
R1992 GND.n710 GND.n709 18.953
R1993 GND.n752 GND.n751 18.953
R1994 GND.n784 GND.n783 18.953
R1995 GND.n828 GND.n827 18.953
R1996 GND.n400 GND.n399 18.953
R1997 GND.n368 GND.n367 18.953
R1998 GND.n323 GND.n322 18.953
R1999 GND.n279 GND.n278 18.953
R2000 GND.n246 GND.n245 18.953
R2001 GND.n204 GND.n203 18.953
R2002 GND.n159 GND.n158 18.953
R2003 GND.n126 GND.n125 18.953
R2004 GND.n19 GND.t4 15.644
R2005 GND.n33 GND.n30 14.864
R2006 GND.n65 GND.n62 14.864
R2007 GND.n97 GND.n94 14.864
R2008 GND.n129 GND.n126 14.864
R2009 GND.n162 GND.n159 14.864
R2010 GND.n207 GND.n204 14.864
R2011 GND.n249 GND.n246 14.864
R2012 GND.n282 GND.n279 14.864
R2013 GND.n326 GND.n323 14.864
R2014 GND.n371 GND.n368 14.864
R2015 GND.n403 GND.n400 14.864
R2016 GND.n829 GND.n828 14.864
R2017 GND.n785 GND.n784 14.864
R2018 GND.n753 GND.n752 14.864
R2019 GND.n711 GND.n710 14.864
R2020 GND.n669 GND.n668 14.864
R2021 GND.n636 GND.n635 14.864
R2022 GND.n594 GND.n593 14.864
R2023 GND.n552 GND.n551 14.864
R2024 GND.n519 GND.n518 14.864
R2025 GND.n474 GND.n473 14.864
R2026 GND.n19 GND.n18 13.541
R2027 GND.n433 GND.n432 9.154
R2028 GND.n440 GND.n435 9.154
R2029 GND.n443 GND.n442 9.154
R2030 GND.n446 GND.n445 9.154
R2031 GND.n449 GND.n448 9.154
R2032 GND.n452 GND.n451 9.154
R2033 GND.n455 GND.n454 9.154
R2034 GND.n458 GND.n457 9.154
R2035 GND.n461 GND.n460 9.154
R2036 GND.n464 GND.n463 9.154
R2037 GND.n467 GND.n466 9.154
R2038 GND.n474 GND.n470 9.154
R2039 GND.n477 GND.n476 9.154
R2040 GND.n485 GND.n479 9.154
R2041 GND.n488 GND.n487 9.154
R2042 GND.n491 GND.n490 9.154
R2043 GND.n494 GND.n493 9.154
R2044 GND.n497 GND.n496 9.154
R2045 GND.n500 GND.n499 9.154
R2046 GND.n503 GND.n502 9.154
R2047 GND.n506 GND.n505 9.154
R2048 GND.n509 GND.n508 9.154
R2049 GND.n512 GND.n511 9.154
R2050 GND.n519 GND.n515 9.154
R2051 GND.n522 GND.n521 9.154
R2052 GND.n530 GND.n529 9.154
R2053 GND.n533 GND.n532 9.154
R2054 GND.n536 GND.n535 9.154
R2055 GND.n539 GND.n538 9.154
R2056 GND.n542 GND.n541 9.154
R2057 GND.n545 GND.n544 9.154
R2058 GND.n552 GND.n548 9.154
R2059 GND.n555 GND.n554 9.154
R2060 GND.n560 GND.n557 9.154
R2061 GND.n563 GND.n562 9.154
R2062 GND.n566 GND.n565 9.154
R2063 GND.n569 GND.n568 9.154
R2064 GND.n572 GND.n571 9.154
R2065 GND.n575 GND.n574 9.154
R2066 GND.n578 GND.n577 9.154
R2067 GND.n581 GND.n580 9.154
R2068 GND.n584 GND.n583 9.154
R2069 GND.n587 GND.n586 9.154
R2070 GND.n594 GND.n590 9.154
R2071 GND.n597 GND.n596 9.154
R2072 GND.n602 GND.n599 9.154
R2073 GND.n605 GND.n604 9.154
R2074 GND.n608 GND.n607 9.154
R2075 GND.n611 GND.n610 9.154
R2076 GND.n614 GND.n613 9.154
R2077 GND.n617 GND.n616 9.154
R2078 GND.n620 GND.n619 9.154
R2079 GND.n623 GND.n622 9.154
R2080 GND.n626 GND.n625 9.154
R2081 GND.n629 GND.n628 9.154
R2082 GND.n636 GND.n632 9.154
R2083 GND.n639 GND.n638 9.154
R2084 GND.n647 GND.n646 9.154
R2085 GND.n650 GND.n649 9.154
R2086 GND.n653 GND.n652 9.154
R2087 GND.n656 GND.n655 9.154
R2088 GND.n659 GND.n658 9.154
R2089 GND.n662 GND.n661 9.154
R2090 GND.n669 GND.n665 9.154
R2091 GND.n672 GND.n671 9.154
R2092 GND.n677 GND.n674 9.154
R2093 GND.n680 GND.n679 9.154
R2094 GND.n683 GND.n682 9.154
R2095 GND.n686 GND.n685 9.154
R2096 GND.n689 GND.n688 9.154
R2097 GND.n692 GND.n691 9.154
R2098 GND.n695 GND.n694 9.154
R2099 GND.n698 GND.n697 9.154
R2100 GND.n701 GND.n700 9.154
R2101 GND.n704 GND.n703 9.154
R2102 GND.n711 GND.n707 9.154
R2103 GND.n714 GND.n713 9.154
R2104 GND.n719 GND.n716 9.154
R2105 GND.n722 GND.n721 9.154
R2106 GND.n725 GND.n724 9.154
R2107 GND.n728 GND.n727 9.154
R2108 GND.n731 GND.n730 9.154
R2109 GND.n734 GND.n733 9.154
R2110 GND.n737 GND.n736 9.154
R2111 GND.n740 GND.n739 9.154
R2112 GND.n743 GND.n742 9.154
R2113 GND.n746 GND.n745 9.154
R2114 GND.n753 GND.n749 9.154
R2115 GND.n756 GND.n755 9.154
R2116 GND.n763 GND.n762 9.154
R2117 GND.n766 GND.n765 9.154
R2118 GND.n769 GND.n768 9.154
R2119 GND.n772 GND.n771 9.154
R2120 GND.n775 GND.n774 9.154
R2121 GND.n778 GND.n777 9.154
R2122 GND.n785 GND.n781 9.154
R2123 GND.n788 GND.n787 9.154
R2124 GND.n795 GND.n790 9.154
R2125 GND.n798 GND.n797 9.154
R2126 GND.n801 GND.n800 9.154
R2127 GND.n804 GND.n803 9.154
R2128 GND.n807 GND.n806 9.154
R2129 GND.n810 GND.n809 9.154
R2130 GND.n813 GND.n812 9.154
R2131 GND.n816 GND.n815 9.154
R2132 GND.n819 GND.n818 9.154
R2133 GND.n822 GND.n821 9.154
R2134 GND.n829 GND.n825 9.154
R2135 GND.n832 GND.n831 9.154
R2136 GND.n837 GND.n834 9.154
R2137 GND.n427 GND.n426 9.154
R2138 GND.n424 GND.n423 9.154
R2139 GND.n421 GND.n420 9.154
R2140 GND.n418 GND.n417 9.154
R2141 GND.n415 GND.n414 9.154
R2142 GND.n412 GND.n411 9.154
R2143 GND.n409 GND.n408 9.154
R2144 GND.n406 GND.n405 9.154
R2145 GND.n403 GND.n402 9.154
R2146 GND.n396 GND.n395 9.154
R2147 GND.n393 GND.n392 9.154
R2148 GND.n390 GND.n389 9.154
R2149 GND.n383 GND.n382 9.154
R2150 GND.n380 GND.n379 9.154
R2151 GND.n377 GND.n376 9.154
R2152 GND.n374 GND.n373 9.154
R2153 GND.n371 GND.n370 9.154
R2154 GND.n364 GND.n363 9.154
R2155 GND.n361 GND.n360 9.154
R2156 GND.n358 GND.n352 9.154
R2157 GND.n350 GND.n349 9.154
R2158 GND.n347 GND.n346 9.154
R2159 GND.n344 GND.n343 9.154
R2160 GND.n341 GND.n340 9.154
R2161 GND.n338 GND.n337 9.154
R2162 GND.n335 GND.n334 9.154
R2163 GND.n332 GND.n331 9.154
R2164 GND.n329 GND.n328 9.154
R2165 GND.n326 GND.n325 9.154
R2166 GND.n319 GND.n318 9.154
R2167 GND.n316 GND.n315 9.154
R2168 GND.n313 GND.n308 9.154
R2169 GND.n306 GND.n305 9.154
R2170 GND.n303 GND.n302 9.154
R2171 GND.n300 GND.n299 9.154
R2172 GND.n297 GND.n296 9.154
R2173 GND.n294 GND.n293 9.154
R2174 GND.n291 GND.n290 9.154
R2175 GND.n288 GND.n287 9.154
R2176 GND.n285 GND.n284 9.154
R2177 GND.n282 GND.n281 9.154
R2178 GND.n275 GND.n274 9.154
R2179 GND.n272 GND.n271 9.154
R2180 GND.n269 GND.n268 9.154
R2181 GND.n261 GND.n260 9.154
R2182 GND.n258 GND.n257 9.154
R2183 GND.n255 GND.n254 9.154
R2184 GND.n252 GND.n251 9.154
R2185 GND.n249 GND.n248 9.154
R2186 GND.n242 GND.n241 9.154
R2187 GND.n239 GND.n238 9.154
R2188 GND.n236 GND.n233 9.154
R2189 GND.n231 GND.n230 9.154
R2190 GND.n228 GND.n227 9.154
R2191 GND.n225 GND.n224 9.154
R2192 GND.n222 GND.n221 9.154
R2193 GND.n219 GND.n218 9.154
R2194 GND.n216 GND.n215 9.154
R2195 GND.n213 GND.n212 9.154
R2196 GND.n210 GND.n209 9.154
R2197 GND.n207 GND.n206 9.154
R2198 GND.n200 GND.n199 9.154
R2199 GND.n197 GND.n196 9.154
R2200 GND.n194 GND.n188 9.154
R2201 GND.n186 GND.n185 9.154
R2202 GND.n183 GND.n182 9.154
R2203 GND.n180 GND.n179 9.154
R2204 GND.n177 GND.n176 9.154
R2205 GND.n174 GND.n173 9.154
R2206 GND.n171 GND.n170 9.154
R2207 GND.n168 GND.n167 9.154
R2208 GND.n165 GND.n164 9.154
R2209 GND.n162 GND.n161 9.154
R2210 GND.n155 GND.n154 9.154
R2211 GND.n152 GND.n151 9.154
R2212 GND.n149 GND.n148 9.154
R2213 GND.n141 GND.n140 9.154
R2214 GND.n138 GND.n137 9.154
R2215 GND.n135 GND.n134 9.154
R2216 GND.n132 GND.n131 9.154
R2217 GND.n129 GND.n128 9.154
R2218 GND.n122 GND.n121 9.154
R2219 GND.n119 GND.n118 9.154
R2220 GND.n116 GND.n115 9.154
R2221 GND.n109 GND.n108 9.154
R2222 GND.n106 GND.n105 9.154
R2223 GND.n103 GND.n102 9.154
R2224 GND.n100 GND.n99 9.154
R2225 GND.n97 GND.n96 9.154
R2226 GND.n90 GND.n89 9.154
R2227 GND.n87 GND.n86 9.154
R2228 GND.n84 GND.n83 9.154
R2229 GND.n77 GND.n76 9.154
R2230 GND.n74 GND.n73 9.154
R2231 GND.n6 GND.n5 9.154
R2232 GND.n12 GND.n11 9.154
R2233 GND.n23 GND.n22 9.154
R2234 GND.n26 GND.n25 9.154
R2235 GND.n33 GND.n32 9.154
R2236 GND.n36 GND.n35 9.154
R2237 GND.n39 GND.n38 9.154
R2238 GND.n42 GND.n41 9.154
R2239 GND.n45 GND.n44 9.154
R2240 GND.n52 GND.n51 9.154
R2241 GND.n55 GND.n54 9.154
R2242 GND.n58 GND.n57 9.154
R2243 GND.n65 GND.n64 9.154
R2244 GND.n68 GND.n67 9.154
R2245 GND.n71 GND.n70 9.154
R2246 GND.n81 GND.n80 8.128
R2247 GND.n113 GND.n112 8.128
R2248 GND.n311 GND.n310 8.128
R2249 GND.n387 GND.n386 8.128
R2250 GND.n793 GND.n792 8.128
R2251 GND.n760 GND.n759 8.128
R2252 GND.n438 GND.n437 8.128
R2253 GND.n49 GND.n48 8.128
R2254 GND.n7 GND.n1 4.795
R2255 GND.n431 GND.n430 4.65
R2256 GND.n75 GND.n74 4.65
R2257 GND.n78 GND.n77 4.65
R2258 GND.n85 GND.n84 4.65
R2259 GND.n88 GND.n87 4.65
R2260 GND.n91 GND.n90 4.65
R2261 GND.n98 GND.n97 4.65
R2262 GND.n101 GND.n100 4.65
R2263 GND.n104 GND.n103 4.65
R2264 GND.n107 GND.n106 4.65
R2265 GND.n110 GND.n109 4.65
R2266 GND.n117 GND.n116 4.65
R2267 GND.n120 GND.n119 4.65
R2268 GND.n123 GND.n122 4.65
R2269 GND.n130 GND.n129 4.65
R2270 GND.n133 GND.n132 4.65
R2271 GND.n136 GND.n135 4.65
R2272 GND.n139 GND.n138 4.65
R2273 GND.n142 GND.n141 4.65
R2274 GND.n150 GND.n149 4.65
R2275 GND.n153 GND.n152 4.65
R2276 GND.n156 GND.n155 4.65
R2277 GND.n163 GND.n162 4.65
R2278 GND.n166 GND.n165 4.65
R2279 GND.n169 GND.n168 4.65
R2280 GND.n172 GND.n171 4.65
R2281 GND.n175 GND.n174 4.65
R2282 GND.n178 GND.n177 4.65
R2283 GND.n181 GND.n180 4.65
R2284 GND.n184 GND.n183 4.65
R2285 GND.n187 GND.n186 4.65
R2286 GND.n195 GND.n194 4.65
R2287 GND.n198 GND.n197 4.65
R2288 GND.n201 GND.n200 4.65
R2289 GND.n208 GND.n207 4.65
R2290 GND.n211 GND.n210 4.65
R2291 GND.n214 GND.n213 4.65
R2292 GND.n217 GND.n216 4.65
R2293 GND.n220 GND.n219 4.65
R2294 GND.n223 GND.n222 4.65
R2295 GND.n226 GND.n225 4.65
R2296 GND.n229 GND.n228 4.65
R2297 GND.n232 GND.n231 4.65
R2298 GND.n237 GND.n236 4.65
R2299 GND.n240 GND.n239 4.65
R2300 GND.n243 GND.n242 4.65
R2301 GND.n250 GND.n249 4.65
R2302 GND.n253 GND.n252 4.65
R2303 GND.n256 GND.n255 4.65
R2304 GND.n259 GND.n258 4.65
R2305 GND.n262 GND.n261 4.65
R2306 GND.n270 GND.n269 4.65
R2307 GND.n273 GND.n272 4.65
R2308 GND.n276 GND.n275 4.65
R2309 GND.n283 GND.n282 4.65
R2310 GND.n286 GND.n285 4.65
R2311 GND.n289 GND.n288 4.65
R2312 GND.n292 GND.n291 4.65
R2313 GND.n295 GND.n294 4.65
R2314 GND.n298 GND.n297 4.65
R2315 GND.n301 GND.n300 4.65
R2316 GND.n304 GND.n303 4.65
R2317 GND.n307 GND.n306 4.65
R2318 GND.n314 GND.n313 4.65
R2319 GND.n317 GND.n316 4.65
R2320 GND.n320 GND.n319 4.65
R2321 GND.n327 GND.n326 4.65
R2322 GND.n330 GND.n329 4.65
R2323 GND.n333 GND.n332 4.65
R2324 GND.n336 GND.n335 4.65
R2325 GND.n339 GND.n338 4.65
R2326 GND.n342 GND.n341 4.65
R2327 GND.n345 GND.n344 4.65
R2328 GND.n348 GND.n347 4.65
R2329 GND.n351 GND.n350 4.65
R2330 GND.n359 GND.n358 4.65
R2331 GND.n362 GND.n361 4.65
R2332 GND.n365 GND.n364 4.65
R2333 GND.n372 GND.n371 4.65
R2334 GND.n375 GND.n374 4.65
R2335 GND.n378 GND.n377 4.65
R2336 GND.n381 GND.n380 4.65
R2337 GND.n384 GND.n383 4.65
R2338 GND.n391 GND.n390 4.65
R2339 GND.n394 GND.n393 4.65
R2340 GND.n397 GND.n396 4.65
R2341 GND.n404 GND.n403 4.65
R2342 GND.n407 GND.n406 4.65
R2343 GND.n410 GND.n409 4.65
R2344 GND.n413 GND.n412 4.65
R2345 GND.n416 GND.n415 4.65
R2346 GND.n419 GND.n418 4.65
R2347 GND.n422 GND.n421 4.65
R2348 GND.n425 GND.n424 4.65
R2349 GND.n428 GND.n427 4.65
R2350 GND.n838 GND.n837 4.65
R2351 GND.n833 GND.n832 4.65
R2352 GND.n830 GND.n829 4.65
R2353 GND.n823 GND.n822 4.65
R2354 GND.n820 GND.n819 4.65
R2355 GND.n817 GND.n816 4.65
R2356 GND.n814 GND.n813 4.65
R2357 GND.n811 GND.n810 4.65
R2358 GND.n808 GND.n807 4.65
R2359 GND.n805 GND.n804 4.65
R2360 GND.n802 GND.n801 4.65
R2361 GND.n799 GND.n798 4.65
R2362 GND.n796 GND.n795 4.65
R2363 GND.n789 GND.n788 4.65
R2364 GND.n786 GND.n785 4.65
R2365 GND.n779 GND.n778 4.65
R2366 GND.n776 GND.n775 4.65
R2367 GND.n773 GND.n772 4.65
R2368 GND.n770 GND.n769 4.65
R2369 GND.n767 GND.n766 4.65
R2370 GND.n764 GND.n763 4.65
R2371 GND.n757 GND.n756 4.65
R2372 GND.n754 GND.n753 4.65
R2373 GND.n747 GND.n746 4.65
R2374 GND.n744 GND.n743 4.65
R2375 GND.n741 GND.n740 4.65
R2376 GND.n738 GND.n737 4.65
R2377 GND.n735 GND.n734 4.65
R2378 GND.n732 GND.n731 4.65
R2379 GND.n729 GND.n728 4.65
R2380 GND.n726 GND.n725 4.65
R2381 GND.n723 GND.n722 4.65
R2382 GND.n720 GND.n719 4.65
R2383 GND.n715 GND.n714 4.65
R2384 GND.n712 GND.n711 4.65
R2385 GND.n705 GND.n704 4.65
R2386 GND.n702 GND.n701 4.65
R2387 GND.n699 GND.n698 4.65
R2388 GND.n696 GND.n695 4.65
R2389 GND.n693 GND.n692 4.65
R2390 GND.n690 GND.n689 4.65
R2391 GND.n687 GND.n686 4.65
R2392 GND.n684 GND.n683 4.65
R2393 GND.n681 GND.n680 4.65
R2394 GND.n678 GND.n677 4.65
R2395 GND.n673 GND.n672 4.65
R2396 GND.n670 GND.n669 4.65
R2397 GND.n663 GND.n662 4.65
R2398 GND.n660 GND.n659 4.65
R2399 GND.n657 GND.n656 4.65
R2400 GND.n654 GND.n653 4.65
R2401 GND.n651 GND.n650 4.65
R2402 GND.n648 GND.n647 4.65
R2403 GND.n640 GND.n639 4.65
R2404 GND.n637 GND.n636 4.65
R2405 GND.n630 GND.n629 4.65
R2406 GND.n627 GND.n626 4.65
R2407 GND.n624 GND.n623 4.65
R2408 GND.n621 GND.n620 4.65
R2409 GND.n618 GND.n617 4.65
R2410 GND.n615 GND.n614 4.65
R2411 GND.n612 GND.n611 4.65
R2412 GND.n609 GND.n608 4.65
R2413 GND.n606 GND.n605 4.65
R2414 GND.n603 GND.n602 4.65
R2415 GND.n598 GND.n597 4.65
R2416 GND.n595 GND.n594 4.65
R2417 GND.n588 GND.n587 4.65
R2418 GND.n585 GND.n584 4.65
R2419 GND.n582 GND.n581 4.65
R2420 GND.n579 GND.n578 4.65
R2421 GND.n576 GND.n575 4.65
R2422 GND.n573 GND.n572 4.65
R2423 GND.n570 GND.n569 4.65
R2424 GND.n567 GND.n566 4.65
R2425 GND.n564 GND.n563 4.65
R2426 GND.n561 GND.n560 4.65
R2427 GND.n556 GND.n555 4.65
R2428 GND.n553 GND.n552 4.65
R2429 GND.n546 GND.n545 4.65
R2430 GND.n543 GND.n542 4.65
R2431 GND.n540 GND.n539 4.65
R2432 GND.n537 GND.n536 4.65
R2433 GND.n534 GND.n533 4.65
R2434 GND.n531 GND.n530 4.65
R2435 GND.n523 GND.n522 4.65
R2436 GND.n520 GND.n519 4.65
R2437 GND.n513 GND.n512 4.65
R2438 GND.n510 GND.n509 4.65
R2439 GND.n507 GND.n506 4.65
R2440 GND.n504 GND.n503 4.65
R2441 GND.n501 GND.n500 4.65
R2442 GND.n498 GND.n497 4.65
R2443 GND.n495 GND.n494 4.65
R2444 GND.n492 GND.n491 4.65
R2445 GND.n489 GND.n488 4.65
R2446 GND.n486 GND.n485 4.65
R2447 GND.n478 GND.n477 4.65
R2448 GND.n475 GND.n474 4.65
R2449 GND.n468 GND.n467 4.65
R2450 GND.n465 GND.n464 4.65
R2451 GND.n462 GND.n461 4.65
R2452 GND.n459 GND.n458 4.65
R2453 GND.n456 GND.n455 4.65
R2454 GND.n453 GND.n452 4.65
R2455 GND.n450 GND.n449 4.65
R2456 GND.n447 GND.n446 4.65
R2457 GND.n444 GND.n443 4.65
R2458 GND.n441 GND.n440 4.65
R2459 GND.n434 GND.n433 4.65
R2460 GND.n7 GND.n6 4.65
R2461 GND.n13 GND.n12 4.65
R2462 GND.n24 GND.n23 4.65
R2463 GND.n27 GND.n26 4.65
R2464 GND.n34 GND.n33 4.65
R2465 GND.n37 GND.n36 4.65
R2466 GND.n40 GND.n39 4.65
R2467 GND.n43 GND.n42 4.65
R2468 GND.n46 GND.n45 4.65
R2469 GND.n53 GND.n52 4.65
R2470 GND.n56 GND.n55 4.65
R2471 GND.n59 GND.n58 4.65
R2472 GND.n66 GND.n65 4.65
R2473 GND.n69 GND.n68 4.65
R2474 GND.n72 GND.n71 4.65
R2475 GND.n15 GND.n14 4.504
R2476 GND.n6 GND.n4 4.129
R2477 GND.n52 GND.n50 4.129
R2478 GND.n84 GND.n82 4.129
R2479 GND.n116 GND.n114 4.129
R2480 GND.n149 GND.n147 4.129
R2481 GND.n269 GND.n267 4.129
R2482 GND.n390 GND.n388 4.129
R2483 GND.n763 GND.n761 4.129
R2484 GND.n647 GND.n645 4.129
R2485 GND.n530 GND.n528 4.129
R2486 GND.n23 GND.n21 3.716
R2487 GND.t4 GND.n15 2.452
R2488 GND.n1 GND.n0 0.475
R2489 GND.n430 GND.n429 0.474
R2490 GND.n9 GND.n8 0.376
R2491 GND.n34 GND.n27 0.29
R2492 GND.n66 GND.n59 0.29
R2493 GND.n98 GND.n91 0.29
R2494 GND.n130 GND.n123 0.29
R2495 GND.n163 GND.n156 0.29
R2496 GND.n208 GND.n201 0.29
R2497 GND.n250 GND.n243 0.29
R2498 GND.n283 GND.n276 0.29
R2499 GND.n327 GND.n320 0.29
R2500 GND.n372 GND.n365 0.29
R2501 GND.n404 GND.n397 0.29
R2502 GND.n830 GND.n823 0.29
R2503 GND.n786 GND.n779 0.29
R2504 GND.n754 GND.n747 0.29
R2505 GND.n712 GND.n705 0.29
R2506 GND.n670 GND.n663 0.29
R2507 GND.n637 GND.n630 0.29
R2508 GND.n595 GND.n588 0.29
R2509 GND.n553 GND.n546 0.29
R2510 GND.n520 GND.n513 0.29
R2511 GND.n475 GND.n468 0.29
R2512 GND.n431 GND 0.207
R2513 GND.n12 GND.n10 0.206
R2514 GND.n194 GND.n193 0.206
R2515 GND.n236 GND.n235 0.206
R2516 GND.n313 GND.n312 0.206
R2517 GND.n358 GND.n357 0.206
R2518 GND.n837 GND.n836 0.206
R2519 GND.n795 GND.n794 0.206
R2520 GND.n719 GND.n718 0.206
R2521 GND.n677 GND.n676 0.206
R2522 GND.n602 GND.n601 0.206
R2523 GND.n560 GND.n559 0.206
R2524 GND.n485 GND.n484 0.206
R2525 GND.n440 GND.n439 0.206
R2526 GND.n181 GND.n178 0.197
R2527 GND.n226 GND.n223 0.197
R2528 GND.n301 GND.n298 0.197
R2529 GND.n345 GND.n342 0.197
R2530 GND.n422 GND.n419 0.197
R2531 GND.n808 GND.n805 0.197
R2532 GND.n732 GND.n729 0.197
R2533 GND.n690 GND.n687 0.197
R2534 GND.n615 GND.n612 0.197
R2535 GND.n573 GND.n570 0.197
R2536 GND.n498 GND.n495 0.197
R2537 GND.n453 GND.n450 0.197
R2538 GND.n46 GND.n43 0.181
R2539 GND.n78 GND.n75 0.181
R2540 GND.n110 GND.n107 0.181
R2541 GND.n142 GND.n139 0.181
R2542 GND.n262 GND.n259 0.181
R2543 GND.n384 GND.n381 0.181
R2544 GND.n770 GND.n767 0.181
R2545 GND.n654 GND.n651 0.181
R2546 GND.n537 GND.n534 0.181
R2547 GND.n13 GND.n7 0.157
R2548 GND.n24 GND.n13 0.157
R2549 GND.n27 GND.n24 0.145
R2550 GND.n37 GND.n34 0.145
R2551 GND.n40 GND.n37 0.145
R2552 GND.n43 GND.n40 0.145
R2553 GND.n53 GND.n46 0.145
R2554 GND.n56 GND.n53 0.145
R2555 GND.n59 GND.n56 0.145
R2556 GND.n69 GND.n66 0.145
R2557 GND.n72 GND.n69 0.145
R2558 GND.n75 GND.n72 0.145
R2559 GND.n85 GND.n78 0.145
R2560 GND.n88 GND.n85 0.145
R2561 GND.n91 GND.n88 0.145
R2562 GND.n101 GND.n98 0.145
R2563 GND.n104 GND.n101 0.145
R2564 GND.n107 GND.n104 0.145
R2565 GND.n117 GND.n110 0.145
R2566 GND.n120 GND.n117 0.145
R2567 GND.n123 GND.n120 0.145
R2568 GND.n133 GND.n130 0.145
R2569 GND.n136 GND.n133 0.145
R2570 GND.n139 GND.n136 0.145
R2571 GND.n150 GND.n142 0.145
R2572 GND.n153 GND.n150 0.145
R2573 GND.n156 GND.n153 0.145
R2574 GND.n166 GND.n163 0.145
R2575 GND.n169 GND.n166 0.145
R2576 GND.n172 GND.n169 0.145
R2577 GND.n175 GND.n172 0.145
R2578 GND.n178 GND.n175 0.145
R2579 GND.n184 GND.n181 0.145
R2580 GND.n187 GND.n184 0.145
R2581 GND.n195 GND.n187 0.145
R2582 GND.n198 GND.n195 0.145
R2583 GND.n201 GND.n198 0.145
R2584 GND.n211 GND.n208 0.145
R2585 GND.n214 GND.n211 0.145
R2586 GND.n217 GND.n214 0.145
R2587 GND.n220 GND.n217 0.145
R2588 GND.n223 GND.n220 0.145
R2589 GND.n229 GND.n226 0.145
R2590 GND.n232 GND.n229 0.145
R2591 GND.n237 GND.n232 0.145
R2592 GND.n240 GND.n237 0.145
R2593 GND.n243 GND.n240 0.145
R2594 GND.n253 GND.n250 0.145
R2595 GND.n256 GND.n253 0.145
R2596 GND.n259 GND.n256 0.145
R2597 GND.n270 GND.n262 0.145
R2598 GND.n273 GND.n270 0.145
R2599 GND.n276 GND.n273 0.145
R2600 GND.n286 GND.n283 0.145
R2601 GND.n289 GND.n286 0.145
R2602 GND.n292 GND.n289 0.145
R2603 GND.n295 GND.n292 0.145
R2604 GND.n298 GND.n295 0.145
R2605 GND.n304 GND.n301 0.145
R2606 GND.n307 GND.n304 0.145
R2607 GND.n314 GND.n307 0.145
R2608 GND.n317 GND.n314 0.145
R2609 GND.n320 GND.n317 0.145
R2610 GND.n330 GND.n327 0.145
R2611 GND.n333 GND.n330 0.145
R2612 GND.n336 GND.n333 0.145
R2613 GND.n339 GND.n336 0.145
R2614 GND.n342 GND.n339 0.145
R2615 GND.n348 GND.n345 0.145
R2616 GND.n351 GND.n348 0.145
R2617 GND.n359 GND.n351 0.145
R2618 GND.n362 GND.n359 0.145
R2619 GND.n365 GND.n362 0.145
R2620 GND.n375 GND.n372 0.145
R2621 GND.n378 GND.n375 0.145
R2622 GND.n381 GND.n378 0.145
R2623 GND.n391 GND.n384 0.145
R2624 GND.n394 GND.n391 0.145
R2625 GND.n397 GND.n394 0.145
R2626 GND.n407 GND.n404 0.145
R2627 GND.n410 GND.n407 0.145
R2628 GND.n413 GND.n410 0.145
R2629 GND.n416 GND.n413 0.145
R2630 GND.n419 GND.n416 0.145
R2631 GND.n425 GND.n422 0.145
R2632 GND.n428 GND.n425 0.145
R2633 GND.n838 GND.n833 0.145
R2634 GND.n833 GND.n830 0.145
R2635 GND.n823 GND.n820 0.145
R2636 GND.n820 GND.n817 0.145
R2637 GND.n817 GND.n814 0.145
R2638 GND.n814 GND.n811 0.145
R2639 GND.n811 GND.n808 0.145
R2640 GND.n805 GND.n802 0.145
R2641 GND.n802 GND.n799 0.145
R2642 GND.n799 GND.n796 0.145
R2643 GND.n796 GND.n789 0.145
R2644 GND.n789 GND.n786 0.145
R2645 GND.n779 GND.n776 0.145
R2646 GND.n776 GND.n773 0.145
R2647 GND.n773 GND.n770 0.145
R2648 GND.n767 GND.n764 0.145
R2649 GND.n764 GND.n757 0.145
R2650 GND.n757 GND.n754 0.145
R2651 GND.n747 GND.n744 0.145
R2652 GND.n744 GND.n741 0.145
R2653 GND.n741 GND.n738 0.145
R2654 GND.n738 GND.n735 0.145
R2655 GND.n735 GND.n732 0.145
R2656 GND.n729 GND.n726 0.145
R2657 GND.n726 GND.n723 0.145
R2658 GND.n723 GND.n720 0.145
R2659 GND.n720 GND.n715 0.145
R2660 GND.n715 GND.n712 0.145
R2661 GND.n705 GND.n702 0.145
R2662 GND.n702 GND.n699 0.145
R2663 GND.n699 GND.n696 0.145
R2664 GND.n696 GND.n693 0.145
R2665 GND.n693 GND.n690 0.145
R2666 GND.n687 GND.n684 0.145
R2667 GND.n684 GND.n681 0.145
R2668 GND.n681 GND.n678 0.145
R2669 GND.n678 GND.n673 0.145
R2670 GND.n673 GND.n670 0.145
R2671 GND.n663 GND.n660 0.145
R2672 GND.n660 GND.n657 0.145
R2673 GND.n657 GND.n654 0.145
R2674 GND.n651 GND.n648 0.145
R2675 GND.n648 GND.n640 0.145
R2676 GND.n640 GND.n637 0.145
R2677 GND.n630 GND.n627 0.145
R2678 GND.n627 GND.n624 0.145
R2679 GND.n624 GND.n621 0.145
R2680 GND.n621 GND.n618 0.145
R2681 GND.n618 GND.n615 0.145
R2682 GND.n612 GND.n609 0.145
R2683 GND.n609 GND.n606 0.145
R2684 GND.n606 GND.n603 0.145
R2685 GND.n603 GND.n598 0.145
R2686 GND.n598 GND.n595 0.145
R2687 GND.n588 GND.n585 0.145
R2688 GND.n585 GND.n582 0.145
R2689 GND.n582 GND.n579 0.145
R2690 GND.n579 GND.n576 0.145
R2691 GND.n576 GND.n573 0.145
R2692 GND.n570 GND.n567 0.145
R2693 GND.n567 GND.n564 0.145
R2694 GND.n564 GND.n561 0.145
R2695 GND.n561 GND.n556 0.145
R2696 GND.n556 GND.n553 0.145
R2697 GND.n546 GND.n543 0.145
R2698 GND.n543 GND.n540 0.145
R2699 GND.n540 GND.n537 0.145
R2700 GND.n534 GND.n531 0.145
R2701 GND.n531 GND.n523 0.145
R2702 GND.n523 GND.n520 0.145
R2703 GND.n513 GND.n510 0.145
R2704 GND.n510 GND.n507 0.145
R2705 GND.n507 GND.n504 0.145
R2706 GND.n504 GND.n501 0.145
R2707 GND.n501 GND.n498 0.145
R2708 GND.n495 GND.n492 0.145
R2709 GND.n492 GND.n489 0.145
R2710 GND.n489 GND.n486 0.145
R2711 GND.n486 GND.n478 0.145
R2712 GND.n478 GND.n475 0.145
R2713 GND.n468 GND.n465 0.145
R2714 GND.n465 GND.n462 0.145
R2715 GND.n462 GND.n459 0.145
R2716 GND.n459 GND.n456 0.145
R2717 GND.n456 GND.n453 0.145
R2718 GND.n450 GND.n447 0.145
R2719 GND.n447 GND.n444 0.145
R2720 GND.n444 GND.n441 0.145
R2721 GND.n441 GND.n434 0.145
R2722 GND.n434 GND.n431 0.145
R2723 GND GND.n838 0.086
R2724 GND GND.n428 0.058
R2725 a_14511_989.n2 a_14511_989.t5 475.572
R2726 a_14511_989.n1 a_14511_989.t6 469.145
R2727 a_14511_989.n6 a_14511_989.t8 454.685
R2728 a_14511_989.n6 a_14511_989.t13 428.979
R2729 a_14511_989.n2 a_14511_989.t11 384.527
R2730 a_14511_989.n1 a_14511_989.t9 384.527
R2731 a_14511_989.n3 a_14511_989.t10 370.613
R2732 a_14511_989.n5 a_14511_989.t7 314.896
R2733 a_14511_989.n7 a_14511_989.t12 311.683
R2734 a_14511_989.n13 a_14511_989.n12 305.581
R2735 a_14511_989.n7 a_14511_989.n6 171.288
R2736 a_14511_989.n14 a_14511_989.n13 159.999
R2737 a_14511_989.n15 a_14511_989.n14 157.963
R2738 a_14511_989.n3 a_14511_989.n2 128.028
R2739 a_14511_989.n4 a_14511_989.n1 126.97
R2740 a_14511_989.n14 a_14511_989.n0 91.706
R2741 a_14511_989.n5 a_14511_989.n4 55.717
R2742 a_14511_989.n12 a_14511_989.n11 30
R2743 a_14511_989.n10 a_14511_989.n9 24.383
R2744 a_14511_989.n12 a_14511_989.n10 23.684
R2745 a_14511_989.n0 a_14511_989.t4 14.282
R2746 a_14511_989.n0 a_14511_989.t3 14.282
R2747 a_14511_989.t1 a_14511_989.n15 14.282
R2748 a_14511_989.n15 a_14511_989.t0 14.282
R2749 a_14511_989.n4 a_14511_989.n3 14.151
R2750 a_14511_989.n8 a_14511_989.n7 7.597
R2751 a_14511_989.n8 a_14511_989.n5 6.509
R2752 a_14511_989.n13 a_14511_989.n8 4.65
R2753 a_15932_209.n4 a_15932_209.t7 512.525
R2754 a_15932_209.n4 a_15932_209.t9 371.139
R2755 a_15932_209.n5 a_15932_209.t8 338.57
R2756 a_15932_209.n10 a_15932_209.n6 227.387
R2757 a_15932_209.n5 a_15932_209.n4 191.629
R2758 a_15932_209.n3 a_15932_209.n2 165.613
R2759 a_15932_209.n6 a_15932_209.n3 132.893
R2760 a_15932_209.n15 a_15932_209.n14 112.771
R2761 a_15932_209.n17 a_15932_209.n15 110.702
R2762 a_15932_209.n10 a_15932_209.n9 106.052
R2763 a_15932_209.n3 a_15932_209.n1 99.355
R2764 a_15932_209.n9 a_15932_209.n7 80.526
R2765 a_15932_209.n18 a_15932_209.n0 55.263
R2766 a_15932_209.n14 a_15932_209.n13 30
R2767 a_15932_209.n9 a_15932_209.n8 30
R2768 a_15932_209.n17 a_15932_209.n16 30
R2769 a_15932_209.n12 a_15932_209.n11 24.383
R2770 a_15932_209.n14 a_15932_209.n12 23.684
R2771 a_15932_209.n18 a_15932_209.n17 23.684
R2772 a_15932_209.n1 a_15932_209.t4 14.282
R2773 a_15932_209.n1 a_15932_209.t3 14.282
R2774 a_15932_209.n2 a_15932_209.t1 14.282
R2775 a_15932_209.n2 a_15932_209.t2 14.282
R2776 a_15932_209.n6 a_15932_209.n5 10.343
R2777 a_15932_209.n15 a_15932_209.n10 7.053
R2778 a_16421_1051.t5 a_16421_1051.n5 179.898
R2779 a_16421_1051.n3 a_16421_1051.n2 165.613
R2780 a_16421_1051.n3 a_16421_1051.n1 142.653
R2781 a_16421_1051.n5 a_16421_1051.n4 106.183
R2782 a_16421_1051.n5 a_16421_1051.n0 99.355
R2783 a_16421_1051.n4 a_16421_1051.n3 82.665
R2784 a_16421_1051.n4 a_16421_1051.t3 73.712
R2785 a_16421_1051.n1 a_16421_1051.t1 14.282
R2786 a_16421_1051.n1 a_16421_1051.t7 14.282
R2787 a_16421_1051.n2 a_16421_1051.t6 14.282
R2788 a_16421_1051.n2 a_16421_1051.t0 14.282
R2789 a_16421_1051.n0 a_16421_1051.t4 14.282
R2790 a_16421_1051.n0 a_16421_1051.t2 14.282
R2791 a_8142_210.n12 a_8142_210.n10 171.558
R2792 a_8142_210.n7 a_8142_210.n6 117.622
R2793 a_8142_210.n5 a_8142_210.n4 92.5
R2794 a_8142_210.n9 a_8142_210.n8 92.5
R2795 a_8142_210.n10 a_8142_210.t1 75.764
R2796 a_8142_210.n5 a_8142_210.n3 65.02
R2797 a_8142_210.n13 a_8142_210.n0 49.6
R2798 a_8142_210.n7 a_8142_210.n5 36.517
R2799 a_8142_210.n3 a_8142_210.n2 35.865
R2800 a_8142_210.n12 a_8142_210.n11 27.2
R2801 a_8142_210.n13 a_8142_210.n12 22.4
R2802 a_8142_210.n9 a_8142_210.n7 19.952
R2803 a_8142_210.t1 a_8142_210.n1 7.04
R2804 a_8142_210.n10 a_8142_210.n9 1.505
R2805 a_5327_187.n4 a_5327_187.t8 512.525
R2806 a_5327_187.n2 a_5327_187.t15 472.359
R2807 a_5327_187.n0 a_5327_187.t12 472.359
R2808 a_5327_187.n5 a_5327_187.t10 417.109
R2809 a_5327_187.n2 a_5327_187.t9 384.527
R2810 a_5327_187.n0 a_5327_187.t7 384.527
R2811 a_5327_187.n11 a_5327_187.n10 379.457
R2812 a_5327_187.n4 a_5327_187.t13 371.139
R2813 a_5327_187.n3 a_5327_187.t14 370.613
R2814 a_5327_187.n1 a_5327_187.t11 370.613
R2815 a_5327_187.n5 a_5327_187.n4 179.837
R2816 a_5327_187.n14 a_5327_187.n13 161.352
R2817 a_5327_187.n3 a_5327_187.n2 127.096
R2818 a_5327_187.n1 a_5327_187.n0 127.096
R2819 a_5327_187.n15 a_5327_187.n11 123.481
R2820 a_5327_187.n14 a_5327_187.n12 95.095
R2821 a_5327_187.n16 a_5327_187.n15 95.094
R2822 a_5327_187.n15 a_5327_187.n14 66.258
R2823 a_5327_187.n10 a_5327_187.n9 22.578
R2824 a_5327_187.n12 a_5327_187.t1 14.282
R2825 a_5327_187.n12 a_5327_187.t3 14.282
R2826 a_5327_187.n13 a_5327_187.t0 14.282
R2827 a_5327_187.n13 a_5327_187.t2 14.282
R2828 a_5327_187.t5 a_5327_187.n16 14.282
R2829 a_5327_187.n16 a_5327_187.t4 14.282
R2830 a_5327_187.n6 a_5327_187.n5 12.222
R2831 a_5327_187.n7 a_5327_187.n1 10.046
R2832 a_5327_187.n10 a_5327_187.n8 8.58
R2833 a_5327_187.n6 a_5327_187.n3 4.65
R2834 a_5327_187.n11 a_5327_187.n7 4.65
R2835 a_5327_187.n7 a_5327_187.n6 4.035
R2836 CLK.n14 CLK.t1 459.505
R2837 CLK.n11 CLK.t14 459.505
R2838 CLK.n8 CLK.t11 459.505
R2839 CLK.n5 CLK.t12 459.505
R2840 CLK.n2 CLK.t2 459.505
R2841 CLK.n0 CLK.t3 459.505
R2842 CLK.n15 CLK.t10 399.181
R2843 CLK.n12 CLK.t17 399.181
R2844 CLK.n9 CLK.t13 399.181
R2845 CLK.n6 CLK.t6 399.181
R2846 CLK.n3 CLK.t5 399.181
R2847 CLK.n1 CLK.t15 399.181
R2848 CLK.n14 CLK.t7 384.527
R2849 CLK.n11 CLK.t4 384.527
R2850 CLK.n8 CLK.t16 384.527
R2851 CLK.n5 CLK.t0 384.527
R2852 CLK.n2 CLK.t8 384.527
R2853 CLK.n0 CLK.t9 384.527
R2854 CLK.n15 CLK.n14 33.832
R2855 CLK.n1 CLK.n0 33.832
R2856 CLK.n3 CLK.n2 33.832
R2857 CLK.n6 CLK.n5 33.832
R2858 CLK.n9 CLK.n8 33.832
R2859 CLK.n12 CLK.n11 33.832
R2860 CLK.n4 CLK.n1 11.555
R2861 CLK.n7 CLK.n4 9.476
R2862 CLK.n10 CLK.n7 9.476
R2863 CLK.n13 CLK.n10 9.476
R2864 CLK.n16 CLK.n13 9.476
R2865 CLK.n4 CLK.n3 2.079
R2866 CLK.n7 CLK.n6 2.079
R2867 CLK.n10 CLK.n9 2.079
R2868 CLK.n13 CLK.n12 2.079
R2869 CLK.n16 CLK.n15 2.079
R2870 CLK.n16 CLK 0.046
R2871 a_2141_1050.n1 a_2141_1050.t5 512.525
R2872 a_2141_1050.n1 a_2141_1050.t6 371.139
R2873 a_2141_1050.n2 a_2141_1050.t7 361.392
R2874 a_2141_1050.n4 a_2141_1050.n3 327.32
R2875 a_2141_1050.n2 a_2141_1050.n1 235.554
R2876 a_2141_1050.n5 a_2141_1050.n4 159.999
R2877 a_2141_1050.n6 a_2141_1050.n5 157.963
R2878 a_2141_1050.n5 a_2141_1050.n0 91.706
R2879 a_2141_1050.n0 a_2141_1050.t1 14.282
R2880 a_2141_1050.n0 a_2141_1050.t0 14.282
R2881 a_2141_1050.t4 a_2141_1050.n6 14.282
R2882 a_2141_1050.n6 a_2141_1050.t3 14.282
R2883 a_2141_1050.n4 a_2141_1050.n2 10.615
R2884 a_9009_1050.n1 a_9009_1050.t8 480.392
R2885 a_9009_1050.n1 a_9009_1050.t7 403.272
R2886 a_9009_1050.n2 a_9009_1050.t9 385.063
R2887 a_9009_1050.n4 a_9009_1050.n3 357.814
R2888 a_9009_1050.n7 a_9009_1050.n6 161.352
R2889 a_9009_1050.n5 a_9009_1050.n4 151.34
R2890 a_9009_1050.n2 a_9009_1050.n1 143.429
R2891 a_9009_1050.n5 a_9009_1050.n0 95.095
R2892 a_9009_1050.n8 a_9009_1050.n7 95.094
R2893 a_9009_1050.n7 a_9009_1050.n5 66.258
R2894 a_9009_1050.n0 a_9009_1050.t5 14.282
R2895 a_9009_1050.n0 a_9009_1050.t6 14.282
R2896 a_9009_1050.n6 a_9009_1050.t0 14.282
R2897 a_9009_1050.n6 a_9009_1050.t1 14.282
R2898 a_9009_1050.t3 a_9009_1050.n8 14.282
R2899 a_9009_1050.n8 a_9009_1050.t2 14.282
R2900 a_9009_1050.n4 a_9009_1050.n2 10.615
R2901 a_9331_989.n2 a_9331_989.t9 512.525
R2902 a_9331_989.n0 a_9331_989.t12 477.179
R2903 a_9331_989.n5 a_9331_989.t10 454.685
R2904 a_9331_989.n1 a_9331_989.t7 440.954
R2905 a_9331_989.n5 a_9331_989.t5 428.979
R2906 a_9331_989.n0 a_9331_989.t8 406.485
R2907 a_9331_989.n2 a_9331_989.t6 371.139
R2908 a_9331_989.n4 a_9331_989.t11 322.918
R2909 a_9331_989.n6 a_9331_989.t13 283.824
R2910 a_9331_989.n12 a_9331_989.n11 277.722
R2911 a_9331_989.n6 a_9331_989.n5 199.147
R2912 a_9331_989.n14 a_9331_989.n12 187.858
R2913 a_9331_989.n14 a_9331_989.n13 157.964
R2914 a_9331_989.n4 a_9331_989.n3 111.608
R2915 a_9331_989.n15 a_9331_989.n14 91.705
R2916 a_9331_989.n3 a_9331_989.n2 77.972
R2917 a_9331_989.n11 a_9331_989.n10 30
R2918 a_9331_989.n7 a_9331_989.n4 24.737
R2919 a_9331_989.n9 a_9331_989.n8 24.383
R2920 a_9331_989.n11 a_9331_989.n9 23.684
R2921 a_9331_989.n1 a_9331_989.n0 21.4
R2922 a_9331_989.n13 a_9331_989.t3 14.282
R2923 a_9331_989.n13 a_9331_989.t4 14.282
R2924 a_9331_989.n15 a_9331_989.t1 14.282
R2925 a_9331_989.t2 a_9331_989.n15 14.282
R2926 a_9331_989.n7 a_9331_989.n6 7.597
R2927 a_9331_989.n3 a_9331_989.n1 6.833
R2928 a_9331_989.n12 a_9331_989.n7 4.65
R2929 a_147_187.n4 a_147_187.t15 512.525
R2930 a_147_187.n2 a_147_187.t9 472.359
R2931 a_147_187.n0 a_147_187.t14 472.359
R2932 a_147_187.n5 a_147_187.t12 417.109
R2933 a_147_187.n2 a_147_187.t13 384.527
R2934 a_147_187.n0 a_147_187.t10 384.527
R2935 a_147_187.n4 a_147_187.t11 371.139
R2936 a_147_187.n3 a_147_187.t8 370.613
R2937 a_147_187.n1 a_147_187.t7 370.613
R2938 a_147_187.n12 a_147_187.n11 363.934
R2939 a_147_187.n5 a_147_187.n4 179.837
R2940 a_147_187.n15 a_147_187.n14 161.352
R2941 a_147_187.n3 a_147_187.n2 127.096
R2942 a_147_187.n1 a_147_187.n0 127.096
R2943 a_147_187.n16 a_147_187.n12 123.481
R2944 a_147_187.n15 a_147_187.n13 95.095
R2945 a_147_187.n17 a_147_187.n16 95.094
R2946 a_147_187.n16 a_147_187.n15 66.258
R2947 a_147_187.n11 a_147_187.n10 30
R2948 a_147_187.n9 a_147_187.n8 24.383
R2949 a_147_187.n11 a_147_187.n9 23.684
R2950 a_147_187.n13 a_147_187.t5 14.282
R2951 a_147_187.n13 a_147_187.t6 14.282
R2952 a_147_187.n14 a_147_187.t4 14.282
R2953 a_147_187.n14 a_147_187.t3 14.282
R2954 a_147_187.n17 a_147_187.t1 14.282
R2955 a_147_187.t2 a_147_187.n17 14.282
R2956 a_147_187.n6 a_147_187.n5 12.222
R2957 a_147_187.n7 a_147_187.n1 10.046
R2958 a_147_187.n6 a_147_187.n3 4.65
R2959 a_147_187.n12 a_147_187.n7 4.65
R2960 a_147_187.n7 a_147_187.n6 4.035
R2961 a_4626_101.n5 a_4626_101.n4 62.817
R2962 a_4626_101.n2 a_4626_101.n0 41.528
R2963 a_4626_101.n5 a_4626_101.n3 26.202
R2964 a_4626_101.t0 a_4626_101.n5 19.737
R2965 a_4626_101.t0 a_4626_101.n6 8.137
R2966 a_4626_101.n2 a_4626_101.n1 3.644
R2967 a_4626_101.t0 a_4626_101.n2 1.093
R2968 a_4151_989.n1 a_4151_989.t11 512.525
R2969 a_4151_989.n0 a_4151_989.t7 512.525
R2970 a_4151_989.n5 a_4151_989.t5 454.685
R2971 a_4151_989.n5 a_4151_989.t8 428.979
R2972 a_4151_989.n1 a_4151_989.t6 371.139
R2973 a_4151_989.n0 a_4151_989.t12 371.139
R2974 a_4151_989.n2 a_4151_989.n1 343.521
R2975 a_4151_989.n4 a_4151_989.n0 287.803
R2976 a_4151_989.n9 a_4151_989.n8 271.602
R2977 a_4151_989.n6 a_4151_989.t9 244.718
R2978 a_4151_989.n6 a_4151_989.n5 227.006
R2979 a_4151_989.n11 a_4151_989.n9 215.717
R2980 a_4151_989.n2 a_4151_989.t13 172.106
R2981 a_4151_989.n3 a_4151_989.t10 165.68
R2982 a_4151_989.n11 a_4151_989.n10 157.964
R2983 a_4151_989.n12 a_4151_989.n11 91.705
R2984 a_4151_989.n4 a_4151_989.n3 55.717
R2985 a_4151_989.n7 a_4151_989.n4 47.59
R2986 a_4151_989.n10 a_4151_989.t0 14.282
R2987 a_4151_989.n10 a_4151_989.t1 14.282
R2988 a_4151_989.n12 a_4151_989.t2 14.282
R2989 a_4151_989.t3 a_4151_989.n12 14.282
R2990 a_4151_989.n3 a_4151_989.n2 10.343
R2991 a_4151_989.n7 a_4151_989.n6 7.597
R2992 a_4151_989.n9 a_4151_989.n7 4.65
R2993 a_1053_103.t0 a_1053_103.n7 59.616
R2994 a_1053_103.n4 a_1053_103.n2 54.496
R2995 a_1053_103.n4 a_1053_103.n3 54.496
R2996 a_1053_103.n1 a_1053_103.n0 24.679
R2997 a_1053_103.n6 a_1053_103.n4 7.859
R2998 a_1053_103.t0 a_1053_103.n1 7.505
R2999 a_1053_103.t0 a_1053_103.n6 3.034
R3000 a_1053_103.n6 a_1053_103.n5 0.443
R3001 a_1334_210.n10 a_1334_210.n8 171.558
R3002 a_1334_210.n8 a_1334_210.t1 75.764
R3003 a_1334_210.n11 a_1334_210.n0 49.6
R3004 a_1334_210.n3 a_1334_210.n2 27.476
R3005 a_1334_210.n10 a_1334_210.n9 27.2
R3006 a_1334_210.n11 a_1334_210.n10 22.4
R3007 a_1334_210.t1 a_1334_210.n5 20.241
R3008 a_1334_210.n7 a_1334_210.n6 19.952
R3009 a_1334_210.t1 a_1334_210.n3 13.984
R3010 a_1334_210.n5 a_1334_210.n4 13.494
R3011 a_1334_210.t1 a_1334_210.n1 7.04
R3012 a_1334_210.n8 a_1334_210.n7 1.505
R3013 a_277_1050.n2 a_277_1050.t8 512.525
R3014 a_277_1050.n0 a_277_1050.t7 512.525
R3015 a_277_1050.n3 a_277_1050.t12 389.251
R3016 a_277_1050.n1 a_277_1050.t11 389.251
R3017 a_277_1050.n2 a_277_1050.t10 371.139
R3018 a_277_1050.n0 a_277_1050.t9 371.139
R3019 a_277_1050.n9 a_277_1050.n8 336.075
R3020 a_277_1050.n3 a_277_1050.n2 207.695
R3021 a_277_1050.n1 a_277_1050.n0 207.695
R3022 a_277_1050.n12 a_277_1050.n11 161.352
R3023 a_277_1050.n13 a_277_1050.n9 151.34
R3024 a_277_1050.n12 a_277_1050.n10 95.095
R3025 a_277_1050.n14 a_277_1050.n13 95.094
R3026 a_277_1050.n13 a_277_1050.n12 66.258
R3027 a_277_1050.n8 a_277_1050.n7 30
R3028 a_277_1050.n6 a_277_1050.n5 24.383
R3029 a_277_1050.n8 a_277_1050.n6 23.684
R3030 a_277_1050.n10 a_277_1050.t6 14.282
R3031 a_277_1050.n10 a_277_1050.t5 14.282
R3032 a_277_1050.n11 a_277_1050.t3 14.282
R3033 a_277_1050.n11 a_277_1050.t4 14.282
R3034 a_277_1050.t2 a_277_1050.n14 14.282
R3035 a_277_1050.n14 a_277_1050.t1 14.282
R3036 a_277_1050.n4 a_277_1050.n1 14.126
R3037 a_277_1050.n9 a_277_1050.n4 5.965
R3038 a_277_1050.n4 a_277_1050.n3 4.65
R3039 a_5457_1050.n4 a_5457_1050.t7 512.525
R3040 a_5457_1050.n2 a_5457_1050.t8 512.525
R3041 a_5457_1050.n5 a_5457_1050.t11 389.251
R3042 a_5457_1050.n3 a_5457_1050.t10 389.251
R3043 a_5457_1050.n4 a_5457_1050.t12 371.139
R3044 a_5457_1050.n2 a_5457_1050.t9 371.139
R3045 a_5457_1050.n8 a_5457_1050.n7 357.814
R3046 a_5457_1050.n5 a_5457_1050.n4 207.695
R3047 a_5457_1050.n3 a_5457_1050.n2 207.695
R3048 a_5457_1050.n11 a_5457_1050.n10 161.352
R3049 a_5457_1050.n9 a_5457_1050.n8 151.34
R3050 a_5457_1050.n9 a_5457_1050.n1 95.095
R3051 a_5457_1050.n10 a_5457_1050.n0 95.095
R3052 a_5457_1050.n10 a_5457_1050.n9 66.258
R3053 a_5457_1050.n1 a_5457_1050.t0 14.282
R3054 a_5457_1050.n1 a_5457_1050.t2 14.282
R3055 a_5457_1050.n0 a_5457_1050.t6 14.282
R3056 a_5457_1050.n0 a_5457_1050.t5 14.282
R3057 a_5457_1050.t4 a_5457_1050.n11 14.282
R3058 a_5457_1050.n11 a_5457_1050.t3 14.282
R3059 a_5457_1050.n6 a_5457_1050.n3 14.126
R3060 a_5457_1050.n8 a_5457_1050.n6 5.965
R3061 a_5457_1050.n6 a_5457_1050.n5 4.65
R3062 a_5779_989.n1 a_5779_989.t11 480.392
R3063 a_5779_989.n3 a_5779_989.t12 454.685
R3064 a_5779_989.n3 a_5779_989.t10 428.979
R3065 a_5779_989.n1 a_5779_989.t9 403.272
R3066 a_5779_989.n2 a_5779_989.t8 357.204
R3067 a_5779_989.n4 a_5779_989.t7 311.683
R3068 a_5779_989.n10 a_5779_989.n9 308.216
R3069 a_5779_989.n11 a_5779_989.n10 179.199
R3070 a_5779_989.n4 a_5779_989.n3 171.288
R3071 a_5779_989.n2 a_5779_989.n1 171.288
R3072 a_5779_989.n13 a_5779_989.n12 161.352
R3073 a_5779_989.n11 a_5779_989.n0 95.095
R3074 a_5779_989.n14 a_5779_989.n13 95.094
R3075 a_5779_989.n13 a_5779_989.n11 66.258
R3076 a_5779_989.n9 a_5779_989.n8 30
R3077 a_5779_989.n7 a_5779_989.n6 24.383
R3078 a_5779_989.n9 a_5779_989.n7 23.684
R3079 a_5779_989.n0 a_5779_989.t3 14.282
R3080 a_5779_989.n0 a_5779_989.t2 14.282
R3081 a_5779_989.n12 a_5779_989.t6 14.282
R3082 a_5779_989.n12 a_5779_989.t5 14.282
R3083 a_5779_989.t1 a_5779_989.n14 14.282
R3084 a_5779_989.n14 a_5779_989.t0 14.282
R3085 a_5779_989.n5 a_5779_989.n4 8.685
R3086 a_5779_989.n5 a_5779_989.n2 5.965
R3087 a_5779_989.n10 a_5779_989.n5 4.65
R3088 a_12396_101.n3 a_12396_101.n1 42.788
R3089 a_12396_101.t0 a_12396_101.n0 8.137
R3090 a_12396_101.n3 a_12396_101.n2 4.665
R3091 a_12396_101.t0 a_12396_101.n3 0.06
R3092 a_3829_1050.n1 a_3829_1050.t9 480.392
R3093 a_3829_1050.n1 a_3829_1050.t7 403.272
R3094 a_3829_1050.n2 a_3829_1050.t8 385.063
R3095 a_3829_1050.n7 a_3829_1050.n6 336.075
R3096 a_3829_1050.n10 a_3829_1050.n9 161.352
R3097 a_3829_1050.n8 a_3829_1050.n7 151.34
R3098 a_3829_1050.n2 a_3829_1050.n1 143.429
R3099 a_3829_1050.n8 a_3829_1050.n0 95.095
R3100 a_3829_1050.n11 a_3829_1050.n10 95.094
R3101 a_3829_1050.n10 a_3829_1050.n8 66.258
R3102 a_3829_1050.n6 a_3829_1050.n5 30
R3103 a_3829_1050.n4 a_3829_1050.n3 24.383
R3104 a_3829_1050.n6 a_3829_1050.n4 23.684
R3105 a_3829_1050.n0 a_3829_1050.t5 14.282
R3106 a_3829_1050.n0 a_3829_1050.t6 14.282
R3107 a_3829_1050.n9 a_3829_1050.t3 14.282
R3108 a_3829_1050.n9 a_3829_1050.t2 14.282
R3109 a_3829_1050.t1 a_3829_1050.n11 14.282
R3110 a_3829_1050.n11 a_3829_1050.t0 14.282
R3111 a_3829_1050.n7 a_3829_1050.n2 10.615
R3112 a_2036_101.n11 a_2036_101.n10 68.43
R3113 a_2036_101.n3 a_2036_101.n2 62.817
R3114 a_2036_101.n7 a_2036_101.n6 38.626
R3115 a_2036_101.n6 a_2036_101.n5 35.955
R3116 a_2036_101.n3 a_2036_101.n1 26.202
R3117 a_2036_101.t0 a_2036_101.n3 19.737
R3118 a_2036_101.t1 a_2036_101.n8 8.137
R3119 a_2036_101.t0 a_2036_101.n4 7.273
R3120 a_2036_101.t0 a_2036_101.n0 6.109
R3121 a_2036_101.t1 a_2036_101.n7 4.864
R3122 a_2036_101.t0 a_2036_101.n12 2.074
R3123 a_2036_101.n12 a_2036_101.t1 0.937
R3124 a_2036_101.t1 a_2036_101.n11 0.763
R3125 a_2036_101.n11 a_2036_101.n9 0.185
R3126 a_10451_103.n5 a_10451_103.n4 66.708
R3127 a_10451_103.n2 a_10451_103.n0 32.662
R3128 a_10451_103.n5 a_10451_103.n3 19.496
R3129 a_10451_103.t0 a_10451_103.n5 13.756
R3130 a_10451_103.t0 a_10451_103.n2 3.034
R3131 a_10451_103.n2 a_10451_103.n1 0.443
R3132 a_15757_1051.n4 a_15757_1051.t0 179.895
R3133 a_15757_1051.n2 a_15757_1051.n1 157.021
R3134 a_15757_1051.n2 a_15757_1051.n0 124.955
R3135 a_15757_1051.n4 a_15757_1051.n3 106.183
R3136 a_15757_1051.n5 a_15757_1051.n4 99.358
R3137 a_15757_1051.n3 a_15757_1051.n2 82.65
R3138 a_15757_1051.n3 a_15757_1051.t7 73.712
R3139 a_15757_1051.n0 a_15757_1051.t3 14.282
R3140 a_15757_1051.n0 a_15757_1051.t2 14.282
R3141 a_15757_1051.n1 a_15757_1051.t4 14.282
R3142 a_15757_1051.n1 a_15757_1051.t5 14.282
R3143 a_15757_1051.t1 a_15757_1051.n5 14.282
R3144 a_15757_1051.n5 a_15757_1051.t6 14.282
R3145 a_15652_101.n4 a_15652_101.n2 41.528
R3146 a_15652_101.n1 a_15652_101.n0 33.123
R3147 a_15652_101.t0 a_15652_101.n1 10.642
R3148 a_15652_101.n6 a_15652_101.n5 7.966
R3149 a_15652_101.n4 a_15652_101.n3 3.644
R3150 a_15652_101.t0 a_15652_101.n4 1.093
R3151 a_15652_101.t0 a_15652_101.n6 0.088
R3152 a_6514_210.n10 a_6514_210.n8 171.558
R3153 a_6514_210.n8 a_6514_210.t1 75.764
R3154 a_6514_210.n3 a_6514_210.n2 27.476
R3155 a_6514_210.n10 a_6514_210.n9 27.2
R3156 a_6514_210.n11 a_6514_210.n0 23.498
R3157 a_6514_210.n11 a_6514_210.n10 22.4
R3158 a_6514_210.t1 a_6514_210.n5 20.241
R3159 a_6514_210.n7 a_6514_210.n6 19.952
R3160 a_6514_210.t1 a_6514_210.n3 13.984
R3161 a_6514_210.n5 a_6514_210.n4 13.494
R3162 a_6514_210.t1 a_6514_210.n1 7.04
R3163 a_6514_210.n8 a_6514_210.n7 1.505
R3164 a_11694_210.n10 a_11694_210.n8 171.558
R3165 a_11694_210.n8 a_11694_210.t1 75.764
R3166 a_11694_210.n11 a_11694_210.n0 49.6
R3167 a_11694_210.n3 a_11694_210.n2 27.476
R3168 a_11694_210.n10 a_11694_210.n9 27.2
R3169 a_11694_210.n11 a_11694_210.n10 22.4
R3170 a_11694_210.t1 a_11694_210.n5 20.241
R3171 a_11694_210.n7 a_11694_210.n6 19.952
R3172 a_11694_210.t1 a_11694_210.n3 13.984
R3173 a_11694_210.n5 a_11694_210.n4 13.494
R3174 a_11694_210.t1 a_11694_210.n1 7.04
R3175 a_11694_210.n8 a_11694_210.n7 1.505
R3176 a_14986_101.n11 a_14986_101.n10 68.43
R3177 a_14986_101.n3 a_14986_101.n2 62.817
R3178 a_14986_101.n7 a_14986_101.n6 38.626
R3179 a_14986_101.n6 a_14986_101.n5 35.955
R3180 a_14986_101.n3 a_14986_101.n1 26.202
R3181 a_14986_101.t0 a_14986_101.n3 19.737
R3182 a_14986_101.t1 a_14986_101.n8 8.137
R3183 a_14986_101.t0 a_14986_101.n4 7.273
R3184 a_14986_101.t0 a_14986_101.n0 6.109
R3185 a_14986_101.t1 a_14986_101.n7 4.864
R3186 a_14986_101.t0 a_14986_101.n12 2.074
R3187 a_14986_101.n12 a_14986_101.t1 0.937
R3188 a_14986_101.t1 a_14986_101.n11 0.763
R3189 a_14986_101.n11 a_14986_101.n9 0.185
R3190 a_12501_1050.n0 a_12501_1050.t7 512.525
R3191 a_12501_1050.n0 a_12501_1050.t5 371.139
R3192 a_12501_1050.n1 a_12501_1050.t6 361.392
R3193 a_12501_1050.n3 a_12501_1050.n2 327.32
R3194 a_12501_1050.n1 a_12501_1050.n0 235.554
R3195 a_12501_1050.n5 a_12501_1050.n3 159.999
R3196 a_12501_1050.n5 a_12501_1050.n4 157.964
R3197 a_12501_1050.n6 a_12501_1050.n5 91.705
R3198 a_12501_1050.n4 a_12501_1050.t4 14.282
R3199 a_12501_1050.n4 a_12501_1050.t3 14.282
R3200 a_12501_1050.t1 a_12501_1050.n6 14.282
R3201 a_12501_1050.n6 a_12501_1050.t0 14.282
R3202 a_12501_1050.n3 a_12501_1050.n1 10.615
R3203 a_7321_1050.n1 a_7321_1050.t5 512.525
R3204 a_7321_1050.n1 a_7321_1050.t7 371.139
R3205 a_7321_1050.n2 a_7321_1050.t6 361.392
R3206 a_7321_1050.n7 a_7321_1050.n6 305.581
R3207 a_7321_1050.n2 a_7321_1050.n1 235.554
R3208 a_7321_1050.n8 a_7321_1050.n7 159.999
R3209 a_7321_1050.n9 a_7321_1050.n8 157.963
R3210 a_7321_1050.n8 a_7321_1050.n0 91.706
R3211 a_7321_1050.n6 a_7321_1050.n5 30
R3212 a_7321_1050.n4 a_7321_1050.n3 24.383
R3213 a_7321_1050.n6 a_7321_1050.n4 23.684
R3214 a_7321_1050.n0 a_7321_1050.t2 14.282
R3215 a_7321_1050.n0 a_7321_1050.t3 14.282
R3216 a_7321_1050.n9 a_7321_1050.t0 14.282
R3217 a_7321_1050.t1 a_7321_1050.n9 14.282
R3218 a_7321_1050.n7 a_7321_1050.n2 10.615
R3219 a_8823_103.t0 a_8823_103.n7 59.616
R3220 a_8823_103.n4 a_8823_103.n2 54.496
R3221 a_8823_103.n4 a_8823_103.n3 54.496
R3222 a_8823_103.n1 a_8823_103.n0 24.679
R3223 a_8823_103.n6 a_8823_103.n4 7.859
R3224 a_8823_103.t0 a_8823_103.n1 7.505
R3225 a_8823_103.t0 a_8823_103.n6 3.034
R3226 a_8823_103.n6 a_8823_103.n5 0.443
R3227 a_9104_210.n10 a_9104_210.n8 171.558
R3228 a_9104_210.n8 a_9104_210.t1 75.764
R3229 a_9104_210.n11 a_9104_210.n0 49.6
R3230 a_9104_210.n3 a_9104_210.n2 27.476
R3231 a_9104_210.n10 a_9104_210.n9 27.2
R3232 a_9104_210.n11 a_9104_210.n10 22.4
R3233 a_9104_210.t1 a_9104_210.n5 20.241
R3234 a_9104_210.n7 a_9104_210.n6 19.952
R3235 a_9104_210.t1 a_9104_210.n3 13.984
R3236 a_9104_210.n5 a_9104_210.n4 13.494
R3237 a_9104_210.t1 a_9104_210.n1 7.04
R3238 a_9104_210.n8 a_9104_210.n7 1.505
R3239 a_16318_101.n2 a_16318_101.n0 42.755
R3240 a_16318_101.n2 a_16318_101.n1 2.198
R3241 a_16318_101.t0 a_16318_101.n2 0.106
R3242 a_372_210.n9 a_372_210.n7 171.558
R3243 a_372_210.t0 a_372_210.n9 75.765
R3244 a_372_210.n3 a_372_210.n1 74.827
R3245 a_372_210.n3 a_372_210.n2 27.476
R3246 a_372_210.n7 a_372_210.n6 27.2
R3247 a_372_210.n5 a_372_210.n4 23.498
R3248 a_372_210.n7 a_372_210.n5 22.4
R3249 a_372_210.t0 a_372_210.n11 20.241
R3250 a_372_210.t0 a_372_210.n3 13.984
R3251 a_372_210.n11 a_372_210.n10 13.494
R3252 a_372_210.t0 a_372_210.n0 8.137
R3253 a_372_210.n9 a_372_210.n8 1.505
R3254 a_10732_210.n8 a_10732_210.n6 185.173
R3255 a_10732_210.t0 a_10732_210.n8 75.765
R3256 a_10732_210.n3 a_10732_210.n1 74.827
R3257 a_10732_210.n3 a_10732_210.n2 27.476
R3258 a_10732_210.n6 a_10732_210.n5 22.349
R3259 a_10732_210.t0 a_10732_210.n10 20.241
R3260 a_10732_210.t0 a_10732_210.n3 13.984
R3261 a_10732_210.n10 a_10732_210.n9 13.494
R3262 a_10732_210.n6 a_10732_210.n4 8.443
R3263 a_10732_210.t0 a_10732_210.n0 8.137
R3264 a_10732_210.n8 a_10732_210.n7 1.505
R3265 a_6233_103.t0 a_6233_103.n7 59.616
R3266 a_6233_103.n4 a_6233_103.n2 54.496
R3267 a_6233_103.n4 a_6233_103.n3 54.496
R3268 a_6233_103.n1 a_6233_103.n0 24.679
R3269 a_6233_103.t0 a_6233_103.n1 7.505
R3270 a_6233_103.n6 a_6233_103.n5 2.455
R3271 a_6233_103.n6 a_6233_103.n4 0.636
R3272 a_6233_103.t0 a_6233_103.n6 0.246
R3273 a_5552_210.n9 a_5552_210.n7 171.558
R3274 a_5552_210.t0 a_5552_210.n9 75.765
R3275 a_5552_210.n3 a_5552_210.n1 74.827
R3276 a_5552_210.n3 a_5552_210.n2 27.476
R3277 a_5552_210.n7 a_5552_210.n6 27.2
R3278 a_5552_210.n5 a_5552_210.n4 23.498
R3279 a_5552_210.n7 a_5552_210.n5 22.4
R3280 a_5552_210.t0 a_5552_210.n11 20.241
R3281 a_5552_210.t0 a_5552_210.n3 13.984
R3282 a_5552_210.n11 a_5552_210.n10 13.494
R3283 a_5552_210.t0 a_5552_210.n0 8.137
R3284 a_5552_210.n9 a_5552_210.n8 1.505
R3285 a_16984_101.n3 a_16984_101.n1 42.788
R3286 a_16984_101.t0 a_16984_101.n0 8.137
R3287 a_16984_101.n3 a_16984_101.n2 4.665
R3288 a_16984_101.t0 a_16984_101.n3 0.06
R3289 a_2962_210.n9 a_2962_210.n7 171.558
R3290 a_2962_210.t0 a_2962_210.n9 75.765
R3291 a_2962_210.n3 a_2962_210.n1 74.827
R3292 a_2962_210.n3 a_2962_210.n2 27.476
R3293 a_2962_210.n7 a_2962_210.n6 27.2
R3294 a_2962_210.n5 a_2962_210.n4 23.498
R3295 a_2962_210.n7 a_2962_210.n5 22.4
R3296 a_2962_210.t0 a_2962_210.n11 20.241
R3297 a_2962_210.t0 a_2962_210.n3 13.984
R3298 a_2962_210.n11 a_2962_210.n10 13.494
R3299 a_2962_210.t0 a_2962_210.n0 8.137
R3300 a_2962_210.n9 a_2962_210.n8 1.505
R3301 a_7861_103.n5 a_7861_103.n4 66.708
R3302 a_7861_103.n2 a_7861_103.n0 25.439
R3303 a_7861_103.n5 a_7861_103.n3 19.496
R3304 a_7861_103.t0 a_7861_103.n5 13.756
R3305 a_7861_103.n2 a_7861_103.n1 2.455
R3306 a_7861_103.t0 a_7861_103.n2 0.246
R3307 Q.n2 Q.n1 349.908
R3308 Q.n2 Q.n0 215.564
R3309 Q.n0 Q.t1 14.282
R3310 Q.n0 Q.t0 14.282
R3311 Q.n3 Q.n2 4.65
R3312 Q.n3 Q 0.046
R3313 a_9806_101.n3 a_9806_101.n1 42.788
R3314 a_9806_101.t0 a_9806_101.n0 8.137
R3315 a_9806_101.n3 a_9806_101.n2 4.665
R3316 a_9806_101.t0 a_9806_101.n3 0.06
R3317 a_7216_101.n11 a_7216_101.n10 68.43
R3318 a_7216_101.n3 a_7216_101.n2 62.817
R3319 a_7216_101.n7 a_7216_101.n6 38.626
R3320 a_7216_101.n6 a_7216_101.n5 35.955
R3321 a_7216_101.n3 a_7216_101.n1 26.202
R3322 a_7216_101.t0 a_7216_101.n3 19.737
R3323 a_7216_101.t1 a_7216_101.n8 8.137
R3324 a_7216_101.t0 a_7216_101.n4 7.273
R3325 a_7216_101.t0 a_7216_101.n0 6.109
R3326 a_7216_101.t1 a_7216_101.n7 4.864
R3327 a_7216_101.t0 a_7216_101.n12 2.074
R3328 a_7216_101.n12 a_7216_101.t1 0.937
R3329 a_7216_101.t1 a_7216_101.n11 0.763
R3330 a_7216_101.n11 a_7216_101.n9 0.185
R3331 a_91_103.n5 a_91_103.n4 66.708
R3332 a_91_103.n2 a_91_103.n0 25.439
R3333 a_91_103.n5 a_91_103.n3 19.496
R3334 a_91_103.t0 a_91_103.n5 13.756
R3335 a_91_103.n2 a_91_103.n1 2.455
R3336 a_91_103.t0 a_91_103.n2 0.246
R3337 a_5271_103.n5 a_5271_103.n4 66.708
R3338 a_5271_103.n2 a_5271_103.n0 25.439
R3339 a_5271_103.n5 a_5271_103.n3 19.496
R3340 a_5271_103.t0 a_5271_103.n5 13.756
R3341 a_5271_103.n2 a_5271_103.n1 2.455
R3342 a_5271_103.t0 a_5271_103.n2 0.246
R3343 a_3924_210.n10 a_3924_210.n8 171.558
R3344 a_3924_210.n8 a_3924_210.t1 75.764
R3345 a_3924_210.n3 a_3924_210.n2 27.476
R3346 a_3924_210.n10 a_3924_210.n9 27.2
R3347 a_3924_210.n11 a_3924_210.n0 23.498
R3348 a_3924_210.n11 a_3924_210.n10 22.4
R3349 a_3924_210.t1 a_3924_210.n5 20.241
R3350 a_3924_210.n7 a_3924_210.n6 19.952
R3351 a_3924_210.t1 a_3924_210.n3 13.984
R3352 a_3924_210.n5 a_3924_210.n4 13.494
R3353 a_3924_210.t1 a_3924_210.n1 7.04
R3354 a_3924_210.n8 a_3924_210.n7 1.505
R3355 a_13322_210.n9 a_13322_210.n7 171.558
R3356 a_13322_210.t0 a_13322_210.n9 75.765
R3357 a_13322_210.n3 a_13322_210.n1 74.827
R3358 a_13322_210.n3 a_13322_210.n2 27.476
R3359 a_13322_210.n7 a_13322_210.n6 27.2
R3360 a_13322_210.n5 a_13322_210.n4 23.498
R3361 a_13322_210.n7 a_13322_210.n5 22.4
R3362 a_13322_210.t0 a_13322_210.n11 20.241
R3363 a_13322_210.t0 a_13322_210.n3 13.984
R3364 a_13322_210.n11 a_13322_210.n10 13.494
R3365 a_13322_210.t0 a_13322_210.n0 8.137
R3366 a_13322_210.n9 a_13322_210.n8 1.505
R3367 a_14284_210.n10 a_14284_210.n8 171.558
R3368 a_14284_210.n8 a_14284_210.t1 75.764
R3369 a_14284_210.n3 a_14284_210.n2 27.476
R3370 a_14284_210.n10 a_14284_210.n9 27.2
R3371 a_14284_210.n11 a_14284_210.n0 23.498
R3372 a_14284_210.n11 a_14284_210.n10 22.4
R3373 a_14284_210.t1 a_14284_210.n5 20.241
R3374 a_14284_210.n7 a_14284_210.n6 19.952
R3375 a_14284_210.t1 a_14284_210.n3 13.984
R3376 a_14284_210.n5 a_14284_210.n4 13.494
R3377 a_14284_210.t1 a_14284_210.n1 7.04
R3378 a_14284_210.n8 a_14284_210.n7 1.505
R3379 a_13041_103.n5 a_13041_103.n4 66.708
R3380 a_13041_103.n2 a_13041_103.n0 25.439
R3381 a_13041_103.n5 a_13041_103.n3 19.496
R3382 a_13041_103.t0 a_13041_103.n5 13.756
R3383 a_13041_103.n2 a_13041_103.n1 2.455
R3384 a_13041_103.t0 a_13041_103.n2 0.246
R3385 a_3643_103.t0 a_3643_103.n7 59.616
R3386 a_3643_103.n4 a_3643_103.n2 54.496
R3387 a_3643_103.n4 a_3643_103.n3 54.496
R3388 a_3643_103.n1 a_3643_103.n0 24.679
R3389 a_3643_103.t0 a_3643_103.n1 7.505
R3390 a_3643_103.n6 a_3643_103.n5 2.455
R3391 a_3643_103.n6 a_3643_103.n4 0.636
R3392 a_3643_103.t0 a_3643_103.n6 0.246
R3393 a_14003_103.n5 a_14003_103.n4 66.708
R3394 a_14003_103.n2 a_14003_103.n0 25.439
R3395 a_14003_103.n5 a_14003_103.n3 19.496
R3396 a_14003_103.t0 a_14003_103.n5 13.756
R3397 a_14003_103.n2 a_14003_103.n1 2.455
R3398 a_14003_103.t0 a_14003_103.n2 0.246
R3399 a_2681_103.n5 a_2681_103.n4 66.708
R3400 a_2681_103.n2 a_2681_103.n0 25.439
R3401 a_2681_103.n5 a_2681_103.n3 19.496
R3402 a_2681_103.t0 a_2681_103.n5 13.756
R3403 a_2681_103.n2 a_2681_103.n1 2.455
R3404 a_2681_103.t0 a_2681_103.n2 0.246
C7 RN GND 7.36fF
C8 VDD GND 29.31fF
C9 a_2681_103.n0 GND 0.11fF
C10 a_2681_103.n1 GND 0.04fF
C11 a_2681_103.n2 GND 0.03fF
C12 a_2681_103.n3 GND 0.07fF
C13 a_2681_103.n4 GND 0.08fF
C14 a_2681_103.n5 GND 0.03fF
C15 a_14003_103.n0 GND 0.11fF
C16 a_14003_103.n1 GND 0.04fF
C17 a_14003_103.n2 GND 0.03fF
C18 a_14003_103.n3 GND 0.07fF
C19 a_14003_103.n4 GND 0.08fF
C20 a_14003_103.n5 GND 0.03fF
C21 a_3643_103.n0 GND 0.08fF
C22 a_3643_103.n1 GND 0.07fF
C23 a_3643_103.n2 GND 0.04fF
C24 a_3643_103.n3 GND 0.06fF
C25 a_3643_103.n4 GND 0.03fF
C26 a_3643_103.n5 GND 0.04fF
C27 a_3643_103.n7 GND 0.08fF
C28 a_13041_103.n0 GND 0.11fF
C29 a_13041_103.n1 GND 0.04fF
C30 a_13041_103.n2 GND 0.03fF
C31 a_13041_103.n3 GND 0.07fF
C32 a_13041_103.n4 GND 0.08fF
C33 a_13041_103.n5 GND 0.03fF
C34 a_14284_210.n0 GND 0.02fF
C35 a_14284_210.n1 GND 0.09fF
C36 a_14284_210.n2 GND 0.12fF
C37 a_14284_210.n3 GND 0.08fF
C38 a_14284_210.n4 GND 0.08fF
C39 a_14284_210.n5 GND 0.02fF
C40 a_14284_210.t1 GND 0.29fF
C41 a_14284_210.n6 GND 0.09fF
C42 a_14284_210.n7 GND 0.02fF
C43 a_14284_210.n8 GND 0.13fF
C44 a_14284_210.n9 GND 0.02fF
C45 a_14284_210.n10 GND 0.03fF
C46 a_14284_210.n11 GND 0.03fF
C47 a_13322_210.n0 GND 0.07fF
C48 a_13322_210.n1 GND 0.09fF
C49 a_13322_210.n2 GND 0.12fF
C50 a_13322_210.n3 GND 0.08fF
C51 a_13322_210.n4 GND 0.02fF
C52 a_13322_210.n5 GND 0.03fF
C53 a_13322_210.n6 GND 0.02fF
C54 a_13322_210.n7 GND 0.03fF
C55 a_13322_210.n8 GND 0.02fF
C56 a_13322_210.n9 GND 0.13fF
C57 a_13322_210.n10 GND 0.08fF
C58 a_13322_210.n11 GND 0.02fF
C59 a_13322_210.t0 GND 0.31fF
C60 a_3924_210.n0 GND 0.02fF
C61 a_3924_210.n1 GND 0.09fF
C62 a_3924_210.n2 GND 0.12fF
C63 a_3924_210.n3 GND 0.08fF
C64 a_3924_210.n4 GND 0.08fF
C65 a_3924_210.n5 GND 0.02fF
C66 a_3924_210.t1 GND 0.29fF
C67 a_3924_210.n6 GND 0.09fF
C68 a_3924_210.n7 GND 0.02fF
C69 a_3924_210.n8 GND 0.13fF
C70 a_3924_210.n9 GND 0.02fF
C71 a_3924_210.n10 GND 0.03fF
C72 a_3924_210.n11 GND 0.03fF
C73 a_5271_103.n0 GND 0.11fF
C74 a_5271_103.n1 GND 0.04fF
C75 a_5271_103.n2 GND 0.03fF
C76 a_5271_103.n3 GND 0.07fF
C77 a_5271_103.n4 GND 0.08fF
C78 a_5271_103.n5 GND 0.03fF
C79 a_91_103.n0 GND 0.10fF
C80 a_91_103.n1 GND 0.03fF
C81 a_91_103.n2 GND 0.03fF
C82 a_91_103.n3 GND 0.07fF
C83 a_91_103.n4 GND 0.08fF
C84 a_91_103.n5 GND 0.03fF
C85 a_7216_101.n0 GND 0.02fF
C86 a_7216_101.n1 GND 0.09fF
C87 a_7216_101.n2 GND 0.08fF
C88 a_7216_101.n3 GND 0.03fF
C89 a_7216_101.n4 GND 0.01fF
C90 a_7216_101.n5 GND 0.04fF
C91 a_7216_101.n6 GND 0.04fF
C92 a_7216_101.n7 GND 0.02fF
C93 a_7216_101.n8 GND 0.05fF
C94 a_7216_101.n9 GND 0.15fF
C95 a_7216_101.n10 GND 0.08fF
C96 a_7216_101.n11 GND 0.08fF
C97 a_7216_101.t1 GND 0.23fF
C98 a_7216_101.n12 GND 0.01fF
C99 a_9806_101.n0 GND 0.05fF
C100 a_9806_101.n1 GND 0.12fF
C101 a_9806_101.n2 GND 0.04fF
C102 a_9806_101.n3 GND 0.17fF
C103 Q.n0 GND 0.58fF
C104 Q.n1 GND 0.36fF
C105 Q.n2 GND 0.66fF
C106 Q.n3 GND 0.01fF
C107 a_7861_103.n0 GND 0.11fF
C108 a_7861_103.n1 GND 0.04fF
C109 a_7861_103.n2 GND 0.03fF
C110 a_7861_103.n3 GND 0.07fF
C111 a_7861_103.n4 GND 0.08fF
C112 a_7861_103.n5 GND 0.03fF
C113 a_2962_210.n0 GND 0.07fF
C114 a_2962_210.n1 GND 0.09fF
C115 a_2962_210.n2 GND 0.12fF
C116 a_2962_210.n3 GND 0.08fF
C117 a_2962_210.n4 GND 0.02fF
C118 a_2962_210.n5 GND 0.03fF
C119 a_2962_210.n6 GND 0.02fF
C120 a_2962_210.n7 GND 0.03fF
C121 a_2962_210.n8 GND 0.02fF
C122 a_2962_210.n9 GND 0.13fF
C123 a_2962_210.n10 GND 0.08fF
C124 a_2962_210.n11 GND 0.02fF
C125 a_2962_210.t0 GND 0.31fF
C126 a_16984_101.n0 GND 0.06fF
C127 a_16984_101.n1 GND 0.13fF
C128 a_16984_101.n2 GND 0.04fF
C129 a_16984_101.n3 GND 0.19fF
C130 a_5552_210.n0 GND 0.07fF
C131 a_5552_210.n1 GND 0.09fF
C132 a_5552_210.n2 GND 0.12fF
C133 a_5552_210.n3 GND 0.08fF
C134 a_5552_210.n4 GND 0.02fF
C135 a_5552_210.n5 GND 0.03fF
C136 a_5552_210.n6 GND 0.02fF
C137 a_5552_210.n7 GND 0.03fF
C138 a_5552_210.n8 GND 0.02fF
C139 a_5552_210.n9 GND 0.13fF
C140 a_5552_210.n10 GND 0.08fF
C141 a_5552_210.n11 GND 0.02fF
C142 a_5552_210.t0 GND 0.31fF
C143 a_6233_103.n0 GND 0.08fF
C144 a_6233_103.n1 GND 0.07fF
C145 a_6233_103.n2 GND 0.04fF
C146 a_6233_103.n3 GND 0.06fF
C147 a_6233_103.n4 GND 0.03fF
C148 a_6233_103.n5 GND 0.04fF
C149 a_6233_103.n7 GND 0.08fF
C150 a_10732_210.n0 GND 0.07fF
C151 a_10732_210.n1 GND 0.09fF
C152 a_10732_210.n2 GND 0.12fF
C153 a_10732_210.n3 GND 0.08fF
C154 a_10732_210.n4 GND 0.02fF
C155 a_10732_210.n5 GND 0.03fF
C156 a_10732_210.n6 GND 0.05fF
C157 a_10732_210.n7 GND 0.02fF
C158 a_10732_210.n8 GND 0.14fF
C159 a_10732_210.n9 GND 0.08fF
C160 a_10732_210.n10 GND 0.02fF
C161 a_10732_210.t0 GND 0.31fF
C162 a_372_210.n0 GND 0.07fF
C163 a_372_210.n1 GND 0.09fF
C164 a_372_210.n2 GND 0.12fF
C165 a_372_210.n3 GND 0.08fF
C166 a_372_210.n4 GND 0.02fF
C167 a_372_210.n5 GND 0.03fF
C168 a_372_210.n6 GND 0.02fF
C169 a_372_210.n7 GND 0.03fF
C170 a_372_210.n8 GND 0.02fF
C171 a_372_210.n9 GND 0.13fF
C172 a_372_210.n10 GND 0.08fF
C173 a_372_210.n11 GND 0.02fF
C174 a_372_210.t0 GND 0.31fF
C175 a_16318_101.n0 GND 0.13fF
C176 a_16318_101.n1 GND 0.14fF
C177 a_16318_101.n2 GND 0.14fF
C178 a_9104_210.n0 GND 0.02fF
C179 a_9104_210.n1 GND 0.09fF
C180 a_9104_210.n2 GND 0.12fF
C181 a_9104_210.n3 GND 0.08fF
C182 a_9104_210.n4 GND 0.08fF
C183 a_9104_210.n5 GND 0.02fF
C184 a_9104_210.t1 GND 0.29fF
C185 a_9104_210.n6 GND 0.09fF
C186 a_9104_210.n7 GND 0.02fF
C187 a_9104_210.n8 GND 0.13fF
C188 a_9104_210.n9 GND 0.02fF
C189 a_9104_210.n10 GND 0.03fF
C190 a_9104_210.n11 GND 0.02fF
C191 a_8823_103.n0 GND 0.08fF
C192 a_8823_103.n1 GND 0.07fF
C193 a_8823_103.n2 GND 0.04fF
C194 a_8823_103.n3 GND 0.06fF
C195 a_8823_103.n4 GND 0.11fF
C196 a_8823_103.n5 GND 0.04fF
C197 a_8823_103.n7 GND 0.08fF
C198 a_7321_1050.n0 GND 0.39fF
C199 a_7321_1050.n1 GND 0.33fF
C200 a_7321_1050.n2 GND 0.67fF
C201 a_7321_1050.n3 GND 0.04fF
C202 a_7321_1050.n4 GND 0.06fF
C203 a_7321_1050.n5 GND 0.03fF
C204 a_7321_1050.n6 GND 0.23fF
C205 a_7321_1050.n7 GND 0.69fF
C206 a_7321_1050.n8 GND 0.59fF
C207 a_7321_1050.n9 GND 0.51fF
C208 a_12501_1050.n0 GND 0.36fF
C209 a_12501_1050.n1 GND 0.72fF
C210 a_12501_1050.n2 GND 0.37fF
C211 a_12501_1050.n3 GND 0.76fF
C212 a_12501_1050.n4 GND 0.54fF
C213 a_12501_1050.n5 GND 0.64fF
C214 a_12501_1050.n6 GND 0.42fF
C215 a_14986_101.n0 GND 0.02fF
C216 a_14986_101.n1 GND 0.09fF
C217 a_14986_101.n2 GND 0.08fF
C218 a_14986_101.n3 GND 0.03fF
C219 a_14986_101.n4 GND 0.01fF
C220 a_14986_101.n5 GND 0.04fF
C221 a_14986_101.n6 GND 0.04fF
C222 a_14986_101.n7 GND 0.02fF
C223 a_14986_101.n8 GND 0.05fF
C224 a_14986_101.n9 GND 0.15fF
C225 a_14986_101.n10 GND 0.08fF
C226 a_14986_101.n11 GND 0.08fF
C227 a_14986_101.t1 GND 0.23fF
C228 a_14986_101.n12 GND 0.01fF
C229 a_11694_210.n0 GND 0.02fF
C230 a_11694_210.n1 GND 0.09fF
C231 a_11694_210.n2 GND 0.12fF
C232 a_11694_210.n3 GND 0.08fF
C233 a_11694_210.n4 GND 0.08fF
C234 a_11694_210.n5 GND 0.02fF
C235 a_11694_210.t1 GND 0.29fF
C236 a_11694_210.n6 GND 0.09fF
C237 a_11694_210.n7 GND 0.02fF
C238 a_11694_210.n8 GND 0.13fF
C239 a_11694_210.n9 GND 0.02fF
C240 a_11694_210.n10 GND 0.03fF
C241 a_11694_210.n11 GND 0.02fF
C242 a_6514_210.n0 GND 0.02fF
C243 a_6514_210.n1 GND 0.09fF
C244 a_6514_210.n2 GND 0.12fF
C245 a_6514_210.n3 GND 0.08fF
C246 a_6514_210.n4 GND 0.08fF
C247 a_6514_210.n5 GND 0.02fF
C248 a_6514_210.t1 GND 0.29fF
C249 a_6514_210.n6 GND 0.09fF
C250 a_6514_210.n7 GND 0.02fF
C251 a_6514_210.n8 GND 0.13fF
C252 a_6514_210.n9 GND 0.02fF
C253 a_6514_210.n10 GND 0.03fF
C254 a_6514_210.n11 GND 0.03fF
C255 a_15652_101.n0 GND 0.09fF
C256 a_15652_101.n1 GND 0.07fF
C257 a_15652_101.n2 GND 0.11fF
C258 a_15652_101.n3 GND 0.02fF
C259 a_15652_101.n4 GND 0.02fF
C260 a_15652_101.n5 GND 0.06fF
C261 a_15652_101.n6 GND 0.21fF
C262 a_15757_1051.n0 GND 0.36fF
C263 a_15757_1051.n1 GND 0.43fF
C264 a_15757_1051.n2 GND 0.80fF
C265 a_15757_1051.n3 GND 0.30fF
C266 a_15757_1051.n4 GND 0.52fF
C267 a_15757_1051.n5 GND 0.32fF
C268 a_10451_103.n0 GND 0.13fF
C269 a_10451_103.n1 GND 0.04fF
C270 a_10451_103.n2 GND 0.09fF
C271 a_10451_103.n3 GND 0.07fF
C272 a_10451_103.n4 GND 0.08fF
C273 a_10451_103.n5 GND 0.03fF
C274 a_2036_101.n0 GND 0.02fF
C275 a_2036_101.n1 GND 0.09fF
C276 a_2036_101.n2 GND 0.08fF
C277 a_2036_101.n3 GND 0.03fF
C278 a_2036_101.n4 GND 0.01fF
C279 a_2036_101.n5 GND 0.04fF
C280 a_2036_101.n6 GND 0.04fF
C281 a_2036_101.n7 GND 0.02fF
C282 a_2036_101.n8 GND 0.05fF
C283 a_2036_101.n9 GND 0.15fF
C284 a_2036_101.n10 GND 0.08fF
C285 a_2036_101.n11 GND 0.08fF
C286 a_2036_101.t1 GND 0.23fF
C287 a_2036_101.n12 GND 0.01fF
C288 a_3829_1050.n0 GND 0.35fF
C289 a_3829_1050.n1 GND 0.28fF
C290 a_3829_1050.n2 GND 0.55fF
C291 a_3829_1050.n3 GND 0.04fF
C292 a_3829_1050.n4 GND 0.05fF
C293 a_3829_1050.n5 GND 0.03fF
C294 a_3829_1050.n6 GND 0.23fF
C295 a_3829_1050.n7 GND 0.63fF
C296 a_3829_1050.n8 GND 0.38fF
C297 a_3829_1050.n9 GND 0.45fF
C298 a_3829_1050.n10 GND 0.43fF
C299 a_3829_1050.n11 GND 0.35fF
C300 a_12396_101.n0 GND 0.05fF
C301 a_12396_101.n1 GND 0.12fF
C302 a_12396_101.n2 GND 0.04fF
C303 a_12396_101.n3 GND 0.17fF
C304 a_5779_989.n0 GND 0.46fF
C305 a_5779_989.n1 GND 0.39fF
C306 a_5779_989.n2 GND 0.56fF
C307 a_5779_989.n3 GND 0.39fF
C308 a_5779_989.t7 GND 0.63fF
C309 a_5779_989.n4 GND 0.75fF
C310 a_5779_989.n5 GND 1.19fF
C311 a_5779_989.n6 GND 0.05fF
C312 a_5779_989.n7 GND 0.06fF
C313 a_5779_989.n8 GND 0.04fF
C314 a_5779_989.n9 GND 0.27fF
C315 a_5779_989.n10 GND 0.62fF
C316 a_5779_989.n11 GND 0.53fF
C317 a_5779_989.n12 GND 0.59fF
C318 a_5779_989.n13 GND 0.56fF
C319 a_5779_989.n14 GND 0.46fF
C320 a_5457_1050.n0 GND 0.60fF
C321 a_5457_1050.n1 GND 0.60fF
C322 a_5457_1050.n2 GND 0.47fF
C323 a_5457_1050.n3 GND 1.86fF
C324 a_5457_1050.n4 GND 0.47fF
C325 a_5457_1050.n5 GND 0.74fF
C326 a_5457_1050.n6 GND 2.64fF
C327 a_5457_1050.n7 GND 0.57fF
C328 a_5457_1050.n8 GND 0.90fF
C329 a_5457_1050.n9 GND 0.65fF
C330 a_5457_1050.n10 GND 0.73fF
C331 a_5457_1050.n11 GND 0.77fF
C332 a_277_1050.n0 GND 0.43fF
C333 a_277_1050.n1 GND 1.71fF
C334 a_277_1050.n2 GND 0.43fF
C335 a_277_1050.n3 GND 0.68fF
C336 a_277_1050.n4 GND 2.43fF
C337 a_277_1050.n5 GND 0.06fF
C338 a_277_1050.n6 GND 0.08fF
C339 a_277_1050.n7 GND 0.05fF
C340 a_277_1050.n8 GND 0.36fF
C341 a_277_1050.n9 GND 0.80fF
C342 a_277_1050.n10 GND 0.56fF
C343 a_277_1050.n11 GND 0.71fF
C344 a_277_1050.n12 GND 0.67fF
C345 a_277_1050.n13 GND 0.59fF
C346 a_277_1050.n14 GND 0.56fF
C347 a_1334_210.n0 GND 0.02fF
C348 a_1334_210.n1 GND 0.09fF
C349 a_1334_210.n2 GND 0.12fF
C350 a_1334_210.n3 GND 0.08fF
C351 a_1334_210.n4 GND 0.08fF
C352 a_1334_210.n5 GND 0.02fF
C353 a_1334_210.t1 GND 0.29fF
C354 a_1334_210.n6 GND 0.09fF
C355 a_1334_210.n7 GND 0.02fF
C356 a_1334_210.n8 GND 0.13fF
C357 a_1334_210.n9 GND 0.02fF
C358 a_1334_210.n10 GND 0.03fF
C359 a_1334_210.n11 GND 0.02fF
C360 a_1053_103.n0 GND 0.08fF
C361 a_1053_103.n1 GND 0.07fF
C362 a_1053_103.n2 GND 0.04fF
C363 a_1053_103.n3 GND 0.06fF
C364 a_1053_103.n4 GND 0.11fF
C365 a_1053_103.n5 GND 0.04fF
C366 a_1053_103.n7 GND 0.08fF
C367 a_4151_989.n0 GND 0.86fF
C368 a_4151_989.n1 GND 0.98fF
C369 a_4151_989.n2 GND 1.36fF
C370 a_4151_989.t10 GND 0.97fF
C371 a_4151_989.n3 GND 0.74fF
C372 a_4151_989.n4 GND 10.33fF
C373 a_4151_989.n5 GND 0.85fF
C374 a_4151_989.t9 GND 1.09fF
C375 a_4151_989.n6 GND 1.19fF
C376 a_4151_989.n7 GND 12.86fF
C377 a_4151_989.n8 GND 0.62fF
C378 a_4151_989.n9 GND 1.14fF
C379 a_4151_989.n10 GND 1.10fF
C380 a_4151_989.n11 GND 1.43fF
C381 a_4151_989.n12 GND 0.86fF
C382 a_4626_101.n0 GND 0.08fF
C383 a_4626_101.n1 GND 0.02fF
C384 a_4626_101.n2 GND 0.02fF
C385 a_4626_101.n3 GND 0.09fF
C386 a_4626_101.n4 GND 0.08fF
C387 a_4626_101.n5 GND 0.03fF
C388 a_4626_101.n6 GND 0.05fF
C389 a_147_187.n0 GND 0.46fF
C390 a_147_187.t7 GND 0.95fF
C391 a_147_187.n1 GND 1.20fF
C392 a_147_187.n2 GND 0.46fF
C393 a_147_187.t8 GND 0.95fF
C394 a_147_187.n3 GND 0.64fF
C395 a_147_187.n4 GND 0.47fF
C396 a_147_187.n5 GND 1.67fF
C397 a_147_187.n6 GND 2.70fF
C398 a_147_187.n7 GND 2.24fF
C399 a_147_187.n8 GND 0.07fF
C400 a_147_187.n9 GND 0.09fF
C401 a_147_187.n10 GND 0.06fF
C402 a_147_187.n11 GND 0.47fF
C403 a_147_187.n12 GND 0.87fF
C404 a_147_187.n13 GND 0.65fF
C405 a_147_187.n14 GND 0.82fF
C406 a_147_187.n15 GND 0.78fF
C407 a_147_187.n16 GND 0.64fF
C408 a_147_187.n17 GND 0.65fF
C409 a_9331_989.n0 GND 0.49fF
C410 a_9331_989.n1 GND 1.52fF
C411 a_9331_989.n2 GND 0.48fF
C412 a_9331_989.n3 GND 1.10fF
C413 a_9331_989.n4 GND 4.30fF
C414 a_9331_989.n5 GND 0.70fF
C415 a_9331_989.t13 GND 1.00fF
C416 a_9331_989.n6 GND 1.08fF
C417 a_9331_989.n7 GND 6.33fF
C418 a_9331_989.n8 GND 0.08fF
C419 a_9331_989.n9 GND 0.11fF
C420 a_9331_989.n10 GND 0.07fF
C421 a_9331_989.n11 GND 0.38fF
C422 a_9331_989.n12 GND 0.98fF
C423 a_9331_989.n13 GND 0.97fF
C424 a_9331_989.n14 GND 1.20fF
C425 a_9331_989.n15 GND 0.76fF
C426 a_9009_1050.n0 GND 0.37fF
C427 a_9009_1050.n1 GND 0.29fF
C428 a_9009_1050.n2 GND 0.58fF
C429 a_9009_1050.n3 GND 0.35fF
C430 a_9009_1050.n4 GND 0.68fF
C431 a_9009_1050.n5 GND 0.40fF
C432 a_9009_1050.n6 GND 0.47fF
C433 a_9009_1050.n7 GND 0.45fF
C434 a_9009_1050.n8 GND 0.37fF
C435 a_2141_1050.n0 GND 0.38fF
C436 a_2141_1050.n1 GND 0.32fF
C437 a_2141_1050.n2 GND 0.64fF
C438 a_2141_1050.n3 GND 0.33fF
C439 a_2141_1050.n4 GND 0.68fF
C440 a_2141_1050.n5 GND 0.57fF
C441 a_2141_1050.n6 GND 0.48fF
C442 a_5327_187.n0 GND 0.49fF
C443 a_5327_187.t11 GND 1.03fF
C444 a_5327_187.n1 GND 1.30fF
C445 a_5327_187.n2 GND 0.49fF
C446 a_5327_187.t14 GND 1.03fF
C447 a_5327_187.n3 GND 0.69fF
C448 a_5327_187.n4 GND 0.51fF
C449 a_5327_187.n5 GND 1.81fF
C450 a_5327_187.n6 GND 2.92fF
C451 a_5327_187.n7 GND 2.42fF
C452 a_5327_187.n8 GND 0.08fF
C453 a_5327_187.n9 GND 0.10fF
C454 a_5327_187.n10 GND 0.54fF
C455 a_5327_187.n11 GND 0.96fF
C456 a_5327_187.n12 GND 0.70fF
C457 a_5327_187.n13 GND 0.89fF
C458 a_5327_187.n14 GND 0.84fF
C459 a_5327_187.n15 GND 0.69fF
C460 a_5327_187.n16 GND 0.70fF
C461 a_8142_210.n0 GND 0.02fF
C462 a_8142_210.n1 GND 0.09fF
C463 a_8142_210.t1 GND 0.23fF
C464 a_8142_210.n2 GND 0.10fF
C465 a_8142_210.n3 GND 0.07fF
C466 a_8142_210.n4 GND 0.04fF
C467 a_8142_210.n5 GND 0.08fF
C468 a_8142_210.n6 GND 0.09fF
C469 a_8142_210.n7 GND 0.04fF
C470 a_8142_210.n8 GND 0.02fF
C471 a_8142_210.n9 GND 0.01fF
C472 a_8142_210.n10 GND 0.13fF
C473 a_8142_210.n11 GND 0.02fF
C474 a_8142_210.n12 GND 0.03fF
C475 a_8142_210.n13 GND 0.02fF
C476 a_16421_1051.n0 GND 0.29fF
C477 a_16421_1051.n1 GND 0.28fF
C478 a_16421_1051.n2 GND 0.37fF
C479 a_16421_1051.n3 GND 0.70fF
C480 a_16421_1051.n4 GND 0.27fF
C481 a_16421_1051.n5 GND 0.45fF
C482 a_15932_209.n0 GND 0.03fF
C483 a_15932_209.n1 GND 0.27fF
C484 a_15932_209.n2 GND 0.34fF
C485 a_15932_209.n3 GND 0.41fF
C486 a_15932_209.n4 GND 0.24fF
C487 a_15932_209.n5 GND 0.47fF
C488 a_15932_209.n6 GND 0.43fF
C489 a_15932_209.n7 GND 0.05fF
C490 a_15932_209.n8 GND 0.03fF
C491 a_15932_209.n9 GND 0.05fF
C492 a_15932_209.n10 GND 0.33fF
C493 a_15932_209.n11 GND 0.03fF
C494 a_15932_209.n12 GND 0.04fF
C495 a_15932_209.n13 GND 0.03fF
C496 a_15932_209.n14 GND 0.04fF
C497 a_15932_209.n15 GND 0.95fF
C498 a_15932_209.n16 GND 0.03fF
C499 a_15932_209.n17 GND 0.03fF
C500 a_15932_209.n18 GND 0.04fF
C501 a_14511_989.n0 GND 0.41fF
C502 a_14511_989.n1 GND 0.30fF
C503 a_14511_989.n2 GND 0.31fF
C504 a_14511_989.t10 GND 0.61fF
C505 a_14511_989.n3 GND 1.06fF
C506 a_14511_989.n4 GND 0.74fF
C507 a_14511_989.t7 GND 0.56fF
C508 a_14511_989.n5 GND 0.41fF
C509 a_14511_989.n6 GND 0.35fF
C510 a_14511_989.t12 GND 0.56fF
C511 a_14511_989.n7 GND 0.59fF
C512 a_14511_989.n8 GND 1.00fF
C513 a_14511_989.n9 GND 0.04fF
C514 a_14511_989.n10 GND 0.06fF
C515 a_14511_989.n11 GND 0.04fF
C516 a_14511_989.n12 GND 0.24fF
C517 a_14511_989.n13 GND 0.53fF
C518 a_14511_989.n14 GND 0.62fF
C519 a_14511_989.n15 GND 0.53fF
C520 a_11413_103.n0 GND 0.03fF
C521 a_11413_103.n1 GND 0.09fF
C522 a_11413_103.n2 GND 0.08fF
C523 a_11413_103.n3 GND 0.04fF
C524 a_11413_103.n4 GND 0.05fF
C525 a_11413_103.n5 GND 0.11fF
C526 a_11413_103.n6 GND 0.04fF
C527 a_11413_103.n8 GND 0.08fF
C528 a_599_989.n0 GND 0.41fF
C529 a_599_989.n1 GND 0.34fF
C530 a_599_989.n2 GND 0.49fF
C531 a_599_989.n3 GND 0.34fF
C532 a_599_989.t9 GND 0.56fF
C533 a_599_989.n4 GND 0.66fF
C534 a_599_989.n5 GND 1.06fF
C535 a_599_989.n6 GND 0.04fF
C536 a_599_989.n7 GND 0.06fF
C537 a_599_989.n8 GND 0.04fF
C538 a_599_989.n9 GND 0.24fF
C539 a_599_989.n10 GND 0.55fF
C540 a_599_989.n11 GND 0.47fF
C541 a_599_989.n12 GND 0.52fF
C542 a_599_989.n13 GND 0.49fF
C543 a_599_989.n14 GND 0.41fF
C544 a_10959_989.n0 GND 0.54fF
C545 a_10959_989.n1 GND 0.54fF
C546 a_10959_989.n2 GND 0.45fF
C547 a_10959_989.n3 GND 0.65fF
C548 a_10959_989.n4 GND 0.45fF
C549 a_10959_989.t11 GND 0.73fF
C550 a_10959_989.n5 GND 0.87fF
C551 a_10959_989.n6 GND 1.38fF
C552 a_10959_989.n7 GND 0.06fF
C553 a_10959_989.n8 GND 0.07fF
C554 a_10959_989.n9 GND 0.05fF
C555 a_10959_989.n10 GND 0.31fF
C556 a_10959_989.n11 GND 0.72fF
C557 a_10959_989.n12 GND 0.62fF
C558 a_10959_989.n13 GND 0.65fF
C559 a_10959_989.n14 GND 0.68fF
C560 a_14189_1050.n0 GND 0.37fF
C561 a_14189_1050.n1 GND 0.37fF
C562 a_14189_1050.n2 GND 0.29fF
C563 a_14189_1050.n3 GND 0.58fF
C564 a_14189_1050.n4 GND 0.35fF
C565 a_14189_1050.n5 GND 0.68fF
C566 a_14189_1050.n6 GND 0.39fF
C567 a_14189_1050.n7 GND 0.44fF
C568 a_14189_1050.n8 GND 0.47fF
C569 a_10637_1050.n0 GND 0.63fF
C570 a_10637_1050.n1 GND 0.63fF
C571 a_10637_1050.n2 GND 0.49fF
C572 a_10637_1050.n3 GND 1.93fF
C573 a_10637_1050.n4 GND 0.49fF
C574 a_10637_1050.n5 GND 0.77fF
C575 a_10637_1050.n6 GND 2.74fF
C576 a_10637_1050.n7 GND 0.59fF
C577 a_10637_1050.n8 GND 0.93fF
C578 a_10637_1050.n9 GND 0.67fF
C579 a_10637_1050.n10 GND 0.75fF
C580 a_10637_1050.n11 GND 0.80fF
C581 VDD.n1 GND 0.03fF
C582 VDD.n2 GND 0.10fF
C583 VDD.n3 GND 0.03fF
C584 VDD.n4 GND 0.02fF
C585 VDD.n5 GND 0.06fF
C586 VDD.n6 GND 0.02fF
C587 VDD.n7 GND 0.02fF
C588 VDD.n8 GND 0.02fF
C589 VDD.n9 GND 0.02fF
C590 VDD.n10 GND 0.02fF
C591 VDD.n11 GND 0.02fF
C592 VDD.n12 GND 0.02fF
C593 VDD.n13 GND 0.02fF
C594 VDD.n14 GND 0.04fF
C595 VDD.n15 GND 0.01fF
C596 VDD.n20 GND 0.48fF
C597 VDD.n21 GND 0.29fF
C598 VDD.n22 GND 0.02fF
C599 VDD.n23 GND 0.03fF
C600 VDD.n24 GND 0.07fF
C601 VDD.n25 GND 0.21fF
C602 VDD.n26 GND 0.01fF
C603 VDD.n27 GND 0.01fF
C604 VDD.n28 GND 0.07fF
C605 VDD.n29 GND 0.18fF
C606 VDD.n30 GND 0.01fF
C607 VDD.n31 GND 0.03fF
C608 VDD.n32 GND 0.03fF
C609 VDD.n33 GND 0.21fF
C610 VDD.n34 GND 0.01fF
C611 VDD.n35 GND 0.07fF
C612 VDD.n36 GND 0.01fF
C613 VDD.n37 GND 0.02fF
C614 VDD.n38 GND 0.29fF
C615 VDD.n39 GND 0.01fF
C616 VDD.n40 GND 0.02fF
C617 VDD.n41 GND 0.04fF
C618 VDD.n42 GND 0.06fF
C619 VDD.n43 GND 0.02fF
C620 VDD.n44 GND 0.02fF
C621 VDD.n45 GND 0.02fF
C622 VDD.n46 GND 0.02fF
C623 VDD.n47 GND 0.02fF
C624 VDD.n48 GND 0.02fF
C625 VDD.n49 GND 0.02fF
C626 VDD.n50 GND 0.02fF
C627 VDD.n51 GND 0.02fF
C628 VDD.n52 GND 0.02fF
C629 VDD.n53 GND 0.02fF
C630 VDD.n54 GND 0.03fF
C631 VDD.n55 GND 0.02fF
C632 VDD.n56 GND 0.19fF
C633 VDD.n57 GND 0.02fF
C634 VDD.n58 GND 0.02fF
C635 VDD.n60 GND 0.02fF
C636 VDD.n64 GND 0.29fF
C637 VDD.n65 GND 0.29fF
C638 VDD.n66 GND 0.01fF
C639 VDD.n67 GND 0.02fF
C640 VDD.n68 GND 0.04fF
C641 VDD.n69 GND 0.26fF
C642 VDD.n70 GND 0.01fF
C643 VDD.n71 GND 0.02fF
C644 VDD.n72 GND 0.02fF
C645 VDD.n73 GND 0.18fF
C646 VDD.n74 GND 0.01fF
C647 VDD.n75 GND 0.02fF
C648 VDD.n76 GND 0.02fF
C649 VDD.n77 GND 0.01fF
C650 VDD.n78 GND 0.03fF
C651 VDD.n79 GND 0.03fF
C652 VDD.n80 GND 0.15fF
C653 VDD.n81 GND 0.01fF
C654 VDD.n82 GND 0.03fF
C655 VDD.n83 GND 0.03fF
C656 VDD.n84 GND 0.17fF
C657 VDD.n85 GND 0.01fF
C658 VDD.n86 GND 0.02fF
C659 VDD.n87 GND 0.02fF
C660 VDD.n88 GND 0.26fF
C661 VDD.n89 GND 0.01fF
C662 VDD.n90 GND 0.02fF
C663 VDD.n91 GND 0.02fF
C664 VDD.n92 GND 0.29fF
C665 VDD.n93 GND 0.01fF
C666 VDD.n94 GND 0.02fF
C667 VDD.n95 GND 0.04fF
C668 VDD.n96 GND 0.22fF
C669 VDD.n97 GND 0.02fF
C670 VDD.n98 GND 0.02fF
C671 VDD.n99 GND 0.02fF
C672 VDD.n100 GND 0.06fF
C673 VDD.n101 GND 0.02fF
C674 VDD.n102 GND 0.02fF
C675 VDD.n103 GND 0.02fF
C676 VDD.n104 GND 0.02fF
C677 VDD.n105 GND 0.02fF
C678 VDD.n106 GND 0.02fF
C679 VDD.n107 GND 0.02fF
C680 VDD.n108 GND 0.02fF
C681 VDD.n109 GND 0.02fF
C682 VDD.n110 GND 0.02fF
C683 VDD.n111 GND 0.03fF
C684 VDD.n112 GND 0.02fF
C685 VDD.n113 GND 0.02fF
C686 VDD.n117 GND 0.29fF
C687 VDD.n118 GND 0.29fF
C688 VDD.n119 GND 0.01fF
C689 VDD.n120 GND 0.02fF
C690 VDD.n121 GND 0.04fF
C691 VDD.n122 GND 0.26fF
C692 VDD.n123 GND 0.01fF
C693 VDD.n124 GND 0.02fF
C694 VDD.n125 GND 0.02fF
C695 VDD.n126 GND 0.17fF
C696 VDD.n127 GND 0.01fF
C697 VDD.n128 GND 0.02fF
C698 VDD.n129 GND 0.02fF
C699 VDD.n130 GND 0.15fF
C700 VDD.n131 GND 0.01fF
C701 VDD.n132 GND 0.03fF
C702 VDD.n133 GND 0.03fF
C703 VDD.n134 GND 0.01fF
C704 VDD.n135 GND 0.03fF
C705 VDD.n136 GND 0.03fF
C706 VDD.n137 GND 0.18fF
C707 VDD.n138 GND 0.01fF
C708 VDD.n139 GND 0.02fF
C709 VDD.n140 GND 0.02fF
C710 VDD.n141 GND 0.26fF
C711 VDD.n142 GND 0.01fF
C712 VDD.n143 GND 0.02fF
C713 VDD.n144 GND 0.02fF
C714 VDD.n145 GND 0.29fF
C715 VDD.n146 GND 0.01fF
C716 VDD.n147 GND 0.02fF
C717 VDD.n148 GND 0.04fF
C718 VDD.n149 GND 0.22fF
C719 VDD.n150 GND 0.02fF
C720 VDD.n151 GND 0.02fF
C721 VDD.n152 GND 0.02fF
C722 VDD.n153 GND 0.06fF
C723 VDD.n154 GND 0.02fF
C724 VDD.n155 GND 0.02fF
C725 VDD.n156 GND 0.02fF
C726 VDD.n157 GND 0.02fF
C727 VDD.n158 GND 0.02fF
C728 VDD.n159 GND 0.02fF
C729 VDD.n160 GND 0.02fF
C730 VDD.n161 GND 0.02fF
C731 VDD.n162 GND 0.02fF
C732 VDD.n163 GND 0.02fF
C733 VDD.n164 GND 0.03fF
C734 VDD.n165 GND 0.02fF
C735 VDD.n166 GND 0.02fF
C736 VDD.n170 GND 0.29fF
C737 VDD.n171 GND 0.29fF
C738 VDD.n172 GND 0.01fF
C739 VDD.n173 GND 0.02fF
C740 VDD.n174 GND 0.04fF
C741 VDD.n175 GND 0.07fF
C742 VDD.n176 GND 0.26fF
C743 VDD.n177 GND 0.01fF
C744 VDD.n178 GND 0.01fF
C745 VDD.n179 GND 0.02fF
C746 VDD.n180 GND 0.18fF
C747 VDD.n181 GND 0.01fF
C748 VDD.n182 GND 0.02fF
C749 VDD.n183 GND 0.02fF
C750 VDD.n184 GND 0.08fF
C751 VDD.n185 GND 0.05fF
C752 VDD.n186 GND 0.01fF
C753 VDD.n187 GND 0.02fF
C754 VDD.n188 GND 0.03fF
C755 VDD.n189 GND 0.15fF
C756 VDD.n190 GND 0.01fF
C757 VDD.n191 GND 0.02fF
C758 VDD.n192 GND 0.03fF
C759 VDD.n193 GND 0.17fF
C760 VDD.n194 GND 0.01fF
C761 VDD.n195 GND 0.02fF
C762 VDD.n196 GND 0.02fF
C763 VDD.n197 GND 0.07fF
C764 VDD.n198 GND 0.26fF
C765 VDD.n199 GND 0.01fF
C766 VDD.n200 GND 0.01fF
C767 VDD.n201 GND 0.02fF
C768 VDD.n202 GND 0.29fF
C769 VDD.n203 GND 0.01fF
C770 VDD.n204 GND 0.02fF
C771 VDD.n205 GND 0.04fF
C772 VDD.n206 GND 0.22fF
C773 VDD.n207 GND 0.02fF
C774 VDD.n208 GND 0.02fF
C775 VDD.n209 GND 0.02fF
C776 VDD.n210 GND 0.06fF
C777 VDD.n211 GND 0.02fF
C778 VDD.n212 GND 0.02fF
C779 VDD.n213 GND 0.02fF
C780 VDD.n214 GND 0.02fF
C781 VDD.n215 GND 0.02fF
C782 VDD.n216 GND 0.02fF
C783 VDD.n217 GND 0.02fF
C784 VDD.n218 GND 0.02fF
C785 VDD.n219 GND 0.02fF
C786 VDD.n220 GND 0.02fF
C787 VDD.n221 GND 0.03fF
C788 VDD.n222 GND 0.02fF
C789 VDD.n223 GND 0.02fF
C790 VDD.n227 GND 0.29fF
C791 VDD.n228 GND 0.29fF
C792 VDD.n229 GND 0.01fF
C793 VDD.n230 GND 0.02fF
C794 VDD.n231 GND 0.04fF
C795 VDD.n232 GND 0.06fF
C796 VDD.n233 GND 0.26fF
C797 VDD.n234 GND 0.01fF
C798 VDD.n235 GND 0.01fF
C799 VDD.n236 GND 0.02fF
C800 VDD.n237 GND 0.18fF
C801 VDD.n238 GND 0.01fF
C802 VDD.n239 GND 0.02fF
C803 VDD.n240 GND 0.02fF
C804 VDD.n241 GND 0.08fF
C805 VDD.n242 GND 0.05fF
C806 VDD.n243 GND 0.01fF
C807 VDD.n244 GND 0.02fF
C808 VDD.n245 GND 0.03fF
C809 VDD.n246 GND 0.15fF
C810 VDD.n247 GND 0.01fF
C811 VDD.n248 GND 0.02fF
C812 VDD.n249 GND 0.03fF
C813 VDD.n250 GND 0.17fF
C814 VDD.n251 GND 0.01fF
C815 VDD.n252 GND 0.02fF
C816 VDD.n253 GND 0.02fF
C817 VDD.n254 GND 0.07fF
C818 VDD.n255 GND 0.26fF
C819 VDD.n256 GND 0.01fF
C820 VDD.n257 GND 0.01fF
C821 VDD.n258 GND 0.02fF
C822 VDD.n259 GND 0.29fF
C823 VDD.n260 GND 0.01fF
C824 VDD.n261 GND 0.02fF
C825 VDD.n262 GND 0.04fF
C826 VDD.n263 GND 0.27fF
C827 VDD.n264 GND 0.02fF
C828 VDD.n265 GND 0.02fF
C829 VDD.n266 GND 0.02fF
C830 VDD.n267 GND 0.06fF
C831 VDD.n268 GND 0.02fF
C832 VDD.n269 GND 0.02fF
C833 VDD.n270 GND 0.02fF
C834 VDD.n271 GND 0.02fF
C835 VDD.n272 GND 0.02fF
C836 VDD.n273 GND 0.02fF
C837 VDD.n274 GND 0.02fF
C838 VDD.n275 GND 0.02fF
C839 VDD.n276 GND 0.02fF
C840 VDD.n277 GND 0.02fF
C841 VDD.n278 GND 0.03fF
C842 VDD.n279 GND 0.02fF
C843 VDD.n280 GND 0.02fF
C844 VDD.n284 GND 0.29fF
C845 VDD.n285 GND 0.29fF
C846 VDD.n286 GND 0.01fF
C847 VDD.n287 GND 0.02fF
C848 VDD.n288 GND 0.04fF
C849 VDD.n289 GND 0.29fF
C850 VDD.n290 GND 0.01fF
C851 VDD.n291 GND 0.02fF
C852 VDD.n292 GND 0.02fF
C853 VDD.n293 GND 0.23fF
C854 VDD.n294 GND 0.01fF
C855 VDD.n295 GND 0.07fF
C856 VDD.n296 GND 0.02fF
C857 VDD.n297 GND 0.18fF
C858 VDD.n298 GND 0.01fF
C859 VDD.n299 GND 0.02fF
C860 VDD.n300 GND 0.02fF
C861 VDD.n301 GND 0.17fF
C862 VDD.n302 GND 0.01fF
C863 VDD.n303 GND 0.08fF
C864 VDD.n304 GND 0.05fF
C865 VDD.n305 GND 0.02fF
C866 VDD.n306 GND 0.02fF
C867 VDD.n307 GND 0.15fF
C868 VDD.n308 GND 0.02fF
C869 VDD.n309 GND 0.02fF
C870 VDD.n310 GND 0.03fF
C871 VDD.n311 GND 0.16fF
C872 VDD.n312 GND 0.02fF
C873 VDD.n313 GND 0.02fF
C874 VDD.n314 GND 0.03fF
C875 VDD.n315 GND 0.08fF
C876 VDD.n316 GND 0.05fF
C877 VDD.n317 GND 0.16fF
C878 VDD.n318 GND 0.01fF
C879 VDD.n319 GND 0.02fF
C880 VDD.n320 GND 0.02fF
C881 VDD.n321 GND 0.18fF
C882 VDD.n322 GND 0.01fF
C883 VDD.n323 GND 0.02fF
C884 VDD.n324 GND 0.02fF
C885 VDD.n325 GND 0.07fF
C886 VDD.n326 GND 0.24fF
C887 VDD.n327 GND 0.01fF
C888 VDD.n328 GND 0.01fF
C889 VDD.n329 GND 0.02fF
C890 VDD.n330 GND 0.29fF
C891 VDD.n331 GND 0.01fF
C892 VDD.n332 GND 0.02fF
C893 VDD.n333 GND 0.02fF
C894 VDD.n334 GND 0.29fF
C895 VDD.n335 GND 0.01fF
C896 VDD.n336 GND 0.02fF
C897 VDD.n337 GND 0.04fF
C898 VDD.n338 GND 0.32fF
C899 VDD.n339 GND 0.02fF
C900 VDD.n340 GND 0.02fF
C901 VDD.n341 GND 0.02fF
C902 VDD.n342 GND 0.06fF
C903 VDD.n343 GND 0.02fF
C904 VDD.n344 GND 0.02fF
C905 VDD.n345 GND 0.02fF
C906 VDD.n346 GND 0.02fF
C907 VDD.n347 GND 0.02fF
C908 VDD.n348 GND 0.02fF
C909 VDD.n349 GND 0.02fF
C910 VDD.n350 GND 0.02fF
C911 VDD.n351 GND 0.02fF
C912 VDD.n352 GND 0.02fF
C913 VDD.n353 GND 0.03fF
C914 VDD.n354 GND 0.02fF
C915 VDD.n355 GND 0.02fF
C916 VDD.n359 GND 0.29fF
C917 VDD.n360 GND 0.29fF
C918 VDD.n361 GND 0.01fF
C919 VDD.n362 GND 0.02fF
C920 VDD.n363 GND 0.04fF
C921 VDD.n364 GND 0.29fF
C922 VDD.n365 GND 0.01fF
C923 VDD.n366 GND 0.02fF
C924 VDD.n367 GND 0.02fF
C925 VDD.n368 GND 0.23fF
C926 VDD.n369 GND 0.01fF
C927 VDD.n370 GND 0.07fF
C928 VDD.n371 GND 0.02fF
C929 VDD.n372 GND 0.18fF
C930 VDD.n373 GND 0.01fF
C931 VDD.n374 GND 0.02fF
C932 VDD.n375 GND 0.02fF
C933 VDD.n376 GND 0.17fF
C934 VDD.n377 GND 0.01fF
C935 VDD.n378 GND 0.08fF
C936 VDD.n379 GND 0.05fF
C937 VDD.n380 GND 0.02fF
C938 VDD.n381 GND 0.02fF
C939 VDD.n382 GND 0.15fF
C940 VDD.n383 GND 0.02fF
C941 VDD.n384 GND 0.02fF
C942 VDD.n385 GND 0.03fF
C943 VDD.n386 GND 0.16fF
C944 VDD.n387 GND 0.02fF
C945 VDD.n388 GND 0.02fF
C946 VDD.n389 GND 0.03fF
C947 VDD.n390 GND 0.08fF
C948 VDD.n391 GND 0.05fF
C949 VDD.n392 GND 0.16fF
C950 VDD.n393 GND 0.01fF
C951 VDD.n394 GND 0.02fF
C952 VDD.n395 GND 0.02fF
C953 VDD.n396 GND 0.18fF
C954 VDD.n397 GND 0.01fF
C955 VDD.n398 GND 0.02fF
C956 VDD.n399 GND 0.02fF
C957 VDD.n400 GND 0.07fF
C958 VDD.n401 GND 0.24fF
C959 VDD.n402 GND 0.01fF
C960 VDD.n403 GND 0.01fF
C961 VDD.n404 GND 0.02fF
C962 VDD.n405 GND 0.29fF
C963 VDD.n406 GND 0.01fF
C964 VDD.n407 GND 0.02fF
C965 VDD.n408 GND 0.02fF
C966 VDD.n409 GND 0.29fF
C967 VDD.n410 GND 0.01fF
C968 VDD.n411 GND 0.02fF
C969 VDD.n412 GND 0.04fF
C970 VDD.n413 GND 0.27fF
C971 VDD.n414 GND 0.02fF
C972 VDD.n415 GND 0.02fF
C973 VDD.n416 GND 0.02fF
C974 VDD.n417 GND 0.06fF
C975 VDD.n418 GND 0.02fF
C976 VDD.n419 GND 0.02fF
C977 VDD.n420 GND 0.02fF
C978 VDD.n421 GND 0.02fF
C979 VDD.n422 GND 0.02fF
C980 VDD.n423 GND 0.02fF
C981 VDD.n424 GND 0.02fF
C982 VDD.n425 GND 0.02fF
C983 VDD.n426 GND 0.02fF
C984 VDD.n427 GND 0.02fF
C985 VDD.n428 GND 0.03fF
C986 VDD.n429 GND 0.02fF
C987 VDD.n430 GND 0.02fF
C988 VDD.n434 GND 0.29fF
C989 VDD.n435 GND 0.29fF
C990 VDD.n436 GND 0.01fF
C991 VDD.n437 GND 0.02fF
C992 VDD.n438 GND 0.04fF
C993 VDD.n439 GND 0.06fF
C994 VDD.n440 GND 0.26fF
C995 VDD.n441 GND 0.01fF
C996 VDD.n442 GND 0.01fF
C997 VDD.n443 GND 0.02fF
C998 VDD.n444 GND 0.18fF
C999 VDD.n445 GND 0.01fF
C1000 VDD.n446 GND 0.02fF
C1001 VDD.n447 GND 0.02fF
C1002 VDD.n448 GND 0.08fF
C1003 VDD.n449 GND 0.05fF
C1004 VDD.n450 GND 0.01fF
C1005 VDD.n451 GND 0.02fF
C1006 VDD.n452 GND 0.03fF
C1007 VDD.n453 GND 0.15fF
C1008 VDD.n454 GND 0.01fF
C1009 VDD.n455 GND 0.02fF
C1010 VDD.n456 GND 0.03fF
C1011 VDD.n457 GND 0.17fF
C1012 VDD.n458 GND 0.01fF
C1013 VDD.n459 GND 0.02fF
C1014 VDD.n460 GND 0.02fF
C1015 VDD.n461 GND 0.07fF
C1016 VDD.n462 GND 0.26fF
C1017 VDD.n463 GND 0.01fF
C1018 VDD.n464 GND 0.01fF
C1019 VDD.n465 GND 0.02fF
C1020 VDD.n466 GND 0.29fF
C1021 VDD.n467 GND 0.01fF
C1022 VDD.n468 GND 0.02fF
C1023 VDD.n469 GND 0.04fF
C1024 VDD.n470 GND 0.27fF
C1025 VDD.n471 GND 0.02fF
C1026 VDD.n472 GND 0.02fF
C1027 VDD.n473 GND 0.02fF
C1028 VDD.n474 GND 0.06fF
C1029 VDD.n475 GND 0.02fF
C1030 VDD.n476 GND 0.02fF
C1031 VDD.n477 GND 0.02fF
C1032 VDD.n478 GND 0.02fF
C1033 VDD.n479 GND 0.02fF
C1034 VDD.n480 GND 0.02fF
C1035 VDD.n481 GND 0.02fF
C1036 VDD.n482 GND 0.02fF
C1037 VDD.n483 GND 0.02fF
C1038 VDD.n484 GND 0.02fF
C1039 VDD.n485 GND 0.03fF
C1040 VDD.n486 GND 0.02fF
C1041 VDD.n487 GND 0.02fF
C1042 VDD.n491 GND 0.29fF
C1043 VDD.n492 GND 0.29fF
C1044 VDD.n493 GND 0.01fF
C1045 VDD.n494 GND 0.02fF
C1046 VDD.n495 GND 0.04fF
C1047 VDD.n496 GND 0.29fF
C1048 VDD.n497 GND 0.01fF
C1049 VDD.n498 GND 0.02fF
C1050 VDD.n499 GND 0.02fF
C1051 VDD.n500 GND 0.23fF
C1052 VDD.n501 GND 0.01fF
C1053 VDD.n502 GND 0.07fF
C1054 VDD.n503 GND 0.02fF
C1055 VDD.n504 GND 0.18fF
C1056 VDD.n505 GND 0.01fF
C1057 VDD.n506 GND 0.02fF
C1058 VDD.n507 GND 0.02fF
C1059 VDD.n508 GND 0.17fF
C1060 VDD.n509 GND 0.01fF
C1061 VDD.n510 GND 0.08fF
C1062 VDD.n511 GND 0.05fF
C1063 VDD.n512 GND 0.02fF
C1064 VDD.n513 GND 0.02fF
C1065 VDD.n514 GND 0.15fF
C1066 VDD.n515 GND 0.02fF
C1067 VDD.n516 GND 0.02fF
C1068 VDD.n517 GND 0.03fF
C1069 VDD.n518 GND 0.16fF
C1070 VDD.n519 GND 0.02fF
C1071 VDD.n520 GND 0.02fF
C1072 VDD.n521 GND 0.03fF
C1073 VDD.n522 GND 0.08fF
C1074 VDD.n523 GND 0.05fF
C1075 VDD.n524 GND 0.16fF
C1076 VDD.n525 GND 0.01fF
C1077 VDD.n526 GND 0.02fF
C1078 VDD.n527 GND 0.02fF
C1079 VDD.n528 GND 0.18fF
C1080 VDD.n529 GND 0.01fF
C1081 VDD.n530 GND 0.02fF
C1082 VDD.n531 GND 0.02fF
C1083 VDD.n532 GND 0.07fF
C1084 VDD.n533 GND 0.24fF
C1085 VDD.n534 GND 0.01fF
C1086 VDD.n535 GND 0.01fF
C1087 VDD.n536 GND 0.02fF
C1088 VDD.n537 GND 0.29fF
C1089 VDD.n538 GND 0.01fF
C1090 VDD.n539 GND 0.02fF
C1091 VDD.n540 GND 0.02fF
C1092 VDD.n541 GND 0.29fF
C1093 VDD.n542 GND 0.01fF
C1094 VDD.n543 GND 0.02fF
C1095 VDD.n544 GND 0.04fF
C1096 VDD.n545 GND 0.32fF
C1097 VDD.n546 GND 0.02fF
C1098 VDD.n547 GND 0.02fF
C1099 VDD.n548 GND 0.02fF
C1100 VDD.n549 GND 0.06fF
C1101 VDD.n550 GND 0.02fF
C1102 VDD.n551 GND 0.02fF
C1103 VDD.n552 GND 0.02fF
C1104 VDD.n553 GND 0.02fF
C1105 VDD.n554 GND 0.02fF
C1106 VDD.n555 GND 0.02fF
C1107 VDD.n556 GND 0.02fF
C1108 VDD.n557 GND 0.02fF
C1109 VDD.n558 GND 0.02fF
C1110 VDD.n559 GND 0.02fF
C1111 VDD.n560 GND 0.03fF
C1112 VDD.n561 GND 0.02fF
C1113 VDD.n562 GND 0.02fF
C1114 VDD.n566 GND 0.29fF
C1115 VDD.n567 GND 0.29fF
C1116 VDD.n568 GND 0.01fF
C1117 VDD.n569 GND 0.02fF
C1118 VDD.n570 GND 0.04fF
C1119 VDD.n571 GND 0.29fF
C1120 VDD.n572 GND 0.01fF
C1121 VDD.n573 GND 0.02fF
C1122 VDD.n574 GND 0.02fF
C1123 VDD.n575 GND 0.23fF
C1124 VDD.n576 GND 0.01fF
C1125 VDD.n577 GND 0.07fF
C1126 VDD.n578 GND 0.02fF
C1127 VDD.n579 GND 0.18fF
C1128 VDD.n580 GND 0.01fF
C1129 VDD.n581 GND 0.02fF
C1130 VDD.n582 GND 0.02fF
C1131 VDD.n583 GND 0.17fF
C1132 VDD.n584 GND 0.01fF
C1133 VDD.n585 GND 0.08fF
C1134 VDD.n586 GND 0.05fF
C1135 VDD.n587 GND 0.02fF
C1136 VDD.n588 GND 0.02fF
C1137 VDD.n589 GND 0.15fF
C1138 VDD.n590 GND 0.02fF
C1139 VDD.n591 GND 0.02fF
C1140 VDD.n592 GND 0.03fF
C1141 VDD.n593 GND 0.16fF
C1142 VDD.n594 GND 0.02fF
C1143 VDD.n595 GND 0.02fF
C1144 VDD.n596 GND 0.03fF
C1145 VDD.n597 GND 0.08fF
C1146 VDD.n598 GND 0.05fF
C1147 VDD.n599 GND 0.16fF
C1148 VDD.n600 GND 0.01fF
C1149 VDD.n601 GND 0.02fF
C1150 VDD.n602 GND 0.02fF
C1151 VDD.n603 GND 0.18fF
C1152 VDD.n604 GND 0.01fF
C1153 VDD.n605 GND 0.02fF
C1154 VDD.n606 GND 0.02fF
C1155 VDD.n607 GND 0.07fF
C1156 VDD.n608 GND 0.24fF
C1157 VDD.n609 GND 0.01fF
C1158 VDD.n610 GND 0.01fF
C1159 VDD.n611 GND 0.02fF
C1160 VDD.n612 GND 0.29fF
C1161 VDD.n613 GND 0.01fF
C1162 VDD.n614 GND 0.02fF
C1163 VDD.n615 GND 0.02fF
C1164 VDD.n616 GND 0.29fF
C1165 VDD.n617 GND 0.01fF
C1166 VDD.n618 GND 0.02fF
C1167 VDD.n619 GND 0.04fF
C1168 VDD.n620 GND 0.27fF
C1169 VDD.n621 GND 0.02fF
C1170 VDD.n622 GND 0.02fF
C1171 VDD.n623 GND 0.02fF
C1172 VDD.n624 GND 0.06fF
C1173 VDD.n625 GND 0.02fF
C1174 VDD.n626 GND 0.02fF
C1175 VDD.n627 GND 0.02fF
C1176 VDD.n628 GND 0.02fF
C1177 VDD.n629 GND 0.02fF
C1178 VDD.n630 GND 0.02fF
C1179 VDD.n631 GND 0.02fF
C1180 VDD.n632 GND 0.02fF
C1181 VDD.n633 GND 0.02fF
C1182 VDD.n634 GND 0.02fF
C1183 VDD.n635 GND 0.03fF
C1184 VDD.n636 GND 0.02fF
C1185 VDD.n637 GND 0.02fF
C1186 VDD.n641 GND 0.29fF
C1187 VDD.n642 GND 0.29fF
C1188 VDD.n643 GND 0.01fF
C1189 VDD.n644 GND 0.02fF
C1190 VDD.n645 GND 0.04fF
C1191 VDD.n646 GND 0.06fF
C1192 VDD.n647 GND 0.26fF
C1193 VDD.n648 GND 0.01fF
C1194 VDD.n649 GND 0.01fF
C1195 VDD.n650 GND 0.02fF
C1196 VDD.n651 GND 0.18fF
C1197 VDD.n652 GND 0.01fF
C1198 VDD.n653 GND 0.02fF
C1199 VDD.n654 GND 0.02fF
C1200 VDD.n655 GND 0.08fF
C1201 VDD.n656 GND 0.05fF
C1202 VDD.n657 GND 0.01fF
C1203 VDD.n658 GND 0.02fF
C1204 VDD.n659 GND 0.03fF
C1205 VDD.n660 GND 0.15fF
C1206 VDD.n661 GND 0.01fF
C1207 VDD.n662 GND 0.02fF
C1208 VDD.n663 GND 0.03fF
C1209 VDD.n664 GND 0.17fF
C1210 VDD.n665 GND 0.01fF
C1211 VDD.n666 GND 0.02fF
C1212 VDD.n667 GND 0.02fF
C1213 VDD.n668 GND 0.07fF
C1214 VDD.n669 GND 0.26fF
C1215 VDD.n670 GND 0.01fF
C1216 VDD.n671 GND 0.01fF
C1217 VDD.n672 GND 0.02fF
C1218 VDD.n673 GND 0.29fF
C1219 VDD.n674 GND 0.01fF
C1220 VDD.n675 GND 0.02fF
C1221 VDD.n676 GND 0.04fF
C1222 VDD.n677 GND 0.27fF
C1223 VDD.n678 GND 0.02fF
C1224 VDD.n679 GND 0.02fF
C1225 VDD.n680 GND 0.02fF
C1226 VDD.n681 GND 0.06fF
C1227 VDD.n682 GND 0.02fF
C1228 VDD.n683 GND 0.02fF
C1229 VDD.n684 GND 0.02fF
C1230 VDD.n685 GND 0.02fF
C1231 VDD.n686 GND 0.02fF
C1232 VDD.n687 GND 0.02fF
C1233 VDD.n688 GND 0.02fF
C1234 VDD.n689 GND 0.02fF
C1235 VDD.n690 GND 0.02fF
C1236 VDD.n691 GND 0.02fF
C1237 VDD.n692 GND 0.03fF
C1238 VDD.n693 GND 0.02fF
C1239 VDD.n694 GND 0.02fF
C1240 VDD.n698 GND 0.29fF
C1241 VDD.n699 GND 0.29fF
C1242 VDD.n700 GND 0.01fF
C1243 VDD.n701 GND 0.02fF
C1244 VDD.n702 GND 0.04fF
C1245 VDD.n703 GND 0.29fF
C1246 VDD.n704 GND 0.01fF
C1247 VDD.n705 GND 0.02fF
C1248 VDD.n706 GND 0.02fF
C1249 VDD.n707 GND 0.23fF
C1250 VDD.n708 GND 0.01fF
C1251 VDD.n709 GND 0.07fF
C1252 VDD.n710 GND 0.02fF
C1253 VDD.n711 GND 0.18fF
C1254 VDD.n712 GND 0.01fF
C1255 VDD.n713 GND 0.02fF
C1256 VDD.n714 GND 0.02fF
C1257 VDD.n715 GND 0.17fF
C1258 VDD.n716 GND 0.01fF
C1259 VDD.n717 GND 0.08fF
C1260 VDD.n718 GND 0.05fF
C1261 VDD.n719 GND 0.02fF
C1262 VDD.n720 GND 0.02fF
C1263 VDD.n721 GND 0.15fF
C1264 VDD.n722 GND 0.02fF
C1265 VDD.n723 GND 0.02fF
C1266 VDD.n724 GND 0.03fF
C1267 VDD.n725 GND 0.16fF
C1268 VDD.n726 GND 0.02fF
C1269 VDD.n727 GND 0.02fF
C1270 VDD.n728 GND 0.03fF
C1271 VDD.n729 GND 0.08fF
C1272 VDD.n730 GND 0.05fF
C1273 VDD.n731 GND 0.16fF
C1274 VDD.n732 GND 0.01fF
C1275 VDD.n733 GND 0.02fF
C1276 VDD.n734 GND 0.02fF
C1277 VDD.n735 GND 0.18fF
C1278 VDD.n736 GND 0.01fF
C1279 VDD.n737 GND 0.02fF
C1280 VDD.n738 GND 0.02fF
C1281 VDD.n739 GND 0.19fF
C1282 VDD.n740 GND 0.02fF
C1283 VDD.n741 GND 0.02fF
C1284 VDD.n742 GND 0.06fF
C1285 VDD.n743 GND 0.02fF
C1286 VDD.n744 GND 0.02fF
C1287 VDD.n745 GND 0.02fF
C1288 VDD.n746 GND 0.02fF
C1289 VDD.n747 GND 0.02fF
C1290 VDD.n748 GND 0.02fF
C1291 VDD.n749 GND 0.02fF
C1292 VDD.n750 GND 0.02fF
C1293 VDD.n751 GND 0.03fF
C1294 VDD.n752 GND 0.04fF
C1295 VDD.n753 GND 0.02fF
C1296 VDD.n757 GND 0.48fF
C1297 VDD.n758 GND 0.29fF
C1298 VDD.n759 GND 0.02fF
C1299 VDD.n760 GND 0.03fF
C1300 VDD.n761 GND 0.03fF
C1301 VDD.n762 GND 0.29fF
C1302 VDD.n763 GND 0.01fF
C1303 VDD.n764 GND 0.02fF
C1304 VDD.n765 GND 0.02fF
C1305 VDD.n766 GND 0.07fF
C1306 VDD.n767 GND 0.24fF
C1307 VDD.n768 GND 0.01fF
C1308 VDD.n769 GND 0.01fF
C1309 VDD.n770 GND 0.02fF
C1310 VDD.n771 GND 0.18fF
C1311 VDD.n772 GND 0.01fF
C1312 VDD.n773 GND 0.02fF
C1313 VDD.n774 GND 0.02fF
C1314 VDD.n775 GND 0.08fF
C1315 VDD.n776 GND 0.05fF
C1316 VDD.n777 GND 0.16fF
C1317 VDD.n778 GND 0.01fF
C1318 VDD.n779 GND 0.02fF
C1319 VDD.n780 GND 0.02fF
C1320 VDD.n781 GND 0.16fF
C1321 VDD.n782 GND 0.02fF
C1322 VDD.n783 GND 0.02fF
C1323 VDD.n784 GND 0.03fF
C1324 VDD.n785 GND 0.15fF
C1325 VDD.n786 GND 0.02fF
C1326 VDD.n787 GND 0.02fF
C1327 VDD.n788 GND 0.03fF
C1328 VDD.n789 GND 0.17fF
C1329 VDD.n790 GND 0.01fF
C1330 VDD.n791 GND 0.08fF
C1331 VDD.n792 GND 0.05fF
C1332 VDD.n793 GND 0.02fF
C1333 VDD.n794 GND 0.02fF
C1334 VDD.n795 GND 0.18fF
C1335 VDD.n796 GND 0.01fF
C1336 VDD.n797 GND 0.02fF
C1337 VDD.n798 GND 0.02fF
C1338 VDD.n799 GND 0.23fF
C1339 VDD.n800 GND 0.01fF
C1340 VDD.n801 GND 0.07fF
C1341 VDD.n802 GND 0.02fF
C1342 VDD.n803 GND 0.29fF
C1343 VDD.n804 GND 0.01fF
C1344 VDD.n805 GND 0.02fF
C1345 VDD.n806 GND 0.02fF
C1346 VDD.n807 GND 0.29fF
C1347 VDD.n808 GND 0.01fF
C1348 VDD.n809 GND 0.02fF
C1349 VDD.n810 GND 0.04fF
C1350 VDD.n811 GND 0.06fF
C1351 VDD.n812 GND 0.02fF
C1352 VDD.n813 GND 0.02fF
C1353 VDD.n814 GND 0.02fF
C1354 VDD.n815 GND 0.02fF
C1355 VDD.n816 GND 0.02fF
C1356 VDD.n817 GND 0.02fF
C1357 VDD.n818 GND 0.02fF
C1358 VDD.n819 GND 0.02fF
C1359 VDD.n820 GND 0.02fF
C1360 VDD.n821 GND 0.02fF
C1361 VDD.n822 GND 0.02fF
C1362 VDD.n823 GND 0.03fF
C1363 VDD.n824 GND 0.02fF
C1364 VDD.n827 GND 0.02fF
C1365 VDD.n829 GND 0.02fF
C1366 VDD.n830 GND 0.33fF
C1367 VDD.n831 GND 0.02fF
C1368 VDD.n833 GND 0.29fF
C1369 VDD.n834 GND 0.29fF
C1370 VDD.n835 GND 0.01fF
C1371 VDD.n836 GND 0.02fF
C1372 VDD.n837 GND 0.04fF
C1373 VDD.n838 GND 0.29fF
C1374 VDD.n839 GND 0.01fF
C1375 VDD.n840 GND 0.02fF
C1376 VDD.n841 GND 0.02fF
C1377 VDD.n842 GND 0.07fF
C1378 VDD.n843 GND 0.24fF
C1379 VDD.n844 GND 0.01fF
C1380 VDD.n845 GND 0.01fF
C1381 VDD.n846 GND 0.02fF
C1382 VDD.n847 GND 0.18fF
C1383 VDD.n848 GND 0.01fF
C1384 VDD.n849 GND 0.02fF
C1385 VDD.n850 GND 0.02fF
C1386 VDD.n851 GND 0.08fF
C1387 VDD.n852 GND 0.05fF
C1388 VDD.n853 GND 0.16fF
C1389 VDD.n854 GND 0.01fF
C1390 VDD.n855 GND 0.02fF
C1391 VDD.n856 GND 0.02fF
C1392 VDD.n857 GND 0.16fF
C1393 VDD.n858 GND 0.02fF
C1394 VDD.n859 GND 0.02fF
C1395 VDD.n860 GND 0.03fF
C1396 VDD.n861 GND 0.15fF
C1397 VDD.n862 GND 0.02fF
C1398 VDD.n863 GND 0.02fF
C1399 VDD.n864 GND 0.03fF
C1400 VDD.n865 GND 0.17fF
C1401 VDD.n866 GND 0.01fF
C1402 VDD.n867 GND 0.08fF
C1403 VDD.n868 GND 0.05fF
C1404 VDD.n869 GND 0.02fF
C1405 VDD.n870 GND 0.02fF
C1406 VDD.n871 GND 0.18fF
C1407 VDD.n872 GND 0.01fF
C1408 VDD.n873 GND 0.02fF
C1409 VDD.n874 GND 0.02fF
C1410 VDD.n875 GND 0.23fF
C1411 VDD.n876 GND 0.01fF
C1412 VDD.n877 GND 0.07fF
C1413 VDD.n878 GND 0.02fF
C1414 VDD.n879 GND 0.29fF
C1415 VDD.n880 GND 0.01fF
C1416 VDD.n881 GND 0.02fF
C1417 VDD.n882 GND 0.02fF
C1418 VDD.n883 GND 0.29fF
C1419 VDD.n884 GND 0.01fF
C1420 VDD.n885 GND 0.02fF
C1421 VDD.n886 GND 0.04fF
C1422 VDD.n887 GND 0.27fF
C1423 VDD.n888 GND 0.02fF
C1424 VDD.n889 GND 0.02fF
C1425 VDD.n890 GND 0.02fF
C1426 VDD.n891 GND 0.06fF
C1427 VDD.n892 GND 0.02fF
C1428 VDD.n893 GND 0.02fF
C1429 VDD.n894 GND 0.02fF
C1430 VDD.n895 GND 0.02fF
C1431 VDD.n896 GND 0.02fF
C1432 VDD.n897 GND 0.02fF
C1433 VDD.n898 GND 0.02fF
C1434 VDD.n899 GND 0.02fF
C1435 VDD.n900 GND 0.02fF
C1436 VDD.n901 GND 0.02fF
C1437 VDD.n902 GND 0.03fF
C1438 VDD.n903 GND 0.02fF
C1439 VDD.n904 GND 0.02fF
C1440 VDD.n908 GND 0.29fF
C1441 VDD.n909 GND 0.29fF
C1442 VDD.n910 GND 0.01fF
C1443 VDD.n911 GND 0.02fF
C1444 VDD.n912 GND 0.04fF
C1445 VDD.n913 GND 0.07fF
C1446 VDD.n914 GND 0.26fF
C1447 VDD.n915 GND 0.01fF
C1448 VDD.n916 GND 0.01fF
C1449 VDD.n917 GND 0.02fF
C1450 VDD.n918 GND 0.17fF
C1451 VDD.n919 GND 0.01fF
C1452 VDD.n920 GND 0.02fF
C1453 VDD.n921 GND 0.02fF
C1454 VDD.n922 GND 0.15fF
C1455 VDD.n923 GND 0.01fF
C1456 VDD.n924 GND 0.02fF
C1457 VDD.n925 GND 0.03fF
C1458 VDD.n926 GND 0.08fF
C1459 VDD.n927 GND 0.05fF
C1460 VDD.n928 GND 0.01fF
C1461 VDD.n929 GND 0.02fF
C1462 VDD.n930 GND 0.03fF
C1463 VDD.n931 GND 0.18fF
C1464 VDD.n932 GND 0.01fF
C1465 VDD.n933 GND 0.02fF
C1466 VDD.n934 GND 0.02fF
C1467 VDD.n935 GND 0.06fF
C1468 VDD.n936 GND 0.26fF
C1469 VDD.n937 GND 0.01fF
C1470 VDD.n938 GND 0.01fF
C1471 VDD.n939 GND 0.02fF
C1472 VDD.n940 GND 0.29fF
C1473 VDD.n941 GND 0.01fF
C1474 VDD.n942 GND 0.02fF
C1475 VDD.n943 GND 0.04fF
C1476 VDD.n944 GND 0.27fF
C1477 VDD.n945 GND 0.02fF
C1478 VDD.n946 GND 0.02fF
C1479 VDD.n947 GND 0.02fF
C1480 VDD.n948 GND 0.06fF
C1481 VDD.n949 GND 0.02fF
C1482 VDD.n950 GND 0.02fF
C1483 VDD.n951 GND 0.02fF
C1484 VDD.n952 GND 0.02fF
C1485 VDD.n953 GND 0.02fF
C1486 VDD.n954 GND 0.02fF
C1487 VDD.n955 GND 0.02fF
C1488 VDD.n956 GND 0.02fF
C1489 VDD.n957 GND 0.02fF
C1490 VDD.n958 GND 0.02fF
C1491 VDD.n959 GND 0.03fF
C1492 VDD.n960 GND 0.02fF
C1493 VDD.n961 GND 0.02fF
C1494 VDD.n965 GND 0.29fF
C1495 VDD.n966 GND 0.29fF
C1496 VDD.n967 GND 0.01fF
C1497 VDD.n968 GND 0.02fF
C1498 VDD.n969 GND 0.04fF
C1499 VDD.n970 GND 0.29fF
C1500 VDD.n971 GND 0.01fF
C1501 VDD.n972 GND 0.02fF
C1502 VDD.n973 GND 0.02fF
C1503 VDD.n974 GND 0.07fF
C1504 VDD.n975 GND 0.24fF
C1505 VDD.n976 GND 0.01fF
C1506 VDD.n977 GND 0.01fF
C1507 VDD.n978 GND 0.02fF
C1508 VDD.n979 GND 0.18fF
C1509 VDD.n980 GND 0.01fF
C1510 VDD.n981 GND 0.02fF
C1511 VDD.n982 GND 0.02fF
C1512 VDD.n983 GND 0.08fF
C1513 VDD.n984 GND 0.05fF
C1514 VDD.n985 GND 0.16fF
C1515 VDD.n986 GND 0.01fF
C1516 VDD.n987 GND 0.02fF
C1517 VDD.n988 GND 0.02fF
C1518 VDD.n989 GND 0.16fF
C1519 VDD.n990 GND 0.02fF
C1520 VDD.n991 GND 0.02fF
C1521 VDD.n992 GND 0.03fF
C1522 VDD.n993 GND 0.15fF
C1523 VDD.n994 GND 0.02fF
C1524 VDD.n995 GND 0.02fF
C1525 VDD.n996 GND 0.03fF
C1526 VDD.n997 GND 0.17fF
C1527 VDD.n998 GND 0.01fF
C1528 VDD.n999 GND 0.08fF
C1529 VDD.n1000 GND 0.05fF
C1530 VDD.n1001 GND 0.02fF
C1531 VDD.n1002 GND 0.02fF
C1532 VDD.n1003 GND 0.18fF
C1533 VDD.n1004 GND 0.01fF
C1534 VDD.n1005 GND 0.02fF
C1535 VDD.n1006 GND 0.02fF
C1536 VDD.n1007 GND 0.23fF
C1537 VDD.n1008 GND 0.01fF
C1538 VDD.n1009 GND 0.07fF
C1539 VDD.n1010 GND 0.02fF
C1540 VDD.n1011 GND 0.29fF
C1541 VDD.n1012 GND 0.01fF
C1542 VDD.n1013 GND 0.02fF
C1543 VDD.n1014 GND 0.02fF
C1544 VDD.n1015 GND 0.29fF
C1545 VDD.n1016 GND 0.01fF
C1546 VDD.n1017 GND 0.02fF
C1547 VDD.n1018 GND 0.04fF
C1548 VDD.n1019 GND 0.32fF
C1549 VDD.n1020 GND 0.02fF
C1550 VDD.n1021 GND 0.02fF
C1551 VDD.n1022 GND 0.02fF
C1552 VDD.n1023 GND 0.06fF
C1553 VDD.n1024 GND 0.02fF
C1554 VDD.n1025 GND 0.02fF
C1555 VDD.n1026 GND 0.02fF
C1556 VDD.n1027 GND 0.02fF
C1557 VDD.n1028 GND 0.02fF
C1558 VDD.n1029 GND 0.02fF
C1559 VDD.n1030 GND 0.02fF
C1560 VDD.n1031 GND 0.02fF
C1561 VDD.n1032 GND 0.02fF
C1562 VDD.n1033 GND 0.02fF
C1563 VDD.n1034 GND 0.03fF
C1564 VDD.n1035 GND 0.02fF
C1565 VDD.n1036 GND 0.02fF
C1566 VDD.n1040 GND 0.29fF
C1567 VDD.n1041 GND 0.29fF
C1568 VDD.n1042 GND 0.01fF
C1569 VDD.n1043 GND 0.02fF
C1570 VDD.n1044 GND 0.04fF
C1571 VDD.n1045 GND 0.29fF
C1572 VDD.n1046 GND 0.01fF
C1573 VDD.n1047 GND 0.02fF
C1574 VDD.n1048 GND 0.02fF
C1575 VDD.n1049 GND 0.07fF
C1576 VDD.n1050 GND 0.24fF
C1577 VDD.n1051 GND 0.01fF
C1578 VDD.n1052 GND 0.01fF
C1579 VDD.n1053 GND 0.02fF
C1580 VDD.n1054 GND 0.18fF
C1581 VDD.n1055 GND 0.01fF
C1582 VDD.n1056 GND 0.02fF
C1583 VDD.n1057 GND 0.02fF
C1584 VDD.n1058 GND 0.08fF
C1585 VDD.n1059 GND 0.05fF
C1586 VDD.n1060 GND 0.16fF
C1587 VDD.n1061 GND 0.01fF
C1588 VDD.n1062 GND 0.02fF
C1589 VDD.n1063 GND 0.02fF
C1590 VDD.n1064 GND 0.16fF
C1591 VDD.n1065 GND 0.02fF
C1592 VDD.n1066 GND 0.02fF
C1593 VDD.n1067 GND 0.03fF
C1594 VDD.n1068 GND 0.15fF
C1595 VDD.n1069 GND 0.02fF
C1596 VDD.n1070 GND 0.02fF
C1597 VDD.n1071 GND 0.03fF
C1598 VDD.n1072 GND 0.17fF
C1599 VDD.n1073 GND 0.01fF
C1600 VDD.n1074 GND 0.08fF
C1601 VDD.n1075 GND 0.05fF
C1602 VDD.n1076 GND 0.02fF
C1603 VDD.n1077 GND 0.02fF
C1604 VDD.n1078 GND 0.18fF
C1605 VDD.n1079 GND 0.01fF
C1606 VDD.n1080 GND 0.02fF
C1607 VDD.n1081 GND 0.02fF
C1608 VDD.n1082 GND 0.23fF
C1609 VDD.n1083 GND 0.01fF
C1610 VDD.n1084 GND 0.07fF
C1611 VDD.n1085 GND 0.02fF
C1612 VDD.n1086 GND 0.29fF
C1613 VDD.n1087 GND 0.01fF
C1614 VDD.n1088 GND 0.02fF
C1615 VDD.n1089 GND 0.02fF
C1616 VDD.n1090 GND 0.29fF
C1617 VDD.n1091 GND 0.01fF
C1618 VDD.n1092 GND 0.02fF
C1619 VDD.n1093 GND 0.04fF
C1620 VDD.n1094 GND 0.27fF
C1621 VDD.n1095 GND 0.02fF
C1622 VDD.n1096 GND 0.02fF
C1623 VDD.n1097 GND 0.02fF
C1624 VDD.n1098 GND 0.06fF
C1625 VDD.n1099 GND 0.02fF
C1626 VDD.n1100 GND 0.02fF
C1627 VDD.n1101 GND 0.02fF
C1628 VDD.n1102 GND 0.02fF
C1629 VDD.n1103 GND 0.02fF
C1630 VDD.n1104 GND 0.02fF
C1631 VDD.n1105 GND 0.02fF
C1632 VDD.n1106 GND 0.02fF
C1633 VDD.n1107 GND 0.02fF
C1634 VDD.n1108 GND 0.02fF
C1635 VDD.n1109 GND 0.03fF
C1636 VDD.n1110 GND 0.02fF
C1637 VDD.n1111 GND 0.02fF
C1638 VDD.n1115 GND 0.29fF
C1639 VDD.n1116 GND 0.29fF
C1640 VDD.n1117 GND 0.01fF
C1641 VDD.n1118 GND 0.02fF
C1642 VDD.n1119 GND 0.04fF
C1643 VDD.n1120 GND 0.07fF
C1644 VDD.n1121 GND 0.26fF
C1645 VDD.n1122 GND 0.01fF
C1646 VDD.n1123 GND 0.01fF
C1647 VDD.n1124 GND 0.02fF
C1648 VDD.n1125 GND 0.17fF
C1649 VDD.n1126 GND 0.01fF
C1650 VDD.n1127 GND 0.02fF
C1651 VDD.n1128 GND 0.02fF
C1652 VDD.n1129 GND 0.15fF
C1653 VDD.n1130 GND 0.01fF
C1654 VDD.n1131 GND 0.02fF
C1655 VDD.n1132 GND 0.03fF
C1656 VDD.n1133 GND 0.08fF
C1657 VDD.n1134 GND 0.05fF
C1658 VDD.n1135 GND 0.01fF
C1659 VDD.n1136 GND 0.02fF
C1660 VDD.n1137 GND 0.03fF
C1661 VDD.n1138 GND 0.18fF
C1662 VDD.n1139 GND 0.01fF
C1663 VDD.n1140 GND 0.02fF
C1664 VDD.n1141 GND 0.02fF
C1665 VDD.n1142 GND 0.06fF
C1666 VDD.n1143 GND 0.26fF
C1667 VDD.n1144 GND 0.01fF
C1668 VDD.n1145 GND 0.01fF
C1669 VDD.n1146 GND 0.02fF
C1670 VDD.n1147 GND 0.29fF
C1671 VDD.n1148 GND 0.01fF
C1672 VDD.n1149 GND 0.02fF
C1673 VDD.n1150 GND 0.04fF
C1674 VDD.n1151 GND 0.27fF
C1675 VDD.n1152 GND 0.02fF
C1676 VDD.n1153 GND 0.02fF
C1677 VDD.n1154 GND 0.02fF
C1678 VDD.n1155 GND 0.06fF
C1679 VDD.n1156 GND 0.02fF
C1680 VDD.n1157 GND 0.02fF
C1681 VDD.n1158 GND 0.02fF
C1682 VDD.n1159 GND 0.02fF
C1683 VDD.n1160 GND 0.02fF
C1684 VDD.n1161 GND 0.02fF
C1685 VDD.n1162 GND 0.02fF
C1686 VDD.n1163 GND 0.02fF
C1687 VDD.n1164 GND 0.02fF
C1688 VDD.n1165 GND 0.02fF
C1689 VDD.n1166 GND 0.03fF
C1690 VDD.n1167 GND 0.02fF
C1691 VDD.n1168 GND 0.02fF
C1692 VDD.n1172 GND 0.29fF
C1693 VDD.n1173 GND 0.29fF
C1694 VDD.n1174 GND 0.01fF
C1695 VDD.n1175 GND 0.02fF
C1696 VDD.n1176 GND 0.04fF
C1697 VDD.n1177 GND 0.29fF
C1698 VDD.n1178 GND 0.01fF
C1699 VDD.n1179 GND 0.02fF
C1700 VDD.n1180 GND 0.02fF
C1701 VDD.n1181 GND 0.07fF
C1702 VDD.n1182 GND 0.24fF
C1703 VDD.n1183 GND 0.01fF
C1704 VDD.n1184 GND 0.01fF
C1705 VDD.n1185 GND 0.02fF
C1706 VDD.n1186 GND 0.18fF
C1707 VDD.n1187 GND 0.01fF
C1708 VDD.n1188 GND 0.02fF
C1709 VDD.n1189 GND 0.02fF
C1710 VDD.n1190 GND 0.08fF
C1711 VDD.n1191 GND 0.05fF
C1712 VDD.n1192 GND 0.16fF
C1713 VDD.n1193 GND 0.01fF
C1714 VDD.n1194 GND 0.02fF
C1715 VDD.n1195 GND 0.02fF
C1716 VDD.n1196 GND 0.16fF
C1717 VDD.n1197 GND 0.02fF
C1718 VDD.n1198 GND 0.02fF
C1719 VDD.n1199 GND 0.03fF
C1720 VDD.n1200 GND 0.15fF
C1721 VDD.n1201 GND 0.02fF
C1722 VDD.n1202 GND 0.02fF
C1723 VDD.n1203 GND 0.03fF
C1724 VDD.n1204 GND 0.17fF
C1725 VDD.n1205 GND 0.01fF
C1726 VDD.n1206 GND 0.08fF
C1727 VDD.n1207 GND 0.05fF
C1728 VDD.n1208 GND 0.02fF
C1729 VDD.n1209 GND 0.02fF
C1730 VDD.n1210 GND 0.18fF
C1731 VDD.n1211 GND 0.01fF
C1732 VDD.n1212 GND 0.02fF
C1733 VDD.n1213 GND 0.02fF
C1734 VDD.n1214 GND 0.23fF
C1735 VDD.n1215 GND 0.01fF
C1736 VDD.n1216 GND 0.07fF
C1737 VDD.n1217 GND 0.02fF
C1738 VDD.n1218 GND 0.29fF
C1739 VDD.n1219 GND 0.01fF
C1740 VDD.n1220 GND 0.02fF
C1741 VDD.n1221 GND 0.02fF
C1742 VDD.n1222 GND 0.29fF
C1743 VDD.n1223 GND 0.01fF
C1744 VDD.n1224 GND 0.02fF
C1745 VDD.n1225 GND 0.04fF
C1746 VDD.n1226 GND 0.32fF
C1747 VDD.n1227 GND 0.02fF
C1748 VDD.n1228 GND 0.02fF
C1749 VDD.n1229 GND 0.02fF
C1750 VDD.n1230 GND 0.06fF
C1751 VDD.n1231 GND 0.02fF
C1752 VDD.n1232 GND 0.02fF
C1753 VDD.n1233 GND 0.02fF
C1754 VDD.n1234 GND 0.02fF
C1755 VDD.n1235 GND 0.02fF
C1756 VDD.n1236 GND 0.02fF
C1757 VDD.n1237 GND 0.02fF
C1758 VDD.n1238 GND 0.02fF
C1759 VDD.n1239 GND 0.02fF
C1760 VDD.n1240 GND 0.02fF
C1761 VDD.n1241 GND 0.03fF
C1762 VDD.n1242 GND 0.02fF
C1763 VDD.n1243 GND 0.02fF
C1764 VDD.n1247 GND 0.29fF
C1765 VDD.n1248 GND 0.29fF
C1766 VDD.n1249 GND 0.01fF
C1767 VDD.n1250 GND 0.02fF
C1768 VDD.n1251 GND 0.04fF
C1769 VDD.n1252 GND 0.29fF
C1770 VDD.n1253 GND 0.01fF
C1771 VDD.n1254 GND 0.02fF
C1772 VDD.n1255 GND 0.02fF
C1773 VDD.n1256 GND 0.07fF
C1774 VDD.n1257 GND 0.24fF
C1775 VDD.n1258 GND 0.01fF
C1776 VDD.n1259 GND 0.01fF
C1777 VDD.n1260 GND 0.02fF
C1778 VDD.n1261 GND 0.18fF
C1779 VDD.n1262 GND 0.01fF
C1780 VDD.n1263 GND 0.02fF
C1781 VDD.n1264 GND 0.02fF
C1782 VDD.n1265 GND 0.08fF
C1783 VDD.n1266 GND 0.05fF
C1784 VDD.n1267 GND 0.16fF
C1785 VDD.n1268 GND 0.01fF
C1786 VDD.n1269 GND 0.02fF
C1787 VDD.n1270 GND 0.02fF
C1788 VDD.n1271 GND 0.16fF
C1789 VDD.n1272 GND 0.02fF
C1790 VDD.n1273 GND 0.02fF
C1791 VDD.n1274 GND 0.03fF
C1792 VDD.n1275 GND 0.15fF
C1793 VDD.n1276 GND 0.02fF
C1794 VDD.n1277 GND 0.02fF
C1795 VDD.n1278 GND 0.03fF
C1796 VDD.n1279 GND 0.17fF
C1797 VDD.n1280 GND 0.01fF
C1798 VDD.n1281 GND 0.08fF
C1799 VDD.n1282 GND 0.05fF
C1800 VDD.n1283 GND 0.02fF
C1801 VDD.n1284 GND 0.02fF
C1802 VDD.n1285 GND 0.18fF
C1803 VDD.n1286 GND 0.01fF
C1804 VDD.n1287 GND 0.02fF
C1805 VDD.n1288 GND 0.02fF
C1806 VDD.n1289 GND 0.23fF
C1807 VDD.n1290 GND 0.01fF
C1808 VDD.n1291 GND 0.07fF
C1809 VDD.n1292 GND 0.02fF
C1810 VDD.n1293 GND 0.29fF
C1811 VDD.n1294 GND 0.01fF
C1812 VDD.n1295 GND 0.02fF
C1813 VDD.n1296 GND 0.02fF
C1814 VDD.n1297 GND 0.29fF
C1815 VDD.n1298 GND 0.01fF
C1816 VDD.n1299 GND 0.02fF
C1817 VDD.n1300 GND 0.04fF
C1818 VDD.n1301 GND 0.27fF
C1819 VDD.n1302 GND 0.02fF
C1820 VDD.n1303 GND 0.02fF
C1821 VDD.n1304 GND 0.02fF
C1822 VDD.n1305 GND 0.06fF
C1823 VDD.n1306 GND 0.02fF
C1824 VDD.n1307 GND 0.02fF
C1825 VDD.n1308 GND 0.02fF
C1826 VDD.n1309 GND 0.02fF
C1827 VDD.n1310 GND 0.02fF
C1828 VDD.n1311 GND 0.02fF
C1829 VDD.n1312 GND 0.02fF
C1830 VDD.n1313 GND 0.02fF
C1831 VDD.n1314 GND 0.02fF
C1832 VDD.n1315 GND 0.02fF
C1833 VDD.n1316 GND 0.03fF
C1834 VDD.n1317 GND 0.02fF
C1835 VDD.n1318 GND 0.02fF
C1836 VDD.n1322 GND 0.29fF
C1837 VDD.n1323 GND 0.29fF
C1838 VDD.n1324 GND 0.01fF
C1839 VDD.n1325 GND 0.02fF
C1840 VDD.n1326 GND 0.04fF
C1841 VDD.n1327 GND 0.07fF
C1842 VDD.n1328 GND 0.26fF
C1843 VDD.n1329 GND 0.01fF
C1844 VDD.n1330 GND 0.01fF
C1845 VDD.n1331 GND 0.02fF
C1846 VDD.n1332 GND 0.17fF
C1847 VDD.n1333 GND 0.01fF
C1848 VDD.n1334 GND 0.02fF
C1849 VDD.n1335 GND 0.02fF
C1850 VDD.n1336 GND 0.15fF
C1851 VDD.n1337 GND 0.01fF
C1852 VDD.n1338 GND 0.02fF
C1853 VDD.n1339 GND 0.03fF
C1854 VDD.n1340 GND 0.08fF
C1855 VDD.n1341 GND 0.05fF
C1856 VDD.n1342 GND 0.01fF
C1857 VDD.n1343 GND 0.02fF
C1858 VDD.n1344 GND 0.03fF
C1859 VDD.n1345 GND 0.18fF
C1860 VDD.n1346 GND 0.01fF
C1861 VDD.n1347 GND 0.02fF
C1862 VDD.n1348 GND 0.02fF
C1863 VDD.n1349 GND 0.06fF
C1864 VDD.n1350 GND 0.26fF
C1865 VDD.n1351 GND 0.01fF
C1866 VDD.n1352 GND 0.01fF
C1867 VDD.n1353 GND 0.02fF
C1868 VDD.n1354 GND 0.29fF
C1869 VDD.n1355 GND 0.01fF
C1870 VDD.n1356 GND 0.02fF
C1871 VDD.n1357 GND 0.04fF
C1872 VDD.n1358 GND 0.27fF
C1873 VDD.n1359 GND 0.02fF
C1874 VDD.n1360 GND 0.02fF
C1875 VDD.n1361 GND 0.02fF
C1876 VDD.n1362 GND 0.06fF
C1877 VDD.n1363 GND 0.02fF
C1878 VDD.n1364 GND 0.02fF
C1879 VDD.n1365 GND 0.02fF
C1880 VDD.n1366 GND 0.02fF
C1881 VDD.n1367 GND 0.02fF
C1882 VDD.n1368 GND 0.02fF
C1883 VDD.n1369 GND 0.02fF
C1884 VDD.n1370 GND 0.02fF
C1885 VDD.n1371 GND 0.02fF
C1886 VDD.n1372 GND 0.02fF
C1887 VDD.n1373 GND 0.03fF
C1888 VDD.n1374 GND 0.02fF
C1889 