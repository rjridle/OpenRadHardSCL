* SPICE3 file created from DLATCH.ext - technology: sky130A

.subckt DLATCH Q D GATE VDD GND
X0 GND a_185_209.t3 a_556_101.t0 GND sky130_fd_pr__nfet_01v8 ad=7.6538p pd=5.332u as=0p ps=0u w=0u l=0u
X1 VDD.t29 a_1771_1050.t5 a_2405_209.t0 ����U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X2 VDD.t20 D.t0 a_1771_1050.t2 ���U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X3 a_185_209.t2 D.t1 VDD.t18 0�N�U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X4 a_1295_209.t2 a_661_1050.t5 VDD.t35  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X5 a_661_1050.t0 GATE.t0 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X6 a_1771_1050.t4 D.t3 VDD.t39  ��B sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X7 Q.t2 a_3007_411.t5 a_2795_1051.t3 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X8 a_3461_1051.t3 a_2405_209.t3 a_3007_411.t1  ��B sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X9 a_661_1050.t3 a_185_209.t4 VDD.t22 ��B sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X10 a_1771_1050.t0 GATE.t1 VDD.t6  ��B sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X11 a_2795_1051.t1 a_1295_209.t3 VDD.t12 ��B sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X12 VDD.t14 Q.t4 a_3461_1051.t1  ��B sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X13 a_2405_209.t2 a_1771_1050.t6 VDD.t27 ��B sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X14 GND GATE.t4 a_1666_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X15 VDD.t10 a_185_209.t5 a_661_1050.t2  ��B sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X16 VDD.t8 GATE.t3 a_1771_1050.t1 ��B sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X17 VDD.t33 D.t5 a_185_209.t1  ��B sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X18 VDD.t25 a_661_1050.t6 a_1295_209.t1 ��B sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X19 a_3007_411.t2 a_2405_209.t4 a_3461_1051.t2  ��B sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X20 Q a_1295_209.t4 GND.t3 GND sky130_fd_pr__nfet_01v8 ad=3.582p pd=3.15u as=0p ps=0u w=0u l=0u
X21 a_2795_1051.t2 a_3007_411.t6 Q.t1 ��B sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X22 a_3461_1051.t0 Q.t6 VDD.t1  ��B sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X23 Q a_3007_411.t4 GND.t5 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X24 VDD.t31 GATE.t5 a_661_1050.t4 ��B sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X25 VDD.t16 a_1295_209.t5 a_2795_1051.t0  ��B sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
C0 Q VDD 0.85fF
C1 GATE D 0.58fF
C2 D VDD 0.73fF
C3 GATE VDD 0.64fF
R0 a_1771_1050.n3 a_1771_1050.t5 512.525
R1 a_1771_1050.n3 a_1771_1050.t6 371.139
R2 a_1771_1050.n7 a_1771_1050.n5 284.244
R3 a_1771_1050.n4 a_1771_1050.t7 282.852
R4 a_1771_1050.n4 a_1771_1050.n3 247.347
R5 a_1771_1050.n5 a_1771_1050.n2 187.858
R6 a_1771_1050.n2 a_1771_1050.n1 157.964
R7 a_1771_1050.n2 a_1771_1050.n0 91.706
R8 a_1771_1050.n7 a_1771_1050.n6 15.218
R9 a_1771_1050.n0 a_1771_1050.t2 14.282
R10 a_1771_1050.n0 a_1771_1050.t4 14.282
R11 a_1771_1050.n1 a_1771_1050.t1 14.282
R12 a_1771_1050.n1 a_1771_1050.t0 14.282
R13 a_1771_1050.n8 a_1771_1050.n7 12.014
R14 a_1771_1050.n5 a_1771_1050.n4 10.343
R15 a_2405_209.n2 a_2405_209.t3 470.752
R16 a_2405_209.n2 a_2405_209.t4 384.527
R17 a_2405_209.n3 a_2405_209.t5 342.755
R18 a_2405_209.n6 a_2405_209.n4 328.169
R19 a_2405_209.n4 a_2405_209.n1 215.564
R20 a_2405_209.n3 a_2405_209.n2 155.073
R21 a_2405_209.n6 a_2405_209.n5 30
R22 a_2405_209.n7 a_2405_209.n0 24.383
R23 a_2405_209.n7 a_2405_209.n6 23.684
R24 a_2405_209.n1 a_2405_209.t0 14.282
R25 a_2405_209.n1 a_2405_209.t2 14.282
R26 a_2405_209.n4 a_2405_209.n3 13.607
R27 VDD.n240 VDD.n229 144.705
R28 VDD.n294 VDD.n287 144.705
R29 VDD.n176 VDD.n169 144.705
R30 VDD.n354 VDD.n347 144.705
R31 VDD.n132 VDD.n125 144.705
R32 VDD.n77 VDD.n66 144.705
R33 VDD.n280 VDD.t31 143.754
R34 VDD.n179 VDD.t20 143.754
R35 VDD.n213 VDD.t18 135.17
R36 VDD.n220 VDD.t33 135.17
R37 VDD.n256 VDD.t22 135.17
R38 VDD.n313 VDD.t35 135.17
R39 VDD.n322 VDD.t25 135.17
R40 VDD.n357 VDD.t6 135.17
R41 VDD.n146 VDD.t27 135.17
R42 VDD.n135 VDD.t29 135.17
R43 VDD.n96 VDD.n95 129.849
R44 VDD.n40 VDD.n39 129.849
R45 VDD.n271 VDD.n270 129.472
R46 VDD.n371 VDD.n370 129.472
R47 VDD.n62 VDD.n61 92.5
R48 VDD.n60 VDD.n59 92.5
R49 VDD.n58 VDD.n57 92.5
R50 VDD.n56 VDD.n55 92.5
R51 VDD.n64 VDD.n63 92.5
R52 VDD.n121 VDD.n120 92.5
R53 VDD.n119 VDD.n118 92.5
R54 VDD.n117 VDD.n116 92.5
R55 VDD.n115 VDD.n114 92.5
R56 VDD.n123 VDD.n122 92.5
R57 VDD.n165 VDD.n164 92.5
R58 VDD.n163 VDD.n162 92.5
R59 VDD.n161 VDD.n160 92.5
R60 VDD.n159 VDD.n158 92.5
R61 VDD.n167 VDD.n166 92.5
R62 VDD.n343 VDD.n342 92.5
R63 VDD.n341 VDD.n340 92.5
R64 VDD.n339 VDD.n338 92.5
R65 VDD.n337 VDD.n336 92.5
R66 VDD.n345 VDD.n344 92.5
R67 VDD.n307 VDD.n306 92.5
R68 VDD.n305 VDD.n304 92.5
R69 VDD.n303 VDD.n302 92.5
R70 VDD.n301 VDD.n300 92.5
R71 VDD.n309 VDD.n308 92.5
R72 VDD.n250 VDD.n249 92.5
R73 VDD.n248 VDD.n247 92.5
R74 VDD.n246 VDD.n245 92.5
R75 VDD.n244 VDD.n243 92.5
R76 VDD.n252 VDD.n251 92.5
R77 VDD.n199 VDD.n198 92.5
R78 VDD.n197 VDD.n196 92.5
R79 VDD.n195 VDD.n194 92.5
R80 VDD.n193 VDD.n192 92.5
R81 VDD.n201 VDD.n200 92.5
R82 VDD.n14 VDD.n1 92.5
R83 VDD.n5 VDD.n4 92.5
R84 VDD.n7 VDD.n6 92.5
R85 VDD.n9 VDD.n8 92.5
R86 VDD.n11 VDD.n10 92.5
R87 VDD.n13 VDD.n12 92.5
R88 VDD.n21 VDD.n20 92.059
R89 VDD.n76 VDD.n75 92.059
R90 VDD.n131 VDD.n130 92.059
R91 VDD.n175 VDD.n174 92.059
R92 VDD.n353 VDD.n352 92.059
R93 VDD.n293 VDD.n292 92.059
R94 VDD.n239 VDD.n238 92.059
R95 VDD.n207 VDD.n206 92.059
R96 VDD.n20 VDD.n16 67.194
R97 VDD.n20 VDD.n17 67.194
R98 VDD.n20 VDD.n18 67.194
R99 VDD.n20 VDD.n19 67.194
R100 VDD.n191 VDD.n190 44.141
R101 VDD.n299 VDD.n298 44.141
R102 VDD.n335 VDD.n334 44.141
R103 VDD.n157 VDD.n156 44.141
R104 VDD.n113 VDD.n112 44.141
R105 VDD.n5 VDD.n3 44.141
R106 VDD.n298 VDD.n296 44.107
R107 VDD.n334 VDD.n332 44.107
R108 VDD.n156 VDD.n154 44.107
R109 VDD.n112 VDD.n110 44.107
R110 VDD.n190 VDD.n188 44.107
R111 VDD.n3 VDD.n2 44.107
R112 VDD.n136 ����U 43.472
R113 VDD.n144 ��B 43.472
R114 VDD.n323 ��B 43.472
R115 VDD.n314 �!��U 43.472
R116 VDD.n221  ��B 43.472
R117 VDD.n211 0�N�U 43.472
R118 VDD.n20 VDD.n15 41.052
R119 VDD.n70 VDD.n68 39.742
R120 VDD.n70 VDD.n69 39.742
R121 VDD.n72 VDD.n71 39.742
R122 VDD.n127 VDD.n126 39.742
R123 VDD.n171 VDD.n170 39.742
R124 VDD.n349 VDD.n348 39.742
R125 VDD.n289 VDD.n288 39.742
R126 VDD.n203 VDD.n202 39.742
R127 VDD.n237 VDD.n234 39.742
R128 VDD.n237 VDD.n236 39.742
R129 VDD.n233 VDD.n232 39.742
R130 VDD.n112 VDD.n111 38
R131 VDD.n156 VDD.n155 38
R132 VDD.n334 VDD.n333 38
R133 VDD.n298 VDD.n297 38
R134 VDD.n190 VDD.n189 38
R135 VDD.n296 VDD.n295 36.774
R136 VDD.n332 VDD.n331 36.774
R137 VDD.n154 VDD.n153 36.774
R138 VDD.n110 VDD.n109 36.774
R139 VDD.n68 VDD.n67 36.774
R140 VDD.n236 VDD.n235 36.774
R141 VDD.n1 VDD.n0 30.923
R142 VDD.n75 VDD.n73 26.38
R143 VDD.n75 VDD.n72 26.38
R144 VDD.n75 VDD.n70 26.38
R145 VDD.n75 VDD.n74 26.38
R146 VDD.n130 VDD.n128 26.38
R147 VDD.n130 VDD.n127 26.38
R148 VDD.n130 VDD.n129 26.38
R149 VDD.n174 VDD.n172 26.38
R150 VDD.n174 VDD.n171 26.38
R151 VDD.n174 VDD.n173 26.38
R152 VDD.n352 VDD.n350 26.38
R153 VDD.n352 VDD.n349 26.38
R154 VDD.n352 VDD.n351 26.38
R155 VDD.n292 VDD.n290 26.38
R156 VDD.n292 VDD.n289 26.38
R157 VDD.n292 VDD.n291 26.38
R158 VDD.n206 VDD.n204 26.38
R159 VDD.n206 VDD.n203 26.38
R160 VDD.n206 VDD.n205 26.38
R161 VDD.n238 VDD.n237 26.38
R162 VDD.n238 VDD.n233 26.38
R163 VDD.n238 VDD.n231 26.38
R164 VDD.n238 VDD.n230 26.38
R165 VDD.n209 VDD.n201 22.915
R166 VDD.n23 VDD.n14 22.915
R167 VDD.n28  ��B 20.457
R168 VDD.n84 ��B 20.457
R169 VDD.n184 ���U 20.457
R170 VDD.n274 ��B 20.457
R171 VDD.n41  ��B 17.9
R172 VDD.n97  ��B 17.9
R173 VDD.n362  ��B 17.9
R174 VDD.n261 ��B 17.9
R175 VDD.n201 VDD.n199 14.864
R176 VDD.n199 VDD.n197 14.864
R177 VDD.n197 VDD.n195 14.864
R178 VDD.n195 VDD.n193 14.864
R179 VDD.n193 VDD.n191 14.864
R180 VDD.n309 VDD.n307 14.864
R181 VDD.n307 VDD.n305 14.864
R182 VDD.n305 VDD.n303 14.864
R183 VDD.n303 VDD.n301 14.864
R184 VDD.n301 VDD.n299 14.864
R185 VDD.n345 VDD.n343 14.864
R186 VDD.n343 VDD.n341 14.864
R187 VDD.n341 VDD.n339 14.864
R188 VDD.n339 VDD.n337 14.864
R189 VDD.n337 VDD.n335 14.864
R190 VDD.n167 VDD.n165 14.864
R191 VDD.n165 VDD.n163 14.864
R192 VDD.n163 VDD.n161 14.864
R193 VDD.n161 VDD.n159 14.864
R194 VDD.n159 VDD.n157 14.864
R195 VDD.n123 VDD.n121 14.864
R196 VDD.n121 VDD.n119 14.864
R197 VDD.n119 VDD.n117 14.864
R198 VDD.n117 VDD.n115 14.864
R199 VDD.n115 VDD.n113 14.864
R200 VDD.n64 VDD.n62 14.864
R201 VDD.n62 VDD.n60 14.864
R202 VDD.n60 VDD.n58 14.864
R203 VDD.n58 VDD.n56 14.864
R204 VDD.n56 VDD.n54 14.864
R205 VDD.n54 VDD.n53 14.864
R206 VDD.n252 VDD.n250 14.864
R207 VDD.n250 VDD.n248 14.864
R208 VDD.n248 VDD.n246 14.864
R209 VDD.n246 VDD.n244 14.864
R210 VDD.n244 VDD.n242 14.864
R211 VDD.n242 VDD.n241 14.864
R212 VDD.n14 VDD.n13 14.864
R213 VDD.n13 VDD.n11 14.864
R214 VDD.n11 VDD.n9 14.864
R215 VDD.n9 VDD.n7 14.864
R216 VDD.n7 VDD.n5 14.864
R217 VDD.n78 VDD.n65 14.864
R218 VDD.n133 VDD.n124 14.864
R219 VDD.n177 VDD.n168 14.864
R220 VDD.n355 VDD.n346 14.864
R221 VDD.n311 VDD.n310 14.864
R222 VDD.n254 VDD.n253 14.864
R223 VDD.n270 VDD.t3 14.282
R224 VDD.n270 VDD.t10 14.282
R225 VDD.n370 VDD.t39 14.282
R226 VDD.n370 VDD.t8 14.282
R227 VDD.n95 VDD.t12 14.282
R228 VDD.n95 VDD.t16 14.282
R229 VDD.n39 VDD.t1 14.282
R230 VDD.n39 VDD.t14 14.282
R231 VDD.n373 VDD.n371 9.083
R232 VDD.n272 VDD.n271 9.083
R233 VDD.n23 VDD.n22 8.855
R234 VDD.n22 VDD.n21 8.855
R235 VDD.n26 VDD.n25 8.855
R236 VDD.n25 VDD.n24 8.855
R237 VDD.n30 VDD.n29 8.855
R238 VDD.n29 VDD.n28 8.855
R239 VDD.n33 VDD.n32 8.855
R240 VDD.n32  ��B 8.855
R241 VDD.n37 VDD.n36 8.855
R242 VDD.n36 VDD.n35 8.855
R243 VDD.n43 VDD.n42 8.855
R244 VDD.n42 VDD.n41 8.855
R245 VDD.n47 VDD.n46 8.855
R246 VDD.n46 VDD.n45 8.855
R247 VDD.n51 VDD.n50 8.855
R248 VDD.n50 VDD.n49 8.855
R249 VDD.n78 VDD.n77 8.855
R250 VDD.n77 VDD.n76 8.855
R251 VDD.n82 VDD.n81 8.855
R252 VDD.n81 VDD.n80 8.855
R253 VDD.n86 VDD.n85 8.855
R254 VDD.n85 VDD.n84 8.855
R255 VDD.n89 VDD.n88 8.855
R256 VDD.n88 VDD.t4 8.855
R257 VDD.n93 VDD.n92 8.855
R258 VDD.n92 VDD.n91 8.855
R259 VDD.n99 VDD.n98 8.855
R260 VDD.n98 VDD.n97 8.855
R261 VDD.n103 VDD.n102 8.855
R262 VDD.n102 VDD.n101 8.855
R263 VDD.n107 VDD.n106 8.855
R264 VDD.n106 VDD.n105 8.855
R265 VDD.n133 VDD.n132 8.855
R266 VDD.n132 VDD.n131 8.855
R267 VDD.n138 VDD.n137 8.855
R268 VDD.n137 VDD.n136 8.855
R269 VDD.n142 VDD.n141 8.855
R270 VDD.n141 VDD.n140 8.855
R271 VDD.n147 VDD.n145 8.855
R272 VDD.n145 VDD.n144 8.855
R273 VDD.n151 VDD.n150 8.855
R274 VDD.n150 VDD.n149 8.855
R275 VDD.n177 VDD.n176 8.855
R276 VDD.n176 VDD.n175 8.855
R277 VDD.n182 VDD.n181 8.855
R278 VDD.n181 VDD.n180 8.855
R279 VDD.n186 VDD.n185 8.855
R280 VDD.n185 VDD.n184 8.855
R281 VDD.n373 VDD.n372 8.855
R282 VDD.n372  ��B 8.855
R283 VDD.n368 VDD.n367 8.855
R284 VDD.n367 VDD.n366 8.855
R285 VDD.n364 VDD.n363 8.855
R286 VDD.n363 VDD.n362 8.855
R287 VDD.n360 VDD.n359 8.855
R288 VDD.n359 VDD.n358 8.855
R289 VDD.n355 VDD.n354 8.855
R290 VDD.n354 VDD.n353 8.855
R291 VDD.n329 VDD.n328 8.855
R292 VDD.n328 VDD.n327 8.855
R293 VDD.n325 VDD.n324 8.855
R294 VDD.n324 VDD.n323 8.855
R295 VDD.n320 VDD.n319 8.855
R296 VDD.n319 VDD.n318 8.855
R297 VDD.n316 VDD.n315 8.855
R298 VDD.n315 VDD.n314 8.855
R299 VDD.n311 VDD.n294 8.855
R300 VDD.n294 VDD.n293 8.855
R301 VDD.n285 VDD.n284 8.855
R302 VDD.n284 VDD.n283 8.855
R303 VDD.n281 VDD.n279 8.855
R304 VDD.n279 VDD.n278 8.855
R305 VDD.n276 VDD.n275 8.855
R306 VDD.n275 VDD.n274 8.855
R307 VDD.n272 VDD.n269 8.855
R308 VDD.n269 VDD.t2 8.855
R309 VDD.n267 VDD.n266 8.855
R310 VDD.n266 VDD.n265 8.855
R311 VDD.n263 VDD.n262 8.855
R312 VDD.n262 VDD.n261 8.855
R313 VDD.n259 VDD.n258 8.855
R314 VDD.n258 VDD.n257 8.855
R315 VDD.n254 VDD.n240 8.855
R316 VDD.n240 VDD.n239 8.855
R317 VDD.n227 VDD.n226 8.855
R318 VDD.n226 VDD.n225 8.855
R319 VDD.n223 VDD.n222 8.855
R320 VDD.n222 VDD.n221 8.855
R321 VDD.n218 VDD.n217 8.855
R322 VDD.n217 VDD.n216 8.855
R323 VDD.n214 VDD.n212 8.855
R324 VDD.n212 VDD.n211 8.855
R325 VDD.n209 VDD.n208 8.855
R326 VDD.n208 VDD.n207 8.855
R327 VDD.n310 VDD.n309 8.051
R328 VDD.n346 VDD.n345 8.051
R329 VDD.n168 VDD.n167 8.051
R330 VDD.n124 VDD.n123 8.051
R331 VDD.n65 VDD.n64 8.051
R332 VDD.n253 VDD.n252 8.051
R333 VDD.n43 VDD.n40 6.193
R334 VDD.n99 VDD.n96 6.193
R335 VDD.n31 VDD.n30 4.65
R336 VDD.n34 VDD.n33 4.65
R337 VDD.n38 VDD.n37 4.65
R338 VDD.n44 VDD.n43 4.65
R339 VDD.n48 VDD.n47 4.65
R340 VDD.n52 VDD.n51 4.65
R341 VDD.n79 VDD.n78 4.65
R342 VDD.n83 VDD.n82 4.65
R343 VDD.n87 VDD.n86 4.65
R344 VDD.n90 VDD.n89 4.65
R345 VDD.n94 VDD.n93 4.65
R346 VDD.n100 VDD.n99 4.65
R347 VDD.n104 VDD.n103 4.65
R348 VDD.n108 VDD.n107 4.65
R349 VDD.n134 VDD.n133 4.65
R350 VDD.n139 VDD.n138 4.65
R351 VDD.n143 VDD.n142 4.65
R352 VDD.n148 VDD.n147 4.65
R353 VDD.n152 VDD.n151 4.65
R354 VDD.n178 VDD.n177 4.65
R355 VDD.n183 VDD.n182 4.65
R356 VDD.n187 VDD.n186 4.65
R357 VDD.n374 VDD.n373 4.65
R358 VDD.n369 VDD.n368 4.65
R359 VDD.n365 VDD.n364 4.65
R360 VDD.n361 VDD.n360 4.65
R361 VDD.n356 VDD.n355 4.65
R362 VDD.n330 VDD.n329 4.65
R363 VDD.n326 VDD.n325 4.65
R364 VDD.n321 VDD.n320 4.65
R365 VDD.n317 VDD.n316 4.65
R366 VDD.n312 VDD.n311 4.65
R367 VDD.n286 VDD.n285 4.65
R368 VDD.n282 VDD.n281 4.65
R369 VDD.n277 VDD.n276 4.65
R370 VDD.n273 VDD.n272 4.65
R371 VDD.n268 VDD.n267 4.65
R372 VDD.n264 VDD.n263 4.65
R373 VDD.n260 VDD.n259 4.65
R374 VDD.n255 VDD.n254 4.65
R375 VDD.n228 VDD.n227 4.65
R376 VDD.n224 VDD.n223 4.65
R377 VDD.n219 VDD.n218 4.65
R378 VDD.n215 VDD.n214 4.65
R379 VDD.n210 VDD.n209 4.65
R380 VDD.n27 VDD.n23 2.933
R381 VDD.n360 VDD.n357 2.89
R382 VDD.n259 VDD.n256 2.89
R383 VDD.n27 VDD.n26 2.844
R384 VDD.n35  ��B 2.557
R385 VDD.n91 ��B 2.557
R386 VDD.n366 ��B 2.557
R387 VDD.n265  ��B 2.557
R388 VDD.n182 VDD.n179 2.477
R389 VDD.n281 VDD.n280 2.477
R390 VDD.n138 VDD.n135 2.064
R391 VDD.n147 VDD.n146 2.064
R392 VDD.n325 VDD.n322 2.064
R393 VDD.n316 VDD.n313 2.064
R394 VDD.n223 VDD.n220 2.064
R395 VDD.n214 VDD.n213 2.064
R396 VDD.n31 VDD.n27 1.063
R397 VDD.n79 VDD.n52 0.29
R398 VDD.n134 VDD.n108 0.29
R399 VDD.n178 VDD.n152 0.29
R400 VDD.n356 VDD.n330 0.29
R401 VDD.n312 VDD.n286 0.29
R402 VDD.n255 VDD.n228 0.29
R403 VDD.n210 VDD 0.207
R404 VDD.n38 VDD.n34 0.181
R405 VDD.n94 VDD.n90 0.181
R406 VDD.n374 VDD.n369 0.181
R407 VDD.n273 VDD.n268 0.181
R408 VDD.n143 VDD.n139 0.157
R409 VDD.n148 VDD.n143 0.157
R410 VDD.n326 VDD.n321 0.157
R411 VDD.n321 VDD.n317 0.157
R412 VDD.n224 VDD.n219 0.157
R413 VDD.n219 VDD.n215 0.157
R414 VDD.n34 VDD.n31 0.145
R415 VDD.n44 VDD.n38 0.145
R416 VDD.n48 VDD.n44 0.145
R417 VDD.n52 VDD.n48 0.145
R418 VDD.n83 VDD.n79 0.145
R419 VDD.n87 VDD.n83 0.145
R420 VDD.n90 VDD.n87 0.145
R421 VDD.n100 VDD.n94 0.145
R422 VDD.n104 VDD.n100 0.145
R423 VDD.n108 VDD.n104 0.145
R424 VDD.n139 VDD.n134 0.145
R425 VDD.n152 VDD.n148 0.145
R426 VDD.n183 VDD.n178 0.145
R427 VDD.n187 VDD.n183 0.145
R428 VDD.n369 VDD.n365 0.145
R429 VDD.n365 VDD.n361 0.145
R430 VDD.n361 VDD.n356 0.145
R431 VDD.n330 VDD.n326 0.145
R432 VDD.n317 VDD.n312 0.145
R433 VDD.n286 VDD.n282 0.145
R434 VDD.n282 VDD.n277 0.145
R435 VDD.n277 VDD.n273 0.145
R436 VDD.n268 VDD.n264 0.145
R437 VDD.n264 VDD.n260 0.145
R438 VDD.n260 VDD.n255 0.145
R439 VDD.n228 VDD.n224 0.145
R440 VDD.n215 VDD.n210 0.145
R441 VDD VDD.n374 0.133
R442 VDD VDD.n187 0.012
R443 a_3007_411.n2 a_3007_411.t6 470.752
R444 a_3007_411.n2 a_3007_411.t5 384.527
R445 a_3007_411.n3 a_3007_411.t4 314.896
R446 a_3007_411.n4 a_3007_411.n1 260.107
R447 a_3007_411.n9 a_3007_411.n8 208.452
R448 a_3007_411.n3 a_3007_411.n2 182.932
R449 a_3007_411.n9 a_3007_411.n4 170.164
R450 a_3007_411.n11 a_3007_411.n9 135.417
R451 a_3007_411.n12 a_3007_411.n0 55.263
R452 a_3007_411.n8 a_3007_411.n7 30
R453 a_3007_411.n11 a_3007_411.n10 30
R454 a_3007_411.n12 a_3007_411.n11 25.263
R455 a_3007_411.n6 a_3007_411.n5 24.383
R456 a_3007_411.n8 a_3007_411.n6 23.684
R457 a_3007_411.n1 a_3007_411.t1 14.282
R458 a_3007_411.n1 a_3007_411.t2 14.282
R459 a_3007_411.n4 a_3007_411.n3 12.247
R460 GND.n162 GND.n161 237.558
R461 GND.n194 GND.n193 237.558
R462 GND.n123 GND.n122 237.558
R463 GND.n227 GND.n226 237.558
R464 GND.n90 GND.n89 237.558
R465 GND.n43 GND.n42 237.558
R466 GND.n40 GND.n39 210.82
R467 GND.n164 GND.n163 210.82
R468 GND.n196 GND.n195 210.82
R469 GND.n229 GND.n228 210.82
R470 GND.n120 GND.n119 210.82
R471 GND.n87 GND.n86 210.82
R472 GND.n174 GND.n173 166.605
R473 GND.n240 GND.n239 151.605
R474 GND.n55 GND.n54 92.5
R475 GND.n71 GND.n70 92.5
R476 GND.n78 GND.t3 45.413
R477 GND.n19 GND.n18 40.431
R478 GND.n65 GND.n64 40.431
R479 GND.n4 GND.n3 40.003
R480 GND.n78 GND.n77 39.307
R481 GND.n32 GND.n31 37.582
R482 GND.n112 GND.n111 37.582
R483 GND.n207 GND.n206 37.582
R484 GND.n142 GND.n141 37.582
R485 GND.n47 GND.n46 35.865
R486 GND.t6 GND.n109 32.601
R487 GND.t4 GND.n204 32.601
R488 GND.t10 GND.n139 32.601
R489 GND.n48 GND.n47 28.503
R490 GND.n239 GND.n238 28.421
R491 GND.n239 GND.n237 25.263
R492 GND.n237 GND.n236 24.383
R493 GND.n79 GND.n78 23.77
R494 GND.n173 GND.n171 23.03
R495 GND.n109 GND.n108 21.734
R496 GND.n204 GND.n203 21.734
R497 GND.n139 GND.n138 21.734
R498 GND.n25 GND.n24 20.705
R499 GND.n20 GND.n19 20.705
R500 GND.n11 GND.n10 20.705
R501 GND.n5 GND.n4 20.705
R502 GND.n33 GND.n32 20.705
R503 GND.n72 GND.n71 20.705
R504 GND.n66 GND.n65 20.705
R505 GND.n56 GND.n55 20.705
R506 GND.n49 GND.n48 20.705
R507 GND.n80 GND.n79 20.705
R508 GND.n95 GND.n94 20.705
R509 GND.n101 GND.n100 20.705
R510 GND.n113 GND.n112 20.705
R511 GND.n219 GND.n218 20.705
R512 GND.n213 GND.n212 20.705
R513 GND.n208 GND.n207 20.705
R514 GND.n154 GND.n153 20.705
R515 GND.n148 GND.n147 20.705
R516 GND.n143 GND.n142 20.705
R517 GND.n94 GND.n93 19.952
R518 GND.n218 GND.n217 19.952
R519 GND.n153 GND.n152 19.952
R520 GND.n41 GND.n40 18.953
R521 GND.n165 GND.n164 18.953
R522 GND.n197 GND.n196 18.953
R523 GND.n230 GND.n229 18.953
R524 GND.n121 GND.n120 18.953
R525 GND.n88 GND.n87 18.953
R526 GND.n3 GND.n2 17.258
R527 GND.n31 GND.t0 15.644
R528 GND.n111 GND.t6 15.644
R529 GND.n206 GND.t4 15.644
R530 GND.n141 GND.t10 15.644
R531 GND.n44 GND.n41 14.864
R532 GND.n91 GND.n88 14.864
R533 GND.n124 GND.n121 14.864
R534 GND.n231 GND.n230 14.864
R535 GND.n198 GND.n197 14.864
R536 GND.n166 GND.n165 14.864
R537 GND.n18 GND.t9 13.654
R538 GND.n64 GND.t5 13.654
R539 GND.n64 GND.n63 13.654
R540 GND.n31 GND.n30 13.541
R541 GND.n111 GND.n110 13.541
R542 GND.n206 GND.n205 13.541
R543 GND.n141 GND.n140 13.541
R544 GND.n22 GND.n20 9.29
R545 GND.n68 GND.n66 9.29
R546 GND.n144 GND.n135 9.154
R547 GND.n150 GND.n149 9.154
R548 GND.n156 GND.n155 9.154
R549 GND.n159 GND.n158 9.154
R550 GND.n166 GND.n162 9.154
R551 GND.n169 GND.n168 9.154
R552 GND.n176 GND.n175 9.154
R553 GND.n179 GND.n178 9.154
R554 GND.n182 GND.n181 9.154
R555 GND.n185 GND.n184 9.154
R556 GND.n188 GND.n187 9.154
R557 GND.n191 GND.n190 9.154
R558 GND.n198 GND.n194 9.154
R559 GND.n209 GND.n200 9.154
R560 GND.n215 GND.n214 9.154
R561 GND.n221 GND.n220 9.154
R562 GND.n224 GND.n223 9.154
R563 GND.n231 GND.n227 9.154
R564 GND.n234 GND.n233 9.154
R565 GND.n242 GND.n241 9.154
R566 GND.n245 GND.n244 9.154
R567 GND.n248 GND.n247 9.154
R568 GND.n130 GND.n129 9.154
R569 GND.n127 GND.n126 9.154
R570 GND.n124 GND.n123 9.154
R571 GND.n117 GND.n116 9.154
R572 GND.n114 GND.n105 9.154
R573 GND.n103 GND.n102 9.154
R574 GND.n97 GND.n96 9.154
R575 GND.n91 GND.n90 9.154
R576 GND.n84 GND.n83 9.154
R577 GND.n81 GND.n76 9.154
R578 GND.n74 GND.n73 9.154
R579 GND.n68 GND.n67 9.154
R580 GND.n60 GND.n59 9.154
R581 GND.n57 GND.n53 9.154
R582 GND.n51 GND.n50 9.154
R583 GND.n44 GND.n43 9.154
R584 GND.n37 GND.n36 9.154
R585 GND.n34 GND.n29 9.154
R586 GND.n27 GND.n26 9.154
R587 GND.n22 GND.n21 9.154
R588 GND.n15 GND.n14 9.154
R589 GND.n12 GND.n9 9.154
R590 GND.n7 GND.n6 9.154
R591 GND.n173 GND.n172 8.128
R592 GND.t9 GND.n17 7.04
R593 GND.t5 GND.n62 7.04
R594 GND.n8 GND.n1 4.795
R595 GND.n134 GND.n133 4.65
R596 GND.n8 GND.n7 4.65
R597 GND.n13 GND.n12 4.65
R598 GND.n16 GND.n15 4.65
R599 GND.n23 GND.n22 4.65
R600 GND.n28 GND.n27 4.65
R601 GND.n35 GND.n34 4.65
R602 GND.n38 GND.n37 4.65
R603 GND.n45 GND.n44 4.65
R604 GND.n52 GND.n51 4.65
R605 GND.n58 GND.n57 4.65
R606 GND.n61 GND.n60 4.65
R607 GND.n69 GND.n68 4.65
R608 GND.n75 GND.n74 4.65
R609 GND.n82 GND.n81 4.65
R610 GND.n85 GND.n84 4.65
R611 GND.n92 GND.n91 4.65
R612 GND.n98 GND.n97 4.65
R613 GND.n104 GND.n103 4.65
R614 GND.n115 GND.n114 4.65
R615 GND.n118 GND.n117 4.65
R616 GND.n125 GND.n124 4.65
R617 GND.n128 GND.n127 4.65
R618 GND.n131 GND.n130 4.65
R619 GND.n249 GND.n248 4.65
R620 GND.n246 GND.n245 4.65
R621 GND.n243 GND.n242 4.65
R622 GND.n235 GND.n234 4.65
R623 GND.n232 GND.n231 4.65
R624 GND.n225 GND.n224 4.65
R625 GND.n222 GND.n221 4.65
R626 GND.n216 GND.n215 4.65
R627 GND.n210 GND.n209 4.65
R628 GND.n199 GND.n198 4.65
R629 GND.n192 GND.n191 4.65
R630 GND.n189 GND.n188 4.65
R631 GND.n186 GND.n185 4.65
R632 GND.n183 GND.n182 4.65
R633 GND.n180 GND.n179 4.65
R634 GND.n177 GND.n176 4.65
R635 GND.n170 GND.n169 4.65
R636 GND.n167 GND.n166 4.65
R637 GND.n160 GND.n159 4.65
R638 GND.n157 GND.n156 4.65
R639 GND.n151 GND.n150 4.65
R640 GND.n145 GND.n144 4.65
R641 GND.n107 GND.n106 4.504
R642 GND.n202 GND.n201 4.504
R643 GND.n137 GND.n136 4.504
R644 GND.n12 GND.n11 4.129
R645 GND.n27 GND.n25 4.129
R646 GND.n57 GND.n56 4.129
R647 GND.n74 GND.n72 4.129
R648 GND.n97 GND.n95 4.129
R649 GND.n242 GND.n240 4.129
R650 GND.n221 GND.n219 4.129
R651 GND.n176 GND.n174 4.129
R652 GND.n156 GND.n154 4.129
R653 GND.n114 GND.n113 3.716
R654 GND.n209 GND.n208 3.716
R655 GND.n144 GND.n143 3.716
R656 GND.t6 GND.n107 2.452
R657 GND.t4 GND.n202 2.452
R658 GND.t10 GND.n137 2.452
R659 GND.n7 GND.n5 1.032
R660 GND.n34 GND.n33 1.032
R661 GND.n51 GND.n49 1.032
R662 GND.n81 GND.n80 1.032
R663 GND.n1 GND.n0 0.474
R664 GND.n133 GND.n132 0.474
R665 GND.n100 GND.n99 0.376
R666 GND.n212 GND.n211 0.376
R667 GND.n147 GND.n146 0.376
R668 GND.n45 GND.n38 0.29
R669 GND.n92 GND.n85 0.29
R670 GND.n125 GND.n118 0.29
R671 GND.n232 GND.n225 0.29
R672 GND.n199 GND.n192 0.29
R673 GND.n167 GND.n160 0.29
R674 GND.n134 GND 0.207
R675 GND.n103 GND.n101 0.206
R676 GND.n215 GND.n213 0.206
R677 GND.n150 GND.n148 0.206
R678 GND.n23 GND.n16 0.181
R679 GND.n69 GND.n61 0.181
R680 GND.n249 GND.n246 0.181
R681 GND.n183 GND.n180 0.181
R682 GND.n104 GND.n98 0.157
R683 GND.n115 GND.n104 0.157
R684 GND.n222 GND.n216 0.157
R685 GND.n216 GND.n210 0.157
R686 GND.n157 GND.n151 0.157
R687 GND.n151 GND.n145 0.157
R688 GND.n13 GND.n8 0.145
R689 GND.n16 GND.n13 0.145
R690 GND.n28 GND.n23 0.145
R691 GND.n35 GND.n28 0.145
R692 GND.n38 GND.n35 0.145
R693 GND.n52 GND.n45 0.145
R694 GND.n58 GND.n52 0.145
R695 GND.n61 GND.n58 0.145
R696 GND.n75 GND.n69 0.145
R697 GND.n82 GND.n75 0.145
R698 GND.n85 GND.n82 0.145
R699 GND.n98 GND.n92 0.145
R700 GND.n118 GND.n115 0.145
R701 GND.n128 GND.n125 0.145
R702 GND.n131 GND.n128 0.145
R703 GND.n246 GND.n243 0.145
R704 GND.n243 GND.n235 0.145
R705 GND.n235 GND.n232 0.145
R706 GND.n225 GND.n222 0.145
R707 GND.n210 GND.n199 0.145
R708 GND.n192 GND.n189 0.145
R709 GND.n189 GND.n186 0.145
R710 GND.n186 GND.n183 0.145
R711 GND.n180 GND.n177 0.145
R712 GND.n177 GND.n170 0.145
R713 GND.n170 GND.n167 0.145
R714 GND.n160 GND.n157 0.145
R715 GND.n145 GND.n134 0.145
R716 GND GND.n249 0.133
R717 GND GND.n131 0.012
R718 Q.n0 Q.t6 486.819
R719 Q.n0 Q.t4 384.527
R720 Q.n1 Q.t5 322.919
R721 Q.n8 Q.n2 287.966
R722 Q.n7 Q.n6 223.975
R723 Q.n1 Q.n0 206.987
R724 Q.n7 Q.n3 157.274
R725 Q.n8 Q.n7 142.305
R726 Q.n6 Q.n5 22.578
R727 Q.n2 Q.t1 14.282
R728 Q.n2 Q.t2 14.282
R729 Q.n6 Q.n4 8.58
R730 Q.n9 Q.n1 5.965
R731 Q.n9 Q.n8 4.65
R732 Q.n9 Q 0.046
R733 D.n2 D.t5 512.525
R734 D.n0 D.t0 472.359
R735 D.n0 D.t3 384.527
R736 D.n2 D.t1 371.139
R737 D.n1 D.t2 342.755
R738 D.n3 D.t4 338.57
R739 D.n3 D.n2 191.629
R740 D.n1 D.n0 154.955
R741 D.n4 D.n1 11.134
R742 D.n4 D.n3 4.65
R743 D.n4 D 0.046
R744 a_185_209.n0 a_185_209.t5 480.392
R745 a_185_209.n0 a_185_209.t4 403.272
R746 a_185_209.n1 a_185_209.t3 357.204
R747 a_185_209.n3 a_185_209.n2 322.049
R748 a_185_209.n4 a_185_209.n3 243.422
R749 a_185_209.n1 a_185_209.n0 171.288
R750 a_185_209.n4 a_185_209.t1 14.282
R751 a_185_209.t2 a_185_209.n4 14.282
R752 a_185_209.n3 a_185_209.n1 10.615
R753 a_661_1050.n1 a_661_1050.t6 512.525
R754 a_661_1050.n1 a_661_1050.t5 371.139
R755 a_661_1050.n4 a_661_1050.n3 299.461
R756 a_661_1050.n2 a_661_1050.t7 282.852
R757 a_661_1050.n2 a_661_1050.n1 247.347
R758 a_661_1050.n5 a_661_1050.n4 187.858
R759 a_661_1050.n6 a_661_1050.n5 157.963
R760 a_661_1050.n5 a_661_1050.n0 91.706
R761 a_661_1050.n0 a_661_1050.t4 14.282
R762 a_661_1050.n0 a_661_1050.t0 14.282
R763 a_661_1050.n6 a_661_1050.t2 14.282
R764 a_661_1050.t3 a_661_1050.n6 14.282
R765 a_661_1050.n4 a_661_1050.n2 10.343
R766 a_1295_209.n0 a_1295_209.t3 486.819
R767 a_1295_209.n0 a_1295_209.t5 384.527
R768 a_1295_209.n1 a_1295_209.t4 350.778
R769 a_1295_209.n3 a_1295_209.n2 322.049
R770 a_1295_209.n4 a_1295_209.n3 243.422
R771 a_1295_209.n1 a_1295_209.n0 179.128
R772 a_1295_209.n3 a_1295_209.n1 14.696
R773 a_1295_209.n4 a_1295_209.t1 14.282
R774 a_1295_209.t2 a_1295_209.n4 14.282
R775 a_1666_101.n3 a_1666_101.n1 42.788
R776 a_1666_101.t0 a_1666_101.n0 8.137
R777 a_1666_101.n3 a_1666_101.n2 4.665
R778 a_1666_101.t0 a_1666_101.n3 0.06
R779 GATE.n0 GATE.t3 480.392
R780 GATE.n2 GATE.t5 472.359
R781 GATE.n0 GATE.t1 403.272
R782 GATE.n2 GATE.t0 384.527
R783 GATE.n1 GATE.t4 301.486
R784 GATE.n3 GATE.t2 259.178
R785 GATE.n3 GATE.n2 238.531
R786 GATE.n1 GATE.n0 227.006
R787 GATE.n4 GATE.n1 8.141
R788 GATE.n4 GATE.n3 4.65
R789 GATE.n4 GATE 0.046
R790 a_556_101.n11 a_556_101.n10 68.43
R791 a_556_101.n3 a_556_101.n2 62.817
R792 a_556_101.n7 a_556_101.n6 38.626
R793 a_556_101.n6 a_556_101.n5 35.955
R794 a_556_101.n3 a_556_101.n1 26.202
R795 a_556_101.t0 a_556_101.n3 19.737
R796 a_556_101.t1 a_556_101.n8 8.137
R797 a_556_101.t0 a_556_101.n4 7.273
R798 a_556_101.t0 a_556_101.n0 6.109
R799 a_556_101.t1 a_556_101.n7 4.864
R800 a_556_101.t0 a_556_101.n12 2.074
R801 a_556_101.n12 a_556_101.t1 0.937
R802 a_556_101.t1 a_556_101.n11 0.763
R803 a_556_101.n11 a_556_101.n9 0.185
R804 a_2795_1051.n0 a_2795_1051.t2 228.369
R805 a_2795_1051.n0 a_2795_1051.t0 219.778
R806 a_2795_1051.n1 a_2795_1051.n0 42.29
R807 a_2795_1051.n1 a_2795_1051.t3 14.282
R808 a_2795_1051.t1 a_2795_1051.n1 14.282
R809 a_3461_1051.n1 a_3461_1051.t3 228.368
R810 a_3461_1051.t1 a_3461_1051.n1 219.777
R811 a_3461_1051.n1 a_3461_1051.n0 42.29
R812 a_3461_1051.n0 a_3461_1051.t2 14.282
R813 a_3461_1051.n0 a_3461_1051.t0 14.282
C4 VDD GND 6.85fF
C5 a_3461_1051.n0 GND 0.21fF
C6 a_3461_1051.n1 GND 0.50fF
C7 a_2795_1051.n0 GND 0.52fF
C8 a_2795_1051.n1 GND 0.22fF
C9 a_556_101.n0 GND 0.02fF
C10 a_556_101.n1 GND 0.09fF
C11 a_556_101.n2 GND 0.08fF
C12 a_556_101.n3 GND 0.03fF
C13 a_556_101.n4 GND 0.01fF
C14 a_556_101.n5 GND 0.04fF
C15 a_556_101.n6 GND 0.04fF
C16 a_556_101.n7 GND 0.02fF
C17 a_556_101.n8 GND 0.05fF
C18 a_556_101.n9 GND 0.15fF
C19 a_556_101.n10 GND 0.08fF
C20 a_556_101.n11 GND 0.08fF
C21 a_556_101.t1 GND 0.23fF
C22 a_556_101.n12 GND 0.01fF
C23 a_1666_101.n0 GND 0.05fF
C24 a_1666_101.n1 GND 0.12fF
C25 a_1666_101.n2 GND 0.04fF
C26 a_1666_101.n3 GND 0.17fF
C27 a_1295_209.n0 GND 0.39fF
C28 a_1295_209.n1 GND 1.25fF
C29 a_1295_209.n2 GND 0.39fF
C30 a_1295_209.n3 GND 1.51fF
C31 a_1295_209.n4 GND 0.72fF
C32 a_661_1050.n0 GND 0.34fF
C33 a_661_1050.n1 GND 0.31fF
C34 a_661_1050.t7 GND 0.45fF
C35 a_661_1050.n2 GND 0.52fF
C36 a_661_1050.n3 GND 0.27fF
C37 a_661_1050.n4 GND 0.58fF
C38 a_661_1050.n5 GND 0.54fF
C39 a_661_1050.n6 GND 0.44fF
C40 a_185_209.n0 GND 0.30fF
C41 a_185_209.n1 GND 0.56fF
C42 a_185_209.n2 GND 0.30fF
C43 a_185_209.n3 GND 0.75fF
C44 a_185_209.n4 GND 0.55fF
C45 Q.n0 GND 0.34fF
C46 Q.t5 GND 0.50fF
C47 Q.n1 GND 0.45fF
C48 Q.n2 GND 0.57fF
C49 Q.n3 GND 0.17fF
C50 Q.n4 GND 0.04fF
C51 Q.n5 GND 0.05fF
C52 Q.n6 GND 0.14fF
C53 Q.n7 GND 0.47fF
C54 Q.n8 GND 0.48fF
C55 Q.n9 GND 0.30fF
C56 a_3007_411.n0 GND 0.05fF
C57 a_3007_411.n1 GND 0.60fF
C58 a_3007_411.n2 GND 0.34fF
C59 a_3007_411.n3 GND 0.83fF
C60 a_3007_411.n4 GND 0.93fF
C61 a_3007_411.n5 GND 0.04fF
C62 a_3007_411.n6 GND 0.06fF
C63 a_3007_411.n7 GND 0.04fF
C64 a_3007_411.n8 GND 0.13fF
C65 a_3007_411.n9 GND 0.54fF
C66 a_3007_411.n10 GND 0.04fF
C67 a_3007_411.n11 GND 0.06fF
C68 a_3007_411.n12 GND 0.05fF
C69 VDD.n1 GND 0.03fF
C70 VDD.n2 GND 0.11fF
C71 VDD.n3 GND 0.02fF
C72 VDD.n4 GND 0.02fF
C73 VDD.n5 GND 0.05fF
C74 VDD.n6 GND 0.02fF
C75 VDD.n7 GND 0.02fF
C76 VDD.n8 GND 0.02fF
C77 VDD.n9 GND 0.02fF
C78 VDD.n10 GND 0.02fF
C79 VDD.n11 GND 0.02fF
C80 VDD.n12 GND 0.02fF
C81 VDD.n13 GND 0.02fF
C82 VDD.n14 GND 0.03fF
C83 VDD.n15 GND 0.01fF
C84 VDD.n20 GND 0.38fF
C85 VDD.n21 GND 0.23fF
C86 VDD.n22 GND 0.02fF
C87 VDD.n23 GND 0.03fF
C88 VDD.n24 GND 0.20fF
C89 VDD.n25 GND 0.01fF
C90 VDD.n26 GND 0.02fF
C91 VDD.n27 GND 0.01fF
C92 VDD.n28 GND 0.14fF
C93 VDD.n29 GND 0.01fF
C94 VDD.n30 GND 0.02fF
C95 VDD.n31 GND 0.07fF
C96 VDD.n32 GND 0.01fF
C97 VDD.n33 GND 0.02fF
C98 VDD.n34 GND 0.02fF
C99 VDD.n35 GND 0.12fF
C100 VDD.n36 GND 0.01fF
C101 VDD.n37 GND 0.02fF
C102 VDD.n38 GND 0.02fF
C103 VDD.n39 GND 0.07fF
C104 VDD.n40 GND 0.04fF
C105 VDD.n41 GND 0.14fF
C106 VDD.n42 GND 0.01fF
C107 VDD.n43 GND 0.01fF
C108 VDD.n44 GND 0.02fF
C109 VDD.n45 GND 0.21fF
C110 VDD.n46 GND 0.01fF
C111 VDD.n47 GND 0.02fF
C112 VDD.n48 GND 0.02fF
C113 VDD.n49 GND 0.23fF
C114 VDD.n50 GND 0.01fF
C115 VDD.n51 GND 0.02fF
C116 VDD.n52 GND 0.03fF
C117 VDD.n53 GND 0.05fF
C118 VDD.n54 GND 0.02fF
C119 VDD.n55 GND 0.02fF
C120 VDD.n56 GND 0.02fF
C121 VDD.n57 GND 0.02fF
C122 VDD.n58 GND 0.02fF
C123 VDD.n59 GND 0.02fF
C124 VDD.n60 GND 0.02fF
C125 VDD.n61 GND 0.02fF
C126 VDD.n62 GND 0.02fF
C127 VDD.n63 GND 0.02fF
C128 VDD.n64 GND 0.01fF
C129 VDD.n65 GND 0.02fF
C130 VDD.n66 GND 0.02fF
C131 VDD.n67 GND 0.18fF
C132 VDD.n68 GND 0.02fF
C133 VDD.n69 GND 0.02fF
C134 VDD.n71 GND 0.02fF
C135 VDD.n75 GND 0.23fF
C136 VDD.n76 GND 0.23fF
C137 VDD.n77 GND 0.01fF
C138 VDD.n78 GND 0.02fF
C139 VDD.n79 GND 0.03fF
C140 VDD.n80 GND 0.20fF
C141 VDD.n81 GND 0.01fF
C142 VDD.n82 GND 0.02fF
C143 VDD.n83 GND 0.02fF
C144 VDD.n84 GND 0.14fF
C145 VDD.n85 GND 0.01fF
C146 VDD.n86 GND 0.02fF
C147 VDD.n87 GND 0.02fF
C148 VDD.n88 GND 0.01fF
C149 VDD.n89 GND 0.02fF
C150 VDD.n90 GND 0.02fF
C151 VDD.n91 GND 0.12fF
C152 VDD.n92 GND 0.01fF
C153 VDD.n93 GND 0.02fF
C154 VDD.n94 GND 0.02fF
C155 VDD.n95 GND 0.07fF
C156 VDD.n96 GND 0.04fF
C157 VDD.n97 GND 0.14fF
C158 VDD.n98 GND 0.01fF
C159 VDD.n99 GND 0.01fF
C160 VDD.n100 GND 0.02fF
C161 VDD.n101 GND 0.21fF
C162 VDD.n102 GND 0.01fF
C163 VDD.n103 GND 0.02fF
C164 VDD.n104 GND 0.02fF
C165 VDD.n105 GND 0.23fF
C166 VDD.n106 GND 0.01fF
C167 VDD.n107 GND 0.02fF
C168 VDD.n108 GND 0.03fF
C169 VDD.n109 GND 0.15fF
C170 VDD.n110 GND 0.02fF
C171 VDD.n111 GND 0.02fF
C172 VDD.n112 GND 0.02fF
C173 VDD.n113 GND 0.05fF
C174 VDD.n114 GND 0.02fF
C175 VDD.n115 GND 0.02fF
C176 VDD.n116 GND 0.02fF
C177 VDD.n117 GND 0.02fF
C178 VDD.n118 GND 0.02fF
C179 VDD.n119 GND 0.02fF
C180 VDD.n120 GND 0.02fF
C181 VDD.n121 GND 0.02fF
C182 VDD.n122 GND 0.02fF
C183 VDD.n123 GND 0.01fF
C184 VDD.n124 GND 0.02fF
C185 VDD.n125 GND 0.02fF
C186 VDD.n126 GND 0.02fF
C187 VDD.n130 GND 0.23fF
C188 VDD.n131 GND 0.23fF
C189 VDD.n132 GND 0.01fF
C190 VDD.n133 GND 0.02fF
C191 VDD.n134 GND 0.03fF
C192 VDD.n135 GND 0.05fF
C193 VDD.n136 GND 0.17fF
C194 VDD.n137 GND 0.01fF
C195 VDD.n138 GND 0.01fF
C196 VDD.n139 GND 0.02fF
C197 VDD.n140 GND 0.14fF
C198 VDD.n141 GND 0.01fF
C199 VDD.n142 GND 0.02fF
C200 VDD.n143 GND 0.02fF
C201 VDD.n144 GND 0.17fF
C202 VDD.n145 GND 0.01fF
C203 VDD.n146 GND 0.05fF
C204 VDD.n147 GND 0.01fF
C205 VDD.n148 GND 0.02fF
C206 VDD.n149 GND 0.23fF
C207 VDD.n150 GND 0.01fF
C208 VDD.n151 GND 0.02fF
C209 VDD.n152 GND 0.03fF
C210 VDD.n153 GND 0.15fF
C211 VDD.n154 GND 0.02fF
C212 VDD.n155 GND 0.02fF
C213 VDD.n156 GND 0.02fF
C214 VDD.n157 GND 0.05fF
C215 VDD.n158 GND 0.02fF
C216 VDD.n159 GND 0.02fF
C217 VDD.n160 GND 0.02fF
C218 VDD.n161 GND 0.02fF
C219 VDD.n162 GND 0.02fF
C220 VDD.n163 GND 0.02fF
C221 VDD.n164 GND 0.02fF
C222 VDD.n165 GND 0.02fF
C223 VDD.n166 GND 0.02fF
C224 VDD.n167 GND 0.01fF
C225 VDD.n168 GND 0.02fF
C226 VDD.n169 GND 0.02fF
C227 VDD.n170 GND 0.02fF
C228 VDD.n174 GND 0.23fF
C229 VDD.n175 GND 0.23fF
C230 VDD.n176 GND 0.01fF
C231 VDD.n177 GND 0.02fF
C232 VDD.n178 GND 0.03fF
C233 VDD.n179 GND 0.05fF
C234 VDD.n180 GND 0.20fF
C235 VDD.n181 GND 0.01fF
C236 VDD.n182 GND 0.01fF
C237 VDD.n183 GND 0.02fF
C238 VDD.n184 GND 0.14fF
C239 VDD.n185 GND 0.01fF
C240 VDD.n186 GND 0.02fF
C241 VDD.n187 GND 0.01fF
C242 VDD.n188 GND 0.08fF
C243 VDD.n189 GND 0.02fF
C244 VDD.n190 GND 0.02fF
C245 VDD.n191 GND 0.05fF
C246 VDD.n192 GND 0.02fF
C247 VDD.n193 GND 0.02fF
C248 VDD.n194 GND 0.02fF
C249 VDD.n195 GND 0.02fF
C250 VDD.n196 GND 0.02fF
C251 VDD.n197 GND 0.02fF
C252 VDD.n198 GND 0.02fF
C253 VDD.n199 GND 0.02fF
C254 VDD.n200 GND 0.03fF
C255 VDD.n201 GND 0.03fF
C256 VDD.n202 GND 0.02fF
C257 VDD.n206 GND 0.38fF
C258 VDD.n207 GND 0.23fF
C259 VDD.n208 GND 0.02fF
C260 VDD.n209 GND 0.03fF
C261 VDD.n210 GND 0.02fF
C262 VDD.n211 GND 0.17fF
C263 VDD.n212 GND 0.01fF
C264 VDD.n213 GND 0.05fF
C265 VDD.n214 GND 0.01fF
C266 VDD.n215 GND 0.02fF
C267 VDD.n216 GND 0.14fF
C268 VDD.n217 GND 0.01fF
C269 VDD.n218 GND 0.02fF
C270 VDD.n219 GND 0.02fF
C271 VDD.n220 GND 0.05fF
C272 VDD.n221 GND 0.17fF
C273 VDD.n222 GND 0.01fF
C274 VDD.n223 GND 0.01fF
C275 VDD.n224 GND 0.02fF
C276 VDD.n225 GND 0.23fF
C277 VDD.n226 GND 0.01fF
C278 VDD.n227 GND 0.02fF
C279 VDD.n228 GND 0.03fF
C280 VDD.n229 GND 0.02fF
C281 VDD.n232 GND 0.02fF
C282 VDD.n234 GND 0.02fF
C283 VDD.n235 GND 0.15fF
C284 VDD.n236 GND 0.02fF
C285 VDD.n238 GND 0.23fF
C286 VDD.n239 GND 0.23fF
C287 VDD.n240 GND 0.01fF
C288 VDD.n241 GND 0.05fF
C289 VDD.n242 GND 0.02fF
C290 VDD.n243 GND 0.02fF
C291 VDD.n244 GND 0.02fF
C292 VDD.n245 GND 0.02fF
C293 VDD.n246 GND 0.02fF
C294 VDD.n247 GND 0.02fF
C295 VDD.n248 GND 0.02fF
C296 VDD.n249 GND 0.02fF
C297 VDD.n250 GND 0.02fF
C298 VDD.n251 GND 0.02fF
C299 VDD.n252 GND 0.01fF
C300 VDD.n253 GND 0.02fF
C301 VDD.n254 GND 0.02fF
C302 VDD.n255 GND 0.03fF
C303 VDD.n256 GND 0.05fF
C304 VDD.n257 GND 0.21fF
C305 VDD.n258 GND 0.01fF
C306 VDD.n259 GND 0.01fF
C307 VDD.n260 GND 0.02fF
C308 VDD.n261 GND 0.14fF
C309 VDD.n262 GND 0.01fF
C310 VDD.n263 GND 0.02fF
C311 VDD.n264 GND 0.02fF
C312 VDD.n265 GND 0.12fF
C313 VDD.n266 GND 0.01fF
C314 VDD.n267 GND 0.02fF
C315 VDD.n268 GND 0.02fF
C316 VDD.n269 GND 0.01fF
C317 VDD.n270 GND 0.07fF
C318 VDD.n271 GND 0.04fF
C319 VDD.n272 GND 0.02fF
C320 VDD.n273 GND 0.02fF
C321 VDD.n274 GND 0.14fF
C322 VDD.n275 GND 0.01fF
C323 VDD.n276 GND 0.02fF
C324 VDD.n277 GND 0.02fF
C325 VDD.n278 GND 0.20fF
C326 VDD.n279 GND 0.01fF
C327 VDD.n280 GND 0.05fF
C328 VDD.n281 GND 0.01fF
C329 VDD.n282 GND 0.02fF
C330 VDD.n283 GND 0.23fF
C331 VDD.n284 GND 0.01fF
C332 VDD.n285 GND 0.02fF
C333 VDD.n286 GND 0.03fF
C334 VDD.n287 GND 0.02fF
C335 VDD.n288 GND 0.02fF
C336 VDD.n292 GND 0.23fF
C337 VDD.n293 GND 0.23fF
C338 VDD.n294 GND 0.01fF
C339 VDD.n295 GND 0.15fF
C340 VDD.n296 GND 0.02fF
C341 VDD.n297 GND 0.02fF
C342 VDD.n298 GND 0.02fF
C343 VDD.n299 GND 0.05fF
C344 VDD.n300 GND 0.02fF
C345 VDD.n301 GND 0.02fF
C346 VDD.n302 GND 0.02fF
C347 VDD.n303 GND 0.02fF
C348 VDD.n304 GND 0.02fF
C349 VDD.n305 GND 0.02fF
C350 VDD.n306 GND 0.02fF
C351 VDD.n307 GND 0.02fF
C352 VDD.n308 GND 0.02fF
C353 VDD.n309 GND 0.01fF
C354 VDD.n310 GND 0.02fF
C355 VDD.n311 GND 0.02fF
C356 VDD.n312 GND 0.03fF
C357 VDD.n313 GND 0.05fF
C358 VDD.n314 GND 0.17fF
C359 VDD.n315 GND 0.01fF
C360 VDD.n316 GND 0.01fF
C361 VDD.n317 GND 0.02fF
C362 VDD.n318 GND 0.14fF
C363 VDD.n319 GND 0.01fF
C364 VDD.n320 GND 0.02fF
C365 VDD.n321 GND 0.02fF
C366 VDD.n322 GND 0.05fF
C367 VDD.n323 GND 0.17fF
C368 VDD.n324 GND 0.01fF
C369 VDD.n325 GND 0.01fF
C370 VDD.n326 GND 0.02fF
C371 VDD.n327 GND 0.23fF
C372 VDD.n328 GND 0.01fF
C373 VDD.n329 GND 0.02fF
C374 VDD.n330 GND 0.03fF
C375 VDD.n331 GND 0.15fF
C376 VDD.n332 GND 0.02fF
C377 VDD.n333 GND 0.02fF
C378 VDD.n334 GND 0.02fF
C379 VDD.n335 GND 0.05fF
C380 VDD.n336 GND 0.02fF
C381 VDD.n337 GND 0.02fF
C382 VDD.n338 GND 0.02fF
C383 VDD.n339 GND 0.02fF
C384 VDD.n340 GND 0.02fF
C385 VDD.n341 GND 0.02fF
C386 VDD.n342 GND 0.02fF
C387 VDD.n343 GND 0.02fF
C388 VDD.n344 GND 0.02fF
C389 VDD.n345 GND 0.01fF
C390 VDD.n346 GND 0.02fF
C391 VDD.n347 GND 0.02fF
C392 VDD.n348 GND 0.02fF
C393 VDD.n352 GND 0.23fF
C394 VDD.n353 GND 0.23fF
C395 VDD.n354 GND 0.01fF
C396 VDD.n355 GND 0.02fF
C397 VDD.n356 GND 0.03fF
C398 VDD.n357 GND 0.05fF
C399 VDD.n358 GND 0.21fF
C400 VDD.n359