* SPICE3 file created from AOI3X1.ext - technology: sky130A

.subckt AOI3X1 YN A B C VDD GND
X0 VDD.t9 A.t0 a_217_1050.t2 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X1 VDD.t5 a_217_1050.t5 a_797_1051.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X2 VDD.t12 B.t0 a_217_1050.t4  ,�X sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X3 YN a_217_1050.t6 GND.t1 GND sky130_fd_pr__nfet_01v8 ad=3.582p pd=3.15u as=0p ps=0u w=0u l=0u
X4 GND A.t1 a_112_101.t0 GND sky130_fd_pr__nfet_01v8 ad=2.1157p pd=1.451u as=0p ps=0u w=0u l=0u
X5 a_797_1051.t3 C.t0 YN.t2 �+�X sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X6 a_217_1050.t3 A.t2 VDD.t7  ,�X sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X7 a_797_1051.t0 a_217_1050.t7 VDD.t3 �+�X sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X8 a_217_1050.t1 B.t1 VDD.t1  ,�X sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X9 YN C.t2 GND.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X10 YN.t1 C.t1 a_797_1051.t2 �+�X sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X11 YN C GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
C0 YN VDD 0.52fF
C1 B VDD 0.32fF
C2 B A 0.27fF
C3 C YN 0.26fF
C4 VDD A 0.32fF
C5 C VDD 0.32fF
R0 A.n0 A.t0 480.392
R1 A.n0 A.t2 403.272
R2 A.n1 A.t1 301.486
R3 A.n1 A.n0 227.006
R4 A.n2 A.n1 4.65
R5 A.n2 A 0.046
R6 a_217_1050.n3 a_217_1050.t7 486.819
R7 a_217_1050.n3 a_217_1050.t5 384.527
R8 a_217_1050.n4 a_217_1050.t6 267.201
R9 a_217_1050.n4 a_217_1050.n3 262.705
R10 a_217_1050.n5 a_217_1050.n2 243.576
R11 a_217_1050.n7 a_217_1050.n5 228.526
R12 a_217_1050.n2 a_217_1050.n1 157.964
R13 a_217_1050.n2 a_217_1050.n0 91.706
R14 a_217_1050.n7 a_217_1050.n6 15.218
R15 a_217_1050.n0 a_217_1050.t4 14.282
R16 a_217_1050.n0 a_217_1050.t1 14.282
R17 a_217_1050.n1 a_217_1050.t2 14.282
R18 a_217_1050.n1 a_217_1050.t3 14.282
R19 a_217_1050.n8 a_217_1050.n7 12.014
R20 a_217_1050.n5 a_217_1050.n4 10.615
R21 VDD.n60 VDD.n49 144.705
R22 VDD.n108 VDD.t12 143.754
R23 VDD.n86 VDD.t7 135.17
R24 VDD.n40 VDD.n39 129.849
R25 VDD.n100 VDD.n99 129.472
R26 VDD.n122 VDD.n121 92.5
R27 VDD.n120 VDD.n119 92.5
R28 VDD.n118 VDD.n117 92.5
R29 VDD.n116 VDD.n115 92.5
R30 VDD.n124 VDD.n123 92.5
R31 VDD.n74 VDD.n73 92.5
R32 VDD.n72 VDD.n71 92.5
R33 VDD.n70 VDD.n69 92.5
R34 VDD.n68 VDD.n67 92.5
R35 VDD.n76 VDD.n75 92.5
R36 VDD.n14 VDD.n1 92.5
R37 VDD.n5 VDD.n4 92.5
R38 VDD.n7 VDD.n6 92.5
R39 VDD.n9 VDD.n8 92.5
R40 VDD.n11 VDD.n10 92.5
R41 VDD.n13 VDD.n12 92.5
R42 VDD.n21 VDD.n20 92.059
R43 VDD.n59 VDD.n58 92.059
R44 VDD.n82 VDD.n81 92.059
R45 VDD.n20 VDD.n16 67.194
R46 VDD.n20 VDD.n17 67.194
R47 VDD.n20 VDD.n18 67.194
R48 VDD.n20 VDD.n19 67.194
R49 VDD.n66 VDD.n65 44.141
R50 VDD.n5 VDD.n3 44.141
R51 VDD.n65 VDD.n63 44.107
R52 VDD.n3 VDD.n2 44.107
R53 VDD.n20 VDD.n15 41.052
R54 VDD.n78 VDD.n77 39.742
R55 VDD.n57 VDD.n54 39.742
R56 VDD.n57 VDD.n56 39.742
R57 VDD.n53 VDD.n52 39.742
R58 VDD.n65 VDD.n64 38
R59 VDD.n56 VDD.n55 36.774
R60 VDD.n1 VDD.n0 30.923
R61 VDD.n81 VDD.n79 26.38
R62 VDD.n81 VDD.n78 26.38
R63 VDD.n81 VDD.n80 26.38
R64 VDD.n58 VDD.n57 26.38
R65 VDD.n58 VDD.n53 26.38
R66 VDD.n58 VDD.n51 26.38
R67 VDD.n58 VDD.n50 26.38
R68 VDD.n84 VDD.n76 22.915
R69 VDD.n23 VDD.n14 22.915
R70 VDD.n28 �+�X 20.457
R71 VDD.n104  ,�X 20.457
R72 VDD.n41  17.9
R73 VDD.n91  ,�X 17.9
R74 VDD.n76 VDD.n74 14.864
R75 VDD.n74 VDD.n72 14.864
R76 VDD.n72 VDD.n70 14.864
R77 VDD.n70 VDD.n68 14.864
R78 VDD.n68 VDD.n66 14.864
R79 VDD.n124 VDD.n122 14.864
R80 VDD.n122 VDD.n120 14.864
R81 VDD.n120 VDD.n118 14.864
R82 VDD.n118 VDD.n116 14.864
R83 VDD.n116 VDD.n114 14.864
R84 VDD.n114 VDD.n113 14.864
R85 VDD.n14 VDD.n13 14.864
R86 VDD.n13 VDD.n11 14.864
R87 VDD.n11 VDD.n9 14.864
R88 VDD.n9 VDD.n7 14.864
R89 VDD.n7 VDD.n5 14.864
R90 VDD.n128 VDD.n125 14.864
R91 VDD.n99 VDD.t1 14.282
R92 VDD.n99 VDD.t9 14.282
R93 VDD.n39 VDD.t3 14.282
R94 VDD.n39 VDD.t5 14.282
R95 VDD.n102 VDD.n100 9.083
R96 VDD.n23 VDD.n22 8.855
R97 VDD.n22 VDD.n21 8.855
R98 VDD.n26 VDD.n25 8.855
R99 VDD.n25 VDD.n24 8.855
R100 VDD.n30 VDD.n29 8.855
R101 VDD.n29 VDD.n28 8.855
R102 VDD.n33 VDD.n32 8.855
R103 VDD.n32 �+�X 8.855
R104 VDD.n37 VDD.n36 8.855
R105 VDD.n36 VDD.n35 8.855
R106 VDD.n43 VDD.n42 8.855
R107 VDD.n42 VDD.n41 8.855
R108 VDD.n47 VDD.n46 8.855
R109 VDD.n46 VDD.n45 8.855
R110 VDD.n61 VDD.n60 8.855
R111 VDD.n60 VDD.n59 8.855
R112 VDD.n128 VDD.n127 8.855
R113 VDD.n127 VDD.n126 8.855
R114 VDD.n111 VDD.n110 8.855
R115 VDD.n110 VDD.n109 8.855
R116 VDD.n106 VDD.n105 8.855
R117 VDD.n105 VDD.n104 8.855
R118 VDD.n102 VDD.n101 8.855
R119 VDD.n101  ,�X 8.855
R120 VDD.n97 VDD.n96 8.855
R121 VDD.n96 VDD.n95 8.855
R122 VDD.n93 VDD.n92 8.855
R123 VDD.n92 VDD.n91 8.855
R124 VDD.n89 VDD.n88 8.855
R125 VDD.n88 VDD.n87 8.855
R126 VDD.n84 VDD.n83 8.855
R127 VDD.n83 VDD.n82 8.855
R128 VDD.n125 VDD.n124 8.051
R129 VDD.n43 VDD.n40 6.193
R130 VDD.n31 VDD.n30 4.65
R131 VDD.n34 VDD.n33 4.65
R132 VDD.n38 VDD.n37 4.65
R133 VDD.n44 VDD.n43 4.65
R134 VDD.n48 VDD.n47 4.65
R135 VDD.n62 VDD.n61 4.65
R136 VDD.n129 VDD.n128 4.65
R137 VDD.n112 VDD.n111 4.65
R138 VDD.n107 VDD.n106 4.65
R139 VDD.n103 VDD.n102 4.65
R140 VDD.n98 VDD.n97 4.65
R141 VDD.n94 VDD.n93 4.65
R142 VDD.n90 VDD.n89 4.65
R143 VDD.n85 VDD.n84 4.65
R144 VDD.n27 VDD.n23 2.933
R145 VDD.n89 VDD.n86 2.89
R146 VDD.n27 VDD.n26 2.844
R147 VDD.n35 �+�X 2.557
R148 VDD.n95 VDD.t8 2.557
R149 VDD.n111 VDD.n108 2.477
R150 VDD.n31 VDD.n27 1.063
R151 VDD.n85 VDD 0.207
R152 VDD.n38 VDD.n34 0.181
R153 VDD.n103 VDD.n98 0.181
R154 VDD.n34 VDD.n31 0.145
R155 VDD.n44 VDD.n38 0.145
R156 VDD.n48 VDD.n44 0.145
R157 VDD.n62 VDD.n48 0.145
R158 VDD VDD.n62 0.145
R159 VDD VDD.n129 0.145
R160 VDD.n129 VDD.n112 0.145
R161 VDD.n112 VDD.n107 0.145
R162 VDD.n107 VDD.n103 0.145
R163 VDD.n98 VDD.n94 0.145
R164 VDD.n94 VDD.n90 0.145
R165 VDD.n90 VDD.n85 0.145
R166 a_797_1051.n1 a_797_1051.t3 228.368
R167 a_797_1051.t1 a_797_1051.n1 219.777
R168 a_797_1051.n1 a_797_1051.n0 42.29
R169 a_797_1051.n0 a_797_1051.t2 14.282
R170 a_797_1051.n0 a_797_1051.t0 14.282
R171 B.n0 B.t0 472.359
R172 B.n0 B.t1 384.527
R173 B.n1 B.t2 287.037
R174 B.n1 B.n0 210.673
R175 B.n2 B.n1 4.65
R176 B.n2 B 0.046
R177 C.n0 C.t0 470.752
R178 C.n0 C.t1 384.527
R179 C.n1 C.t2 314.896
R180 C.n1 C.n0 182.932
R181 C.n2 C.n1 4.65
R182 C.n2 C 0.046
R183 YN.n9 YN.n0 232.248
R184 YN.n8 YN.n7 208.452
R185 YN.n9 YN.n8 198.023
R186 YN.n8 YN.n3 135.417
R187 YN.n3 YN.n1 80.526
R188 YN.n7 YN.n6 30
R189 YN.n3 YN.n2 30
R190 YN.n5 YN.n4 24.383
R191 YN.n7 YN.n5 23.684
R192 YN.n0 YN.t2 14.282
R193 YN.n0 YN.t1 14.282
R194 YN.n10 YN.n9 4.65
R195 YN.n10 YN 0.046
R196 a_112_101.t0 a_112_101.n1 93.333
R197 a_112_101.n4 a_112_101.n2 79.092
R198 a_112_101.t0 a_112_101.n0 8.137
R199 a_112_101.n4 a_112_101.n3 4.614
R200 a_112_101.t0 a_112_101.n4 0.111
R201 GND.n37 GND.n36 237.558
R202 GND.n39 GND.n38 210.82
R203 GND.n52 GND.n51 166.605
R204 GND.n19 GND.n18 40.431
R205 GND.n4 GND.n3 40.003
R206 GND.n32 GND.n31 37.582
R207 GND.n51 GND.n49 23.03
R208 GND.n25 GND.n24 20.705
R209 GND.n20 GND.n19 20.705
R210 GND.n11 GND.n10 20.705
R211 GND.n5 GND.n4 20.705
R212 GND.n33 GND.n32 20.705
R213 GND.n40 GND.n39 18.953
R214 GND.n3 GND.n2 17.258
R215 GND.n31 GND.t1 15.644
R216 GND.n41 GND.n40 14.864
R217 GND.n18 GND.t0 13.654
R218 GND.n31 GND.n30 13.541
R219 GND.n22 GND.n20 9.29
R220 GND.n47 GND.n46 9.154
R221 GND.n54 GND.n53 9.154
R222 GND.n57 GND.n56 9.154
R223 GND.n60 GND.n59 9.154
R224 GND.n63 GND.n62 9.154
R225 GND.n66 GND.n65 9.154
R226 GND.n69 GND.n68 9.154
R227 GND.n41 GND.n37 9.154
R228 GND.n34 GND.n29 9.154
R229 GND.n27 GND.n26 9.154
R230 GND.n22 GND.n21 9.154
R231 GND.n15 GND.n14 9.154
R232 GND.n12 GND.n9 9.154
R233 GND.n7 GND.n6 9.154
R234 GND.n51 GND.n50 8.128
R235 GND.t0 GND.n17 7.04
R236 GND.n8 GND.n1 4.795
R237 GND.n45 GND.n44 4.65
R238 GND.n8 GND.n7 4.65
R239 GND.n13 GND.n12 4.65
R240 GND.n16 GND.n15 4.65
R241 GND.n23 GND.n22 4.65
R242 GND.n28 GND.n27 4.65
R243 GND.n35 GND.n34 4.65
R244 GND.n42 GND.n41 4.65
R245 GND.n70 GND.n69 4.65
R246 GND.n67 GND.n66 4.65
R247 GND.n64 GND.n63 4.65
R248 GND.n61 GND.n60 4.65
R249 GND.n58 GND.n57 4.65
R250 GND.n55 GND.n54 4.65
R251 GND.n48 GND.n47 4.65
R252 GND.n12 GND.n11 4.129
R253 GND.n27 GND.n25 4.129
R254 GND.n54 GND.n52 4.129
R255 GND.n7 GND.n5 1.032
R256 GND.n34 GND.n33 1.032
R257 GND.n1 GND.n0 0.474
R258 GND.n44 GND.n43 0.474
R259 GND.n45 GND 0.207
R260 GND.n23 GND.n16 0.181
R261 GND.n61 GND.n58 0.181
R262 GND.n13 GND.n8 0.145
R263 GND.n16 GND.n13 0.145
R264 GND.n28 GND.n23 0.145
R265 GND.n35 GND.n28 0.145
R266 GND.n42 GND.n35 0.145
R267 GND GND.n42 0.145
R268 GND GND.n70 0.145
R269 GND.n70 GND.n67 0.145
R270 GND.n67 GND.n64 0.145
R271 GND.n64 GND.n61 0.145
R272 GND.n58 GND.n55 0.145
R273 GND.n55 GND.n48 0.145
R274 GND.n48 GND.n45 0.145
C6 VDD GND 2.70fF
C7 a_112_101.n0 GND 0.05fF
C8 a_112_101.n1 GND 0.02fF
C9 a_112_101.n2 GND 0.11fF
C10 a_112_101.n3 GND 0.03fF
C11 a_112_101.n4 GND 0.16fF
C12 YN.n0 GND 0.49fF
C13 YN.n1 GND 0.06fF
C14 YN.n2 GND 0.03fF
C15 YN.n3 GND 0.08fF
C16 YN.n4 GND 0.04fF
C17 YN.n5 GND 0.05fF
C18 YN.n6 GND 0.03fF
C19 YN.n7 GND 0.11fF
C20 YN.n8 GND 0.49fF
C21 YN.n9 GND 0.47fF
C22 YN.n10 GND 0.01fF
C23 a_797_1051.n0 GND 0.21fF
C24 a_797_1051.n1 GND 0.50fF
C25 VDD.n1 GND 0.03fF
C26 VDD.n2 GND 0.12fF
C27 VDD.n3 GND 0.02fF
C28 VDD.n4 GND 0.02fF
C29 VDD.n5 GND 0.05fF
C30 VDD.n6 GND 0.02fF
C31 VDD.n7 GND 0.02fF
C32 VDD.n8 GND 0.02fF
C33 VDD.n9 GND 0.02fF
C34 VDD.n10 GND 0.02fF
C35 VDD.n11 GND 0.02fF
C36 VDD.n12 GND 0.02fF
C37 VDD.n13 GND 0.02fF
C38 VDD.n14 GND 0.03fF
C39 VDD.n15 GND 0.01fF
C40 VDD.n20 GND 0.39fF
C41 VDD.n21 GND 0.23fF
C42 VDD.n22 GND 0.02fF
C43 VDD.n23 GND 0.03fF
C44 VDD.n24 GND 0.21fF
C45 VDD.n25 GND 0.01fF
C46 VDD.n26 GND 0.02fF
C47 VDD.n27 GND 0.01fF
C48 VDD.n28 GND 0.14fF
C49 VDD.n29 GND 0.01fF
C50 VDD.n30 GND 0.02fF
C51 VDD.n31 GND 0.07fF
C52 VDD.n32 GND 0.01fF
C53 VDD.n33 GND 0.02fF
C54 VDD.n34 GND 0.02fF
C55 VDD.n35 GND 0.12fF
C56 VDD.n36 GND 0.01fF
C57 VDD.n37 GND 0.02fF
C58 VDD.n38 GND 0.02fF
C59 VDD.n39 GND 0.07fF
C60 VDD.n40 GND 0.04fF
C61 VDD.n41 GND 0.14fF
C62 VDD.n42 GND 0.01fF
C63 VDD.n43 GND 0.01fF
C64 VDD.n44 GND 0.02fF
C65 VDD.n45 GND 0.21fF
C66 VDD.n46 GND 0.01fF
C67 VDD.n47 GND 0.02fF
C68 VDD.n48 GND 0.02fF
C69 VDD.n49 GND 0.02fF
C70 VDD.n52 GND 0.02fF
C71 VDD.n54 GND 0.02fF
C72 VDD.n55 GND 0.19fF
C73 VDD.n56 GND 0.02fF
C74 VDD.n58 GND 0.23fF
C75 VDD.n59 GND 0.23fF
C76 VDD.n60 GND 0.01fF
C77 VDD.n61 GND 0.02fF
C78 VDD.n62 GND 0.02fF
C79 VDD.n63 GND 0.12fF
C80 VDD.n64 GND 0.02fF
C81 VDD.n65 GND 0.02fF
C82 VDD.n66 GND 0.05fF
C83 VDD.n67 GND 0.02fF
C84 VDD.n68 GND 0.02fF
C85 VDD.n69 GND 0.02fF
C86 VDD.n70 GND 0.02fF
C87 VDD.n71 GND 0.02fF
C88 VDD.n72 GND 0.02fF
C89 VDD.n73 GND 0.02fF
C90 VDD.n74 GND 0.02fF
C91 VDD.n75 GND 0.03fF
C92 VDD.n76 GND 0.03fF
C93 VDD.n77 GND 0.02fF
C94 VDD.n81 GND 0.39fF
C95 VDD.n82 GND 0.23fF
C96 VDD.n83 GND 0.02fF
C97 VDD.n84 GND 0.03fF
C98 VDD.n85 GND 0.02fF
C99 VDD.n86 GND 0.05fF
C100 VDD.n87 GND 0.21fF
C101 VDD.n88 GND 0.01fF
C102 VDD.n89 GND 0.01fF
C103 VDD.n90 GND 0.02fF
C104 VDD.n91 GND 0.14fF
C105 VDD.n92 GND 0.01fF
C106 VDD.n93 GND 0.02fF
C107 VDD.n94 GND 0.02fF
C108 VDD.n95 GND 0.12fF
C109 VDD.n96 GND 0.01fF
C110 VDD.n97 GND 0.02fF
C111 VDD.n98 GND 0.02fF
C112 VDD.n99 GND 0.07fF
C113 VDD.n100 GND 0.04fF
C114 VDD.n101 GND 0.01fF
C115 VDD.n102 GND 0.02fF
C116 VDD.n103 GND 0.02fF
C117 VDD.n104 GND 0.14fF
C118 VDD.n105 GND 0.01fF
C119 VDD.n106 GND 0.02fF
C120 VDD.n107 GND 0.02fF
C121 VDD.n108 GND 0.05fF
C122 VDD.n109 GND 0.21fF
C123 VDD.n110 GND 0.01fF
C124 VDD.n111 GND 0.01fF
C125 VDD.n112 GND 0.02fF
C126 VDD.n113 GND 0.05fF
C127 VDD.n114 GND 0.02fF
C128 VDD.n115 GND 0.02fF
C129 VDD.n116 GND 0.02fF
C130 VDD.n117 GND 0.02fF
C131 VDD.n118 GND 0.02fF
C132 VDD.n119 GND 0.02fF
C133 VDD.n120 GND 0.02fF
C134 VDD.n121 GND 0.02fF
C135 VDD.n122 GND 0.02fF
C136 VDD.n123 GND 0.02fF
C137 VDD.n124 GND 0.02fF
C138 VDD.n125 GND 0.02fF
C139 VDD.n126 GND 0.23fF
C140 VDD.n127 GND 0.01fF
C141 VDD.n128 GND 0.02fF
C142 VDD.n129 GND 0.02fF
C143 a_217_1050.n0 GND 0.29fF
C144 a_217_1050.n1 GND 0.37fF
C145 a_217_1050.n2 GND 0.51fF
C146 a_217_1050.n3 GND 0.31fF
C147 a_217_1050.n4 GND 0.44fF
C148 a_217_1050.n5 GND 0.