* NGSPICE file created from NOR2X1.ext - technology: sky130A

.subckt pmos2_1 a_144_n460# a_262_n399# a_88_n399# w_52_n435# a_174_n399#
X0 a_174_n399# a_144_n460# a_88_n399# w_52_n435# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.6e+11p ps=4.56e+06u w=2e+06u l=150000u
X1 a_262_n399# a_144_n460# a_174_n399# w_52_n435# sky130_fd_pr__pfet_01v8 ad=5.4e+11p pd=4.54e+06u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt nmos_top_trim1 a_56_92# a_86_108# a_0_0# VSUBS
X0 a_86_108# a_56_92# a_0_0# VSUBS sky130_fd_pr__nfet_01v8 ad=1.772e+11p pd=1.56e+06u as=1.15725e+12p ps=8.12e+06u w=3e+06u l=150000u
.ends

.subckt nmos_top_trim2 a_56_92# a_86_108# a_0_0# VSUBS
X0 a_86_108# a_56_92# a_0_0# VSUBS sky130_fd_pr__nfet_01v8 ad=1.772e+11p pd=1.56e+06u as=1.15725e+12p ps=8.12e+06u w=3e+06u l=150000u
.ends

.subckt nor2x1_pcell VDD VSS a_168_403# a_362_410# a_405_1105#
Xpmos2_1_0 a_168_403# a_317_1377# a_317_1377# VDD VDD pmos2_1
Xpmos2_1_1 a_362_410# a_317_1377# a_317_1377# VDD a_405_1105# pmos2_1
Xnmos_top_trim1_1 a_168_403# a_405_1105# VSS VSS nmos_top_trim1
Xnmos_top_trim2_0 a_362_410# a_405_1105# VSS VSS nmos_top_trim2
.ends

.subckt NOR2X1 A B Y VSS VDD
Xnor2x1_pcell_0 VDD VSS A B Y nor2x1_pcell
.ends

