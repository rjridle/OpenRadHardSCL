* SPICE3 file created from DFFSNQNX1.ext - technology: sky130A

.subckt DFFSNQNX1 QN D CLK SN VDD VSS
X0 VDD D a_217_1050 VDD sky130_fd_pr__pfet_01v8 ad=1.182p pd=9.582u as=0p ps=0u w=2u l=0.15u M=2
X1 VDD a_1265_989 a_1905_1050 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X2 a_3599_411 a_1265_989 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X3 a_1265_989 CLK a_2702_101 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X4 a_1905_1050 a_217_1050 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X5 a_4294_210 SN a_4013_103 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X6 VDD a_343_411 a_217_1050 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X7 VDD a_217_1050 a_343_411 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X8 QN a_3599_411 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.16p pd=9.16u as=0p ps=0u w=2u l=0.15u M=2
X9 a_1905_1050 a_1265_989 a_2000_210 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X10 VDD CLK a_343_411 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X11 QN a_343_411 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X12 VDD a_1905_1050 a_1265_989 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X13 a_343_411 a_1265_989 a_1038_210 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X14 VDD QN a_3599_411 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X15 VSS a_217_1050 a_757_103 VSS sky130_fd_pr__nfet_01v8 ad=1.0746p pd=9.42u as=0p ps=0u w=3u l=0.15u
X16 VDD a_1265_989 a_343_411 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X17 VSS D a_112_101 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X18 VSS a_343_411 a_3368_101 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X19 VDD SN a_3599_411 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X20 a_1905_1050 SN VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X21 VSS a_217_1050 a_1719_103 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X22 a_1038_210 CLK a_757_103 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X23 VSS a_1905_1050 a_2702_101 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X24 a_217_1050 a_343_411 a_112_101 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X25 VDD CLK a_1265_989 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X26 a_2000_210 SN a_1719_103 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X27 a_3599_411 a_1265_989 a_4294_210 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X28 QN a_3599_411 a_3368_101 VSS sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=0p ps=0u w=3u l=0.15u
X29 VSS QN a_4013_103 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
C0 a_217_1050 VDD 2.52fF
C1 a_343_411 CLK 2.41fF
C2 a_343_411 VDD 6.03fF
C3 a_1265_989 a_343_411 3.02fF
C4 QN VDD 2.20fF
C5 a_3599_411 VDD 2.82fF
C6 a_1265_989 VDD 2.79fF
C7 a_1905_1050 VDD 2.82fF
C8 VDD VSS 7.98fF
.ends
