magic
tech sky130A
magscale 1 2
timestamp 1645050624
<< locali >>
rect -33 -17 -17 17
rect 17 -17 33 17
<< viali >>
rect -17 -17 17 17
<< metal1 >>
rect -17 23 17 53
rect -23 17 23 23
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -23 23 -17
rect -17 -29 17 -23
<< end >>
