* SPICE3 file created from BUFX1.ext - technology: sky130A

.subckt BUFX1 Y A VDD GND
X0 a_185_209.t2 A.t0 VDD.t5  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X1 VDD.t7 a_185_209.t3 Y.t2 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X2 Y a_185_209.t5 GND.t0 GND sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=0p ps=0u w=0u l=0u
X3 VDD.t3 A.t2 a_185_209.t1  �.�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X4 Y.t1 a_185_209.t4 VDD.t1 �.�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
C0 VDD A 0.38fF
C1 Y VDD 1.08fF
R0 A.n0 A.t2 512.525
R1 A.n0 A.t0 371.139
R2 A.n1 A.t1 282.852
R3 A.n1 A.n0 247.347
R4 A.n2 A.n1 4.65
R5 A.n2 A 0.046
R6 VDD.n103 VDD.n101 144.705
R7 VDD.n76 VDD.t5 135.17
R8 VDD.n83 VDD.t3 135.17
R9 VDD.n33 VDD.t1 135.17
R10 VDD.n24 VDD.t7 135.17
R11 VDD.n97 VDD.n96 92.5
R12 VDD.n95 VDD.n94 92.5
R13 VDD.n93 VDD.n92 92.5
R14 VDD.n91 VDD.n90 92.5
R15 VDD.n99 VDD.n98 92.5
R16 VDD.n62 VDD.n61 92.5
R17 VDD.n60 VDD.n59 92.5
R18 VDD.n58 VDD.n57 92.5
R19 VDD.n56 VDD.n55 92.5
R20 VDD.n64 VDD.n63 92.5
R21 VDD.n14 VDD.n1 92.5
R22 VDD.n5 VDD.n4 92.5
R23 VDD.n7 VDD.n6 92.5
R24 VDD.n9 VDD.n8 92.5
R25 VDD.n11 VDD.n10 92.5
R26 VDD.n13 VDD.n12 92.5
R27 VDD.n21 VDD.n20 92.059
R28 VDD.n47 VDD.n46 92.059
R29 VDD.n70 VDD.n69 92.059
R30 VDD.n20 VDD.n16 67.194
R31 VDD.n20 VDD.n17 67.194
R32 VDD.n20 VDD.n18 67.194
R33 VDD.n20 VDD.n19 67.194
R34 VDD.n54 VDD.n53 44.141
R35 VDD.n5 VDD.n3 44.141
R36 VDD.n53 VDD.n51 44.107
R37 VDD.n3 VDD.n2 44.107
R38 VDD.n25 VDD.t6 43.472
R39 VDD.n34 �.�� 43.472
R40 VDD.n84  �.�� 43.472
R41 VDD.n74 ���+V 43.472
R42 VDD.n20 VDD.n15 41.052
R43 VDD.n66 VDD.n65 39.742
R44 VDD.n45 VDD.n42 39.742
R45 VDD.n45 VDD.n44 39.742
R46 VDD.n41 VDD.n40 39.742
R47 VDD.n53 VDD.n52 38
R48 VDD.n44 VDD.n43 36.774
R49 VDD.n1 VDD.n0 30.923
R50 VDD.n69 VDD.n67 26.38
R51 VDD.n69 VDD.n66 26.38
R52 VDD.n69 VDD.n68 26.38
R53 VDD.n46 VDD.n45 26.38
R54 VDD.n46 VDD.n41 26.38
R55 VDD.n46 VDD.n39 26.38
R56 VDD.n46 VDD.n38 26.38
R57 VDD.n72 VDD.n64 22.915
R58 VDD.n23 VDD.n14 22.915
R59 VDD.n64 VDD.n62 14.864
R60 VDD.n62 VDD.n60 14.864
R61 VDD.n60 VDD.n58 14.864
R62 VDD.n58 VDD.n56 14.864
R63 VDD.n56 VDD.n54 14.864
R64 VDD.n99 VDD.n97 14.864
R65 VDD.n97 VDD.n95 14.864
R66 VDD.n95 VDD.n93 14.864
R67 VDD.n93 VDD.n91 14.864
R68 VDD.n91 VDD.n89 14.864
R69 VDD.n89 VDD.n88 14.864
R70 VDD.n14 VDD.n13 14.864
R71 VDD.n13 VDD.n11 14.864
R72 VDD.n11 VDD.n9 14.864
R73 VDD.n9 VDD.n7 14.864
R74 VDD.n7 VDD.n5 14.864
R75 VDD.n104 VDD.n100 14.864
R76 VDD.n23 VDD.n22 8.855
R77 VDD.n22 VDD.n21 8.855
R78 VDD.n27 VDD.n26 8.855
R79 VDD.n26 VDD.n25 8.855
R80 VDD.n31 VDD.n30 8.855
R81 VDD.n30 VDD.n29 8.855
R82 VDD.n36 VDD.n35 8.855
R83 VDD.n35 VDD.n34 8.855
R84 VDD.n49 VDD.n48 8.855
R85 VDD.n48 VDD.n47 8.855
R86 VDD.n104 VDD.n103 8.855
R87 VDD.n103 VDD.n102 8.855
R88 VDD.n86 VDD.n85 8.855
R89 VDD.n85 VDD.n84 8.855
R90 VDD.n81 VDD.n80 8.855
R91 VDD.n80 VDD.n79 8.855
R92 VDD.n77 VDD.n75 8.855
R93 VDD.n75 VDD.n74 8.855
R94 VDD.n72 VDD.n71 8.855
R95 VDD.n71 VDD.n70 8.855
R96 VDD.n100 VDD.n99 8.051
R97 VDD.n28 VDD.n23 4.795
R98 VDD.n28 VDD.n27 4.65
R99 VDD.n32 VDD.n31 4.65
R100 VDD.n37 VDD.n36 4.65
R101 VDD.n50 VDD.n49 4.65
R102 VDD.n105 VDD.n104 4.65
R103 VDD.n87 VDD.n86 4.65
R104 VDD.n82 VDD.n81 4.65
R105 VDD.n78 VDD.n77 4.65
R106 VDD.n73 VDD.n72 4.65
R107 VDD.n27 VDD.n24 2.064
R108 VDD.n36 VDD.n33 2.064
R109 VDD.n86 VDD.n83 2.064
R110 VDD.n77 VDD.n76 2.064
R111 VDD.n73 VDD 0.207
R112 VDD.n32 VDD.n28 0.157
R113 VDD.n37 VDD.n32 0.157
R114 VDD.n87 VDD.n82 0.157
R115 VDD.n82 VDD.n78 0.157
R116 VDD.n50 VDD.n37 0.145
R117 VDD VDD.n50 0.145
R118 VDD VDD.n105 0.145
R119 VDD.n105 VDD.n87 0.145
R120 VDD.n78 VDD.n73 0.145
R121 a_185_209.n0 a_185_209.t3 512.525
R122 a_185_209.n0 a_185_209.t4 371.139
R123 a_185_209.n7 a_185_209.n6 326.998
R124 a_185_209.n1 a_185_209.n0 303.065
R125 a_185_209.n1 a_185_209.t5 227.134
R126 a_185_209.n6 a_185_209.n5 216.733
R127 a_185_209.n5 a_185_209.n4 30
R128 a_185_209.n3 a_185_209.n2 24.383
R129 a_185_209.n5 a_185_209.n3 23.684
R130 a_185_209.n7 a_185_209.t1 14.282
R131 a_185_209.t2 a_185_209.n7 14.282
R132 a_185_209.n6 a_185_209.n1 10.343
R133 GND.n60 GND.n59 237.558
R134 GND.n29 GND.n28 210.82
R135 GND.n5 GND.n4 120.01
R136 GND.n3 GND.n2 92.5
R137 GND.n12 GND.n11 92.5
R138 GND.n22 GND.t0 45.413
R139 GND.n22 GND.n21 39.307
R140 GND.n43 GND.n42 37.582
R141 GND.t1 GND.n40 32.601
R142 GND.n23 GND.n22 23.77
R143 GND.n40 GND.n39 21.734
R144 GND.n6 GND.n5 20.705
R145 GND.n14 GND.n13 20.705
R146 GND.n24 GND.n23 20.705
R147 GND.n55 GND.n54 20.705
R148 GND.n49 GND.n48 20.705
R149 GND.n44 GND.n43 20.705
R150 GND.n5 GND.n3 19.952
R151 GND.n54 GND.n53 19.952
R152 GND.n30 GND.n29 18.953
R153 GND.n42 GND.t1 15.644
R154 GND.n31 GND.n30 14.864
R155 GND.n42 GND.n41 13.541
R156 GND.n45 GND.n36 9.154
R157 GND.n51 GND.n50 9.154
R158 GND.n57 GND.n56 9.154
R159 GND.n61 GND.n60 9.154
R160 GND.n31 GND.n27 9.154
R161 GND.n25 GND.n18 9.154
R162 GND.n16 GND.n15 9.154
R163 GND.n8 GND.n7 9.154
R164 GND.n9 GND.n1 4.795
R165 GND.n35 GND.n34 4.65
R166 GND.n9 GND.n8 4.65
R167 GND.n17 GND.n16 4.65
R168 GND.n26 GND.n25 4.65
R169 GND.n32 GND.n31 4.65
R170 GND.n62 GND.n61 4.65
R171 GND.n58 GND.n57 4.65
R172 GND.n52 GND.n51 4.65
R173 GND.n46 GND.n45 4.65
R174 GND.n20 GND.n19 4.504
R175 GND.n38 GND.n37 4.504
R176 GND.n8 GND.n6 4.129
R177 GND.n57 GND.n55 4.129
R178 GND.n25 GND.n24 3.716
R179 GND.n45 GND.n44 3.716
R180 GND.t0 GND.n20 2.452
R181 GND.t1 GND.n38 2.452
R182 GND.n11 GND.n10 1.935
R183 GND.n1 GND.n0 0.474
R184 GND.n34 GND.n33 0.474
R185 GND.n13 GND.n12 0.376
R186 GND.n48 GND.n47 0.376
R187 GND.n35 GND 0.207
R188 GND.n16 GND.n14 0.206
R189 GND.n51 GND.n49 0.206
R190 GND.n17 GND.n9 0.157
R191 GND.n26 GND.n17 0.157
R192 GND.n58 GND.n52 0.157
R193 GND.n52 GND.n46 0.157
R194 GND.n32 GND.n26 0.145
R195 GND GND.n32 0.145
R196 GND GND.n62 0.145
R197 GND.n62 GND.n58 0.145
R198 GND.n46 GND.n35 0.145
R199 Y.n2 Y.n1 294.19
R200 Y.n2 Y.n0 271.281
R201 Y.n0 Y.t2 14.282
R202 Y.n0 Y.t1 14.282
R203 Y.n3 Y.n2 4.65
R204 Y.n3 Y 0.046
C2 VDD GND 1.62fF
C3 Y.n0 GND 0.64fF
C4 Y.n1 GND 0.30fF
C5 Y.n2 GND 0.64fF
C6 Y.n3 GND 0.01fF
C7 a_185_209.n0 GND 0.31fF
C8 a_185_209.n1 GND 0.44fF
C9 a_185_209.n2 GND 0.03fF
C10 a_185_209.n3 GND 0.04fF
C11 a_185_209.n4 GND 0.03fF
C12 a_185_209.n5 GND 0.10fF
C13 a_185_209.n6 GND 0.59fF
C14 a_185_209.n7 GND 0.55fF
C15 VDD.n1 GND 0.02fF
C16 VDD.n2 GND 0.06fF
C17 VDD.n3 GND 0.02fF
C18 VDD.n4 GND 0.01fF
C19 VDD.n5 GND 0.04fF
C20 VDD.n6 GND 0.01fF
C21 VDD.n7 GND 0.01fF
C22 VDD.n8 GND 0.01fF
C23 VDD.n9 GND 0.01fF
C24 VDD.n10 GND 0.01fF
C25 VDD.n11 GND 0.01fF
C26 VDD.n12 GND 0.01fF
C27 VDD.n13 GND 0.01fF
C28 VDD.n14 GND 0.02fF
C29 VDD.n15 GND 0.01fF
C30 VDD.n20 GND 0.30fF
C31 VDD.n21 GND 0.18fF
C32 VDD.n22 GND 0.01fF
C33 VDD.n23 GND 0.02fF
C34 VDD.n24 GND 0.04fF
C35 VDD.n25 GND 0.13fF
C36 VDD.n26 GND 0.01fF
C37 VDD.n27 GND 0.01fF
C38 VDD.n28 GND 0.04fF
C39 VDD.n29 GND 0.11fF
C40 VDD.n30 GND 0.01fF
C41 VDD.n31 GND 0.02fF
C42 VDD.n32 GND 0.02fF
C43 VDD.n33 GND 0.04fF
C44 VDD.n34 GND 0.13fF
C45 VDD.n35 GND 0.01fF
C46 VDD.n36 GND 0.01fF
C47 VDD.n37 GND 0.02fF
C48 VDD.n40 GND 0.01fF
C49 VDD.n42 GND 0.01fF
C50 VDD.n43 GND 0.10fF
C51 VDD.n44 GND 0.01fF
C52 VDD.n46 GND 0.18fF
C53 VDD.n47 GND 0.18fF
C54 VDD.n48 GND 0.01fF
C55 VDD.n49 GND 0.01fF
C56 VDD.n50 GND 0.01fF
C57 VDD.n51 GND 0.06fF
C58 VDD.n52 GND 0.01fF
C59 VDD.n53 GND 0.01fF
C60 VDD.n54 GND 0.04fF
C61 VDD.n55 GND 0.01fF
C62 VDD.n56 GND 0.01fF
C63 VDD.n57 GND 0.01fF
C64 VDD.n58 GND 0.01fF
C65 VDD.n59 GND 0.01fF
C66 VDD.n60 GND 0.01fF
C67 VDD.n61 GND 0.01fF
C68 VDD.n62 GND 0.01fF
C69 VDD.n63 GND 0.02fF
C70 VDD.n64 GND 0.02fF
C71 VDD.n65 GND 0.01fF
C72 VDD.n69 GND 0.30fF
C73 VDD.n70 GND 0.18fF
C74 VDD.n71 GND 0.01fF
C75 VDD.n72 GND 0.02fF
C76 VDD.n73 GND 0.02fF
C77 VDD.n74 GND 0.13fF
C78 VDD.n75 GND 0.01fF
C79 VDD.n76 GND 0.04fF
C80 VDD.n77 GND 0.01fF
C81 VDD.n78 GND 0.02fF
C82 VDD.n79 GND 0.11fF
C83 VDD.n80 GND 0.01fF
C84 VDD.n81 GND 0.02fF
C85 VDD.n82 GND 0.02fF
C86 VDD.n83 GND 0.04fF
C87 VDD.n84 GND 0.13fF
C88 VDD.n85 GND 0.01fF
C89 VDD.n86 GND 0.01fF
C90 VDD.n87 GND 0.02fF
C91 VDD.n88 GND 0.04fF
C92 VDD.n89 GND 0.01fF
C93 VDD.n9