magic
tech sky130A
magscale 1 2
timestamp 1642379819
<< error_p >>
rect 85 322 86 323
rect 269 322 270 323
rect 86 321 87 322
rect 270 321 271 322
rect 101 291 102 292
rect 136 291 137 292
rect 285 291 286 292
rect 320 291 321 292
rect 101 188 102 189
rect 136 188 137 189
rect 285 188 286 189
rect 320 188 321 189
<< nwell >>
rect -36 591 464 1353
<< nmos >>
rect 56 322 86 375
rect 240 322 270 375
rect 56 292 152 322
tri 152 292 182 322 sw
rect 56 188 86 292
tri 86 276 102 292 nw
tri 136 276 152 292 ne
tri 86 188 102 204 sw
tri 136 188 152 204 se
rect 152 188 182 292
rect 240 292 336 322
tri 336 292 366 322 sw
tri 56 158 86 188 ne
rect 86 158 152 188
tri 152 158 182 188 nw
rect 240 188 270 292
tri 270 276 286 292 nw
tri 320 276 336 292 ne
tri 270 188 286 204 sw
tri 320 188 336 204 se
rect 336 188 366 292
tri 240 158 270 188 ne
rect 270 158 336 188
tri 336 158 366 188 nw
<< pmos >>
rect 64 629 94 1229
rect 152 629 182 1229
rect 240 629 270 1229
rect 328 629 358 1229
<< ndiff >>
rect 0 298 56 375
rect 86 322 240 375
rect 270 322 420 375
rect 0 264 10 298
rect 44 264 56 298
tri 152 292 182 322 ne
rect 182 298 240 322
rect 0 215 56 264
rect 0 181 10 215
rect 44 181 56 215
tri 86 276 102 292 se
rect 102 276 136 292
tri 136 276 152 292 sw
rect 86 242 152 276
rect 86 208 98 242
rect 132 208 152 242
rect 86 204 152 208
tri 86 188 102 204 ne
rect 102 188 136 204
tri 136 188 152 204 nw
rect 182 264 194 298
rect 228 264 240 298
tri 336 292 366 322 ne
rect 366 298 420 322
rect 182 215 240 264
rect 0 158 56 181
tri 56 158 86 188 sw
tri 152 158 182 188 se
rect 182 181 194 215
rect 228 181 240 215
tri 270 276 286 292 se
rect 286 276 320 292
tri 320 276 336 292 sw
rect 270 242 336 276
rect 270 208 282 242
rect 316 208 336 242
rect 270 204 336 208
tri 270 188 286 204 ne
rect 286 188 320 204
tri 320 188 336 204 nw
rect 366 264 378 298
rect 412 264 420 298
rect 366 215 420 264
rect 182 158 240 181
tri 240 158 270 188 sw
tri 336 158 366 188 se
rect 366 181 378 215
rect 412 181 420 215
rect 366 158 420 181
rect 0 147 420 158
rect 0 113 10 147
rect 44 113 98 147
rect 132 113 194 147
rect 228 113 282 147
rect 316 113 378 147
rect 412 113 420 147
rect 0 101 420 113
<< pdiff >>
rect 10 1213 64 1229
rect 10 1179 18 1213
rect 52 1179 64 1213
rect 10 1145 64 1179
rect 10 1111 18 1145
rect 52 1111 64 1145
rect 10 1077 64 1111
rect 10 1043 18 1077
rect 52 1043 64 1077
rect 10 1009 64 1043
rect 10 975 18 1009
rect 52 975 64 1009
rect 10 941 64 975
rect 10 907 18 941
rect 52 907 64 941
rect 10 873 64 907
rect 10 839 18 873
rect 52 839 64 873
rect 10 805 64 839
rect 10 771 18 805
rect 52 771 64 805
rect 10 737 64 771
rect 10 703 18 737
rect 52 703 64 737
rect 10 629 64 703
rect 94 1213 152 1229
rect 94 1179 106 1213
rect 140 1179 152 1213
rect 94 1145 152 1179
rect 94 1111 106 1145
rect 140 1111 152 1145
rect 94 1077 152 1111
rect 94 1043 106 1077
rect 140 1043 152 1077
rect 94 1009 152 1043
rect 94 975 106 1009
rect 140 975 152 1009
rect 94 941 152 975
rect 94 907 106 941
rect 140 907 152 941
rect 94 873 152 907
rect 94 839 106 873
rect 140 839 152 873
rect 94 805 152 839
rect 94 771 106 805
rect 140 771 152 805
rect 94 737 152 771
rect 94 703 106 737
rect 140 703 152 737
rect 94 629 152 703
rect 182 1213 240 1229
rect 182 1179 194 1213
rect 228 1179 240 1213
rect 182 1145 240 1179
rect 182 1111 194 1145
rect 228 1111 240 1145
rect 182 1077 240 1111
rect 182 1043 194 1077
rect 228 1043 240 1077
rect 182 1009 240 1043
rect 182 975 194 1009
rect 228 975 240 1009
rect 182 941 240 975
rect 182 907 194 941
rect 228 907 240 941
rect 182 873 240 907
rect 182 839 194 873
rect 228 839 240 873
rect 182 805 240 839
rect 182 771 194 805
rect 228 771 240 805
rect 182 737 240 771
rect 182 703 194 737
rect 228 703 240 737
rect 182 629 240 703
rect 270 1213 328 1229
rect 270 1179 282 1213
rect 316 1179 328 1213
rect 270 1145 328 1179
rect 270 1111 282 1145
rect 316 1111 328 1145
rect 270 1077 328 1111
rect 270 1043 282 1077
rect 316 1043 328 1077
rect 270 1009 328 1043
rect 270 975 282 1009
rect 316 975 328 1009
rect 270 941 328 975
rect 270 907 282 941
rect 316 907 328 941
rect 270 873 328 907
rect 270 839 282 873
rect 316 839 328 873
rect 270 805 328 839
rect 270 771 282 805
rect 316 771 328 805
rect 270 737 328 771
rect 270 703 282 737
rect 316 703 328 737
rect 270 629 328 703
rect 358 1213 412 1229
rect 358 1179 370 1213
rect 404 1179 412 1213
rect 358 1145 412 1179
rect 358 1111 370 1145
rect 404 1111 412 1145
rect 358 1077 412 1111
rect 358 1043 370 1077
rect 404 1043 412 1077
rect 358 1009 412 1043
rect 358 975 370 1009
rect 404 975 412 1009
rect 358 941 412 975
rect 358 907 370 941
rect 404 907 412 941
rect 358 873 412 907
rect 358 839 370 873
rect 404 839 412 873
rect 358 805 412 839
rect 358 771 370 805
rect 404 771 412 805
rect 358 737 412 771
rect 358 703 370 737
rect 404 703 412 737
rect 358 629 412 703
<< ndiffc >>
rect 10 264 44 298
rect 10 181 44 215
rect 98 208 132 242
rect 194 264 228 298
rect 194 181 228 215
rect 282 208 316 242
rect 378 264 412 298
rect 378 181 412 215
rect 10 113 44 147
rect 98 113 132 147
rect 194 113 228 147
rect 282 113 316 147
rect 378 113 412 147
<< pdiffc >>
rect 18 1179 52 1213
rect 18 1111 52 1145
rect 18 1043 52 1077
rect 18 975 52 1009
rect 18 907 52 941
rect 18 839 52 873
rect 18 771 52 805
rect 18 703 52 737
rect 106 1179 140 1213
rect 106 1111 140 1145
rect 106 1043 140 1077
rect 106 975 140 1009
rect 106 907 140 941
rect 106 839 140 873
rect 106 771 140 805
rect 106 703 140 737
rect 194 1179 228 1213
rect 194 1111 228 1145
rect 194 1043 228 1077
rect 194 975 228 1009
rect 194 907 228 941
rect 194 839 228 873
rect 194 771 228 805
rect 194 703 228 737
rect 282 1179 316 1213
rect 282 1111 316 1145
rect 282 1043 316 1077
rect 282 975 316 1009
rect 282 907 316 941
rect 282 839 316 873
rect 282 771 316 805
rect 282 703 316 737
rect 370 1179 404 1213
rect 370 1111 404 1145
rect 370 1043 404 1077
rect 370 975 404 1009
rect 370 907 404 941
rect 370 839 404 873
rect 370 771 404 805
rect 370 703 404 737
<< psubdiff >>
rect 0 13 24 47
rect 58 13 92 47
rect 126 13 160 47
rect 194 13 228 47
rect 262 13 296 47
rect 330 13 364 47
rect 398 13 428 47
<< nsubdiff >>
rect 0 1283 24 1317
rect 58 1283 92 1317
rect 126 1283 160 1317
rect 195 1283 229 1317
rect 263 1283 297 1317
rect 331 1283 365 1317
rect 399 1283 428 1317
<< psubdiffcont >>
rect 24 13 58 47
rect 92 13 126 47
rect 160 13 194 47
rect 228 13 262 47
rect 296 13 330 47
rect 364 13 398 47
<< nsubdiffcont >>
rect 24 1283 58 1317
rect 92 1283 126 1317
rect 160 1283 195 1317
rect 229 1283 263 1317
rect 297 1283 331 1317
rect 365 1283 399 1317
<< poly >>
rect 64 1229 94 1255
rect 152 1229 182 1255
rect 240 1229 270 1255
rect 328 1229 358 1255
rect 64 612 94 629
rect 152 612 182 629
rect 240 612 270 629
rect 328 612 358 629
rect 64 582 358 612
rect 240 540 270 582
rect 204 524 270 540
rect 204 490 214 524
rect 248 490 270 524
rect 204 474 270 490
rect 240 429 270 474
rect 56 399 270 429
rect 56 375 86 399
rect 240 375 270 399
<< polycont >>
rect 214 490 248 524
<< locali >>
rect 0 1317 428 1332
rect 0 1283 24 1317
rect 58 1283 92 1317
rect 126 1283 160 1317
rect 195 1283 229 1317
rect 263 1283 297 1317
rect 331 1283 365 1317
rect 399 1283 428 1317
rect 0 1270 428 1283
rect 18 1213 52 1270
rect 18 1145 52 1179
rect 18 1077 52 1111
rect 18 1009 52 1043
rect 18 941 52 975
rect 18 873 52 907
rect 18 805 52 839
rect 18 737 52 771
rect 18 627 52 703
rect 106 1213 140 1229
rect 106 1145 140 1179
rect 106 1077 140 1111
rect 106 1009 140 1043
rect 106 941 140 975
rect 106 873 140 907
rect 106 805 140 839
rect 106 737 140 771
rect 106 672 140 703
rect 194 1213 228 1270
rect 194 1145 228 1179
rect 194 1077 228 1111
rect 194 1009 228 1043
rect 194 941 228 975
rect 194 873 228 907
rect 194 805 228 839
rect 194 737 228 771
rect 194 627 228 703
rect 282 1213 316 1229
rect 282 1145 316 1179
rect 282 1077 316 1111
rect 282 1009 316 1043
rect 282 941 316 975
rect 282 873 316 907
rect 282 805 316 839
rect 282 737 316 771
rect 282 673 316 703
rect 214 524 248 540
rect 214 474 248 490
rect 10 298 44 343
rect 194 298 228 343
rect 10 215 44 264
rect 98 278 132 287
rect 98 242 132 244
rect 98 192 132 208
rect 194 215 228 264
rect 10 147 44 181
rect 282 278 316 638
rect 370 1213 404 1270
rect 370 1145 404 1179
rect 370 1077 404 1111
rect 370 1009 404 1043
rect 370 941 404 975
rect 370 873 404 907
rect 370 805 404 839
rect 370 737 404 771
rect 370 627 404 703
rect 282 242 316 244
rect 282 192 316 208
rect 378 298 412 343
rect 378 215 412 264
rect 194 147 228 181
rect 378 147 412 181
rect 44 113 98 147
rect 132 113 194 147
rect 228 113 282 147
rect 316 113 378 147
rect 10 62 44 113
rect 194 62 228 113
rect 378 62 412 113
rect 0 47 428 62
rect 0 13 24 47
rect 58 13 92 47
rect 126 13 160 47
rect 194 13 228 47
rect 262 13 296 47
rect 330 13 364 47
rect 398 13 428 47
rect 0 0 428 13
<< viali >>
rect 24 1283 58 1317
rect 92 1283 126 1317
rect 160 1283 195 1317
rect 229 1283 263 1317
rect 297 1283 331 1317
rect 365 1283 399 1317
rect 106 638 140 672
rect 282 638 316 673
rect 214 490 248 524
rect 98 244 132 278
rect 282 244 316 278
rect 24 13 58 47
rect 92 13 126 47
rect 160 13 194 47
rect 228 13 262 47
rect 296 13 330 47
rect 364 13 398 47
<< metal1 >>
rect 0 1317 428 1332
rect 0 1283 24 1317
rect 58 1283 92 1317
rect 126 1283 160 1317
rect 195 1283 229 1317
rect 263 1283 297 1317
rect 331 1283 365 1317
rect 399 1283 428 1317
rect 0 1270 428 1283
rect 94 672 151 678
rect 270 673 328 679
rect 270 672 282 673
rect 94 638 106 672
rect 140 638 282 672
rect 316 638 328 673
rect 94 632 151 638
rect 270 632 328 638
rect 282 629 316 632
rect 214 531 248 548
rect 208 524 254 531
rect 208 490 214 524
rect 248 490 254 524
rect 208 483 254 490
rect 214 467 248 483
rect 98 285 132 290
rect 282 285 316 290
rect 92 278 138 285
rect 276 278 322 285
rect 92 244 98 278
rect 132 244 282 278
rect 316 244 322 278
rect 92 237 138 244
rect 276 237 322 244
rect 98 232 132 237
rect 282 232 316 237
rect 0 47 428 62
rect 0 13 24 47
rect 58 13 92 47
rect 126 13 160 47
rect 194 13 228 47
rect 262 13 296 47
rect 330 13 364 47
rect 398 13 428 47
rect 0 0 428 13
<< labels >>
rlabel metal1 281 1301 281 1301 1 VDD
port 1 n
rlabel metal1 229 503 229 503 1 A
port 2 n
rlabel metal1 297 653 297 653 1 Y
port 3 n
rlabel metal1 278 26 278 26 1 VSS
port 4 n
<< end >>
