* HSPICE file created from tmp.ext - technology: sky130A

.option scale=5000u

.subckt tmp Y A B VDD VSS
X0 a_131_1051 A VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=33600 ps=1368 w=400 l=30 M=2
X1 Y a_198_209 VDD VDD sky130_fd_pr__pfet_01v8 ad=11600 pd=458 as=0 ps=0 w=400 l=30 M=2
X2 a_198_209 A VSS VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=123966 ps=4212 w=598 l=30
X3 a_131_1051 B a_198_209 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=400 l=30 M=2
X4 a_198_209 B VSS VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=598 l=30
X5 Y a_198_209 VSS VSS sky130_fd_pr__nfet_01v8 ad=7088 pd=312 as=0 ps=0 w=598 l=30
.ends

** hspice subcircuit dictionary
