magic
tech sky130A
magscale 1 2
timestamp 1648048189
<< nwell >>
rect 55 1505 89 1539
<< psubdiffcont >>
rect 55 13 89 47
<< nsubdiffcont >>
rect 55 1505 89 1539
<< viali >>
rect 55 1505 89 1539
rect 55 13 89 47
<< metal1 >>
rect 907 871 2780 905
rect 205 797 239 831
rect 537 797 1822 831
rect 2313 797 3429 831
rect 3941 797 4684 831
rect 4719 797 4753 831
rect 1351 723 3683 757
rect 4053 723 4087 757
rect 4123 723 4569 757
rect 2461 649 2909 683
rect 406 575 4398 609
use nand3x1_pcell  nand3x1_pcell_0 pcells
timestamp 1647328266
transform 1 0 666 0 1 0
box -84 0 1046 1575
use nand2x1_pcell  nand2x1_pcell_5 pcells
timestamp 1647328257
transform 1 0 0 0 1 0
box -84 0 750 1575
use li1_M1_contact  li1_M1_contact_20 pcells
timestamp 1646004885
transform 1 0 222 0 1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_5
timestamp 1646004885
transform -1 0 888 0 -1 888
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_3
timestamp 1646004885
transform -1 0 518 0 -1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_1
timestamp 1646004885
transform -1 0 370 0 -1 592
box -53 -33 29 33
use nand3x1_pcell  nand3x1_pcell_2
timestamp 1647328266
transform 1 0 1628 0 1 0
box -84 0 1046 1575
use li1_M1_contact  li1_M1_contact_13
timestamp 1646004885
transform 1 0 2072 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1646004885
transform -1 0 1332 0 -1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_14
timestamp 1646004885
transform 1 0 1850 0 1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_15
timestamp 1646004885
transform -1 0 1110 0 -1 813
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_16
timestamp 1646004885
transform -1 0 1479 0 -1 592
box -53 -33 29 33
use nand3x1_pcell  nand3x1_pcell_1
timestamp 1647328266
transform 1 0 3256 0 1 0
box -84 0 1046 1575
use nand2x1_pcell  nand2x1_pcell_0
timestamp 1647328257
transform 1 0 2590 0 1 0
box -84 0 750 1575
use li1_M1_contact  li1_M1_contact_12
timestamp 1646004885
transform 1 0 3108 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_10
timestamp 1646004885
transform 1 0 2812 0 1 888
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_18
timestamp 1646004885
transform 1 0 2960 0 1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_17
timestamp 1646004885
transform -1 0 2442 0 -1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_8
timestamp 1646004885
transform -1 0 2294 0 -1 814
box -53 -33 29 33
use nand2x1_pcell  nand2x1_pcell_1
timestamp 1647328257
transform 1 0 4218 0 1 0
box -84 0 750 1575
use li1_M1_contact  li1_M1_contact_11
timestamp 1646004885
transform 1 0 3700 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_9
timestamp 1646004885
transform 1 0 3478 0 1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_6
timestamp 1646004885
transform -1 0 4070 0 -1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_4
timestamp 1646004885
transform -1 0 3922 0 -1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_19
timestamp 1646004885
transform 1 0 4440 0 1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_7
timestamp 1646004885
transform 1 0 4588 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_2
timestamp 1646004885
transform 1 0 4736 0 1 814
box -53 -33 29 33
<< labels >>
rlabel metal1 871 871 905 905 1 CLK
port 1 n
rlabel metal1 2277 797 2311 831 1 SN
port 2 n
rlabel metal1 4053 723 4087 757 1 Q
port 3 n
rlabel metal1 4719 797 4753 831 1 QN
port 4 n
rlabel metal1 205 797 239 831 1 D
port 5 n
rlabel metal1 55 1505 89 1539 1 VDD
port 6 n
rlabel metal1 55 13 89 47 1 VSS
port 7 n
<< end >>
