magic
tech sky130A
magscale 1 2
timestamp 1648740352
<< metal1 >>
rect 1867 797 2108 831
use votern3x1_pcell  votern3x1_pcell_0
timestamp 1648740297
transform 1 0 0 0 1 0
box -84 0 2082 1575
use invx1_pcell  invx1_pcell_0
timestamp 1648064504
transform 1 0 1998 0 1 0
box -84 0 528 1575
use li1_M1_contact  li1_M1_contact_16
timestamp 1648061256
transform -1 0 1850 0 -1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform 1 0 2146 0 1 814
box -53 -33 29 33
<< labels >>
rlabel space 2277 427 2311 979 1 Y
<< end >>
