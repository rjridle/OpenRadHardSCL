magic
tech sky130A
magscale 1 2
timestamp 1645915072
<< nmos >>
rect 161 215 191 276
tri 56 185 86 215 se
rect 86 185 191 215
rect 56 103 86 185
tri 86 169 102 185 nw
tri 145 169 161 185 ne
tri 86 103 90 107 sw
rect 56 91 90 103
tri 90 91 102 103 sw
tri 145 91 161 107 se
rect 161 91 191 185
tri 56 61 86 91 ne
rect 86 61 161 91
tri 161 61 191 91 nw
<< ndiff >>
rect 0 260 161 276
rect 0 226 10 260
rect 44 226 100 260
rect 134 226 161 260
rect 0 215 161 226
rect 191 260 248 276
rect 191 226 204 260
rect 238 226 248 260
rect 0 189 56 215
rect 0 155 10 189
rect 44 155 56 189
tri 56 185 86 215 nw
rect 0 121 56 155
rect 0 87 10 121
rect 44 87 56 121
tri 86 169 102 185 se
rect 102 169 145 185
tri 145 169 161 185 sw
rect 86 141 161 169
rect 86 107 107 141
rect 141 107 161 141
tri 86 103 90 107 ne
rect 90 103 145 107
tri 90 91 102 103 ne
rect 102 91 145 103
tri 145 91 161 107 nw
rect 0 61 56 87
tri 56 61 86 91 sw
tri 161 61 191 91 se
rect 191 61 248 226
rect 0 50 248 61
rect 0 16 10 50
rect 44 16 107 50
rect 141 16 204 50
rect 238 16 248 50
rect 0 0 248 16
<< ndiffc >>
rect 10 226 44 260
rect 100 226 134 260
rect 204 226 238 260
rect 10 155 44 189
rect 10 87 44 121
rect 107 107 141 141
rect 10 16 44 50
rect 107 16 141 50
rect 204 16 238 50
<< poly >>
rect 161 276 191 302
<< locali >>
rect 10 260 44 276
rect 204 260 238 276
rect 44 226 100 260
rect 134 226 204 260
rect 10 189 44 226
rect 204 210 238 226
rect 10 121 44 155
rect 107 141 141 143
rect 107 91 141 107
rect 10 50 44 87
rect 204 50 238 66
rect 44 16 107 50
rect 141 16 204 50
rect 10 0 44 16
rect 204 0 238 16
<< viali >>
rect 107 143 141 177
<< metal1 >>
rect 101 177 147 183
rect 95 143 107 177
rect 141 143 230 177
rect 101 137 147 143
<< end >>
