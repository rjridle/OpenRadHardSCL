magic
tech sky130A
magscale 1 2
timestamp 1645918728
<< nmos >>
rect 125 182 155 243
tri 20 152 50 182 se
rect 50 152 155 182
rect 20 58 50 152
tri 50 136 66 152 nw
tri 109 136 125 152 ne
tri 50 58 66 74 sw
tri 109 58 125 74 se
rect 125 58 155 152
tri 20 28 50 58 ne
rect 50 28 125 58
tri 125 28 155 58 nw
<< ndiff >>
rect -37 227 125 243
rect -37 193 -27 227
rect 7 193 70 227
rect 104 193 125 227
rect -37 182 125 193
rect 155 227 211 243
rect 155 193 167 227
rect 201 193 211 227
rect -37 28 20 182
tri 20 152 50 182 nw
rect 155 156 211 193
tri 50 136 66 152 se
rect 66 136 109 152
tri 109 136 125 152 sw
rect 50 108 125 136
rect 50 74 70 108
rect 104 74 125 108
tri 50 58 66 74 ne
rect 66 58 109 74
tri 109 58 125 74 nw
rect 155 122 167 156
rect 201 122 211 156
rect 155 88 211 122
tri 20 28 50 58 sw
tri 125 28 155 58 se
rect 155 54 167 88
rect 201 54 211 88
rect 155 28 211 54
rect -37 17 211 28
rect -37 -17 -27 17
rect 7 -17 70 17
rect 104 -17 167 17
rect 201 -17 211 17
rect -37 -33 211 -17
<< ndiffc >>
rect -27 193 7 227
rect 70 193 104 227
rect 167 193 201 227
rect 70 74 104 108
rect 167 122 201 156
rect 167 54 201 88
rect -27 -17 7 17
rect 70 -17 104 17
rect 167 -17 201 17
<< poly >>
rect 125 243 155 269
<< locali >>
rect -27 227 7 243
rect 167 227 201 243
rect 7 193 70 227
rect 104 193 167 227
rect -27 175 7 193
rect 167 156 201 193
rect 70 108 104 143
rect 70 58 104 74
rect 167 88 201 122
rect -27 17 7 35
rect 167 17 201 54
rect 7 -17 70 17
rect 104 -17 167 17
rect -27 -33 7 -17
rect 167 -33 201 -17
<< end >>
