* SPICE3 file created from TIELO.ext - technology: sky130A

.subckt TIELO YN VDD VSS
X0 a_121_411 a_121_411 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.1p ps=9.1u w=2u l=0.15u M=2
X1 YN a_121_411 VSS VSS sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=1.1408p ps=8.1u w=3u l=0.15u
.ends
