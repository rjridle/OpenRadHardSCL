magic
tech sky130
magscale 1 2
timestamp 1651259505
<< metal1 >>
rect 315 501 569 535
use invx1_pcell  invx1_pcell_1
timestamp 1651259471
transform 1 0 444 0 1 0
box -84 0 528 1575
use invx1_pcell  invx1_pcell_0
timestamp 1651259471
transform 1 0 0 0 1 0
box -84 0 528 1575
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform -1 0 296 0 -1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform 1 0 592 0 1 518
box -53 -33 29 33
<< end >>
