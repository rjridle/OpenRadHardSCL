* SPICE3 file created from TMRDFFSNRNQX1.ext - technology: sky130A

.subckt TMRDFFSNRNQX1 Q D CLK SN RN VDD GND
X0 GND a_6049_1050.t8 a_6825_103.t0 GND sky130_fd_pr__nfet_01v8 ad=4.9019p pd=4.107u as=0p ps=0u w=0u l=0u
X1 VDD.t176 RN.t1 a_15669_1050.t3 ��{�9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X2 GND a_4125_1050.t7 a_4901_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X3 a_599_989.t6 CLK.t0 VDD.t69 ��h�9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X4 VDD.t174 RN.t2 a_9897_1050.t4  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X5 VDD.t46 CLK.t1 a_1561_989.t6 VDD.t45 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X6 a_11821_1050.t4 a_12143_989.t7 VDD.t102 �+�إ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X7 VDD.t235 a_13105_989.t7 a_13745_1050.t6 ��ў9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X8 VDD.t188 a_277_1050.t7 a_2201_1050.t3  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X9 a_7333_989.t6 CLK.t2 VDD.t67 VDD.t66 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X10 a_10219_989.t1 SN.t0 VDD.t93 �+�إ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X11 VDD.t104 a_7333_989.t7 a_6371_989.t3 �WȞ9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X12 VDD.t24 CLK.t3 a_12143_989.t3  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X13 GND a_4447_989.t8 a_18760_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X14 GND a_15991_989.t9 a_18094_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X15 a_13105_989.t3 RN.t4 VDD.t172 VDD.t171 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X16 GND D.t0 a_11635_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X17 VDD.t170 RN.t5 a_277_1050.t6 �+�إ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X18 a_6371_989.t4 a_6049_1050.t7 VDD.t221 �}ߝ9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X19 GND a_6049_1050.t9 a_7787_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X20 VDD.t128 a_7973_1050.t7 a_7333_989.t1 ��˞9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X21 VDD.t215 a_9897_1050.t7 a_10219_989.t6 `�i�9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X22 a_17533_1051.t5 a_15991_989.t8 VDD.t44 �eh�9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X23 a_12143_989.t2 CLK.t7 VDD.t65  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X24 GND a_6371_989.t9 a_9711_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X25 a_599_989.t3 a_1561_989.t7 VDD.t73 VDD.t72 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X26 a_15991_989.t3 a_15669_1050.t7 VDD.t140 �+�إ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X27 GND D.t1 a_5863_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X28 VDD.t168 RN.t6 a_1561_989.t4 P��9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X29 a_9897_1050.t2 a_6371_989.t7 VDD.t79 P��9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X30 a_4125_1050.t3 a_599_989.t8 VDD.t48 ��b�9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X31 VDD.t108 SN.t2 a_2201_1050.t1 @{�9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X32 a_4125_1050.t1 a_4447_989.t7 VDD.t110 0�ǝ9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X33 VDD.t184 a_6371_989.t8 a_6049_1050.t4  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X34 a_18197_1051.t5 a_15991_989.t10 a_17533_1051.t2 VDD.t94 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X35 a_1561_989.t5 CLK.t8 VDD.t180 �+�إ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X36 GND a_11821_1050.t8 a_12597_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X37 VDD.t199 a_599_989.t9 a_277_1050.t4 ����9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X38 a_13745_1050.t0 SN.t4 VDD.t1 ��x�9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X39 GND a_13745_1050.t8 a_14521_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X40 GND a_9897_1050.t8 a_10673_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X41 a_17533_1051.t7 a_10219_989.t7 VDD.t182 �+��9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X42 GND a_7973_1050.t9 a_8749_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X43 a_12143_989.t0 a_11821_1050.t7 VDD.t54 P�ԝ9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X44 VDD.t40 a_13745_1050.t7 a_13105_989.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X45 Q a_17708_209.t8 GND.t8 GND sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=0p ps=0u w=0u l=0u
X46 a_15991_989.t1 SN.t5 VDD.t209  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X47 a_15669_1050.t2 a_12143_989.t8 VDD.t75 VDD.t74 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X48 GND D.t4 a_91_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X49 a_4125_1050.t5 RN.t8 VDD.t166 �+�إ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X50 VDD.t11 a_17708_209.t7 Q.t1 �3h�9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X51 VDD.t194 a_1561_989.t8 a_2201_1050.t6 `b��9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X52 VDD.t164 RN.t9 a_6049_1050.t6  w��9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X53 a_7333_989.t0 a_7973_1050.t8 VDD.t112  �ɝ9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X54 a_7973_1050.t6 a_7333_989.t8 VDD.t38 �M��9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X55 a_9897_1050.t1 a_10219_989.t9 VDD.t42  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X56 VDD.t233 a_13105_989.t10 a_15991_989.t6 VDD.t232 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X57 a_1561_989.t1 a_2201_1050.t7 VDD.t30 �+�إ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X58 a_18197_1051.t1 a_4447_989.t9 a_17533_1051.t1 �F�9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X59 VDD.t126 a_4125_1050.t8 a_4447_989.t1 `h�9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X60 GND a_15991_989.t12 a_17428_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X61 a_6371_989.t6 CLK.t10 VDD.t32  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X62 VDD.t120 CLK.t11 a_7333_989.t5 0�l�9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X63 a_6049_1050.t0 D.t2 VDD.t132 ���9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X64 GND a_11821_1050.t10 a_13559_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X65 a_17708_209.t4 a_10219_989.t10 a_18197_1051.t7  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X66 GND a_12143_989.t9 a_15483_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X67 a_277_1050.t1 D.t3 VDD.t130 VDD.t129 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X68 VDD.t96 CLK.t12 a_13105_989.t2 �+�إ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X69 a_15991_989.t5 a_13105_989.t11 VDD.t231 ����9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X70 VDD.t203 a_11821_1050.t9 a_13745_1050.t3 ��i�9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X71 a_10219_989.t4 a_7333_989.t9 VDD.t56 ��9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X72 VDD.t229 a_13105_989.t12 a_12143_989.t6 @�9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X73 a_15669_1050.t4 RN.t10 VDD.t162 �b��9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X74 VDD.t5 a_277_1050.t8 a_599_989.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X75 a_9897_1050.t3 RN.t11 VDD.t160 VDD.t159 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X76 VDD.t158 RN.t13 a_11821_1050.t6 �+�إ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X77 VDD.t16 a_1561_989.t9 a_599_989.t2 ���9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X78 a_13745_1050.t5 a_13105_989.t13 VDD.t227 ���9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X79 VDD.t223 SN.t6 a_4447_989.t3  "��9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X80 a_18197_1051.t3 a_4447_989.t10 a_17708_209.t1 �䛝9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X81 VDD.t211 a_15991_989.t11 a_15669_1050.t6 ���9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X82 a_6371_989.t2 a_7333_989.t10 VDD.t50  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X83 GND a_15669_1050.t8 a_16445_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X84 VDD.t156 RN.t15 a_7333_989.t4 VDD.t155 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X85 VDD.t85 SN.t7 a_7973_1050.t3 �+�إ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X86 a_277_1050.t5 RN.t16 VDD.t152 ���9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X87 a_11821_1050.t5 RN.t17 VDD.t154 ��I�9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X88 VDD.t61 SN.t8 a_13745_1050.t1 �J�9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X89 a_10219_989.t5 a_9897_1050.t9 VDD.t34 �J�9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X90 VDD.t213 CLK.t14 a_599_989.t5 �AK�9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X91 VDD.t36 a_12143_989.t10 a_11821_1050.t3  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X92 a_1561_989.t3 RN.t18 VDD.t150 VDD.t149 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X93 VDD.t22 a_1561_989.t10 a_4447_989.t6 �+�إ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X94 a_2201_1050.t0 SN.t11 VDD.t26 ���9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X95 GND a_277_1050.t11 a_2015_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X96 VDD.t148 RN.t19 a_4125_1050.t4 �L�9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X97 a_12143_989.t5 a_13105_989.t14 VDD.t225 ��ϝ9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X98 a_599_989.t1 a_277_1050.t9 VDD.t7 ��ѝ9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X99 VDD.t98 a_6049_1050.t10 a_7973_1050.t1 P[��9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X100 VDD.t146 RN.t21 a_13105_989.t4  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X101 a_277_1050.t3 a_599_989.t11 VDD.t71 VDD.t70 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X102 a_11821_1050.t1 D.t5 VDD.t134 �+�إ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X103 a_13105_989.t6 a_13745_1050.t9 VDD.t207 @��9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X104 VDD.t138 a_15669_1050.t9 a_15991_989.t2 �Ӵ�9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X105 a_7973_1050.t0 a_6049_1050.t11 VDD.t118 @Q��9V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X106 VDD.t9 a_6371_989.t10 a_9897_1050.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X107 a_2201_1050.t2 a_277_1050.t10 VDD.t106 VDD.t105 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X108 VDD.t205 a_7333_989.t11 a_10219_989.t3  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X109 Q.t0 a_17708_209.t9 VDD.t28  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X110 a_2201_1050.t5 a_1561_989.t12 VDD.t100  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X111 VDD.t14 a_599_989.t12 a_4125_1050.t2  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X112 GND a_2201_1050.t8 a_2977_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X113 VDD.t190 a_4447_989.t13 a_4125_1050.t6  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X114 a_6049_1050.t5 RN.t23 VDD.t144  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X115 a_17533_1051.t3 a_15991_989.t13 a_18197_1051.t4  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X116 a_4447_989.t0 a_4125_1050.t9 VDD.t124  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X117 VDD.t52 a_6049_1050.t12 a_6371_989.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X118 GND a_277_1050.t12 a_1053_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X119 a_4447_989.t5 a_1561_989.t15 VDD.t192  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X120 a_15669_1050.t1 a_15991_989.t14 VDD.t20  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X121 VDD.t77 a_11821_1050.t11 a_12143_989.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X122 VDD.t91 a_10219_989.t11 a_17533_1051.t6  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X123 a_13105_989.t1 CLK.t16 VDD.t63  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X124 VDD.t219 SN.t13 a_15991_989.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X125 VDD.t59 SN.t14 a_10219_989.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X126 a_13745_1050.t2 a_11821_1050.t12 VDD.t18  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X127 VDD.t201 a_12143_989.t12 a_15669_1050.t5  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X128 GND a_599_989.t7 a_3939_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X129 a_6049_1050.t3 a_6371_989.t12 VDD.t88  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X130 VDD.t196 a_7333_989.t14 a_7973_1050.t5  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X131 VDD.t217 a_10219_989.t14 a_9897_1050.t6  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X132 VDD.t3 a_2201_1050.t9 a_1561_989.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X133 a_4447_989.t2 SN.t15 VDD.t81  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X134 a_17708_209.t0 a_4447_989.t14 a_18197_1051.t2  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X135 a_17533_1051.t0 a_4447_989.t15 a_18197_1051.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X136 VDD.t178 CLK.t17 a_6371_989.t5  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X137 a_7333_989.t3 RN.t25 VDD.t142  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X138 VDD.t136 D.t6 a_6049_1050.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X139 a_7973_1050.t2 SN.t16 VDD.t186  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X140 a_18197_1051.t6 a_10219_989.t15 a_17708_209.t3  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X141 VDD.t83 a_15991_989.t15 a_17533_1051.t4  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X142 VDD.t114 D.t7 a_277_1050.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X143 VDD.t116 D.t8 a_11821_1050.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
C0 VDD RN 2.65fF
C1 CLK VDD 8.69fF
C2 D RN 2.36fF
C3 SN VDD 1.76fF
C4 CLK D 12.06fF
C5 SN D 0.31fF
C6 CLK RN 1.11fF
C7 Q VDD 1.05fF
C8 SN RN 16.07fF
C9 CLK SN 0.63fF
C10 VDD D 11.48fF
R0 RN.n23 RN.t5 479.223
R1 RN.n17 RN.t19 479.223
R2 RN.n14 RN.t9 479.223
R3 RN.n8 RN.t2 479.223
R4 RN.n5 RN.t13 479.223
R5 RN.n0 RN.t1 479.223
R6 RN.n20 RN.t18 454.685
R7 RN.n11 RN.t25 454.685
R8 RN.n2 RN.t4 454.685
R9 RN.n20 RN.t6 428.979
R10 RN.n11 RN.t15 428.979
R11 RN.n2 RN.t21 428.979
R12 RN.n23 RN.t16 375.52
R13 RN.n17 RN.t8 375.52
R14 RN.n14 RN.t23 375.52
R15 RN.n8 RN.t11 375.52
R16 RN.n5 RN.t17 375.52
R17 RN.n0 RN.t10 375.52
R18 RN.n21 RN.n20 254.865
R19 RN.n12 RN.n11 254.865
R20 RN.n3 RN.n2 254.865
R21 RN.n24 RN.n23 252.188
R22 RN.n18 RN.n17 252.188
R23 RN.n15 RN.n14 252.188
R24 RN.n9 RN.n8 252.188
R25 RN.n6 RN.n5 252.188
R26 RN.n1 RN.n0 252.188
R27 RN.n24 RN.t20 231.854
R28 RN.n18 RN.t26 231.854
R29 RN.n15 RN.t7 231.854
R30 RN.n9 RN.t14 231.854
R31 RN.n6 RN.t12 231.854
R32 RN.n1 RN.t22 231.854
R33 RN.n21 RN.t24 228.106
R34 RN.n12 RN.t3 228.106
R35 RN.n3 RN.t0 228.106
R36 RN.n7 RN.n4 11.381
R37 RN.n16 RN.n13 11.381
R38 RN.n25 RN.n22 11.381
R39 RN.n4 RN.n1 7.325
R40 RN.n10 RN.n7 7.028
R41 RN.n19 RN.n16 7.028
R42 RN.n4 RN.n3 4.65
R43 RN.n7 RN.n6 4.65
R44 RN.n10 RN.n9 4.65
R45 RN.n13 RN.n12 4.65
R46 RN.n16 RN.n15 4.65
R47 RN.n19 RN.n18 4.65
R48 RN.n22 RN.n21 4.65
R49 RN.n25 RN.n24 4.65
R50 RN.n13 RN.n10 2.675
R51 RN.n22 RN.n19 2.675
R52 RN.n25 RN 0.046
R53 a_14802_210.n10 a_14802_210.n7 185.173
R54 a_14802_210.n1 a_14802_210.n0 102.58
R55 a_14802_210.t0 a_14802_210.n12 83.571
R56 a_14802_210.t0 a_14802_210.n10 75.765
R57 a_14802_210.n3 a_14802_210.n2 65.02
R58 a_14802_210.t0 a_14802_210.n3 58.043
R59 a_14802_210.n12 a_14802_210.n11 55.714
R60 a_14802_210.n3 a_14802_210.n1 35.865
R61 a_14802_210.n7 a_14802_210.n6 22.349
R62 a_14802_210.n9 a_14802_210.n8 19.952
R63 a_14802_210.n7 a_14802_210.n5 8.443
R64 a_14802_210.t0 a_14802_210.n4 8.137
R65 a_14802_210.n10 a_14802_210.n9 1.505
R66 a_13105_989.n7 a_13105_989.t13 454.685
R67 a_13105_989.n9 a_13105_989.t14 454.685
R68 a_13105_989.n5 a_13105_989.t11 454.685
R69 a_13105_989.n7 a_13105_989.t7 428.979
R70 a_13105_989.n9 a_13105_989.t12 428.979
R71 a_13105_989.n5 a_13105_989.t10 428.979
R72 a_13105_989.n15 a_13105_989.n13 342.597
R73 a_13105_989.n8 a_13105_989.t8 339.542
R74 a_13105_989.n6 a_13105_989.t9 339.542
R75 a_13105_989.n10 a_13105_989.t15 339.186
R76 a_13105_989.n3 a_13105_989.n2 161.352
R77 a_13105_989.n13 a_13105_989.n4 151.34
R78 a_13105_989.n8 a_13105_989.n7 143.429
R79 a_13105_989.n6 a_13105_989.n5 143.429
R80 a_13105_989.n10 a_13105_989.n9 143.074
R81 a_13105_989.n4 a_13105_989.n0 95.095
R82 a_13105_989.n3 a_13105_989.n1 95.095
R83 a_13105_989.n4 a_13105_989.n3 66.258
R84 a_13105_989.n15 a_13105_989.n14 15.218
R85 a_13105_989.n0 a_13105_989.t4 14.282
R86 a_13105_989.n0 a_13105_989.t3 14.282
R87 a_13105_989.n1 a_13105_989.t2 14.282
R88 a_13105_989.n1 a_13105_989.t1 14.282
R89 a_13105_989.n2 a_13105_989.t0 14.282
R90 a_13105_989.n2 a_13105_989.t6 14.282
R91 a_13105_989.n16 a_13105_989.n15 12.014
R92 a_13105_989.n12 a_13105_989.n6 11.134
R93 a_13105_989.n11 a_13105_989.n10 8.145
R94 a_13105_989.n11 a_13105_989.n8 4.65
R95 a_13105_989.n13 a_13105_989.n12 4.65
R96 a_13105_989.n12 a_13105_989.n11 4.035
R97 GND.n32 GND.n31 237.558
R98 GND.n64 GND.n63 237.558
R99 GND.n498 GND.n497 237.558
R100 GND.n540 GND.n539 237.558
R101 GND.n582 GND.n581 237.558
R102 GND.n626 GND.n625 237.558
R103 GND.n670 GND.n669 237.558
R104 GND.n715 GND.n714 237.558
R105 GND.n760 GND.n759 237.558
R106 GND.n805 GND.n804 237.558
R107 GND.n847 GND.n846 237.558
R108 GND.n432 GND.n431 237.558
R109 GND.n889 GND.n888 237.558
R110 GND.n388 GND.n387 237.558
R111 GND.n344 GND.n343 237.558
R112 GND.n302 GND.n301 237.558
R113 GND.n258 GND.n257 237.558
R114 GND.n216 GND.n215 237.558
R115 GND.n172 GND.n171 237.558
R116 GND.n128 GND.n127 237.558
R117 GND.n96 GND.n95 237.558
R118 GND.n29 GND.n28 210.82
R119 GND.n61 GND.n60 210.82
R120 GND.n93 GND.n92 210.82
R121 GND.n500 GND.n499 210.82
R122 GND.n542 GND.n541 210.82
R123 GND.n584 GND.n583 210.82
R124 GND.n628 GND.n627 210.82
R125 GND.n672 GND.n671 210.82
R126 GND.n717 GND.n716 210.82
R127 GND.n762 GND.n761 210.82
R128 GND.n807 GND.n806 210.82
R129 GND.n849 GND.n848 210.82
R130 GND.n891 GND.n890 210.82
R131 GND.n429 GND.n428 210.82
R132 GND.n385 GND.n384 210.82
R133 GND.n341 GND.n340 210.82
R134 GND.n299 GND.n298 210.82
R135 GND.n255 GND.n254 210.82
R136 GND.n213 GND.n212 210.82
R137 GND.n169 GND.n168 210.82
R138 GND.n125 GND.n124 210.82
R139 GND.n245 GND.n244 173.365
R140 GND.n331 GND.n330 173.365
R141 GND.n900 GND.n899 173.365
R142 GND.n858 GND.n857 173.365
R143 GND.n816 GND.n815 173.365
R144 GND.n551 GND.n550 173.365
R145 GND.n509 GND.n508 173.365
R146 GND.n467 GND.n466 173.365
R147 GND.n159 GND.n158 167.358
R148 GND.n203 GND.n202 167.358
R149 GND.n289 GND.n288 167.358
R150 GND.n375 GND.n374 167.358
R151 GND.n419 GND.n418 167.358
R152 GND.n639 GND.n638 167.358
R153 GND.n595 GND.n594 167.358
R154 GND.n82 GND.n81 166.605
R155 GND.n114 GND.n113 166.605
R156 GND.n50 GND.n49 166.605
R157 GND.n774 GND.n773 152.358
R158 GND.n729 GND.n728 152.358
R159 GND.n684 GND.n683 152.358
R160 GND.n20 GND.n19 37.582
R161 GND.t8 GND.n17 32.601
R162 GND.n773 GND.n772 28.421
R163 GND.n728 GND.n727 28.421
R164 GND.n683 GND.n682 28.421
R165 GND.n773 GND.n771 25.263
R166 GND.n728 GND.n726 25.263
R167 GND.n683 GND.n681 25.263
R168 GND.n771 GND.n770 24.383
R169 GND.n726 GND.n725 24.383
R170 GND.n681 GND.n680 24.383
R171 GND.n81 GND.n79 23.03
R172 GND.n113 GND.n111 23.03
R173 GND.n158 GND.n156 23.03
R174 GND.n202 GND.n200 23.03
R175 GND.n288 GND.n286 23.03
R176 GND.n374 GND.n372 23.03
R177 GND.n418 GND.n416 23.03
R178 GND.n638 GND.n636 23.03
R179 GND.n594 GND.n592 23.03
R180 GND.n49 GND.n47 23.03
R181 GND.n17 GND.n16 21.734
R182 GND.n4 GND.n3 20.705
R183 GND.n10 GND.n9 20.705
R184 GND.n21 GND.n20 20.705
R185 GND.n3 GND.n2 19.952
R186 GND.n30 GND.n29 18.953
R187 GND.n62 GND.n61 18.953
R188 GND.n94 GND.n93 18.953
R189 GND.n501 GND.n500 18.953
R190 GND.n543 GND.n542 18.953
R191 GND.n585 GND.n584 18.953
R192 GND.n629 GND.n628 18.953
R193 GND.n673 GND.n672 18.953
R194 GND.n718 GND.n717 18.953
R195 GND.n763 GND.n762 18.953
R196 GND.n808 GND.n807 18.953
R197 GND.n850 GND.n849 18.953
R198 GND.n892 GND.n891 18.953
R199 GND.n430 GND.n429 18.953
R200 GND.n386 GND.n385 18.953
R201 GND.n342 GND.n341 18.953
R202 GND.n300 GND.n299 18.953
R203 GND.n256 GND.n255 18.953
R204 GND.n214 GND.n213 18.953
R205 GND.n170 GND.n169 18.953
R206 GND.n126 GND.n125 18.953
R207 GND.n19 GND.t8 15.644
R208 GND.n33 GND.n30 14.864
R209 GND.n65 GND.n62 14.864
R210 GND.n97 GND.n94 14.864
R211 GND.n129 GND.n126 14.864
R212 GND.n173 GND.n170 14.864
R213 GND.n217 GND.n214 14.864
R214 GND.n259 GND.n256 14.864
R215 GND.n303 GND.n300 14.864
R216 GND.n345 GND.n342 14.864
R217 GND.n389 GND.n386 14.864
R218 GND.n433 GND.n430 14.864
R219 GND.n893 GND.n892 14.864
R220 GND.n851 GND.n850 14.864
R221 GND.n809 GND.n808 14.864
R222 GND.n764 GND.n763 14.864
R223 GND.n719 GND.n718 14.864
R224 GND.n674 GND.n673 14.864
R225 GND.n630 GND.n629 14.864
R226 GND.n586 GND.n585 14.864
R227 GND.n544 GND.n543 14.864
R228 GND.n502 GND.n501 14.864
R229 GND.n19 GND.n18 13.541
R230 GND.n463 GND.n462 9.154
R231 GND.n468 GND.n465 9.154
R232 GND.n471 GND.n470 9.154
R233 GND.n474 GND.n473 9.154
R234 GND.n477 GND.n476 9.154
R235 GND.n480 GND.n479 9.154
R236 GND.n483 GND.n482 9.154
R237 GND.n486 GND.n485 9.154
R238 GND.n489 GND.n488 9.154
R239 GND.n492 GND.n491 9.154
R240 GND.n495 GND.n494 9.154
R241 GND.n502 GND.n498 9.154
R242 GND.n505 GND.n504 9.154
R243 GND.n510 GND.n507 9.154
R244 GND.n513 GND.n512 9.154
R245 GND.n516 GND.n515 9.154
R246 GND.n519 GND.n518 9.154
R247 GND.n522 GND.n521 9.154
R248 GND.n525 GND.n524 9.154
R249 GND.n528 GND.n527 9.154
R250 GND.n531 GND.n530 9.154
R251 GND.n534 GND.n533 9.154
R252 GND.n537 GND.n536 9.154
R253 GND.n544 GND.n540 9.154
R254 GND.n547 GND.n546 9.154
R255 GND.n552 GND.n549 9.154
R256 GND.n555 GND.n554 9.154
R257 GND.n558 GND.n557 9.154
R258 GND.n561 GND.n560 9.154
R259 GND.n564 GND.n563 9.154
R260 GND.n567 GND.n566 9.154
R261 GND.n570 GND.n569 9.154
R262 GND.n573 GND.n572 9.154
R263 GND.n576 GND.n575 9.154
R264 GND.n579 GND.n578 9.154
R265 GND.n586 GND.n582 9.154
R266 GND.n589 GND.n588 9.154
R267 GND.n596 GND.n591 9.154
R268 GND.n599 GND.n598 9.154
R269 GND.n602 GND.n601 9.154
R270 GND.n605 GND.n604 9.154
R271 GND.n608 GND.n607 9.154
R272 GND.n611 GND.n610 9.154
R273 GND.n614 GND.n613 9.154
R274 GND.n617 GND.n616 9.154
R275 GND.n620 GND.n619 9.154
R276 GND.n623 GND.n622 9.154
R277 GND.n630 GND.n626 9.154
R278 GND.n633 GND.n632 9.154
R279 GND.n640 GND.n635 9.154
R280 GND.n643 GND.n642 9.154
R281 GND.n646 GND.n645 9.154
R282 GND.n649 GND.n648 9.154
R283 GND.n652 GND.n651 9.154
R284 GND.n655 GND.n654 9.154
R285 GND.n658 GND.n657 9.154
R286 GND.n661 GND.n660 9.154
R287 GND.n664 GND.n663 9.154
R288 GND.n667 GND.n666 9.154
R289 GND.n674 GND.n670 9.154
R290 GND.n677 GND.n676 9.154
R291 GND.n685 GND.n679 9.154
R292 GND.n688 GND.n687 9.154
R293 GND.n691 GND.n690 9.154
R294 GND.n694 GND.n693 9.154
R295 GND.n697 GND.n696 9.154
R296 GND.n700 GND.n699 9.154
R297 GND.n703 GND.n702 9.154
R298 GND.n706 GND.n705 9.154
R299 GND.n709 GND.n708 9.154
R300 GND.n712 GND.n711 9.154
R301 GND.n719 GND.n715 9.154
R302 GND.n722 GND.n721 9.154
R303 GND.n730 GND.n724 9.154
R304 GND.n733 GND.n732 9.154
R305 GND.n736 GND.n735 9.154
R306 GND.n739 GND.n738 9.154
R307 GND.n742 GND.n741 9.154
R308 GND.n745 GND.n744 9.154
R309 GND.n748 GND.n747 9.154
R310 GND.n751 GND.n750 9.154
R311 GND.n754 GND.n753 9.154
R312 GND.n757 GND.n756 9.154
R313 GND.n764 GND.n760 9.154
R314 GND.n767 GND.n766 9.154
R315 GND.n775 GND.n769 9.154
R316 GND.n778 GND.n777 9.154
R317 GND.n781 GND.n780 9.154
R318 GND.n784 GND.n783 9.154
R319 GND.n787 GND.n786 9.154
R320 GND.n790 GND.n789 9.154
R321 GND.n793 GND.n792 9.154
R322 GND.n796 GND.n795 9.154
R323 GND.n799 GND.n798 9.154
R324 GND.n802 GND.n801 9.154
R325 GND.n809 GND.n805 9.154
R326 GND.n812 GND.n811 9.154
R327 GND.n817 GND.n814 9.154
R328 GND.n820 GND.n819 9.154
R329 GND.n823 GND.n822 9.154
R330 GND.n826 GND.n825 9.154
R331 GND.n829 GND.n828 9.154
R332 GND.n832 GND.n831 9.154
R333 GND.n835 GND.n834 9.154
R334 GND.n838 GND.n837 9.154
R335 GND.n841 GND.n840 9.154
R336 GND.n844 GND.n843 9.154
R337 GND.n851 GND.n847 9.154
R338 GND.n854 GND.n853 9.154
R339 GND.n859 GND.n856 9.154
R340 GND.n862 GND.n861 9.154
R341 GND.n865 GND.n864 9.154
R342 GND.n868 GND.n867 9.154
R343 GND.n871 GND.n870 9.154
R344 GND.n874 GND.n873 9.154
R345 GND.n877 GND.n876 9.154
R346 GND.n880 GND.n879 9.154
R347 GND.n883 GND.n882 9.154
R348 GND.n886 GND.n885 9.154
R349 GND.n893 GND.n889 9.154
R350 GND.n896 GND.n895 9.154
R351 GND.n901 GND.n898 9.154
R352 GND.n457 GND.n456 9.154
R353 GND.n454 GND.n453 9.154
R354 GND.n451 GND.n450 9.154
R355 GND.n448 GND.n447 9.154
R356 GND.n445 GND.n444 9.154
R357 GND.n442 GND.n441 9.154
R358 GND.n439 GND.n438 9.154
R359 GND.n436 GND.n435 9.154
R360 GND.n433 GND.n432 9.154
R361 GND.n426 GND.n425 9.154
R362 GND.n423 GND.n422 9.154
R363 GND.n420 GND.n415 9.154
R364 GND.n413 GND.n412 9.154
R365 GND.n410 GND.n409 9.154
R366 GND.n407 GND.n406 9.154
R367 GND.n404 GND.n403 9.154
R368 GND.n401 GND.n400 9.154
R369 GND.n398 GND.n397 9.154
R370 GND.n395 GND.n394 9.154
R371 GND.n392 GND.n391 9.154
R372 GND.n389 GND.n388 9.154
R373 GND.n382 GND.n381 9.154
R374 GND.n379 GND.n378 9.154
R375 GND.n376 GND.n371 9.154
R376 GND.n369 GND.n368 9.154
R377 GND.n366 GND.n365 9.154
R378 GND.n363 GND.n362 9.154
R379 GND.n360 GND.n359 9.154
R380 GND.n357 GND.n356 9.154
R381 GND.n354 GND.n353 9.154
R382 GND.n351 GND.n350 9.154
R383 GND.n348 GND.n347 9.154
R384 GND.n345 GND.n344 9.154
R385 GND.n338 GND.n337 9.154
R386 GND.n335 GND.n334 9.154
R387 GND.n332 GND.n329 9.154
R388 GND.n327 GND.n326 9.154
R389 GND.n324 GND.n323 9.154
R390 GND.n321 GND.n320 9.154
R391 GND.n318 GND.n317 9.154
R392 GND.n315 GND.n314 9.154
R393 GND.n312 GND.n311 9.154
R394 GND.n309 GND.n308 9.154
R395 GND.n306 GND.n305 9.154
R396 GND.n303 GND.n302 9.154
R397 GND.n296 GND.n295 9.154
R398 GND.n293 GND.n292 9.154
R399 GND.n290 GND.n285 9.154
R400 GND.n283 GND.n282 9.154
R401 GND.n280 GND.n279 9.154
R402 GND.n277 GND.n276 9.154
R403 GND.n274 GND.n273 9.154
R404 GND.n271 GND.n270 9.154
R405 GND.n268 GND.n267 9.154
R406 GND.n265 GND.n264 9.154
R407 GND.n262 GND.n261 9.154
R408 GND.n259 GND.n258 9.154
R409 GND.n252 GND.n251 9.154
R410 GND.n249 GND.n248 9.154
R411 GND.n246 GND.n243 9.154
R412 GND.n241 GND.n240 9.154
R413 GND.n238 GND.n237 9.154
R414 GND.n235 GND.n234 9.154
R415 GND.n232 GND.n231 9.154
R416 GND.n229 GND.n228 9.154
R417 GND.n226 GND.n225 9.154
R418 GND.n223 GND.n222 9.154
R419 GND.n220 GND.n219 9.154
R420 GND.n217 GND.n216 9.154
R421 GND.n210 GND.n209 9.154
R422 GND.n207 GND.n206 9.154
R423 GND.n204 GND.n199 9.154
R424 GND.n197 GND.n196 9.154
R425 GND.n194 GND.n193 9.154
R426 GND.n191 GND.n190 9.154
R427 GND.n188 GND.n187 9.154
R428 GND.n185 GND.n184 9.154
R429 GND.n182 GND.n181 9.154
R430 GND.n179 GND.n178 9.154
R431 GND.n176 GND.n175 9.154
R432 GND.n173 GND.n172 9.154
R433 GND.n166 GND.n165 9.154
R434 GND.n163 GND.n162 9.154
R435 GND.n160 GND.n155 9.154
R436 GND.n153 GND.n152 9.154
R437 GND.n150 GND.n149 9.154
R438 GND.n147 GND.n146 9.154
R439 GND.n144 GND.n143 9.154
R440 GND.n141 GND.n140 9.154
R441 GND.n138 GND.n137 9.154
R442 GND.n135 GND.n134 9.154
R443 GND.n132 GND.n131 9.154
R444 GND.n129 GND.n128 9.154
R445 GND.n122 GND.n121 9.154
R446 GND.n119 GND.n118 9.154
R447 GND.n116 GND.n115 9.154
R448 GND.n109 GND.n108 9.154
R449 GND.n106 GND.n105 9.154
R450 GND.n103 GND.n102 9.154
R451 GND.n100 GND.n99 9.154
R452 GND.n97 GND.n96 9.154
R453 GND.n90 GND.n89 9.154
R454 GND.n87 GND.n86 9.154
R455 GND.n84 GND.n83 9.154
R456 GND.n77 GND.n76 9.154
R457 GND.n74 GND.n73 9.154
R458 GND.n6 GND.n5 9.154
R459 GND.n12 GND.n11 9.154
R460 GND.n23 GND.n22 9.154
R461 GND.n26 GND.n25 9.154
R462 GND.n33 GND.n32 9.154
R463 GND.n36 GND.n35 9.154
R464 GND.n39 GND.n38 9.154
R465 GND.n42 GND.n41 9.154
R466 GND.n45 GND.n44 9.154
R467 GND.n52 GND.n51 9.154
R468 GND.n55 GND.n54 9.154
R469 GND.n58 GND.n57 9.154
R470 GND.n65 GND.n64 9.154
R471 GND.n68 GND.n67 9.154
R472 GND.n71 GND.n70 9.154
R473 GND.n81 GND.n80 8.128
R474 GND.n113 GND.n112 8.128
R475 GND.n158 GND.n157 8.128
R476 GND.n202 GND.n201 8.128
R477 GND.n288 GND.n287 8.128
R478 GND.n374 GND.n373 8.128
R479 GND.n418 GND.n417 8.128
R480 GND.n638 GND.n637 8.128
R481 GND.n594 GND.n593 8.128
R482 GND.n49 GND.n48 8.128
R483 GND.n7 GND.n1 4.795
R484 GND.n461 GND.n460 4.65
R485 GND.n75 GND.n74 4.65
R486 GND.n78 GND.n77 4.65
R487 GND.n85 GND.n84 4.65
R488 GND.n88 GND.n87 4.65
R489 GND.n91 GND.n90 4.65
R490 GND.n98 GND.n97 4.65
R491 GND.n101 GND.n100 4.65
R492 GND.n104 GND.n103 4.65
R493 GND.n107 GND.n106 4.65
R494 GND.n110 GND.n109 4.65
R495 GND.n117 GND.n116 4.65
R496 GND.n120 GND.n119 4.65
R497 GND.n123 GND.n122 4.65
R498 GND.n130 GND.n129 4.65
R499 GND.n133 GND.n132 4.65
R500 GND.n136 GND.n135 4.65
R501 GND.n139 GND.n138 4.65
R502 GND.n142 GND.n141 4.65
R503 GND.n145 GND.n144 4.65
R504 GND.n148 GND.n147 4.65
R505 GND.n151 GND.n150 4.65
R506 GND.n154 GND.n153 4.65
R507 GND.n161 GND.n160 4.65
R508 GND.n164 GND.n163 4.65
R509 GND.n167 GND.n166 4.65
R510 GND.n174 GND.n173 4.65
R511 GND.n177 GND.n176 4.65
R512 GND.n180 GND.n179 4.65
R513 GND.n183 GND.n182 4.65
R514 GND.n186 GND.n185 4.65
R515 GND.n189 GND.n188 4.65
R516 GND.n192 GND.n191 4.65
R517 GND.n195 GND.n194 4.65
R518 GND.n198 GND.n197 4.65
R519 GND.n205 GND.n204 4.65
R520 GND.n208 GND.n207 4.65
R521 GND.n211 GND.n210 4.65
R522 GND.n218 GND.n217 4.65
R523 GND.n221 GND.n220 4.65
R524 GND.n224 GND.n223 4.65
R525 GND.n227 GND.n226 4.65
R526 GND.n230 GND.n229 4.65
R527 GND.n233 GND.n232 4.65
R528 GND.n236 GND.n235 4.65
R529 GND.n239 GND.n238 4.65
R530 GND.n242 GND.n241 4.65
R531 GND.n247 GND.n246 4.65
R532 GND.n250 GND.n249 4.65
R533 GND.n253 GND.n252 4.65
R534 GND.n260 GND.n259 4.65
R535 GND.n263 GND.n262 4.65
R536 GND.n266 GND.n265 4.65
R537 GND.n269 GND.n268 4.65
R538 GND.n272 GND.n271 4.65
R539 GND.n275 GND.n274 4.65
R540 GND.n278 GND.n277 4.65
R541 GND.n281 GND.n280 4.65
R542 GND.n284 GND.n283 4.65
R543 GND.n291 GND.n290 4.65
R544 GND.n294 GND.n293 4.65
R545 GND.n297 GND.n296 4.65
R546 GND.n304 GND.n303 4.65
R547 GND.n307 GND.n306 4.65
R548 GND.n310 GND.n309 4.65
R549 GND.n313 GND.n312 4.65
R550 GND.n316 GND.n315 4.65
R551 GND.n319 GND.n318 4.65
R552 GND.n322 GND.n321 4.65
R553 GND.n325 GND.n324 4.65
R554 GND.n328 GND.n327 4.65
R555 GND.n333 GND.n332 4.65
R556 GND.n336 GND.n335 4.65
R557 GND.n339 GND.n338 4.65
R558 GND.n346 GND.n345 4.65
R559 GND.n349 GND.n348 4.65
R560 GND.n352 GND.n351 4.65
R561 GND.n355 GND.n354 4.65
R562 GND.n358 GND.n357 4.65
R563 GND.n361 GND.n360 4.65
R564 GND.n364 GND.n363 4.65
R565 GND.n367 GND.n366 4.65
R566 GND.n370 GND.n369 4.65
R567 GND.n377 GND.n376 4.65
R568 GND.n380 GND.n379 4.65
R569 GND.n383 GND.n382 4.65
R570 GND.n390 GND.n389 4.65
R571 GND.n393 GND.n392 4.65
R572 GND.n396 GND.n395 4.65
R573 GND.n399 GND.n398 4.65
R574 GND.n402 GND.n401 4.65
R575 GND.n405 GND.n404 4.65
R576 GND.n408 GND.n407 4.65
R577 GND.n411 GND.n410 4.65
R578 GND.n414 GND.n413 4.65
R579 GND.n421 GND.n420 4.65
R580 GND.n424 GND.n423 4.65
R581 GND.n427 GND.n426 4.65
R582 GND.n434 GND.n433 4.65
R583 GND.n437 GND.n436 4.65
R584 GND.n440 GND.n439 4.65
R585 GND.n443 GND.n442 4.65
R586 GND.n446 GND.n445 4.65
R587 GND.n449 GND.n448 4.65
R588 GND.n452 GND.n451 4.65
R589 GND.n455 GND.n454 4.65
R590 GND.n458 GND.n457 4.65
R591 GND.n902 GND.n901 4.65
R592 GND.n897 GND.n896 4.65
R593 GND.n894 GND.n893 4.65
R594 GND.n887 GND.n886 4.65
R595 GND.n884 GND.n883 4.65
R596 GND.n881 GND.n880 4.65
R597 GND.n878 GND.n877 4.65
R598 GND.n875 GND.n874 4.65
R599 GND.n872 GND.n871 4.65
R600 GND.n869 GND.n868 4.65
R601 GND.n866 GND.n865 4.65
R602 GND.n863 GND.n862 4.65
R603 GND.n860 GND.n859 4.65
R604 GND.n855 GND.n854 4.65
R605 GND.n852 GND.n851 4.65
R606 GND.n845 GND.n844 4.65
R607 GND.n842 GND.n841 4.65
R608 GND.n839 GND.n838 4.65
R609 GND.n836 GND.n835 4.65
R610 GND.n833 GND.n832 4.65
R611 GND.n830 GND.n829 4.65
R612 GND.n827 GND.n826 4.65
R613 GND.n824 GND.n823 4.65
R614 GND.n821 GND.n820 4.65
R615 GND.n818 GND.n817 4.65
R616 GND.n813 GND.n812 4.65
R617 GND.n810 GND.n809 4.65
R618 GND.n803 GND.n802 4.65
R619 GND.n800 GND.n799 4.65
R620 GND.n797 GND.n796 4.65
R621 GND.n794 GND.n793 4.65
R622 GND.n791 GND.n790 4.65
R623 GND.n788 GND.n787 4.65
R624 GND.n785 GND.n784 4.65
R625 GND.n782 GND.n781 4.65
R626 GND.n779 GND.n778 4.65
R627 GND.n776 GND.n775 4.65
R628 GND.n768 GND.n767 4.65
R629 GND.n765 GND.n764 4.65
R630 GND.n758 GND.n757 4.65
R631 GND.n755 GND.n754 4.65
R632 GND.n752 GND.n751 4.65
R633 GND.n749 GND.n748 4.65
R634 GND.n746 GND.n745 4.65
R635 GND.n743 GND.n742 4.65
R636 GND.n740 GND.n739 4.65
R637 GND.n737 GND.n736 4.65
R638 GND.n734 GND.n733 4.65
R639 GND.n731 GND.n730 4.65
R640 GND.n723 GND.n722 4.65
R641 GND.n720 GND.n719 4.65
R642 GND.n713 GND.n712 4.65
R643 GND.n710 GND.n709 4.65
R644 GND.n707 GND.n706 4.65
R645 GND.n704 GND.n703 4.65
R646 GND.n701 GND.n700 4.65
R647 GND.n698 GND.n697 4.65
R648 GND.n695 GND.n694 4.65
R649 GND.n692 GND.n691 4.65
R650 GND.n689 GND.n688 4.65
R651 GND.n686 GND.n685 4.65
R652 GND.n678 GND.n677 4.65
R653 GND.n675 GND.n674 4.65
R654 GND.n668 GND.n667 4.65
R655 GND.n665 GND.n664 4.65
R656 GND.n662 GND.n661 4.65
R657 GND.n659 GND.n658 4.65
R658 GND.n656 GND.n655 4.65
R659 GND.n653 GND.n652 4.65
R660 GND.n650 GND.n649 4.65
R661 GND.n647 GND.n646 4.65
R662 GND.n644 GND.n643 4.65
R663 GND.n641 GND.n640 4.65
R664 GND.n634 GND.n633 4.65
R665 GND.n631 GND.n630 4.65
R666 GND.n624 GND.n623 4.65
R667 GND.n621 GND.n620 4.65
R668 GND.n618 GND.n617 4.65
R669 GND.n615 GND.n614 4.65
R670 GND.n612 GND.n611 4.65
R671 GND.n609 GND.n608 4.65
R672 GND.n606 GND.n605 4.65
R673 GND.n603 GND.n602 4.65
R674 GND.n600 GND.n599 4.65
R675 GND.n597 GND.n596 4.65
R676 GND.n590 GND.n589 4.65
R677 GND.n587 GND.n586 4.65
R678 GND.n580 GND.n579 4.65
R679 GND.n577 GND.n576 4.65
R680 GND.n574 GND.n573 4.65
R681 GND.n571 GND.n570 4.65
R682 GND.n568 GND.n567 4.65
R683 GND.n565 GND.n564 4.65
R684 GND.n562 GND.n561 4.65
R685 GND.n559 GND.n558 4.65
R686 GND.n556 GND.n555 4.65
R687 GND.n553 GND.n552 4.65
R688 GND.n548 GND.n547 4.65
R689 GND.n545 GND.n544 4.65
R690 GND.n538 GND.n537 4.65
R691 GND.n535 GND.n534 4.65
R692 GND.n532 GND.n531 4.65
R693 GND.n529 GND.n528 4.65
R694 GND.n526 GND.n525 4.65
R695 GND.n523 GND.n522 4.65
R696 GND.n520 GND.n519 4.65
R697 GND.n517 GND.n516 4.65
R698 GND.n514 GND.n513 4.65
R699 GND.n511 GND.n510 4.65
R700 GND.n506 GND.n505 4.65
R701 GND.n503 GND.n502 4.65
R702 GND.n496 GND.n495 4.65
R703 GND.n493 GND.n492 4.65
R704 GND.n490 GND.n489 4.65
R705 GND.n487 GND.n486 4.65
R706 GND.n484 GND.n483 4.65
R707 GND.n481 GND.n480 4.65
R708 GND.n478 GND.n477 4.65
R709 GND.n475 GND.n474 4.65
R710 GND.n472 GND.n471 4.65
R711 GND.n469 GND.n468 4.65
R712 GND.n464 GND.n463 4.65
R713 GND.n7 GND.n6 4.65
R714 GND.n13 GND.n12 4.65
R715 GND.n24 GND.n23 4.65
R716 GND.n27 GND.n26 4.65
R717 GND.n34 GND.n33 4.65
R718 GND.n37 GND.n36 4.65
R719 GND.n40 GND.n39 4.65
R720 GND.n43 GND.n42 4.65
R721 GND.n46 GND.n45 4.65
R722 GND.n53 GND.n52 4.65
R723 GND.n56 GND.n55 4.65
R724 GND.n59 GND.n58 4.65
R725 GND.n66 GND.n65 4.65
R726 GND.n69 GND.n68 4.65
R727 GND.n72 GND.n71 4.65
R728 GND.n15 GND.n14 4.504
R729 GND.n6 GND.n4 4.129
R730 GND.n52 GND.n50 4.129
R731 GND.n84 GND.n82 4.129
R732 GND.n116 GND.n114 4.129
R733 GND.n23 GND.n21 3.716
R734 GND.t8 GND.n15 2.452
R735 GND.n1 GND.n0 0.475
R736 GND.n460 GND.n459 0.474
R737 GND.n9 GND.n8 0.376
R738 GND.n34 GND.n27 0.29
R739 GND.n66 GND.n59 0.29
R740 GND.n98 GND.n91 0.29
R741 GND.n130 GND.n123 0.29
R742 GND.n174 GND.n167 0.29
R743 GND.n218 GND.n211 0.29
R744 GND.n260 GND.n253 0.29
R745 GND.n304 GND.n297 0.29
R746 GND.n346 GND.n339 0.29
R747 GND.n390 GND.n383 0.29
R748 GND.n434 GND.n427 0.29
R749 GND.n894 GND.n887 0.29
R750 GND.n852 GND.n845 0.29
R751 GND.n810 GND.n803 0.29
R752 GND.n765 GND.n758 0.29
R753 GND.n720 GND.n713 0.29
R754 GND.n675 GND.n668 0.29
R755 GND.n631 GND.n624 0.29
R756 GND.n587 GND.n580 0.29
R757 GND.n545 GND.n538 0.29
R758 GND.n503 GND.n496 0.29
R759 GND.n461 GND 0.207
R760 GND.n12 GND.n10 0.206
R761 GND.n160 GND.n159 0.206
R762 GND.n204 GND.n203 0.206
R763 GND.n246 GND.n245 0.206
R764 GND.n290 GND.n289 0.206
R765 GND.n332 GND.n331 0.206
R766 GND.n376 GND.n375 0.206
R767 GND.n420 GND.n419 0.206
R768 GND.n901 GND.n900 0.206
R769 GND.n859 GND.n858 0.206
R770 GND.n817 GND.n816 0.206
R771 GND.n775 GND.n774 0.206
R772 GND.n730 GND.n729 0.206
R773 GND.n685 GND.n684 0.206
R774 GND.n640 GND.n639 0.206
R775 GND.n596 GND.n595 0.206
R776 GND.n552 GND.n551 0.206
R777 GND.n510 GND.n509 0.206
R778 GND.n468 GND.n467 0.206
R779 GND.n148 GND.n145 0.197
R780 GND.n192 GND.n189 0.197
R781 GND.n236 GND.n233 0.197
R782 GND.n278 GND.n275 0.197
R783 GND.n322 GND.n319 0.197
R784 GND.n364 GND.n361 0.197
R785 GND.n408 GND.n405 0.197
R786 GND.n452 GND.n449 0.197
R787 GND.n872 GND.n869 0.197
R788 GND.n830 GND.n827 0.197
R789 GND.n788 GND.n785 0.197
R790 GND.n743 GND.n740 0.197
R791 GND.n698 GND.n695 0.197
R792 GND.n653 GND.n650 0.197
R793 GND.n609 GND.n606 0.197
R794 GND.n565 GND.n562 0.197
R795 GND.n523 GND.n520 0.197
R796 GND.n481 GND.n478 0.197
R797 GND.n46 GND.n43 0.181
R798 GND.n78 GND.n75 0.181
R799 GND.n110 GND.n107 0.181
R800 GND.n13 GND.n7 0.157
R801 GND.n24 GND.n13 0.157
R802 GND.n27 GND.n24 0.145
R803 GND.n37 GND.n34 0.145
R804 GND.n40 GND.n37 0.145
R805 GND.n43 GND.n40 0.145
R806 GND.n53 GND.n46 0.145
R807 GND.n56 GND.n53 0.145
R808 GND.n59 GND.n56 0.145
R809 GND.n69 GND.n66 0.145
R810 GND.n72 GND.n69 0.145
R811 GND.n75 GND.n72 0.145
R812 GND.n85 GND.n78 0.145
R813 GND.n88 GND.n85 0.145
R814 GND.n91 GND.n88 0.145
R815 GND.n101 GND.n98 0.145
R816 GND.n104 GND.n101 0.145
R817 GND.n107 GND.n104 0.145
R818 GND.n117 GND.n110 0.145
R819 GND.n120 GND.n117 0.145
R820 GND.n123 GND.n120 0.145
R821 GND.n133 GND.n130 0.145
R822 GND.n136 GND.n133 0.145
R823 GND.n139 GND.n136 0.145
R824 GND.n142 GND.n139 0.145
R825 GND.n145 GND.n142 0.145
R826 GND.n151 GND.n148 0.145
R827 GND.n154 GND.n151 0.145
R828 GND.n161 GND.n154 0.145
R829 GND.n164 GND.n161 0.145
R830 GND.n167 GND.n164 0.145
R831 GND.n177 GND.n174 0.145
R832 GND.n180 GND.n177 0.145
R833 GND.n183 GND.n180 0.145
R834 GND.n186 GND.n183 0.145
R835 GND.n189 GND.n186 0.145
R836 GND.n195 GND.n192 0.145
R837 GND.n198 GND.n195 0.145
R838 GND.n205 GND.n198 0.145
R839 GND.n208 GND.n205 0.145
R840 GND.n211 GND.n208 0.145
R841 GND.n221 GND.n218 0.145
R842 GND.n224 GND.n221 0.145
R843 GND.n227 GND.n224 0.145
R844 GND.n230 GND.n227 0.145
R845 GND.n233 GND.n230 0.145
R846 GND.n239 GND.n236 0.145
R847 GND.n242 GND.n239 0.145
R848 GND.n247 GND.n242 0.145
R849 GND.n250 GND.n247 0.145
R850 GND.n253 GND.n250 0.145
R851 GND.n263 GND.n260 0.145
R852 GND.n266 GND.n263 0.145
R853 GND.n269 GND.n266 0.145
R854 GND.n272 GND.n269 0.145
R855 GND.n275 GND.n272 0.145
R856 GND.n281 GND.n278 0.145
R857 GND.n284 GND.n281 0.145
R858 GND.n291 GND.n284 0.145
R859 GND.n294 GND.n291 0.145
R860 GND.n297 GND.n294 0.145
R861 GND.n307 GND.n304 0.145
R862 GND.n310 GND.n307 0.145
R863 GND.n313 GND.n310 0.145
R864 GND.n316 GND.n313 0.145
R865 GND.n319 GND.n316 0.145
R866 GND.n325 GND.n322 0.145
R867 GND.n328 GND.n325 0.145
R868 GND.n333 GND.n328 0.145
R869 GND.n336 GND.n333 0.145
R870 GND.n339 GND.n336 0.145
R871 GND.n349 GND.n346 0.145
R872 GND.n352 GND.n349 0.145
R873 GND.n355 GND.n352 0.145
R874 GND.n358 GND.n355 0.145
R875 GND.n361 GND.n358 0.145
R876 GND.n367 GND.n364 0.145
R877 GND.n370 GND.n367 0.145
R878 GND.n377 GND.n370 0.145
R879 GND.n380 GND.n377 0.145
R880 GND.n383 GND.n380 0.145
R881 GND.n393 GND.n390 0.145
R882 GND.n396 GND.n393 0.145
R883 GND.n399 GND.n396 0.145
R884 GND.n402 GND.n399 0.145
R885 GND.n405 GND.n402 0.145
R886 GND.n411 GND.n408 0.145
R887 GND.n414 GND.n411 0.145
R888 GND.n421 GND.n414 0.145
R889 GND.n424 GND.n421 0.145
R890 GND.n427 GND.n424 0.145
R891 GND.n437 GND.n434 0.145
R892 GND.n440 GND.n437 0.145
R893 GND.n443 GND.n440 0.145
R894 GND.n446 GND.n443 0.145
R895 GND.n449 GND.n446 0.145
R896 GND.n455 GND.n452 0.145
R897 GND.n458 GND.n455 0.145
R898 GND.n902 GND.n897 0.145
R899 GND.n897 GND.n894 0.145
R900 GND.n887 GND.n884 0.145
R901 GND.n884 GND.n881 0.145
R902 GND.n881 GND.n878 0.145
R903 GND.n878 GND.n875 0.145
R904 GND.n875 GND.n872 0.145
R905 GND.n869 GND.n866 0.145
R906 GND.n866 GND.n863 0.145
R907 GND.n863 GND.n860 0.145
R908 GND.n860 GND.n855 0.145
R909 GND.n855 GND.n852 0.145
R910 GND.n845 GND.n842 0.145
R911 GND.n842 GND.n839 0.145
R912 GND.n839 GND.n836 0.145
R913 GND.n836 GND.n833 0.145
R914 GND.n833 GND.n830 0.145
R915 GND.n827 GND.n824 0.145
R916 GND.n824 GND.n821 0.145
R917 GND.n821 GND.n818 0.145
R918 GND.n818 GND.n813 0.145
R919 GND.n813 GND.n810 0.145
R920 GND.n803 GND.n800 0.145
R921 GND.n800 GND.n797 0.145
R922 GND.n797 GND.n794 0.145
R923 GND.n794 GND.n791 0.145
R924 GND.n791 GND.n788 0.145
R925 GND.n785 GND.n782 0.145
R926 GND.n782 GND.n779 0.145
R927 GND.n779 GND.n776 0.145
R928 GND.n776 GND.n768 0.145
R929 GND.n768 GND.n765 0.145
R930 GND.n758 GND.n755 0.145
R931 GND.n755 GND.n752 0.145
R932 GND.n752 GND.n749 0.145
R933 GND.n749 GND.n746 0.145
R934 GND.n746 GND.n743 0.145
R935 GND.n740 GND.n737 0.145
R936 GND.n737 GND.n734 0.145
R937 GND.n734 GND.n731 0.145
R938 GND.n731 GND.n723 0.145
R939 GND.n723 GND.n720 0.145
R940 GND.n713 GND.n710 0.145
R941 GND.n710 GND.n707 0.145
R942 GND.n707 GND.n704 0.145
R943 GND.n704 GND.n701 0.145
R944 GND.n701 GND.n698 0.145
R945 GND.n695 GND.n692 0.145
R946 GND.n692 GND.n689 0.145
R947 GND.n689 GND.n686 0.145
R948 GND.n686 GND.n678 0.145
R949 GND.n678 GND.n675 0.145
R950 GND.n668 GND.n665 0.145
R951 GND.n665 GND.n662 0.145
R952 GND.n662 GND.n659 0.145
R953 GND.n659 GND.n656 0.145
R954 GND.n656 GND.n653 0.145
R955 GND.n650 GND.n647 0.145
R956 GND.n647 GND.n644 0.145
R957 GND.n644 GND.n641 0.145
R958 GND.n641 GND.n634 0.145
R959 GND.n634 GND.n631 0.145
R960 GND.n624 GND.n621 0.145
R961 GND.n621 GND.n618 0.145
R962 GND.n618 GND.n615 0.145
R963 GND.n615 GND.n612 0.145
R964 GND.n612 GND.n609 0.145
R965 GND.n606 GND.n603 0.145
R966 GND.n603 GND.n600 0.145
R967 GND.n600 GND.n597 0.145
R968 GND.n597 GND.n590 0.145
R969 GND.n590 GND.n587 0.145
R970 GND.n580 GND.n577 0.145
R971 GND.n577 GND.n574 0.145
R972 GND.n574 GND.n571 0.145
R973 GND.n571 GND.n568 0.145
R974 GND.n568 GND.n565 0.145
R975 GND.n562 GND.n559 0.145
R976 GND.n559 GND.n556 0.145
R977 GND.n556 GND.n553 0.145
R978 GND.n553 GND.n548 0.145
R979 GND.n548 GND.n545 0.145
R980 GND.n538 GND.n535 0.145
R981 GND.n535 GND.n532 0.145
R982 GND.n532 GND.n529 0.145
R983 GND.n529 GND.n526 0.145
R984 GND.n526 GND.n523 0.145
R985 GND.n520 GND.n517 0.145
R986 GND.n517 GND.n514 0.145
R987 GND.n514 GND.n511 0.145
R988 GND.n511 GND.n506 0.145
R989 GND.n506 GND.n503 0.145
R990 GND.n496 GND.n493 0.145
R991 GND.n493 GND.n490 0.145
R992 GND.n490 GND.n487 0.145
R993 GND.n487 GND.n484 0.145
R994 GND.n484 GND.n481 0.145
R995 GND.n478 GND.n475 0.145
R996 GND.n475 GND.n472 0.145
R997 GND.n472 GND.n469 0.145
R998 GND.n469 GND.n464 0.145
R999 GND.n464 GND.n461 0.145
R1000 GND GND.n902 0.086
R1001 GND GND.n458 0.058
R1002 a_15669_1050.n5 a_15669_1050.t9 512.525
R1003 a_15669_1050.n5 a_15669_1050.t7 371.139
R1004 a_15669_1050.n6 a_15669_1050.t8 361.392
R1005 a_15669_1050.n9 a_15669_1050.n7 314.738
R1006 a_15669_1050.n6 a_15669_1050.n5 235.554
R1007 a_15669_1050.n7 a_15669_1050.n4 179.199
R1008 a_15669_1050.n3 a_15669_1050.n2 161.352
R1009 a_15669_1050.n4 a_15669_1050.n0 95.095
R1010 a_15669_1050.n3 a_15669_1050.n1 95.095
R1011 a_15669_1050.n4 a_15669_1050.n3 66.258
R1012 a_15669_1050.n9 a_15669_1050.n8 15.218
R1013 a_15669_1050.n0 a_15669_1050.t6 14.282
R1014 a_15669_1050.n0 a_15669_1050.t1 14.282
R1015 a_15669_1050.n1 a_15669_1050.t3 14.282
R1016 a_15669_1050.n1 a_15669_1050.t4 14.282
R1017 a_15669_1050.n2 a_15669_1050.t5 14.282
R1018 a_15669_1050.n2 a_15669_1050.t2 14.282
R1019 a_15669_1050.n10 a_15669_1050.n9 12.014
R1020 a_15669_1050.n7 a_15669_1050.n6 10.615
R1021 VDD.n889 VDD.n878 144.705
R1022 VDD.n964 VDD.n957 144.705
R1023 VDD.n1039 VDD.n1032 144.705
R1024 VDD.n1114 VDD.n1107 144.705
R1025 VDD.n1189 VDD.n1182 144.705
R1026 VDD.n1264 VDD.n1257 144.705
R1027 VDD.n1339 VDD.n1332 144.705
R1028 VDD.n1414 VDD.n1407 144.705
R1029 VDD.n1489 VDD.n1482 144.705
R1030 VDD.n754 VDD.n747 144.705
R1031 VDD.n1564 VDD.n1557 144.705
R1032 VDD.n679 VDD.n672 144.705
R1033 VDD.n604 VDD.n597 144.705
R1034 VDD.n529 VDD.n522 144.705
R1035 VDD.n454 VDD.n447 144.705
R1036 VDD.n379 VDD.n372 144.705
R1037 VDD.n304 VDD.n297 144.705
R1038 VDD.n229 VDD.n222 144.705
R1039 VDD.n172 VDD.n165 144.705
R1040 VDD.n119 VDD.n112 144.705
R1041 VDD.n66 VDD.n55 144.705
R1042 VDD.n855 VDD.t199 143.754
R1043 VDD.n931 VDD.t16 143.754
R1044 VDD.n1006 VDD.t194 143.754
R1045 VDD.n1081 VDD.t168 143.754
R1046 VDD.n1156 VDD.t190 143.754
R1047 VDD.n1231 VDD.t22 143.754
R1048 VDD.n1306 VDD.t184 143.754
R1049 VDD.n1381 VDD.t104 143.754
R1050 VDD.n1456 VDD.t196 143.754
R1051 VDD.n1531 VDD.t156 143.754
R1052 VDD.n763 VDD.t217 143.754
R1053 VDD.n688 VDD.t205 143.754
R1054 VDD.n613 VDD.t36 143.754
R1055 VDD.n538 VDD.t229 143.754
R1056 VDD.n463 VDD.t235 143.754
R1057 VDD.n388 VDD.t146 143.754
R1058 VDD.n313 VDD.t211 143.754
R1059 VDD.n238 VDD.t233 143.754
R1060 VDD.n197 VDD.t44 135.539
R1061 VDD.n175 VDD.t91 135.539
R1062 VDD.n820 VDD.t130 135.17
R1063 VDD.n896 VDD.t7 135.17
R1064 VDD.n971 VDD.t106 135.17
R1065 VDD.n1046 VDD.t30 135.17
R1066 VDD.n1121 VDD.t48 135.17
R1067 VDD.n1196 VDD.t124 135.17
R1068 VDD.n1271 VDD.t132 135.17
R1069 VDD.n1346 VDD.t221 135.17
R1070 VDD.n1421 VDD.t118 135.17
R1071 VDD.n1496 VDD.t112 135.17
R1072 VDD.n1571 VDD.t79 135.17
R1073 VDD.n718 VDD.t34 135.17
R1074 VDD.n643 VDD.t134 135.17
R1075 VDD.n568 VDD.t54 135.17
R1076 VDD.n493 VDD.t18 135.17
R1077 VDD.n418 VDD.t207 135.17
R1078 VDD.n343 VDD.t75 135.17
R1079 VDD.n268 VDD.t140 135.17
R1080 VDD.n35 VDD.t28 135.17
R1081 VDD.n24 VDD.t11 135.17
R1082 VDD.n185 VDD.n184 129.849
R1083 VDD.n830 VDD.n829 129.472
R1084 VDD.n846 VDD.n845 129.472
R1085 VDD.n906 VDD.n905 129.472
R1086 VDD.n922 VDD.n921 129.472
R1087 VDD.n981 VDD.n980 129.472
R1088 VDD.n997 VDD.n996 129.472
R1089 VDD.n1056 VDD.n1055 129.472
R1090 VDD.n1072 VDD.n1071 129.472
R1091 VDD.n1131 VDD.n1130 129.472
R1092 VDD.n1147 VDD.n1146 129.472
R1093 VDD.n1206 VDD.n1205 129.472
R1094 VDD.n1222 VDD.n1221 129.472
R1095 VDD.n1281 VDD.n1280 129.472
R1096 VDD.n1297 VDD.n1296 129.472
R1097 VDD.n1356 VDD.n1355 129.472
R1098 VDD.n1372 VDD.n1371 129.472
R1099 VDD.n1431 VDD.n1430 129.472
R1100 VDD.n1447 VDD.n1446 129.472
R1101 VDD.n1506 VDD.n1505 129.472
R1102 VDD.n1522 VDD.n1521 129.472
R1103 VDD.n784 VDD.n783 129.472
R1104 VDD.n772 VDD.n771 129.472
R1105 VDD.n709 VDD.n708 129.472
R1106 VDD.n697 VDD.n696 129.472
R1107 VDD.n634 VDD.n633 129.472
R1108 VDD.n622 VDD.n621 129.472
R1109 VDD.n559 VDD.n558 129.472
R1110 VDD.n547 VDD.n546 129.472
R1111 VDD.n484 VDD.n483 129.472
R1112 VDD.n472 VDD.n471 129.472
R1113 VDD.n409 VDD.n408 129.472
R1114 VDD.n397 VDD.n396 129.472
R1115 VDD.n334 VDD.n333 129.472
R1116 VDD.n322 VDD.n321 129.472
R1117 VDD.n259 VDD.n258 129.472
R1118 VDD.n247 VDD.n246 129.472
R1119 VDD.n51 VDD.n50 92.5
R1120 VDD.n49 VDD.n48 92.5
R1121 VDD.n47 VDD.n46 92.5
R1122 VDD.n45 VDD.n44 92.5
R1123 VDD.n53 VDD.n52 92.5
R1124 VDD.n108 VDD.n107 92.5
R1125 VDD.n106 VDD.n105 92.5
R1126 VDD.n104 VDD.n103 92.5
R1127 VDD.n102 VDD.n101 92.5
R1128 VDD.n110 VDD.n109 92.5
R1129 VDD.n161 VDD.n160 92.5
R1130 VDD.n159 VDD.n158 92.5
R1131 VDD.n157 VDD.n156 92.5
R1132 VDD.n155 VDD.n154 92.5
R1133 VDD.n163 VDD.n162 92.5
R1134 VDD.n218 VDD.n217 92.5
R1135 VDD.n216 VDD.n215 92.5
R1136 VDD.n214 VDD.n213 92.5
R1137 VDD.n212 VDD.n211 92.5
R1138 VDD.n220 VDD.n219 92.5
R1139 VDD.n293 VDD.n292 92.5
R1140 VDD.n291 VDD.n290 92.5
R1141 VDD.n289 VDD.n288 92.5
R1142 VDD.n287 VDD.n286 92.5
R1143 VDD.n295 VDD.n294 92.5
R1144 VDD.n368 VDD.n367 92.5
R1145 VDD.n366 VDD.n365 92.5
R1146 VDD.n364 VDD.n363 92.5
R1147 VDD.n362 VDD.n361 92.5
R1148 VDD.n370 VDD.n369 92.5
R1149 VDD.n443 VDD.n442 92.5
R1150 VDD.n441 VDD.n440 92.5
R1151 VDD.n439 VDD.n438 92.5
R1152 VDD.n437 VDD.n436 92.5
R1153 VDD.n445 VDD.n444 92.5
R1154 VDD.n518 VDD.n517 92.5
R1155 VDD.n516 VDD.n515 92.5
R1156 VDD.n514 VDD.n513 92.5
R1157 VDD.n512 VDD.n511 92.5
R1158 VDD.n520 VDD.n519 92.5
R1159 VDD.n593 VDD.n592 92.5
R1160 VDD.n591 VDD.n590 92.5
R1161 VDD.n589 VDD.n588 92.5
R1162 VDD.n587 VDD.n586 92.5
R1163 VDD.n595 VDD.n594 92.5
R1164 VDD.n668 VDD.n667 92.5
R1165 VDD.n666 VDD.n665 92.5
R1166 VDD.n664 VDD.n663 92.5
R1167 VDD.n662 VDD.n661 92.5
R1168 VDD.n670 VDD.n669 92.5
R1169 VDD.n743 VDD.n742 92.5
R1170 VDD.n741 VDD.n740 92.5
R1171 VDD.n739 VDD.n738 92.5
R1172 VDD.n737 VDD.n736 92.5
R1173 VDD.n745 VDD.n744 92.5
R1174 VDD.n1553 VDD.n1552 92.5
R1175 VDD.n1551 VDD.n1550 92.5
R1176 VDD.n1549 VDD.n1548 92.5
R1177 VDD.n1547 VDD.n1546 92.5
R1178 VDD.n1555 VDD.n1554 92.5
R1179 VDD.n1478 VDD.n1477 92.5
R1180 VDD.n1476 VDD.n1475 92.5
R1181 VDD.n1474 VDD.n1473 92.5
R1182 VDD.n1472 VDD.n1471 92.5
R1183 VDD.n1480 VDD.n1479 92.5
R1184 VDD.n1403 VDD.n1402 92.5
R1185 VDD.n1401 VDD.n1400 92.5
R1186 VDD.n1399 VDD.n1398 92.5
R1187 VDD.n1397 VDD.n1396 92.5
R1188 VDD.n1405 VDD.n1404 92.5
R1189 VDD.n1328 VDD.n1327 92.5
R1190 VDD.n1326 VDD.n1325 92.5
R1191 VDD.n1324 VDD.n1323 92.5
R1192 VDD.n1322 VDD.n1321 92.5
R1193 VDD.n1330 VDD.n1329 92.5
R1194 VDD.n1253 VDD.n1252 92.5
R1195 VDD.n1251 VDD.n1250 92.5
R1196 VDD.n1249 VDD.n1248 92.5
R1197 VDD.n1247 VDD.n1246 92.5
R1198 VDD.n1255 VDD.n1254 92.5
R1199 VDD.n1178 VDD.n1177 92.5
R1200 VDD.n1176 VDD.n1175 92.5
R1201 VDD.n1174 VDD.n1173 92.5
R1202 VDD.n1172 VDD.n1171 92.5
R1203 VDD.n1180 VDD.n1179 92.5
R1204 VDD.n1103 VDD.n1102 92.5
R1205 VDD.n1101 VDD.n1100 92.5
R1206 VDD.n1099 VDD.n1098 92.5
R1207 VDD.n1097 VDD.n1096 92.5
R1208 VDD.n1105 VDD.n1104 92.5
R1209 VDD.n1028 VDD.n1027 92.5
R1210 VDD.n1026 VDD.n1025 92.5
R1211 VDD.n1024 VDD.n1023 92.5
R1212 VDD.n1022 VDD.n1021 92.5
R1213 VDD.n1030 VDD.n1029 92.5
R1214 VDD.n953 VDD.n952 92.5
R1215 VDD.n951 VDD.n950 92.5
R1216 VDD.n949 VDD.n948 92.5
R1217 VDD.n947 VDD.n946 92.5
R1218 VDD.n955 VDD.n954 92.5
R1219 VDD.n874 VDD.n873 92.5
R1220 VDD.n872 VDD.n871 92.5
R1221 VDD.n870 VDD.n869 92.5
R1222 VDD.n868 VDD.n867 92.5
R1223 VDD.n876 VDD.n875 92.5
R1224 VDD.n804 VDD.n803 92.5
R1225 VDD.n802 VDD.n801 92.5
R1226 VDD.n800 VDD.n799 92.5
R1227 VDD.n798 VDD.n797 92.5
R1228 VDD.n806 VDD.n805 92.5
R1229 VDD.n14 VDD.n1 92.5
R1230 VDD.n5 VDD.n4 92.5
R1231 VDD.n7 VDD.n6 92.5
R1232 VDD.n9 VDD.n8 92.5
R1233 VDD.n11 VDD.n10 92.5
R1234 VDD.n13 VDD.n12 92.5
R1235 VDD.n21 VDD.n20 92.059
R1236 VDD.n65 VDD.n64 92.059
R1237 VDD.n118 VDD.n117 92.059
R1238 VDD.n171 VDD.n170 92.059
R1239 VDD.n228 VDD.n227 92.059
R1240 VDD.n303 VDD.n302 92.059
R1241 VDD.n378 VDD.n377 92.059
R1242 VDD.n453 VDD.n452 92.059
R1243 VDD.n528 VDD.n527 92.059
R1244 VDD.n603 VDD.n602 92.059
R1245 VDD.n678 VDD.n677 92.059
R1246 VDD.n753 VDD.n752 92.059
R1247 VDD.n1563 VDD.n1562 92.059
R1248 VDD.n1488 VDD.n1487 92.059
R1249 VDD.n1413 VDD.n1412 92.059
R1250 VDD.n1338 VDD.n1337 92.059
R1251 VDD.n1263 VDD.n1262 92.059
R1252 VDD.n1188 VDD.n1187 92.059
R1253 VDD.n1113 VDD.n1112 92.059
R1254 VDD.n1038 VDD.n1037 92.059
R1255 VDD.n963 VDD.n962 92.059
R1256 VDD.n888 VDD.n887 92.059
R1257 VDD.n812 VDD.n811 92.059
R1258 VDD.n20 VDD.n16 67.194
R1259 VDD.n20 VDD.n17 67.194
R1260 VDD.n20 VDD.n18 67.194
R1261 VDD.n20 VDD.n19 67.194
R1262 VDD.n796 VDD.n795 44.141
R1263 VDD.n945 VDD.n944 44.141
R1264 VDD.n1020 VDD.n1019 44.141
R1265 VDD.n1095 VDD.n1094 44.141
R1266 VDD.n1170 VDD.n1169 44.141
R1267 VDD.n1245 VDD.n1244 44.141
R1268 VDD.n1320 VDD.n1319 44.141
R1269 VDD.n1395 VDD.n1394 44.141
R1270 VDD.n1470 VDD.n1469 44.141
R1271 VDD.n1545 VDD.n1544 44.141
R1272 VDD.n735 VDD.n734 44.141
R1273 VDD.n660 VDD.n659 44.141
R1274 VDD.n585 VDD.n584 44.141
R1275 VDD.n510 VDD.n509 44.141
R1276 VDD.n435 VDD.n434 44.141
R1277 VDD.n360 VDD.n359 44.141
R1278 VDD.n285 VDD.n284 44.141
R1279 VDD.n210 VDD.n209 44.141
R1280 VDD.n153 VDD.n152 44.141
R1281 VDD.n100 VDD.n99 44.141
R1282 VDD.n5 VDD.n3 44.141
R1283 VDD.n944 VDD.n942 44.107
R1284 VDD.n1019 VDD.n1017 44.107
R1285 VDD.n1094 VDD.n1092 44.107
R1286 VDD.n1169 VDD.n1167 44.107
R1287 VDD.n1244 VDD.n1242 44.107
R1288 VDD.n1319 VDD.n1317 44.107
R1289 VDD.n1394 VDD.n1392 44.107
R1290 VDD.n1469 VDD.n1467 44.107
R1291 VDD.n1544 VDD.n1542 44.107
R1292 VDD.n734 VDD.n732 44.107
R1293 VDD.n659 VDD.n657 44.107
R1294 VDD.n584 VDD.n582 44.107
R1295 VDD.n509 VDD.n507 44.107
R1296 VDD.n434 VDD.n432 44.107
R1297 VDD.n359 VDD.n357 44.107
R1298 VDD.n284 VDD.n282 44.107
R1299 VDD.n209 VDD.n207 44.107
R1300 VDD.n152 VDD.n150 44.107
R1301 VDD.n99 VDD.n97 44.107
R1302 VDD.n795 VDD.n793 44.107
R1303 VDD.n3 VDD.n2 44.107
R1304 VDD.n25 �3h�9V 43.472
R1305 VDD.n33  43.472
R1306 VDD.n20 VDD.n15 41.052
R1307 VDD.n59 VDD.n57 39.742
R1308 VDD.n59 VDD.n58 39.742
R1309 VDD.n61 VDD.n60 39.742
R1310 VDD.n114 VDD.n113 39.742
R1311 VDD.n167 VDD.n166 39.742
R1312 VDD.n224 VDD.n223 39.742
R1313 VDD.n299 VDD.n298 39.742
R1314 VDD.n374 VDD.n373 39.742
R1315 VDD.n449 VDD.n448 39.742
R1316 VDD.n524 VDD.n523 39.742
R1317 VDD.n599 VDD.n598 39.742
R1318 VDD.n674 VDD.n673 39.742
R1319 VDD.n749 VDD.n748 39.742
R1320 VDD.n1559 VDD.n1558 39.742
R1321 VDD.n1484 VDD.n1483 39.742
R1322 VDD.n1409 VDD.n1408 39.742
R1323 VDD.n1334 VDD.n1333 39.742
R1324 VDD.n1259 VDD.n1258 39.742
R1325 VDD.n1184 VDD.n1183 39.742
R1326 VDD.n1109 VDD.n1108 39.742
R1327 VDD.n1034 VDD.n1033 39.742
R1328 VDD.n959 VDD.n958 39.742
R1329 VDD.n808 VDD.n807 39.742
R1330 VDD.n886 VDD.n883 39.742
R1331 VDD.n886 VDD.n885 39.742
R1332 VDD.n882 VDD.n881 39.742
R1333 VDD.n99 VDD.n98 38
R1334 VDD.n152 VDD.n151 38
R1335 VDD.n209 VDD.n208 38
R1336 VDD.n284 VDD.n283 38
R1337 VDD.n359 VDD.n358 38
R1338 VDD.n434 VDD.n433 38
R1339 VDD.n509 VDD.n508 38
R1340 VDD.n584 VDD.n583 38
R1341 VDD.n659 VDD.n658 38
R1342 VDD.n734 VDD.n733 38
R1343 VDD.n1544 VDD.n1543 38
R1344 VDD.n1469 VDD.n1468 38
R1345 VDD.n1394 VDD.n1393 38
R1346 VDD.n1319 VDD.n1318 38
R1347 VDD.n1244 VDD.n1243 38
R1348 VDD.n1169 VDD.n1168 38
R1349 VDD.n1094 VDD.n1093 38
R1350 VDD.n1019 VDD.n1018 38
R1351 VDD.n944 VDD.n943 38
R1352 VDD.n795 VDD.n794 38
R1353 VDD.n942 VDD.n941 36.774
R1354 VDD.n1017 VDD.n1016 36.774
R1355 VDD.n1092 VDD.n1091 36.774
R1356 VDD.n1167 VDD.n1166 36.774
R1357 VDD.n1242 VDD.n1241 36.774
R1358 VDD.n1317 VDD.n1316 36.774
R1359 VDD.n1392 VDD.n1391 36.774
R1360 VDD.n1467 VDD.n1466 36.774
R1361 VDD.n1542 VDD.n1541 36.774
R1362 VDD.n732 VDD.n731 36.774
R1363 VDD.n657 VDD.n656 36.774
R1364 VDD.n582 VDD.n581 36.774
R1365 VDD.n507 VDD.n506 36.774
R1366 VDD.n432 VDD.n431 36.774
R1367 VDD.n357 VDD.n356 36.774
R1368 VDD.n282 VDD.n281 36.774
R1369 VDD.n207 VDD.n206 36.774
R1370 VDD.n150 VDD.n149 36.774
R1371 VDD.n97 VDD.n96 36.774
R1372 VDD.n57 VDD.n56 36.774
R1373 VDD.n885 VDD.n884 36.774
R1374 VDD.n240 VDD.t232 35.8
R1375 VDD.n315 ���9V 35.8
R1376 VDD.n390  W�9V 35.8
R1377 VDD.n465 ��ў9V 35.8
R1378 VDD.n540 @�9V 35.8
R1379 VDD.n615 �fb�9V 35.8
R1380 VDD.n690  35.8
R1381 VDD.n765  35.8
R1382 VDD.n1525 VDD.t155 35.8
R1383 VDD.n1450  35.8
R1384 VDD.n1375 �WȞ9V 35.8
R1385 VDD.n1300  35.8
R1386 VDD.n1225 `>H�9V 35.8
R1387 VDD.n1150  35.8
R1388 VDD.n1075 P��9V 35.8
R1389 VDD.n1000 `b��9V 35.8
R1390 VDD.n925 ���9V 35.8
R1391 VDD.n849 ����9V 35.8
R1392 VDD.n264 �+�إ 33.243
R1393 VDD.n339 VDD.t74 33.243
R1394 VDD.n414 @��9V 33.243
R1395 VDD.n489  33.243
R1396 VDD.n564 P�ԝ9V 33.243
R1397 VDD.n639 �H�9V 33.243
R1398 VDD.n714 �J�9V 33.243
R1399 VDD.n789 P��9V 33.243
R1400 VDD.n1501  �ɝ9V 33.243
R1401 VDD.n1426 @Q��9V 33.243
R1402 VDD.n1351 �}ߝ9V 33.243
R1403 VDD.n1276 ���9V 33.243
R1404 VDD.n1201  33.243
R1405 VDD.n1126 ��b�9V 33.243
R1406 VDD.n1051 �+�إ 33.243
R1407 VDD.n976 VDD.t105 33.243
R1408 VDD.n901 ��ѝ9V 33.243
R1409 VDD.n825 VDD.t129 33.243
R1410 VDD.n1 VDD.n0 30.923
R1411 VDD.n64 VDD.n62 26.38
R1412 VDD.n64 VDD.n61 26.38
R1413 VDD.n64 VDD.n59 26.38
R1414 VDD.n64 VDD.n63 26.38
R1415 VDD.n117 VDD.n115 26.38
R1416 VDD.n117 VDD.n114 26.38
R1417 VDD.n117 VDD.n116 26.38
R1418 VDD.n170 VDD.n168 26.38
R1419 VDD.n170 VDD.n167 26.38
R1420 VDD.n170 VDD.n169 26.38
R1421 VDD.n227 VDD.n225 26.38
R1422 VDD.n227 VDD.n224 26.38
R1423 VDD.n227 VDD.n226 26.38
R1424 VDD.n302 VDD.n300 26.38
R1425 VDD.n302 VDD.n299 26.38
R1426 VDD.n302 VDD.n301 26.38
R1427 VDD.n377 VDD.n375 26.38
R1428 VDD.n377 VDD.n374 26.38
R1429 VDD.n377 VDD.n376 26.38
R1430 VDD.n452 VDD.n450 26.38
R1431 VDD.n452 VDD.n449 26.38
R1432 VDD.n452 VDD.n451 26.38
R1433 VDD.n527 VDD.n525 26.38
R1434 VDD.n527 VDD.n524 26.38
R1435 VDD.n527 VDD.n526 26.38
R1436 VDD.n602 VDD.n600 26.38
R1437 VDD.n602 VDD.n599 26.38
R1438 VDD.n602 VDD.n601 26.38
R1439 VDD.n677 VDD.n675 26.38
R1440 VDD.n677 VDD.n674 26.38
R1441 VDD.n677 VDD.n676 26.38
R1442 VDD.n752 VDD.n750 26.38
R1443 VDD.n752 VDD.n749 26.38
R1444 VDD.n752 VDD.n751 26.38
R1445 VDD.n1562 VDD.n1560 26.38
R1446 VDD.n1562 VDD.n1559 26.38
R1447 VDD.n1562 VDD.n1561 26.38
R1448 VDD.n1487 VDD.n1485 26.38
R1449 VDD.n1487 VDD.n1484 26.38
R1450 VDD.n1487 VDD.n1486 26.38
R1451 VDD.n1412 VDD.n1410 26.38
R1452 VDD.n1412 VDD.n1409 26.38
R1453 VDD.n1412 VDD.n1411 26.38
R1454 VDD.n1337 VDD.n1335 26.38
R1455 VDD.n1337 VDD.n1334 26.38
R1456 VDD.n1337 VDD.n1336 26.38
R1457 VDD.n1262 VDD.n1260 26.38
R1458 VDD.n1262 VDD.n1259 26.38
R1459 VDD.n1262 VDD.n1261 26.38
R1460 VDD.n1187 VDD.n1185 26.38
R1461 VDD.n1187 VDD.n1184 26.38
R1462 VDD.n1187 VDD.n1186 26.38
R1463 VDD.n1112 VDD.n1110 26.38
R1464 VDD.n1112 VDD.n1109 26.38
R1465 VDD.n1112 VDD.n1111 26.38
R1466 VDD.n1037 VDD.n1035 26.38
R1467 VDD.n1037 VDD.n1034 26.38
R1468 VDD.n1037 VDD.n1036 26.38
R1469 VDD.n962 VDD.n960 26.38
R1470 VDD.n962 VDD.n959 26.38
R1471 VDD.n962 VDD.n961 26.38
R1472 VDD.n811 VDD.n809 26.38
R1473 VDD.n811 VDD.n808 26.38
R1474 VDD.n811 VDD.n810 26.38
R1475 VDD.n887 VDD.n886 26.38
R1476 VDD.n887 VDD.n882 26.38
R1477 VDD.n887 VDD.n880 26.38
R1478 VDD.n887 VDD.n879 26.38
R1479 VDD.n814 VDD.n806 22.915
R1480 VDD.n23 VDD.n14 22.915
R1481 VDD.n73  20.457
R1482 VDD.n137 VDD.t94 20.457
R1483 VDD.n180  20.457
R1484 VDD.n84  17.9
R1485 VDD.n126  17.9
R1486 VDD.n193 �eh�9V 17.9
R1487 VDD.n244 ����9V 15.343
R1488 VDD.n319  15.343
R1489 VDD.n394 VDD.t171 15.343
R1490 VDD.n469 ���9V 15.343
R1491 VDD.n544 ��ϝ9V 15.343
R1492 VDD.n619 �+�إ 15.343
R1493 VDD.n694 ��9V 15.343
R1494 VDD.n769 б��9V 15.343
R1495 VDD.n1519  15.343
R1496 VDD.n1444 �M��9V 15.343
R1497 VDD.n1369  15.343
R1498 VDD.n1294  15.343
R1499 VDD.n1219  15.343
R1500 VDD.n1144 0�ǝ9V 15.343
R1501 VDD.n1069 VDD.t149 15.343
R1502 VDD.n994  15.343
R1503 VDD.n919 VDD.t72 15.343
R1504 VDD.n843 VDD.t70 15.343
R1505 VDD.n806 VDD.n804 14.864
R1506 VDD.n804 VDD.n802 14.864
R1507 VDD.n802 VDD.n800 14.864
R1508 VDD.n800 VDD.n798 14.864
R1509 VDD.n798 VDD.n796 14.864
R1510 VDD.n955 VDD.n953 14.864
R1511 VDD.n953 VDD.n951 14.864
R1512 VDD.n951 VDD.n949 14.864
R1513 VDD.n949 VDD.n947 14.864
R1514 VDD.n947 VDD.n945 14.864
R1515 VDD.n1030 VDD.n1028 14.864
R1516 VDD.n1028 VDD.n1026 14.864
R1517 VDD.n1026 VDD.n1024 14.864
R1518 VDD.n1024 VDD.n1022 14.864
R1519 VDD.n1022 VDD.n1020 14.864
R1520 VDD.n1105 VDD.n1103 14.864
R1521 VDD.n1103 VDD.n1101 14.864
R1522 VDD.n1101 VDD.n1099 14.864
R1523 VDD.n1099 VDD.n1097 14.864
R1524 VDD.n1097 VDD.n1095 14.864
R1525 VDD.n1180 VDD.n1178 14.864
R1526 VDD.n1178 VDD.n1176 14.864
R1527 VDD.n1176 VDD.n1174 14.864
R1528 VDD.n1174 VDD.n1172 14.864
R1529 VDD.n1172 VDD.n1170 14.864
R1530 VDD.n1255 VDD.n1253 14.864
R1531 VDD.n1253 VDD.n1251 14.864
R1532 VDD.n1251 VDD.n1249 14.864
R1533 VDD.n1249 VDD.n1247 14.864
R1534 VDD.n1247 VDD.n1245 14.864
R1535 VDD.n1330 VDD.n1328 14.864
R1536 VDD.n1328 VDD.n1326 14.864
R1537 VDD.n1326 VDD.n1324 14.864
R1538 VDD.n1324 VDD.n1322 14.864
R1539 VDD.n1322 VDD.n1320 14.864
R1540 VDD.n1405 VDD.n1403 14.864
R1541 VDD.n1403 VDD.n1401 14.864
R1542 VDD.n1401 VDD.n1399 14.864
R1543 VDD.n1399 VDD.n1397 14.864
R1544 VDD.n1397 VDD.n1395 14.864
R1545 VDD.n1480 VDD.n1478 14.864
R1546 VDD.n1478 VDD.n1476 14.864
R1547 VDD.n1476 VDD.n1474 14.864
R1548 VDD.n1474 VDD.n1472 14.864
R1549 VDD.n1472 VDD.n1470 14.864
R1550 VDD.n1555 VDD.n1553 14.864
R1551 VDD.n1553 VDD.n1551 14.864
R1552 VDD.n1551 VDD.n1549 14.864
R1553 VDD.n1549 VDD.n1547 14.864
R1554 VDD.n1547 VDD.n1545 14.864
R1555 VDD.n745 VDD.n743 14.864
R1556 VDD.n743 VDD.n741 14.864
R1557 VDD.n741 VDD.n739 14.864
R1558 VDD.n739 VDD.n737 14.864
R1559 VDD.n737 VDD.n735 14.864
R1560 VDD.n670 VDD.n668 14.864
R1561 VDD.n668 VDD.n666 14.864
R1562 VDD.n666 VDD.n664 14.864
R1563 VDD.n664 VDD.n662 14.864
R1564 VDD.n662 VDD.n660 14.864
R1565 VDD.n595 VDD.n593 14.864
R1566 VDD.n593 VDD.n591 14.864
R1567 VDD.n591 VDD.n589 14.864
R1568 VDD.n589 VDD.n587 14.864
R1569 VDD.n587 VDD.n585 14.864
R1570 VDD.n520 VDD.n518 14.864
R1571 VDD.n518 VDD.n516 14.864
R1572 VDD.n516 VDD.n514 14.864
R1573 VDD.n514 VDD.n512 14.864
R1574 VDD.n512 VDD.n510 14.864
R1575 VDD.n445 VDD.n443 14.864
R1576 VDD.n443 VDD.n441 14.864
R1577 VDD.n441 VDD.n439 14.864
R1578 VDD.n439 VDD.n437 14.864
R1579 VDD.n437 VDD.n435 14.864
R1580 VDD.n370 VDD.n368 14.864
R1581 VDD.n368 VDD.n366 14.864
R1582 VDD.n366 VDD.n364 14.864
R1583 VDD.n364 VDD.n362 14.864
R1584 VDD.n362 VDD.n360 14.864
R1585 VDD.n295 VDD.n293 14.864
R1586 VDD.n293 VDD.n291 14.864
R1587 VDD.n291 VDD.n289 14.864
R1588 VDD.n289 VDD.n287 14.864
R1589 VDD.n287 VDD.n285 14.864
R1590 VDD.n220 VDD.n218 14.864
R1591 VDD.n218 VDD.n216 14.864
R1592 VDD.n216 VDD.n214 14.864
R1593 VDD.n214 VDD.n212 14.864
R1594 VDD.n212 VDD.n210 14.864
R1595 VDD.n163 VDD.n161 14.864
R1596 VDD.n161 VDD.n159 14.864
R1597 VDD.n159 VDD.n157 14.864
R1598 VDD.n157 VDD.n155 14.864
R1599 VDD.n155 VDD.n153 14.864
R1600 VDD.n110 VDD.n108 14.864
R1601 VDD.n108 VDD.n106 14.864
R1602 VDD.n106 VDD.n104 14.864
R1603 VDD.n104 VDD.n102 14.864
R1604 VDD.n102 VDD.n100 14.864
R1605 VDD.n53 VDD.n51 14.864
R1606 VDD.n51 VDD.n49 14.864
R1607 VDD.n49 VDD.n47 14.864
R1608 VDD.n47 VDD.n45 14.864
R1609 VDD.n45 VDD.n43 14.864
R1610 VDD.n43 VDD.n42 14.864
R1611 VDD.n876 VDD.n874 14.864
R1612 VDD.n874 VDD.n872 14.864
R1613 VDD.n872 VDD.n870 14.864
R1614 VDD.n870 VDD.n868 14.864
R1615 VDD.n868 VDD.n866 14.864
R1616 VDD.n866 VDD.n865 14.864
R1617 VDD.n14 VDD.n13 14.864
R1618 VDD.n13 VDD.n11 14.864
R1619 VDD.n11 VDD.n9 14.864
R1620 VDD.n9 VDD.n7 14.864
R1621 VDD.n7 VDD.n5 14.864
R1622 VDD.n67 VDD.n54 14.864
R1623 VDD.n120 VDD.n111 14.864
R1624 VDD.n173 VDD.n164 14.864
R1625 VDD.n230 VDD.n221 14.864
R1626 VDD.n305 VDD.n296 14.864
R1627 VDD.n380 VDD.n371 14.864
R1628 VDD.n455 VDD.n446 14.864
R1629 VDD.n530 VDD.n521 14.864
R1630 VDD.n605 VDD.n596 14.864
R1631 VDD.n680 VDD.n671 14.864
R1632 VDD.n755 VDD.n746 14.864
R1633 VDD.n1565 VDD.n1556 14.864
R1634 VDD.n1490 VDD.n1481 14.864
R1635 VDD.n1415 VDD.n1406 14.864
R1636 VDD.n1340 VDD.n1331 14.864
R1637 VDD.n1265 VDD.n1256 14.864
R1638 VDD.n1190 VDD.n1181 14.864
R1639 VDD.n1115 VDD.n1106 14.864
R1640 VDD.n1040 VDD.n1031 14.864
R1641 VDD.n965 VDD.n956 14.864
R1642 VDD.n890 VDD.n877 14.864
R1643 VDD.n829 VDD.t152 14.282
R1644 VDD.n829 VDD.t114 14.282
R1645 VDD.n845 VDD.t71 14.282
R1646 VDD.n845 VDD.t170 14.282
R1647 VDD.n905 VDD.t69 14.282
R1648 VDD.n905 VDD.t5 14.282
R1649 VDD.n921 VDD.t73 14.282
R1650 VDD.n921 VDD.t213 14.282
R1651 VDD.n980 VDD.t26 14.282
R1652 VDD.n980 VDD.t188 14.282
R1653 VDD.n996 VDD.t100 14.282
R1654 VDD.n996 VDD.t108 14.282
R1655 VDD.n1055 VDD.t180 14.282
R1656 VDD.n1055 VDD.t3 14.282
R1657 VDD.n1071 VDD.t150 14.282
R1658 VDD.n1071 VDD.t46 14.282
R1659 VDD.n1130 VDD.t166 14.282
R1660 VDD.n1130 VDD.t14 14.282
R1661 VDD.n1146 VDD.t110 14.282
R1662 VDD.n1146 VDD.t148 14.282
R1663 VDD.n1205 VDD.t81 14.282
R1664 VDD.n1205 VDD.t126 14.282
R1665 VDD.n1221 VDD.t192 14.282
R1666 VDD.n1221 VDD.t223 14.282
R1667 VDD.n1280 VDD.t144 14.282
R1668 VDD.n1280 VDD.t136 14.282
R1669 VDD.n1296 VDD.t88 14.282
R1670 VDD.n1296 VDD.t164 14.282
R1671 VDD.n1355 VDD.t32 14.282
R1672 VDD.n1355 VDD.t52 14.282
R1673 VDD.n1371 VDD.t50 14.282
R1674 VDD.n1371 VDD.t178 14.282
R1675 VDD.n1430 VDD.t186 14.282
R1676 VDD.n1430 VDD.t98 14.282
R1677 VDD.n1446 VDD.t38 14.282
R1678 VDD.n1446 VDD.t85 14.282
R1679 VDD.n1505 VDD.t67 14.282
R1680 VDD.n1505 VDD.t128 14.282
R1681 VDD.n1521 VDD.t142 14.282
R1682 VDD.n1521 VDD.t120 14.282
R1683 VDD.n783 VDD.t160 14.282
R1684 VDD.n783 VDD.t9 14.282
R1685 VDD.n771 VDD.t42 14.282
R1686 VDD.n771 VDD.t174 14.282
R1687 VDD.n708 VDD.t93 14.282
R1688 VDD.n708 VDD.t215 14.282
R1689 VDD.n696 VDD.t56 14.282
R1690 VDD.n696 VDD.t59 14.282
R1691 VDD.n633 VDD.t154 14.282
R1692 VDD.n633 VDD.t116 14.282
R1693 VDD.n621 VDD.t102 14.282
R1694 VDD.n621 VDD.t158 14.282
R1695 VDD.n558 VDD.t65 14.282
R1696 VDD.n558 VDD.t77 14.282
R1697 VDD.n546 VDD.t225 14.282
R1698 VDD.n546 VDD.t24 14.282
R1699 VDD.n483 VDD.t1 14.282
R1700 VDD.n483 VDD.t203 14.282
R1701 VDD.n471 VDD.t227 14.282
R1702 VDD.n471 VDD.t61 14.282
R1703 VDD.n408 VDD.t63 14.282
R1704 VDD.n408 VDD.t40 14.282
R1705 VDD.n396 VDD.t172 14.282
R1706 VDD.n396 VDD.t96 14.282
R1707 VDD.n333 VDD.t162 14.282
R1708 VDD.n333 VDD.t201 14.282
R1709 VDD.n321 VDD.t20 14.282
R1710 VDD.n321 VDD.t176 14.282
R1711 VDD.n258 VDD.t209 14.282
R1712 VDD.n258 VDD.t138 14.282
R1713 VDD.n246 VDD.t231 14.282
R1714 VDD.n246 VDD.t219 14.282
R1715 VDD.n184 VDD.t182 14.282
R1716 VDD.n184 VDD.t83 14.282
R1717 VDD.n260 �Ӵ�9V 12.786
R1718 VDD.n335  12.786
R1719 VDD.n410  12.786
R1720 VDD.n485 ��i�9V 12.786
R1721 VDD.n560  12.786
R1722 VDD.n635  12.786
R1723 VDD.n710 `�i�9V 12.786
R1724 VDD.n785 �ઝ9V 12.786
R1725 VDD.n1507 ��˞9V 12.786
R1726 VDD.n1432 P[��9V 12.786
R1727 VDD.n1357  12.786
R1728 VDD.n1282  12.786
R1729 VDD.n1207 `h�9V 12.786
R1730 VDD.n1132  12.786
R1731 VDD.n1057  12.786
R1732 VDD.n982 ��ѝ9V 12.786
R1733 VDD.n907 �i�9V 12.786
R1734 VDD.n831  12.786
R1735 VDD.n187 VDD.n185 9.083
R1736 VDD.n23 VDD.n22 8.855
R1737 VDD.n22 VDD.n21 8.855
R1738 VDD.n27 VDD.n26 8.855
R1739 VDD.n26 VDD.n25 8.855
R1740 VDD.n31 VDD.n30 8.855
R1741 VDD.n30 VDD.n29 8.855
R1742 VDD.n36 VDD.n34 8.855
R1743 VDD.n34 VDD.n33 8.855
R1744 VDD.n40 VDD.n39 8.855
R1745 VDD.n39 VDD.n38 8.855
R1746 VDD.n67 VDD.n66 8.855
R1747 VDD.n66 VDD.n65 8.855
R1748 VDD.n71 VDD.n70 8.855
R1749 VDD.n70 VDD.n69 8.855
R1750 VDD.n75 VDD.n74 8.855
R1751 VDD.n74 VDD.n73 8.855
R1752 VDD.n78 VDD.n77 8.855
R1753 VDD.n77 ��x�9V 8.855
R1754 VDD.n82 VDD.n81 8.855
R1755 VDD.n81 VDD.n80 8.855
R1756 VDD.n86 VDD.n85 8.855
R1757 VDD.n85 VDD.n84 8.855
R1758 VDD.n90 VDD.n89 8.855
R1759 VDD.n89 VDD.n88 8.855
R1760 VDD.n94 VDD.n93 8.855
R1761 VDD.n93 VDD.n92 8.855
R1762 VDD.n120 VDD.n119 8.855
R1763 VDD.n119 VDD.n118 8.855
R1764 VDD.n124 VDD.n123 8.855
R1765 VDD.n123 VDD.n122 8.855
R1766 VDD.n128 VDD.n127 8.855
R1767 VDD.n127 VDD.n126 8.855
R1768 VDD.n132 VDD.n131 8.855
R1769 VDD.n131 VDD.n130 8.855
R1770 VDD.n135 VDD.n134 8.855
R1771 VDD.n134  8.855
R1772 VDD.n139 VDD.n138 8.855
R1773 VDD.n138 VDD.n137 8.855
R1774 VDD.n143 VDD.n142 8.855
R1775 VDD.n142 VDD.n141 8.855
R1776 VDD.n147 VDD.n146 8.855
R1777 VDD.n146 VDD.n145 8.855
R1778 VDD.n173 VDD.n172 8.855
R1779 VDD.n172 VDD.n171 8.855
R1780 VDD.n178 VDD.n177 8.855
R1781 VDD.n177 VDD.n176 8.855
R1782 VDD.n182 VDD.n181 8.855
R1783 VDD.n181 VDD.n180 8.855
R1784 VDD.n187 VDD.n186 8.855
R1785 VDD.n186 �+��9V 8.855
R1786 VDD.n191 VDD.n190 8.855
R1787 VDD.n190 VDD.n189 8.855
R1788 VDD.n195 VDD.n194 8.855
R1789 VDD.n194 VDD.n193 8.855
R1790 VDD.n200 VDD.n199 8.855
R1791 VDD.n199 VDD.n198 8.855
R1792 VDD.n204 VDD.n203 8.855
R1793 VDD.n203 VDD.n202 8.855
R1794 VDD.n230 VDD.n229 8.855
R1795 VDD.n229 VDD.n228 8.855
R1796 VDD.n234 VDD.n233 8.855
R1797 VDD.n233 VDD.n232 8.855
R1798 VDD.n238 VDD.n237 8.855
R1799 VDD.n237 VDD.n236 8.855
R1800 VDD.n242 VDD.n241 8.855
R1801 VDD.n241 VDD.n240 8.855
R1802 VDD.n248 VDD.n245 8.855
R1803 VDD.n245 VDD.n244 8.855
R1804 VDD.n252 VDD.n251 8.855
R1805 VDD.n251 VDD.n250 8.855
R1806 VDD.n256 VDD.n255 8.855
R1807 VDD.n255 VDD.n254 8.855
R1808 VDD.n262 VDD.n261 8.855
R1809 VDD.n261 VDD.n260 8.855
R1810 VDD.n266 VDD.n265 8.855
R1811 VDD.n265 VDD.n264 8.855
R1812 VDD.n271 VDD.n270 8.855
R1813 VDD.n270 VDD.n269 8.855
R1814 VDD.n275 VDD.n274 8.855
R1815 VDD.n274 VDD.n273 8.855
R1816 VDD.n279 VDD.n278 8.855
R1817 VDD.n278 VDD.n277 8.855
R1818 VDD.n305 VDD.n304 8.855
R1819 VDD.n304 VDD.n303 8.855
R1820 VDD.n309 VDD.n308 8.855
R1821 VDD.n308 VDD.n307 8.855
R1822 VDD.n313 VDD.n312 8.855
R1823 VDD.n312 VDD.n311 8.855
R1824 VDD.n317 VDD.n316 8.855
R1825 VDD.n316 VDD.n315 8.855
R1826 VDD.n323 VDD.n320 8.855
R1827 VDD.n320 VDD.n319 8.855
R1828 VDD.n327 VDD.n326 8.855
R1829 VDD.n326 VDD.n325 8.855
R1830 VDD.n331 VDD.n330 8.855
R1831 VDD.n330 VDD.n329 8.855
R1832 VDD.n337 VDD.n336 8.855
R1833 VDD.n336 VDD.n335 8.855
R1834 VDD.n341 VDD.n340 8.855
R1835 VDD.n340 VDD.n339 8.855
R1836 VDD.n346 VDD.n345 8.855
R1837 VDD.n345 VDD.n344 8.855
R1838 VDD.n350 VDD.n349 8.855
R1839 VDD.n349 VDD.n348 8.855
R1840 VDD.n354 VDD.n353 8.855
R1841 VDD.n353 VDD.n352 8.855
R1842 VDD.n380 VDD.n379 8.855
R1843 VDD.n379 VDD.n378 8.855
R1844 VDD.n384 VDD.n383 8.855
R1845 VDD.n383 VDD.n382 8.855
R1846 VDD.n388 VDD.n387 8.855
R1847 VDD.n387 VDD.n386 8.855
R1848 VDD.n392 VDD.n391 8.855
R1849 VDD.n391 VDD.n390 8.855
R1850 VDD.n398 VDD.n395 8.855
R1851 VDD.n395 VDD.n394 8.855
R1852 VDD.n402 VDD.n401 8.855
R1853 VDD.n401 VDD.n400 8.855
R1854 VDD.n406 VDD.n405 8.855
R1855 VDD.n405 VDD.n404 8.855
R1856 VDD.n412 VDD.n411 8.855
R1857 VDD.n411 VDD.n410 8.855
R1858 VDD.n416 VDD.n415 8.855
R1859 VDD.n415 VDD.n414 8.855
R1860 VDD.n421 VDD.n420 8.855
R1861 VDD.n420 VDD.n419 8.855
R1862 VDD.n425 VDD.n424 8.855
R1863 VDD.n424 VDD.n423 8.855
R1864 VDD.n429 VDD.n428 8.855
R1865 VDD.n428 VDD.n427 8.855
R1866 VDD.n455 VDD.n454 8.855
R1867 VDD.n454 VDD.n453 8.855
R1868 VDD.n459 VDD.n458 8.855
R1869 VDD.n458 VDD.n457 8.855
R1870 VDD.n463 VDD.n462 8.855
R1871 VDD.n462 VDD.n461 8.855
R1872 VDD.n467 VDD.n466 8.855
R1873 VDD.n466 VDD.n465 8.855
R1874 VDD.n473 VDD.n470 8.855
R1875 VDD.n470 VDD.n469 8.855
R1876 VDD.n477 VDD.n476 8.855
R1877 VDD.n476 VDD.n475 8.855
R1878 VDD.n481 VDD.n480 8.855
R1879 VDD.n480 VDD.n479 8.855
R1880 VDD.n487 VDD.n486 8.855
R1881 VDD.n486 VDD.n485 8.855
R1882 VDD.n491 VDD.n490 8.855
R1883 VDD.n490 VDD.n489 8.855
R1884 VDD.n496 VDD.n495 8.855
R1885 VDD.n495 VDD.n494 8.855
R1886 VDD.n500 VDD.n499 8.855
R1887 VDD.n499 VDD.n498 8.855
R1888 VDD.n504 VDD.n503 8.855
R1889 VDD.n503 VDD.n502 8.855
R1890 VDD.n530 VDD.n529 8.855
R1891 VDD.n529 VDD.n528 8.855
R1892 VDD.n534 VDD.n533 8.855
R1893 VDD.n533 VDD.n532 8.855
R1894 VDD.n538 VDD.n537 8.855
R1895 VDD.n537 VDD.n536 8.855
R1896 VDD.n542 VDD.n541 8.855
R1897 VDD.n541 VDD.n540 8.855
R1898 VDD.n548 VDD.n545 8.855
R1899 VDD.n545 VDD.n544 8.855
R1900 VDD.n552 VDD.n551 8.855
R1901 VDD.n551 VDD.n550 8.855
R1902 VDD.n556 VDD.n555 8.855
R1903 VDD.n555 VDD.n554 8.855
R1904 VDD.n562 VDD.n561 8.855
R1905 VDD.n561 VDD.n560 8.855
R1906 VDD.n566 VDD.n565 8.855
R1907 VDD.n565 VDD.n564 8.855
R1908 VDD.n571 VDD.n570 8.855
R1909 VDD.n570 VDD.n569 8.855
R1910 VDD.n575 VDD.n574 8.855
R1911 VDD.n574 VDD.n573 8.855
R1912 VDD.n579 VDD.n578 8.855
R1913 VDD.n578 VDD.n577 8.855
R1914 VDD.n605 VDD.n604 8.855
R1915 VDD.n604 VDD.n603 8.855
R1916 VDD.n609 VDD.n608 8.855
R1917 VDD.n608 VDD.n607 8.855
R1918 VDD.n613 VDD.n612 8.855
R1919 VDD.n612 VDD.n611 8.855
R1920 VDD.n617 VDD.n616 8.855
R1921 VDD.n616 VDD.n615 8.855
R1922 VDD.n623 VDD.n620 8.855
R1923 VDD.n620 VDD.n619 8.855
R1924 VDD.n627 VDD.n626 8.855
R1925 VDD.n626 VDD.n625 8.855
R1926 VDD.n631 VDD.n630 8.855
R1927 VDD.n630 VDD.n629 8.855
R1928 VDD.n637 VDD.n636 8.855
R1929 VDD.n636 VDD.n635 8.855
R1930 VDD.n641 VDD.n640 8.855
R1931 VDD.n640 VDD.n639 8.855
R1932 VDD.n646 VDD.n645 8.855
R1933 VDD.n645 VDD.n644 8.855
R1934 VDD.n650 VDD.n649 8.855
R1935 VDD.n649 VDD.n648 8.855
R1936 VDD.n654 VDD.n653 8.855
R1937 VDD.n653 VDD.n652 8.855
R1938 VDD.n680 VDD.n679 8.855
R1939 VDD.n679 VDD.n678 8.855
R1940 VDD.n684 VDD.n683 8.855
R1941 VDD.n683 VDD.n682 8.855
R1942 VDD.n688 VDD.n687 8.855
R1943 VDD.n687 VDD.n686 8.855
R1944 VDD.n692 VDD.n691 8.855
R1945 VDD.n691 VDD.n690 8.855
R1946 VDD.n698 VDD.n695 8.855
R1947 VDD.n695 VDD.n694 8.855
R1948 VDD.n702 VDD.n701 8.855
R1949 VDD.n701 VDD.n700 8.855
R1950 VDD.n706 VDD.n705 8.855
R1951 VDD.n705 VDD.n704 8.855
R1952 VDD.n712 VDD.n711 8.855
R1953 VDD.n711 VDD.n710 8.855
R1954 VDD.n716 VDD.n715 8.855
R1955 VDD.n715 VDD.n714 8.855
R1956 VDD.n721 VDD.n720 8.855
R1957 VDD.n720 VDD.n719 8.855
R1958 VDD.n725 VDD.n724 8.855
R1959 VDD.n724 VDD.n723 8.855
R1960 VDD.n729 VDD.n728 8.855
R1961 VDD.n728 VDD.n727 8.855
R1962 VDD.n755 VDD.n754 8.855
R1963 VDD.n754 VDD.n753 8.855
R1964 VDD.n759 VDD.n758 8.855
R1965 VDD.n758 VDD.n757 8.855
R1966 VDD.n763 VDD.n762 8.855
R1967 VDD.n762 VDD.n761 8.855
R1968 VDD.n767 VDD.n766 8.855
R1969 VDD.n766 VDD.n765 8.855
R1970 VDD.n773 VDD.n770 8.855
R1971 VDD.n770 VDD.n769 8.855
R1972 VDD.n777 VDD.n776 8.855
R1973 VDD.n776 VDD.n775 8.855
R1974 VDD.n781 VDD.n780 8.855
R1975 VDD.n780 VDD.n779 8.855
R1976 VDD.n787 VDD.n786 8.855
R1977 VDD.n786 VDD.n785 8.855
R1978 VDD.n791 VDD.n790 8.855
R1979 VDD.n790 VDD.n789 8.855
R1980 VDD.n1574 VDD.n1573 8.855
R1981 VDD.n1573 VDD.n1572 8.855
R1982 VDD.n1569 VDD.n1568 8.855
R1983 VDD.n1568 VDD.n1567 8.855
R1984 VDD.n1565 VDD.n1564 8.855
R1985 VDD.n1564 VDD.n1563 8.855
R1986 VDD.n1539 VDD.n1538 8.855
R1987 VDD.n1538 VDD.n1537 8.855
R1988 VDD.n1535 VDD.n1534 8.855
R1989 VDD.n1534 VDD.n1533 8.855
R1990 VDD.n1531 VDD.n1530 8.855
R1991 VDD.n1530 VDD.n1529 8.855
R1992 VDD.n1527 VDD.n1526 8.855
R1993 VDD.n1526 VDD.n1525 8.855
R1994 VDD.n1523 VDD.n1520 8.855
R1995 VDD.n1520 VDD.n1519 8.855
R1996 VDD.n1517 VDD.n1516 8.855
R1997 VDD.n1516 VDD.n1515 8.855
R1998 VDD.n1513 VDD.n1512 8.855
R1999 VDD.n1512 VDD.n1511 8.855
R2000 VDD.n1509 VDD.n1508 8.855
R2001 VDD.n1508 VDD.n1507 8.855
R2002 VDD.n1503 VDD.n1502 8.855
R2003 VDD.n1502 VDD.n1501 8.855
R2004 VDD.n1499 VDD.n1498 8.855
R2005 VDD.n1498 VDD.n1497 8.855
R2006 VDD.n1494 VDD.n1493 8.855
R2007 VDD.n1493 VDD.n1492 8.855
R2008 VDD.n1490 VDD.n1489 8.855
R2009 VDD.n1489 VDD.n1488 8.855
R2010 VDD.n1464 VDD.n1463 8.855
R2011 VDD.n1463 VDD.n1462 8.855
R2012 VDD.n1460 VDD.n1459 8.855
R2013 VDD.n1459 VDD.n1458 8.855
R2014 VDD.n1456 VDD.n1455 8.855
R2015 VDD.n1455 VDD.n1454 8.855
R2016 VDD.n1452 VDD.n1451 8.855
R2017 VDD.n1451 VDD.n1450 8.855
R2018 VDD.n1448 VDD.n1445 8.855
R2019 VDD.n1445 VDD.n1444 8.855
R2020 VDD.n1442 VDD.n1441 8.855
R2021 VDD.n1441 VDD.n1440 8.855
R2022 VDD.n1438 VDD.n1437 8.855
R2023 VDD.n1437 VDD.n1436 8.855
R2024 VDD.n1434 VDD.n1433 8.855
R2025 VDD.n1433 VDD.n1432 8.855
R2026 VDD.n1428 VDD.n1427 8.855
R2027 VDD.n1427 VDD.n1426 8.855
R2028 VDD.n1424 VDD.n1423 8.855
R2029 VDD.n1423 VDD.n1422 8.855
R2030 VDD.n1419 VDD.n1418 8.855
R2031 VDD.n1418 VDD.n1417 8.855
R2032 VDD.n1415 VDD.n1414 8.855
R2033 VDD.n1414 VDD.n1413 8.855
R2034 VDD.n1389 VDD.n1388 8.855
R2035 VDD.n1388 VDD.n1387 8.855
R2036 VDD.n1385 VDD.n1384 8.855
R2037 VDD.n1384 VDD.n1383 8.855
R2038 VDD.n1381 VDD.n1380 8.855
R2039 VDD.n1380 VDD.n1379 8.855
R2040 VDD.n1377 VDD.n1376 8.855
R2041 VDD.n1376 VDD.n1375 8.855
R2042 VDD.n1373 VDD.n1370 8.855
R2043 VDD.n1370 VDD.n1369 8.855
R2044 VDD.n1367 VDD.n1366 8.855
R2045 VDD.n1366 VDD.n1365 8.855
R2046 VDD.n1363 VDD.n1362 8.855
R2047 VDD.n1362 VDD.n1361 8.855
R2048 VDD.n1359 VDD.n1358 8.855
R2049 VDD.n1358 VDD.n1357 8.855
R2050 VDD.n1353 VDD.n1352 8.855
R2051 VDD.n1352 VDD.n1351 8.855
R2052 VDD.n1349 VDD.n1348 8.855
R2053 VDD.n1348 VDD.n1347 8.855
R2054 VDD.n1344 VDD.n1343 8.855
R2055 VDD.n1343 VDD.n1342 8.855
R2056 VDD.n1340 VDD.n1339 8.855
R2057 VDD.n1339 VDD.n1338 8.855
R2058 VDD.n1314 VDD.n1313 8.855
R2059 VDD.n1313 VDD.n1312 8.855
R2060 VDD.n1310 VDD.n1309 8.855
R2061 VDD.n1309 VDD.n1308 8.855
R2062 VDD.n1306 VDD.n1305 8.855
R2063 VDD.n1305 VDD.n1304 8.855
R2064 VDD.n1302 VDD.n1301 8.855
R2065 VDD.n1301 VDD.n1300 8.855
R2066 VDD.n1298 VDD.n1295 8.855
R2067 VDD.n1295 VDD.n1294 8.855
R2068 VDD.n1292 VDD.n1291 8.855
R2069 VDD.n1291 VDD.n1290 8.855
R2070 VDD.n1288 VDD.n1287 8.855
R2071 VDD.n1287 VDD.n1286 8.855
R2072 VDD.n1284 VDD.n1283 8.855
R2073 VDD.n1283 VDD.n1282 8.855
R2074 VDD.n1278 VDD.n1277 8.855
R2075 VDD.n1277 VDD.n1276 8.855
R2076 VDD.n1274 VDD.n1273 8.855
R2077 VDD.n1273 VDD.n1272 8.855
R2078 VDD.n1269 VDD.n1268 8.855
R2079 VDD.n1268 VDD.n1267 8.855
R2080 VDD.n1265 VDD.n1264 8.855
R2081 VDD.n1264 VDD.n1263 8.855
R2082 VDD.n1239 VDD.n1238 8.855
R2083 VDD.n1238 VDD.n1237 8.855
R2084 VDD.n1235 VDD.n1234 8.855
R2085 VDD.n1234 VDD.n1233 8.855
R2086 VDD.n1231 VDD.n1230 8.855
R2087 VDD.n1230 VDD.n1229 8.855
R2088 VDD.n1227 VDD.n1226 8.855
R2089 VDD.n1226 VDD.n1225 8.855
R2090 VDD.n1223 VDD.n1220 8.855
R2091 VDD.n1220 VDD.n1219 8.855
R2092 VDD.n1217 VDD.n1216 8.855
R2093 VDD.n1216 VDD.n1215 8.855
R2094 VDD.n1213 VDD.n1212 8.855
R2095 VDD.n1212 VDD.n1211 8.855
R2096 VDD.n1209 VDD.n1208 8.855
R2097 VDD.n1208 VDD.n1207 8.855
R2098 VDD.n1203 VDD.n1202 8.855
R2099 VDD.n1202 VDD.n1201 8.855
R2100 VDD.n1199 VDD.n1198 8.855
R2101 VDD.n1198 VDD.n1197 8.855
R2102 VDD.n1194 VDD.n1193 8.855
R2103 VDD.n1193 VDD.n1192 8.855
R2104 VDD.n1190 VDD.n1189 8.855
R2105 VDD.n1189 VDD.n1188 8.855
R2106 VDD.n1164 VDD.n1163 8.855
R2107 VDD.n1163 VDD.n1162 8.855
R2108 VDD.n1160 VDD.n1159 8.855
R2109 VDD.n1159 VDD.n1158 8.855
R2110 VDD.n1156 VDD.n1155 8.855
R2111 VDD.n1155 VDD.n1154 8.855
R2112 VDD.n1152 VDD.n1151 8.855
R2113 VDD.n1151 VDD.n1150 8.855
R2114 VDD.n1148 VDD.n1145 8.855
R2115 VDD.n1145 VDD.n1144 8.855
R2116 VDD.n1142 VDD.n1141 8.855
R2117 VDD.n1141 VDD.n1140 8.855
R2118 VDD.n1138 VDD.n1137 8.855
R2119 VDD.n1137 VDD.n1136 8.855
R2120 VDD.n1134 VDD.n1133 8.855
R2121 VDD.n1133 VDD.n1132 8.855
R2122 VDD.n1128 VDD.n1127 8.855
R2123 VDD.n1127 VDD.n1126 8.855
R2124 VDD.n1124 VDD.n1123 8.855
R2125 VDD.n1123 VDD.n1122 8.855
R2126 VDD.n1119 VDD.n1118 8.855
R2127 VDD.n1118 VDD.n1117 8.855
R2128 VDD.n1115 VDD.n1114 8.855
R2129 VDD.n1114 VDD.n1113 8.855
R2130 VDD.n1089 VDD.n1088 8.855
R2131 VDD.n1088 VDD.n1087 8.855
R2132 VDD.n1085 VDD.n1084 8.855
R2133 VDD.n1084 VDD.n1083 8.855
R2134 VDD.n1081 VDD.n1080 8.855
R2135 VDD.n1080 VDD.n1079 8.855
R2136 VDD.n1077 VDD.n1076 8.855
R2137 VDD.n1076 VDD.n1075 8.855
R2138 VDD.n1073 VDD.n1070 8.855
R2139 VDD.n1070 VDD.n1069 8.855
R2140 VDD.n1067 VDD.n1066 8.855
R2141 VDD.n1066 VDD.n1065 8.855
R2142 VDD.n1063 VDD.n1062 8.855
R2143 VDD.n1062 VDD.n1061 8.855
R2144 VDD.n1059 VDD.n1058 8.855
R2145 VDD.n1058 VDD.n1057 8.855
R2146 VDD.n1053 VDD.n1052 8.855
R2147 VDD.n1052 VDD.n1051 8.855
R2148 VDD.n1049 VDD.n1048 8.855
R2149 VDD.n1048 VDD.n1047 8.855
R2150 VDD.n1044 VDD.n1043 8.855
R2151 VDD.n1043 VDD.n1042 8.855
R2152 VDD.n1040 VDD.n1039 8.855
R2153 VDD.n1039 VDD.n1038 8.855
R2154 VDD.n1014 VDD.n1013 8.855
R2155 VDD.n1013 VDD.n1012 8.855
R2156 VDD.n1010 VDD.n1009 8.855
R2157 VDD.n1009 VDD.n1008 8.855
R2158 VDD.n1006 VDD.n1005 8.855
R2159 VDD.n1005 VDD.n1004 8.855
R2160 VDD.n1002 VDD.n1001 8.855
R2161 VDD.n1001 VDD.n1000 8.855
R2162 VDD.n998 VDD.n995 8.855
R2163 VDD.n995 VDD.n994 8.855
R2164 VDD.n992 VDD.n991 8.855
R2165 VDD.n991 VDD.n990 8.855
R2166 VDD.n988 VDD.n987 8.855
R2167 VDD.n987 VDD.n986 8.855
R2168 VDD.n984 VDD.n983 8.855
R2169 VDD.n983 VDD.n982 8.855
R2170 VDD.n978 VDD.n977 8.855
R2171 VDD.n977 VDD.n976 8.855
R2172 VDD.n974 VDD.n973 8.855
R2173 VDD.n973 VDD.n972 8.855
R2174 VDD.n969 VDD.n968 8.855
R2175 VDD.n968 VDD.n967 8.855
R2176 VDD.n965 VDD.n964 8.855
R2177 VDD.n964 VDD.n963 8.855
R2178 VDD.n939 VDD.n938 8.855
R2179 VDD.n938 VDD.n937 8.855
R2180 VDD.n935 VDD.n934 8.855
R2181 VDD.n934 VDD.n933 8.855
R2182 VDD.n931 VDD.n930 8.855
R2183 VDD.n930 VDD.n929 8.855
R2184 VDD.n927 VDD.n926 8.855
R2185 VDD.n926 VDD.n925 8.855
R2186 VDD.n923 VDD.n920 8.855
R2187 VDD.n920 VDD.n919 8.855
R2188 VDD.n917 VDD.n916 8.855
R2189 VDD.n916 VDD.n915 8.855
R2190 VDD.n913 VDD.n912 8.855
R2191 VDD.n912 VDD.n911 8.855
R2192 VDD.n909 VDD.n908 8.855
R2193 VDD.n908 VDD.n907 8.855
R2194 VDD.n903 VDD.n902 8.855
R2195 VDD.n902 VDD.n901 8.855
R2196 VDD.n899 VDD.n898 8.855
R2197 VDD.n898 VDD.n897 8.855
R2198 VDD.n894 VDD.n893 8.855
R2199 VDD.n893 VDD.n892 8.855
R2200 VDD.n890 VDD.n889 8.855
R2201 VDD.n889 VDD.n888 8.855
R2202 VDD.n863 VDD.n862 8.855
R2203 VDD.n862 VDD.n861 8.855
R2204 VDD.n859 VDD.n858 8.855
R2205 VDD.n858 VDD.n857 8.855
R2206 VDD.n855 VDD.n854 8.855
R2207 VDD.n854 VDD.n853 8.855
R2208 VDD.n851 VDD.n850 8.855
R2209 VDD.n850 VDD.n849 8.855
R2210 VDD.n847 VDD.n844 8.855
R2211 VDD.n844 VDD.n843 8.855
R2212 VDD.n841 VDD.n840 8.855
R2213 VDD.n840 VDD.n839 8.855
R2214 VDD.n837 VDD.n836 8.855
R2215 VDD.n836 VDD.n835 8.855
R2216 VDD.n833 VDD.n832 8.855
R2217 VDD.n832 VDD.n831 8.855
R2218 VDD.n827 VDD.n826 8.855
R2219 VDD.n826 VDD.n825 8.855
R2220 VDD.n823 VDD.n822 8.855
R2221 VDD.n822 VDD.n821 8.855
R2222 VDD.n818 VDD.n817 8.855
R2223 VDD.n817 VDD.n816 8.855
R2224 VDD.n814 VDD.n813 8.855
R2225 VDD.n813 VDD.n812 8.855
R2226 VDD.n956 VDD.n955 8.051
R2227 VDD.n1031 VDD.n1030 8.051
R2228 VDD.n1106 VDD.n1105 8.051
R2229 VDD.n1181 VDD.n1180 8.051
R2230 VDD.n1256 VDD.n1255 8.051
R2231 VDD.n1331 VDD.n1330 8.051
R2232 VDD.n1406 VDD.n1405 8.051
R2233 VDD.n1481 VDD.n1480 8.051
R2234 VDD.n1556 VDD.n1555 8.051
R2235 VDD.n746 VDD.n745 8.051
R2236 VDD.n671 VDD.n670 8.051
R2237 VDD.n596 VDD.n595 8.051
R2238 VDD.n521 VDD.n520 8.051
R2239 VDD.n446 VDD.n445 8.051
R2240 VDD.n371 VDD.n370 8.051
R2241 VDD.n296 VDD.n295 8.051
R2242 VDD.n221 VDD.n220 8.051
R2243 VDD.n164 VDD.n163 8.051
R2244 VDD.n111 VDD.n110 8.051
R2245 VDD.n54 VDD.n53 8.051
R2246 VDD.n877 VDD.n876 8.051
R2247 VDD.n254 ��9V 7.671
R2248 VDD.n329 �b��9V 7.671
R2249 VDD.n404  7.671
R2250 VDD.n479 ��x�9V 7.671
R2251 VDD.n554  ���9V 7.671
R2252 VDD.n629 ��I�9V 7.671
R2253 VDD.n704 �+�إ 7.671
R2254 VDD.n779 VDD.t159 7.671
R2255 VDD.n1511 VDD.t66 7.671
R2256 VDD.n1436  7.671
R2257 VDD.n1361  7.671
R2258 VDD.n1286  7.671
R2259 VDD.n1211  7.671
R2260 VDD.n1136 �+�إ 7.671
R2261 VDD.n1061 �+�إ 7.671
R2262 VDD.n986 ���9V 7.671
R2263 VDD.n911 ��h�9V 7.671
R2264 VDD.n835 ���9V 7.671
R2265 VDD.n262 VDD.n259 7.019
R2266 VDD.n337 VDD.n334 7.019
R2267 VDD.n412 VDD.n409 7.019
R2268 VDD.n487 VDD.n484 7.019
R2269 VDD.n562 VDD.n559 7.019
R2270 VDD.n637 VDD.n634 7.019
R2271 VDD.n712 VDD.n709 7.019
R2272 VDD.n787 VDD.n784 7.019
R2273 VDD.n1509 VDD.n1506 7.019
R2274 VDD.n1434 VDD.n1431 7.019
R2275 VDD.n1359 VDD.n1356 7.019
R2276 VDD.n1284 VDD.n1281 7.019
R2277 VDD.n1209 VDD.n1206 7.019
R2278 VDD.n1134 VDD.n1131 7.019
R2279 VDD.n1059 VDD.n1056 7.019
R2280 VDD.n984 VDD.n981 7.019
R2281 VDD.n909 VDD.n906 7.019
R2282 VDD.n833 VDD.n830 7.019
R2283 VDD.n248 VDD.n247 6.606
R2284 VDD.n323 VDD.n322 6.606
R2285 VDD.n398 VDD.n397 6.606
R2286 VDD.n473 VDD.n472 6.606
R2287 VDD.n548 VDD.n547 6.606
R2288 VDD.n623 VDD.n622 6.606
R2289 VDD.n698 VDD.n697 6.606
R2290 VDD.n773 VDD.n772 6.606
R2291 VDD.n1523 VDD.n1522 6.606
R2292 VDD.n1448 VDD.n1447 6.606
R2293 VDD.n1373 VDD.n1372 6.606
R2294 VDD.n1298 VDD.n1297 6.606
R2295 VDD.n1223 VDD.n1222 6.606
R2296 VDD.n1148 VDD.n1147 6.606
R2297 VDD.n1073 VDD.n1072 6.606
R2298 VDD.n998 VDD.n997 6.606
R2299 VDD.n923 VDD.n922 6.606
R2300 VDD.n847 VDD.n846 6.606
R2301 VDD.n250  5.114
R2302 VDD.n325 ��{�9V 5.114
R2303 VDD.n400 �+�إ 5.114
R2304 VDD.n475 �J�9V 5.114
R2305 VDD.n550 p���9V 5.114
R2306 VDD.n625 �+�إ 5.114
R2307 VDD.n700  5.114
R2308 VDD.n775 �	6�9V 5.114
R2309 VDD.n1515 0�l�9V 5.114
R2310 VDD.n1440 �+�إ 5.114
R2311 VDD.n1365  5.114
R2312 VDD.n1290  w��9V 5.114
R2313 VDD.n1215  "��9V 5.114
R2314 VDD.n1140 �L�9V 5.114
R2315 VDD.n1065 VDD.t45 5.114
R2316 VDD.n990 @{�9V 5.114
R2317 VDD.n915 �AK�9V 5.114
R2318 VDD.n839 �+�إ 5.114
R2319 VDD.n28 VDD.n23 4.795
R2320 VDD.n28 VDD.n27 4.65
R2321 VDD.n32 VDD.n31 4.65
R2322 VDD.n37 VDD.n36 4.65
R2323 VDD.n41 VDD.n40 4.65
R2324 VDD.n68 VDD.n67 4.65
R2325 VDD.n72 VDD.n71 4.65
R2326 VDD.n76 VDD.n75 4.65
R2327 VDD.n79 VDD.n78 4.65
R2328 VDD.n83 VDD.n82 4.65
R2329 VDD.n87 VDD.n86 4.65
R2330 VDD.n91 VDD.n90 4.65
R2331 VDD.n95 VDD.n94 4.65
R2332 VDD.n121 VDD.n120 4.65
R2333 VDD.n125 VDD.n124 4.65
R2334 VDD.n129 VDD.n128 4.65
R2335 VDD.n133 VDD.n132 4.65
R2336 VDD.n136 VDD.n135 4.65
R2337 VDD.n140 VDD.n139 4.65
R2338 VDD.n144 VDD.n143 4.65
R2339 VDD.n148 VDD.n147 4.65
R2340 VDD.n174 VDD.n173 4.65
R2341 VDD.n179 VDD.n178 4.65
R2342 VDD.n183 VDD.n182 4.65
R2343 VDD.n188 VDD.n187 4.65
R2344 VDD.n192 VDD.n191 4.65
R2345 VDD.n196 VDD.n195 4.65
R2346 VDD.n201 VDD.n200 4.65
R2347 VDD.n205 VDD.n204 4.65
R2348 VDD.n231 VDD.n230 4.65
R2349 VDD.n235 VDD.n234 4.65
R2350 VDD.n239 VDD.n238 4.65
R2351 VDD.n243 VDD.n242 4.65
R2352 VDD.n249 VDD.n248 4.65
R2353 VDD.n253 VDD.n252 4.65
R2354 VDD.n257 VDD.n256 4.65
R2355 VDD.n263 VDD.n262 4.65
R2356 VDD.n267 VDD.n266 4.65
R2357 VDD.n272 VDD.n271 4.65
R2358 VDD.n276 VDD.n275 4.65
R2359 VDD.n280 VDD.n279 4.65
R2360 VDD.n306 VDD.n305 4.65
R2361 VDD.n310 VDD.n309 4.65
R2362 VDD.n314 VDD.n313 4.65
R2363 VDD.n318 VDD.n317 4.65
R2364 VDD.n324 VDD.n323 4.65
R2365 VDD.n328 VDD.n327 4.65
R2366 VDD.n332 VDD.n331 4.65
R2367 VDD.n338 VDD.n337 4.65
R2368 VDD.n342 VDD.n341 4.65
R2369 VDD.n347 VDD.n346 4.65
R2370 VDD.n351 VDD.n350 4.65
R2371 VDD.n355 VDD.n354 4.65
R2372 VDD.n381 VDD.n380 4.65
R2373 VDD.n385 VDD.n384 4.65
R2374 VDD.n389 VDD.n388 4.65
R2375 VDD.n393 VDD.n392 4.65
R2376 VDD.n399 VDD.n398 4.65
R2377 VDD.n403 VDD.n402 4.65
R2378 VDD.n407 VDD.n406 4.65
R2379 VDD.n413 VDD.n412 4.65
R2380 VDD.n417 VDD.n416 4.65
R2381 VDD.n422 VDD.n421 4.65
R2382 VDD.n426 VDD.n425 4.65
R2383 VDD.n430 VDD.n429 4.65
R2384 VDD.n456 VDD.n455 4.65
R2385 VDD.n460 VDD.n459 4.65
R2386 VDD.n464 VDD.n463 4.65
R2387 VDD.n468 VDD.n467 4.65
R2388 VDD.n474 VDD.n473 4.65
R2389 VDD.n478 VDD.n477 4.65
R2390 VDD.n482 VDD.n481 4.65
R2391 VDD.n488 VDD.n487 4.65
R2392 VDD.n492 VDD.n491 4.65
R2393 VDD.n497 VDD.n496 4.65
R2394 VDD.n501 VDD.n500 4.65
R2395 VDD.n505 VDD.n504 4.65
R2396 VDD.n531 VDD.n530 4.65
R2397 VDD.n535 VDD.n534 4.65
R2398 VDD.n539 VDD.n538 4.65
R2399 VDD.n543 VDD.n542 4.65
R2400 VDD.n549 VDD.n548 4.65
R2401 VDD.n553 VDD.n552 4.65
R2402 VDD.n557 VDD.n556 4.65
R2403 VDD.n563 VDD.n562 4.65
R2404 VDD.n567 VDD.n566 4.65
R2405 VDD.n572 VDD.n571 4.65
R2406 VDD.n576 VDD.n575 4.65
R2407 VDD.n580 VDD.n579 4.65
R2408 VDD.n606 VDD.n605 4.65
R2409 VDD.n610 VDD.n609 4.65
R2410 VDD.n614 VDD.n613 4.65
R2411 VDD.n618 VDD.n617 4.65
R2412 VDD.n624 VDD.n623 4.65
R2413 VDD.n628 VDD.n627 4.65
R2414 VDD.n632 VDD.n631 4.65
R2415 VDD.n638 VDD.n637 4.65
R2416 VDD.n642 VDD.n641 4.65
R2417 VDD.n647 VDD.n646 4.65
R2418 VDD.n651 VDD.n650 4.65
R2419 VDD.n655 VDD.n654 4.65
R2420 VDD.n681 VDD.n680 4.65
R2421 VDD.n685 VDD.n684 4.65
R2422 VDD.n689 VDD.n688 4.65
R2423 VDD.n693 VDD.n692 4.65
R2424 VDD.n699 VDD.n698 4.65
R2425 VDD.n703 VDD.n702 4.65
R2426 VDD.n707 VDD.n706 4.65
R2427 VDD.n713 VDD.n712 4.65
R2428 VDD.n717 VDD.n716 4.65
R2429 VDD.n722 VDD.n721 4.65
R2430 VDD.n726 VDD.n725 4.65
R2431 VDD.n730 VDD.n729 4.65
R2432 VDD.n756 VDD.n755 4.65
R2433 VDD.n760 VDD.n759 4.65
R2434 VDD.n764 VDD.n763 4.65
R2435 VDD.n768 VDD.n767 4.65
R2436 VDD.n774 VDD.n773 4.65
R2437 VDD.n778 VDD.n777 4.65
R2438 VDD.n782 VDD.n781 4.65
R2439 VDD.n788 VDD.n787 4.65
R2440 VDD.n792 VDD.n791 4.65
R2441 VDD.n1575 VDD.n1574 4.65
R2442 VDD.n1570 VDD.n1569 4.65
R2443 VDD.n1566 VDD.n1565 4.65
R2444 VDD.n1540 VDD.n1539 4.65
R2445 VDD.n1536 VDD.n1535 4.65
R2446 VDD.n1532 VDD.n1531 4.65
R2447 VDD.n1528 VDD.n1527 4.65
R2448 VDD.n1524 VDD.n1523 4.65
R2449 VDD.n1518 VDD.n1517 4.65
R2450 VDD.n1514 VDD.n1513 4.65
R2451 VDD.n1510 VDD.n1509 4.65
R2452 VDD.n1504 VDD.n1503 4.65
R2453 VDD.n1500 VDD.n1499 4.65
R2454 VDD.n1495 VDD.n1494 4.65
R2455 VDD.n1491 VDD.n1490 4.65
R2456 VDD.n1465 VDD.n1464 4.65
R2457 VDD.n1461 VDD.n1460 4.65
R2458 VDD.n1457 VDD.n1456 4.65
R2459 VDD.n1453 VDD.n1452 4.65
R2460 VDD.n1449 VDD.n1448 4.65
R2461 VDD.n1443 VDD.n1442 4.65
R2462 VDD.n1439 VDD.n1438 4.65
R2463 VDD.n1435 VDD.n1434 4.65
R2464 VDD.n1429 VDD.n1428 4.65
R2465 VDD.n1425 VDD.n1424 4.65
R2466 VDD.n1420 VDD.n1419 4.65
R2467 VDD.n1416 VDD.n1415 4.65
R2468 VDD.n1390 VDD.n1389 4.65
R2469 VDD.n1386 VDD.n1385 4.65
R2470 VDD.n1382 VDD.n1381 4.65
R2471 VDD.n1378 VDD.n1377 4.65
R2472 VDD.n1374 VDD.n1373 4.65
R2473 VDD.n1368 VDD.n1367 4.65
R2474 VDD.n1364 VDD.n1363 4.65
R2475 VDD.n1360 VDD.n1359 4.65
R2476 VDD.n1354 VDD.n1353 4.65
R2477 VDD.n1350 VDD.n1349 4.65
R2478 VDD.n1345 VDD.n1344 4.65
R2479 VDD.n1341 VDD.n1340 4.65
R2480 VDD.n1315 VDD.n1314 4.65
R2481 VDD.n1311 VDD.n1310 4.65
R2482 VDD.n1307 VDD.n1306 4.65
R2483 VDD.n1303 VDD.n1302 4.65
R2484 VDD.n1299 VDD.n1298 4.65
R2485 VDD.n1293 VDD.n1292 4.65
R2486 VDD.n1289 VDD.n1288 4.65
R2487 VDD.n1285 VDD.n1284 4.65
R2488 VDD.n1279 VDD.n1278 4.65
R2489 VDD.n1275 VDD.n1274 4.65
R2490 VDD.n1270 VDD.n1269 4.65
R2491 VDD.n1266 VDD.n1265 4.65
R2492 VDD.n1240 VDD.n1239 4.65
R2493 VDD.n1236 VDD.n1235 4.65
R2494 VDD.n1232 VDD.n1231 4.65
R2495 VDD.n1228 VDD.n1227 4.65
R2496 VDD.n1224 VDD.n1223 4.65
R2497 VDD.n1218 VDD.n1217 4.65
R2498 VDD.n1214 VDD.n1213 4.65
R2499 VDD.n1210 VDD.n1209 4.65
R2500 VDD.n1204 VDD.n1203 4.65
R2501 VDD.n1200 VDD.n1199 4.65
R2502 VDD.n1195 VDD.n1194 4.65
R2503 VDD.n1191 VDD.n1190 4.65
R2504 VDD.n1165 VDD.n1164 4.65
R2505 VDD.n1161 VDD.n1160 4.65
R2506 VDD.n1157 VDD.n1156 4.65
R2507 VDD.n1153 VDD.n1152 4.65
R2508 VDD.n1149 VDD.n1148 4.65
R2509 VDD.n1143 VDD.n1142 4.65
R2510 VDD.n1139 VDD.n1138 4.65
R2511 VDD.n1135 VDD.n1134 4.65
R2512 VDD.n1129 VDD.n1128 4.65
R2513 VDD.n1125 VDD.n1124 4.65
R2514 VDD.n1120 VDD.n1119 4.65
R2515 VDD.n1116 VDD.n1115 4.65
R2516 VDD.n1090 VDD.n1089 4.65
R2517 VDD.n1086 VDD.n1085 4.65
R2518 VDD.n1082 VDD.n1081 4.65
R2519 VDD.n1078 VDD.n1077 4.65
R2520 VDD.n1074 VDD.n1073 4.65
R2521 VDD.n1068 VDD.n1067 4.65
R2522 VDD.n1064 VDD.n1063 4.65
R2523 VDD.n1060 VDD.n1059 4.65
R2524 VDD.n1054 VDD.n1053 4.65
R2525 VDD.n1050 VDD.n1049 4.65
R2526 VDD.n1045 VDD.n1044 4.65
R2527 VDD.n1041 VDD.n1040 4.65
R2528 VDD.n1015 VDD.n1014 4.65
R2529 VDD.n1011 VDD.n1010 4.65
R2530 VDD.n1007 VDD.n1006 4.65
R2531 VDD.n1003 VDD.n1002 4.65
R2532 VDD.n999 VDD.n998 4.65
R2533 VDD.n993 VDD.n992 4.65
R2534 VDD.n989 VDD.n988 4.65
R2535 VDD.n985 VDD.n984 4.65
R2536 VDD.n979 VDD.n978 4.65
R2537 VDD.n975 VDD.n974 4.65
R2538 VDD.n970 VDD.n969 4.65
R2539 VDD.n966 VDD.n965 4.65
R2540 VDD.n940 VDD.n939 4.65
R2541 VDD.n936 VDD.n935 4.65
R2542 VDD.n932 VDD.n931 4.65
R2543 VDD.n928 VDD.n927 4.65
R2544 VDD.n924 VDD.n923 4.65
R2545 VDD.n918 VDD.n917 4.65
R2546 VDD.n914 VDD.n913 4.65
R2547 VDD.n910 VDD.n909 4.65
R2548 VDD.n904 VDD.n903 4.65
R2549 VDD.n900 VDD.n899 4.65
R2550 VDD.n895 VDD.n894 4.65
R2551 VDD.n891 VDD.n890 4.65
R2552 VDD.n864 VDD.n863 4.65
R2553 VDD.n860 VDD.n859 4.65
R2554 VDD.n856 VDD.n855 4.65
R2555 VDD.n852 VDD.n851 4.65
R2556 VDD.n848 VDD.n847 4.65
R2557 VDD.n842 VDD.n841 4.65
R2558 VDD.n838 VDD.n837 4.65
R2559 VDD.n834 VDD.n833 4.65
R2560 VDD.n828 VDD.n827 4.65
R2561 VDD.n824 VDD.n823 4.65
R2562 VDD.n819 VDD.n818 4.65
R2563 VDD.n815 VDD.n814 4.65
R2564 VDD.n200 VDD.n197 2.89
R2565 VDD.n80 �䛝9V 2.557
R2566 VDD.n130 �F�9V 2.557
R2567 VDD.n189  2.557
R2568 VDD.n178 VDD.n175 2.477
R2569 VDD.n27 VDD.n24 2.064
R2570 VDD.n36 VDD.n35 2.064
R2571 VDD.n271 VDD.n268 0.412
R2572 VDD.n346 VDD.n343 0.412
R2573 VDD.n421 VDD.n418 0.412
R2574 VDD.n496 VDD.n493 0.412
R2575 VDD.n571 VDD.n568 0.412
R2576 VDD.n646 VDD.n643 0.412
R2577 VDD.n721 VDD.n718 0.412
R2578 VDD.n1574 VDD.n1571 0.412
R2579 VDD.n1499 VDD.n1496 0.412
R2580 VDD.n1424 VDD.n1421 0.412
R2581 VDD.n1349 VDD.n1346 0.412
R2582 VDD.n1274 VDD.n1271 0.412
R2583 VDD.n1199 VDD.n1196 0.412
R2584 VDD.n1124 VDD.n1121 0.412
R2585 VDD.n1049 VDD.n1046 0.412
R2586 VDD.n974 VDD.n971 0.412
R2587 VDD.n899 VDD.n896 0.412
R2588 VDD.n823 VDD.n820 0.412
R2589 VDD.n68 VDD.n41 0.29
R2590 VDD.n121 VDD.n95 0.29
R2591 VDD.n174 VDD.n148 0.29
R2592 VDD.n231 VDD.n205 0.29
R2593 VDD.n306 VDD.n280 0.29
R2594 VDD.n381 VDD.n355 0.29
R2595 VDD.n456 VDD.n430 0.29
R2596 VDD.n531 VDD.n505 0.29
R2597 VDD.n606 VDD.n580 0.29
R2598 VDD.n681 VDD.n655 0.29
R2599 VDD.n756 VDD.n730 0.29
R2600 VDD.n1566 VDD.n1540 0.29
R2601 VDD.n1491 VDD.n1465 0.29
R2602 VDD.n1416 VDD.n1390 0.29
R2603 VDD.n1341 VDD.n1315 0.29
R2604 VDD.n1266 VDD.n1240 0.29
R2605 VDD.n1191 VDD.n1165 0.29
R2606 VDD.n1116 VDD.n1090 0.29
R2607 VDD.n1041 VDD.n1015 0.29
R2608 VDD.n966 VDD.n940 0.29
R2609 VDD.n891 VDD.n864 0.29
R2610 VDD.n815 VDD 0.207
R2611 VDD.n257 VDD.n253 0.197
R2612 VDD.n332 VDD.n328 0.197
R2613 VDD.n407 VDD.n403 0.197
R2614 VDD.n482 VDD.n478 0.197
R2615 VDD.n557 VDD.n553 0.197
R2616 VDD.n632 VDD.n628 0.197
R2617 VDD.n707 VDD.n703 0.197
R2618 VDD.n782 VDD.n778 0.197
R2619 VDD.n1518 VDD.n1514 0.197
R2620 VDD.n1443 VDD.n1439 0.197
R2621 VDD.n1368 VDD.n1364 0.197
R2622 VDD.n1293 VDD.n1289 0.197
R2623 VDD.n1218 VDD.n1214 0.197
R2624 VDD.n1143 VDD.n1139 0.197
R2625 VDD.n1068 VDD.n1064 0.197
R2626 VDD.n993 VDD.n989 0.197
R2627 VDD.n918 VDD.n914 0.197
R2628 VDD.n842 VDD.n838 0.197
R2629 VDD.n83 VDD.n79 0.181
R2630 VDD.n136 VDD.n133 0.181
R2631 VDD.n192 VDD.n188 0.181
R2632 VDD.n32 VDD.n28 0.157
R2633 VDD.n37 VDD.n32 0.157
R2634 VDD.n41 VDD.n37 0.145
R2635 VDD.n72 VDD.n68 0.145
R2636 VDD.n76 VDD.n72 0.145
R2637 VDD.n79 VDD.n76 0.145
R2638 VDD.n87 VDD.n83 0.145
R2639 VDD.n91 VDD.n87 0.145
R2640 VDD.n95 VDD.n91 0.145
R2641 VDD.n125 VDD.n121 0.145
R2642 VDD.n129 VDD.n125 0.145
R2643 VDD.n133 VDD.n129 0.145
R2644 VDD.n140 VDD.n136 0.145
R2645 VDD.n144 VDD.n140 0.145
R2646 VDD.n148 VDD.n144 0.145
R2647 VDD.n179 VDD.n174 0.145
R2648 VDD.n183 VDD.n179 0.145
R2649 VDD.n188 VDD.n183 0.145
R2650 VDD.n196 VDD.n192 0.145
R2651 VDD.n201 VDD.n196 0.145
R2652 VDD.n205 VDD.n201 0.145
R2653 VDD.n235 VDD.n231 0.145
R2654 VDD.n239 VDD.n235 0.145
R2655 VDD.n243 VDD.n239 0.145
R2656 VDD.n249 VDD.n243 0.145
R2657 VDD.n253 VDD.n249 0.145
R2658 VDD.n263 VDD.n257 0.145
R2659 VDD.n267 VDD.n263 0.145
R2660 VDD.n272 VDD.n267 0.145
R2661 VDD.n276 VDD.n272 0.145
R2662 VDD.n280 VDD.n276 0.145
R2663 VDD.n310 VDD.n306 0.145
R2664 VDD.n314 VDD.n310 0.145
R2665 VDD.n318 VDD.n314 0.145
R2666 VDD.n324 VDD.n318 0.145
R2667 VDD.n328 VDD.n324 0.145
R2668 VDD.n338 VDD.n332 0.145
R2669 VDD.n342 VDD.n338 0.145
R2670 VDD.n347 VDD.n342 0.145
R2671 VDD.n351 VDD.n347 0.145
R2672 VDD.n355 VDD.n351 0.145
R2673 VDD.n385 VDD.n381 0.145
R2674 VDD.n389 VDD.n385 0.145
R2675 VDD.n393 VDD.n389 0.145
R2676 VDD.n399 VDD.n393 0.145
R2677 VDD.n403 VDD.n399 0.145
R2678 VDD.n413 VDD.n407 0.145
R2679 VDD.n417 VDD.n413 0.145
R2680 VDD.n422 VDD.n417 0.145
R2681 VDD.n426 VDD.n422 0.145
R2682 VDD.n430 VDD.n426 0.145
R2683 VDD.n460 VDD.n456 0.145
R2684 VDD.n464 VDD.n460 0.145
R2685 VDD.n468 VDD.n464 0.145
R2686 VDD.n474 VDD.n468 0.145
R2687 VDD.n478 VDD.n474 0.145
R2688 VDD.n488 VDD.n482 0.145
R2689 VDD.n492 VDD.n488 0.145
R2690 VDD.n497 VDD.n492 0.145
R2691 VDD.n501 VDD.n497 0.145
R2692 VDD.n505 VDD.n501 0.145
R2693 VDD.n535 VDD.n531 0.145
R2694 VDD.n539 VDD.n535 0.145
R2695 VDD.n543 VDD.n539 0.145
R2696 VDD.n549 VDD.n543 0.145
R2697 VDD.n553 VDD.n549 0.145
R2698 VDD.n563 VDD.n557 0.145
R2699 VDD.n567 VDD.n563 0.145
R2700 VDD.n572 VDD.n567 0.145
R2701 VDD.n576 VDD.n572 0.145
R2702 VDD.n580 VDD.n576 0.145
R2703 VDD.n610 VDD.n606 0.145
R2704 VDD.n614 VDD.n610 0.145
R2705 VDD.n618 VDD.n614 0.145
R2706 VDD.n624 VDD.n618 0.145
R2707 VDD.n628 VDD.n624 0.145
R2708 VDD.n638 VDD.n632 0.145
R2709 VDD.n642 VDD.n638 0.145
R2710 VDD.n647 VDD.n642 0.145
R2711 VDD.n651 VDD.n647 0.145
R2712 VDD.n655 VDD.n651 0.145
R2713 VDD.n685 VDD.n681 0.145
R2714 VDD.n689 VDD.n685 0.145
R2715 VDD.n693 VDD.n689 0.145
R2716 VDD.n699 VDD.n693 0.145
R2717 VDD.n703 VDD.n699 0.145
R2718 VDD.n713 VDD.n707 0.145
R2719 VDD.n717 VDD.n713 0.145
R2720 VDD.n722 VDD.n717 0.145
R2721 VDD.n726 VDD.n722 0.145
R2722 VDD.n730 VDD.n726 0.145
R2723 VDD.n760 VDD.n756 0.145
R2724 VDD.n764 VDD.n760 0.145
R2725 VDD.n768 VDD.n764 0.145
R2726 VDD.n774 VDD.n768 0.145
R2727 VDD.n778 VDD.n774 0.145
R2728 VDD.n788 VDD.n782 0.145
R2729 VDD.n792 VDD.n788 0.145
R2730 VDD.n1575 VDD.n1570 0.145
R2731 VDD.n1570 VDD.n1566 0.145
R2732 VDD.n1540 VDD.n1536 0.145
R2733 VDD.n1536 VDD.n1532 0.145
R2734 VDD.n1532 VDD.n1528 0.145
R2735 VDD.n1528 VDD.n1524 0.145
R2736 VDD.n1524 VDD.n1518 0.145
R2737 VDD.n1514 VDD.n1510 0.145
R2738 VDD.n1510 VDD.n1504 0.145
R2739 VDD.n1504 VDD.n1500 0.145
R2740 VDD.n1500 VDD.n1495 0.145
R2741 VDD.n1495 VDD.n1491 0.145
R2742 VDD.n1465 VDD.n1461 0.145
R2743 VDD.n1461 VDD.n1457 0.145
R2744 VDD.n1457 VDD.n1453 0.145
R2745 VDD.n1453 VDD.n1449 0.145
R2746 VDD.n1449 VDD.n1443 0.145
R2747 VDD.n1439 VDD.n1435 0.145
R2748 VDD.n1435 VDD.n1429 0.145
R2749 VDD.n1429 VDD.n1425 0.145
R2750 VDD.n1425 VDD.n1420 0.145
R2751 VDD.n1420 VDD.n1416 0.145
R2752 VDD.n1390 VDD.n1386 0.145
R2753 VDD.n1386 VDD.n1382 0.145
R2754 VDD.n1382 VDD.n1378 0.145
R2755 VDD.n1378 VDD.n1374 0.145
R2756 VDD.n1374 VDD.n1368 0.145
R2757 VDD.n1364 VDD.n1360 0.145
R2758 VDD.n1360 VDD.n1354 0.145
R2759 VDD.n1354 VDD.n1350 0.145
R2760 VDD.n1350 VDD.n1345 0.145
R2761 VDD.n1345 VDD.n1341 0.145
R2762 VDD.n1315 VDD.n1311 0.145
R2763 VDD.n1311 VDD.n1307 0.145
R2764 VDD.n1307 VDD.n1303 0.145
R2765 VDD.n1303 VDD.n1299 0.145
R2766 VDD.n1299 VDD.n1293 0.145
R2767 VDD.n1289 VDD.n1285 0.145
R2768 VDD.n1285 VDD.n1279 0.145
R2769 VDD.n1279 VDD.n1275 0.145
R2770 VDD.n1275 VDD.n1270 0.145
R2771 VDD.n1270 VDD.n1266 0.145
R2772 VDD.n1240 VDD.n1236 0.145
R2773 VDD.n1236 VDD.n1232 0.145
R2774 VDD.n1232 VDD.n1228 0.145
R2775 VDD.n1228 VDD.n1224 0.145
R2776 VDD.n1224 VDD.n1218 0.145
R2777 VDD.n1214 VDD.n1210 0.145
R2778 VDD.n1210 VDD.n1204 0.145
R2779 VDD.n1204 VDD.n1200 0.145
R2780 VDD.n1200 VDD.n1195 0.145
R2781 VDD.n1195 VDD.n1191 0.145
R2782 VDD.n1165 VDD.n1161 0.145
R2783 VDD.n1161 VDD.n1157 0.145
R2784 VDD.n1157 VDD.n1153 0.145
R2785 VDD.n1153 VDD.n1149 0.145
R2786 VDD.n1149 VDD.n1143 0.145
R2787 VDD.n1139 VDD.n1135 0.145
R2788 VDD.n1135 VDD.n1129 0.145
R2789 VDD.n1129 VDD.n1125 0.145
R2790 VDD.n1125 VDD.n1120 0.145
R2791 VDD.n1120 VDD.n1116 0.145
R2792 VDD.n1090 VDD.n1086 0.145
R2793 VDD.n1086 VDD.n1082 0.145
R2794 VDD.n1082 VDD.n1078 0.145
R2795 VDD.n1078 VDD.n1074 0.145
R2796 VDD.n1074 VDD.n1068 0.145
R2797 VDD.n1064 VDD.n1060 0.145
R2798 VDD.n1060 VDD.n1054 0.145
R2799 VDD.n1054 VDD.n1050 0.145
R2800 VDD.n1050 VDD.n1045 0.145
R2801 VDD.n1045 VDD.n1041 0.145
R2802 VDD.n1015 VDD.n1011 0.145
R2803 VDD.n1011 VDD.n1007 0.145
R2804 VDD.n1007 VDD.n1003 0.145
R2805 VDD.n1003 VDD.n999 0.145
R2806 VDD.n999 VDD.n993 0.145
R2807 VDD.n989 VDD.n985 0.145
R2808 VDD.n985 VDD.n979 0.145
R2809 VDD.n979 VDD.n975 0.145
R2810 VDD.n975 VDD.n970 0.145
R2811 VDD.n970 VDD.n966 0.145
R2812 VDD.n940 VDD.n936 0.145
R2813 VDD.n936 VDD.n932 0.145
R2814 VDD.n932 VDD.n928 0.145
R2815 VDD.n928 VDD.n924 0.145
R2816 VDD.n924 VDD.n918 0.145
R2817 VDD.n914 VDD.n910 0.145
R2818 VDD.n910 VDD.n904 0.145
R2819 VDD.n904 VDD.n900 0.145
R2820 VDD.n900 VDD.n895 0.145
R2821 VDD.n895 VDD.n891 0.145
R2822 VDD.n864 VDD.n860 0.145
R2823 VDD.n860 VDD.n856 0.145
R2824 VDD.n856 VDD.n852 0.145
R2825 VDD.n852 VDD.n848 0.145
R2826 VDD.n848 VDD.n842 0.145
R2827 VDD.n838 VDD.n834 0.145
R2828 VDD.n834 VDD.n828 0.145
R2829 VDD.n828 VDD.n824 0.145
R2830 VDD.n824 VDD.n819 0.145
R2831 VDD.n819 VDD.n815 0.145
R2832 VDD VDD.n1575 0.086
R2833 VDD VDD.n792 0.058
R2834 CLK.n18 CLK.t14 459.505
R2835 CLK.n15 CLK.t1 459.505
R2836 CLK.n12 CLK.t17 459.505
R2837 CLK.n7 CLK.t11 459.505
R2838 CLK.n4 CLK.t3 459.505
R2839 CLK.n0 CLK.t12 459.505
R2840 CLK.n16 CLK.t6 399.181
R2841 CLK.n8 CLK.t9 399.181
R2842 CLK.n1 CLK.t13 399.181
R2843 CLK.n20 CLK.t5 398.835
R2844 CLK.n10 CLK.t4 397.657
R2845 CLK.n2 CLK.t15 397.657
R2846 CLK.n18 CLK.t0 384.527
R2847 CLK.n15 CLK.t8 384.527
R2848 CLK.n12 CLK.t10 384.527
R2849 CLK.n7 CLK.t2 384.527
R2850 CLK.n4 CLK.t7 384.527
R2851 CLK.n0 CLK.t16 384.527
R2852 CLK.n1 CLK.n0 33.832
R2853 CLK.n8 CLK.n7 33.832
R2854 CLK.n16 CLK.n15 33.832
R2855 CLK.n19 CLK.n18 30.851
R2856 CLK.n13 CLK.n12 30.851
R2857 CLK.n5 CLK.n4 30.851
R2858 CLK.n9 CLK.n6 14.075
R2859 CLK.n17 CLK.n14 14.075
R2860 CLK.n19 CLK 9.3
R2861 CLK.n3 CLK.n1 9.111
R2862 CLK.n11 CLK.n9 7.032
R2863 CLK.n21 CLK.n17 7.032
R2864 CLK.n6 CLK.n5 4.639
R2865 CLK.n14 CLK.n13 4.639
R2866 CLK.n3 CLK.n2 4.234
R2867 CLK.n11 CLK.n10 4.234
R2868 CLK.n20 CLK.n19 2.59
R2869 CLK.n21 CLK.n20 2.1
R2870 CLK.n9 CLK.n8 2.079
R2871 CLK.n17 CLK.n16 2.079
R2872 CLK.n21 CLK 0.046
R2873 CLK.n6 CLK.n3 0.023
R2874 CLK.n14 CLK.n11 0.023
R2875 a_599_989.n1 a_599_989.t12 512.525
R2876 a_599_989.n3 a_599_989.t11 454.685
R2877 a_599_989.n3 a_599_989.t9 428.979
R2878 a_599_989.n1 a_599_989.t8 371.139
R2879 a_599_989.n2 a_599_989.t7 361.392
R2880 a_599_989.n7 a_599_989.n6 329.955
R2881 a_599_989.n4 a_599_989.t10 311.683
R2882 a_599_989.n2 a_599_989.n1 235.554
R2883 a_599_989.n8 a_599_989.n7 179.199
R2884 a_599_989.n4 a_599_989.n3 171.288
R2885 a_599_989.n10 a_599_989.n9 161.352
R2886 a_599_989.n8 a_599_989.n0 95.095
R2887 a_599_989.n11 a_599_989.n10 95.094
R2888 a_599_989.n10 a_599_989.n8 66.258
R2889 a_599_989.n0 a_599_989.t2 14.282
R2890 a_599_989.n0 a_599_989.t3 14.282
R2891 a_599_989.n9 a_599_989.t0 14.282
R2892 a_599_989.n9 a_599_989.t1 14.282
R2893 a_599_989.n11 a_599_989.t5 14.282
R2894 a_599_989.t6 a_599_989.n11 14.282
R2895 a_599_989.n5 a_599_989.n2 13.038
R2896 a_599_989.n5 a_599_989.n4 8.685
R2897 a_599_989.n7 a_599_989.n5 4.65
R2898 a_9897_1050.n1 a_9897_1050.t7 512.525
R2899 a_9897_1050.n1 a_9897_1050.t9 371.139
R2900 a_9897_1050.n2 a_9897_1050.t8 361.392
R2901 a_9897_1050.n4 a_9897_1050.n3 329.955
R2902 a_9897_1050.n2 a_9897_1050.n1 235.554
R2903 a_9897_1050.n5 a_9897_1050.n4 179.199
R2904 a_9897_1050.n7 a_9897_1050.n6 161.352
R2905 a_9897_1050.n5 a_9897_1050.n0 95.095
R2906 a_9897_1050.n8 a_9897_1050.n7 95.094
R2907 a_9897_1050.n7 a_9897_1050.n5 66.258
R2908 a_9897_1050.n0 a_9897_1050.t6 14.282
R2909 a_9897_1050.n0 a_9897_1050.t1 14.282
R2910 a_9897_1050.n6 a_9897_1050.t0 14.282
R2911 a_9897_1050.n6 a_9897_1050.t2 14.282
R2912 a_9897_1050.t4 a_9897_1050.n8 14.282
R2913 a_9897_1050.n8 a_9897_1050.t3 14.282
R2914 a_9897_1050.n4 a_9897_1050.n2 10.615
R2915 a_3939_103.n5 a_3939_103.n4 66.708
R2916 a_3939_103.n2 a_3939_103.n0 32.662
R2917 a_3939_103.n5 a_3939_103.n3 19.496
R2918 a_3939_103.t0 a_3939_103.n5 13.756
R2919 a_3939_103.t0 a_3939_103.n2 3.034
R2920 a_3939_103.n2 a_3939_103.n1 0.443
R2921 a_1561_989.n2 a_1561_989.t12 454.685
R2922 a_1561_989.n4 a_1561_989.t7 454.685
R2923 a_1561_989.n0 a_1561_989.t15 454.685
R2924 a_1561_989.n2 a_1561_989.t8 428.979
R2925 a_1561_989.n4 a_1561_989.t9 428.979
R2926 a_1561_989.n0 a_1561_989.t10 428.979
R2927 a_1561_989.n3 a_1561_989.t11 339.542
R2928 a_1561_989.n1 a_1561_989.t14 339.542
R2929 a_1561_989.n5 a_1561_989.t13 339.186
R2930 a_1561_989.n12 a_1561_989.n11 336.075
R2931 a_1561_989.n15 a_1561_989.n14 161.352
R2932 a_1561_989.n16 a_1561_989.n12 151.34
R2933 a_1561_989.n3 a_1561_989.n2 143.429
R2934 a_1561_989.n1 a_1561_989.n0 143.429
R2935 a_1561_989.n5 a_1561_989.n4 143.074
R2936 a_1561_989.n15 a_1561_989.n13 95.095
R2937 a_1561_989.n17 a_1561_989.n16 95.094
R2938 a_1561_989.n16 a_1561_989.n15 66.258
R2939 a_1561_989.n11 a_1561_989.n10 30
R2940 a_1561_989.n9 a_1561_989.n8 24.383
R2941 a_1561_989.n11 a_1561_989.n9 23.684
R2942 a_1561_989.n13 a_1561_989.t6 14.282
R2943 a_1561_989.n13 a_1561_989.t5 14.282
R2944 a_1561_989.n14 a_1561_989.t0 14.282
R2945 a_1561_989.n14 a_1561_989.t1 14.282
R2946 a_1561_989.t4 a_1561_989.n17 14.282
R2947 a_1561_989.n17 a_1561_989.t3 14.282
R2948 a_1561_989.n7 a_1561_989.n1 11.134
R2949 a_1561_989.n6 a_1561_989.n5 8.145
R2950 a_1561_989.n6 a_1561_989.n3 4.65
R2951 a_1561_989.n12 a_1561_989.n7 4.65
R2952 a_1561_989.n7 a_1561_989.n6 4.035
R2953 a_12143_989.n1 a_12143_989.t12 512.525
R2954 a_12143_989.n3 a_12143_989.t7 454.685
R2955 a_12143_989.n3 a_12143_989.t10 428.979
R2956 a_12143_989.n1 a_12143_989.t8 371.139
R2957 a_12143_989.n2 a_12143_989.t9 361.392
R2958 a_12143_989.n4 a_12143_989.t11 311.683
R2959 a_12143_989.n10 a_12143_989.n9 308.216
R2960 a_12143_989.n2 a_12143_989.n1 235.554
R2961 a_12143_989.n11 a_12143_989.n10 179.199
R2962 a_12143_989.n4 a_12143_989.n3 171.288
R2963 a_12143_989.n13 a_12143_989.n12 161.352
R2964 a_12143_989.n11 a_12143_989.n0 95.095
R2965 a_12143_989.n14 a_12143_989.n13 95.094
R2966 a_12143_989.n13 a_12143_989.n11 66.258
R2967 a_12143_989.n9 a_12143_989.n8 30
R2968 a_12143_989.n7 a_12143_989.n6 24.383
R2969 a_12143_989.n9 a_12143_989.n7 23.684
R2970 a_12143_989.n0 a_12143_989.t6 14.282
R2971 a_12143_989.n0 a_12143_989.t5 14.282
R2972 a_12143_989.n12 a_12143_989.t1 14.282
R2973 a_12143_989.n12 a_12143_989.t0 14.282
R2974 a_12143_989.t3 a_12143_989.n14 14.282
R2975 a_12143_989.n14 a_12143_989.t2 14.282
R2976 a_12143_989.n5 a_12143_989.n2 13.038
R2977 a_12143_989.n5 a_12143_989.n4 8.685
R2978 a_12143_989.n10 a_12143_989.n5 4.65
R2979 a_11821_1050.n2 a_11821_1050.t11 512.525
R2980 a_11821_1050.n0 a_11821_1050.t9 512.525
R2981 a_11821_1050.n2 a_11821_1050.t7 371.139
R2982 a_11821_1050.n0 a_11821_1050.t12 371.139
R2983 a_11821_1050.n3 a_11821_1050.t8 306.051
R2984 a_11821_1050.n1 a_11821_1050.t10 306.051
R2985 a_11821_1050.n3 a_11821_1050.n2 290.895
R2986 a_11821_1050.n1 a_11821_1050.n0 290.895
R2987 a_11821_1050.n9 a_11821_1050.n8 252.875
R2988 a_11821_1050.n13 a_11821_1050.n9 234.54
R2989 a_11821_1050.n12 a_11821_1050.n11 161.352
R2990 a_11821_1050.n12 a_11821_1050.n10 95.095
R2991 a_11821_1050.n14 a_11821_1050.n13 95.094
R2992 a_11821_1050.n13 a_11821_1050.n12 66.258
R2993 a_11821_1050.n8 a_11821_1050.n7 30
R2994 a_11821_1050.n6 a_11821_1050.n5 24.383
R2995 a_11821_1050.n8 a_11821_1050.n6 23.684
R2996 a_11821_1050.n10 a_11821_1050.t6 14.282
R2997 a_11821_1050.n10 a_11821_1050.t5 14.282
R2998 a_11821_1050.n11 a_11821_1050.t0 14.282
R2999 a_11821_1050.n11 a_11821_1050.t1 14.282
R3000 a_11821_1050.n14 a_11821_1050.t3 14.282
R3001 a_11821_1050.t4 a_11821_1050.n14 14.282
R3002 a_11821_1050.n4 a_11821_1050.n1 8.141
R3003 a_11821_1050.n9 a_11821_1050.n4 5.965
R3004 a_11821_1050.n4 a_11821_1050.n3 4.65
R3005 a_9030_210.n11 a_9030_210.n8 171.558
R3006 a_9030_210.n1 a_9030_210.n0 102.58
R3007 a_9030_210.t0 a_9030_210.n13 83.571
R3008 a_9030_210.t0 a_9030_210.n11 75.765
R3009 a_9030_210.n3 a_9030_210.n2 65.02
R3010 a_9030_210.t0 a_9030_210.n3 58.043
R3011 a_9030_210.n13 a_9030_210.n12 55.714
R3012 a_9030_210.n3 a_9030_210.n1 35.865
R3013 a_9030_210.n8 a_9030_210.n7 27.2
R3014 a_9030_210.n6 a_9030_210.n5 23.498
R3015 a_9030_210.n8 a_9030_210.n6 22.4
R3016 a_9030_210.n10 a_9030_210.n9 19.952
R3017 a_9030_210.t0 a_9030_210.n4 8.137
R3018 a_9030_210.n11 a_9030_210.n10 1.505
R3019 a_7333_989.n2 a_7333_989.t8 454.685
R3020 a_7333_989.n4 a_7333_989.t10 454.685
R3021 a_7333_989.n0 a_7333_989.t9 454.685
R3022 a_7333_989.n2 a_7333_989.t14 428.979
R3023 a_7333_989.n4 a_7333_989.t7 428.979
R3024 a_7333_989.n0 a_7333_989.t11 428.979
R3025 a_7333_989.n9 a_7333_989.n8 357.814
R3026 a_7333_989.n3 a_7333_989.t13 339.542
R3027 a_7333_989.n1 a_7333_989.t15 339.542
R3028 a_7333_989.n5 a_7333_989.t12 339.186
R3029 a_7333_989.n12 a_7333_989.n11 161.352
R3030 a_7333_989.n13 a_7333_989.n9 151.34
R3031 a_7333_989.n3 a_7333_989.n2 143.429
R3032 a_7333_989.n1 a_7333_989.n0 143.429
R3033 a_7333_989.n5 a_7333_989.n4 143.074
R3034 a_7333_989.n12 a_7333_989.n10 95.095
R3035 a_7333_989.n14 a_7333_989.n13 95.094
R3036 a_7333_989.n13 a_7333_989.n12 66.258
R3037 a_7333_989.n10 a_7333_989.t5 14.282
R3038 a_7333_989.n10 a_7333_989.t6 14.282
R3039 a_7333_989.n11 a_7333_989.t1 14.282
R3040 a_7333_989.n11 a_7333_989.t0 14.282
R3041 a_7333_989.t4 a_7333_989.n14 14.282
R3042 a_7333_989.n14 a_7333_989.t3 14.282
R3043 a_7333_989.n7 a_7333_989.n1 11.134
R3044 a_7333_989.n6 a_7333_989.n5 8.145
R3045 a_7333_989.n6 a_7333_989.n3 4.65
R3046 a_7333_989.n9 a_7333_989.n7 4.65
R3047 a_7333_989.n7 a_7333_989.n6 4.035
R3048 a_13745_1050.n2 a_13745_1050.t7 512.525
R3049 a_13745_1050.n2 a_13745_1050.t9 371.139
R3050 a_13745_1050.n3 a_13745_1050.t8 305.674
R3051 a_13745_1050.n3 a_13745_1050.n2 291.272
R3052 a_13745_1050.n8 a_13745_1050.n7 252.498
R3053 a_13745_1050.n9 a_13745_1050.n8 234.917
R3054 a_13745_1050.n11 a_13745_1050.n10 161.352
R3055 a_13745_1050.n9 a_13745_1050.n1 95.095
R3056 a_13745_1050.n10 a_13745_1050.n0 95.095
R3057 a_13745_1050.n10 a_13745_1050.n9 66.258
R3058 a_13745_1050.n7 a_13745_1050.n6 30
R3059 a_13745_1050.n5 a_13745_1050.n4 24.383
R3060 a_13745_1050.n7 a_13745_1050.n5 23.684
R3061 a_13745_1050.n1 a_13745_1050.t6 14.282
R3062 a_13745_1050.n1 a_13745_1050.t5 14.282
R3063 a_13745_1050.n0 a_13745_1050.t1 14.282
R3064 a_13745_1050.n0 a_13745_1050.t0 14.282
R3065 a_13745_1050.t3 a_13745_1050.n11 14.282
R3066 a_13745_1050.n11 a_13745_1050.t2 14.282
R3067 a_13745_1050.n8 a_13745_1050.n3 10.615
R3068 a_277_1050.n2 a_277_1050.t8 512.525
R3069 a_277_1050.n0 a_277_1050.t7 512.525
R3070 a_277_1050.n2 a_277_1050.t9 371.139
R3071 a_277_1050.n0 a_277_1050.t10 371.139
R3072 a_277_1050.n3 a_277_1050.t12 306.051
R3073 a_277_1050.n1 a_277_1050.t11 306.051
R3074 a_277_1050.n3 a_277_1050.n2 290.895
R3075 a_277_1050.n1 a_277_1050.n0 290.895
R3076 a_277_1050.n9 a_277_1050.n8 252.875
R3077 a_277_1050.n13 a_277_1050.n9 234.54
R3078 a_277_1050.n12 a_277_1050.n11 161.352
R3079 a_277_1050.n12 a_277_1050.n10 95.095
R3080 a_277_1050.n14 a_277_1050.n13 95.094
R3081 a_277_1050.n13 a_277_1050.n12 66.258
R3082 a_277_1050.n8 a_277_1050.n7 30
R3083 a_277_1050.n6 a_277_1050.n5 24.383
R3084 a_277_1050.n8 a_277_1050.n6 23.684
R3085 a_277_1050.n10 a_277_1050.t6 14.282
R3086 a_277_1050.n10 a_277_1050.t5 14.282
R3087 a_277_1050.n11 a_277_1050.t0 14.282
R3088 a_277_1050.n11 a_277_1050.t1 14.282
R3089 a_277_1050.t4 a_277_1050.n14 14.282
R3090 a_277_1050.n14 a_277_1050.t3 14.282
R3091 a_277_1050.n4 a_277_1050.n1 8.141
R3092 a_277_1050.n9 a_277_1050.n4 5.965
R3093 a_277_1050.n4 a_277_1050.n3 4.65
R3094 a_2201_1050.n2 a_2201_1050.t9 512.525
R3095 a_2201_1050.n2 a_2201_1050.t7 371.139
R3096 a_2201_1050.n3 a_2201_1050.t8 305.674
R3097 a_2201_1050.n3 a_2201_1050.n2 291.272
R3098 a_2201_1050.n8 a_2201_1050.n7 252.498
R3099 a_2201_1050.n9 a_2201_1050.n8 234.917
R3100 a_2201_1050.n11 a_2201_1050.n10 161.352
R3101 a_2201_1050.n9 a_2201_1050.n1 95.095
R3102 a_2201_1050.n10 a_2201_1050.n0 95.095
R3103 a_2201_1050.n10 a_2201_1050.n9 66.258
R3104 a_2201_1050.n7 a_2201_1050.n6 30
R3105 a_2201_1050.n5 a_2201_1050.n4 24.383
R3106 a_2201_1050.n7 a_2201_1050.n5 23.684
R3107 a_2201_1050.n1 a_2201_1050.t6 14.282
R3108 a_2201_1050.n1 a_2201_1050.t5 14.282
R3109 a_2201_1050.n0 a_2201_1050.t1 14.282
R3110 a_2201_1050.n0 a_2201_1050.t0 14.282
R3111 a_2201_1050.t3 a_2201_1050.n11 14.282
R3112 a_2201_1050.n11 a_2201_1050.t2 14.282
R3113 a_2201_1050.n8 a_2201_1050.n3 10.615
R3114 SN.n14 SN.t2 479.223
R3115 SN.n11 SN.t6 479.223
R3116 SN.n8 SN.t7 479.223
R3117 SN.n5 SN.t14 479.223
R3118 SN.n2 SN.t8 479.223
R3119 SN.n0 SN.t13 479.223
R3120 SN.n14 SN.t11 375.52
R3121 SN.n11 SN.t15 375.52
R3122 SN.n8 SN.t16 375.52
R3123 SN.n5 SN.t0 375.52
R3124 SN.n2 SN.t4 375.52
R3125 SN.n0 SN.t5 375.52
R3126 SN.n12 SN.n11 280.047
R3127 SN.n6 SN.n5 280.047
R3128 SN.n1 SN.n0 280.047
R3129 SN.n3 SN.n2 276.525
R3130 SN.n9 SN.n8 276.525
R3131 SN.n15 SN.n14 276.525
R3132 SN.n12 SN.t1 136.76
R3133 SN.n6 SN.t9 136.76
R3134 SN.n1 SN.t10 136.76
R3135 SN.n15 SN.t17 135.513
R3136 SN.n9 SN.t3 135.513
R3137 SN.n3 SN.t12 135.513
R3138 SN.n4 SN.n1 15.211
R3139 SN.n7 SN.n4 10.564
R3140 SN.n13 SN.n10 10.564
R3141 SN.n10 SN.n7 10.561
R3142 SN.n16 SN.n13 10.561
R3143 SN.n7 SN.n6 4.65
R3144 SN.n13 SN.n12 4.65
R3145 SN.n4 SN.n3 2.113
R3146 SN.n10 SN.n9 2.113
R3147 SN.n16 SN.n15 2.113
R3148 SN.n16 SN 0.046
R3149 a_10219_989.n1 a_10219_989.t15 475.572
R3150 a_10219_989.n3 a_10219_989.t11 469.145
R3151 a_10219_989.n6 a_10219_989.t9 454.685
R3152 a_10219_989.n6 a_10219_989.t14 428.979
R3153 a_10219_989.n3 a_10219_989.t7 384.527
R3154 a_10219_989.n1 a_10219_989.t10 384.527
R3155 a_10219_989.n4 a_10219_989.t12 370.613
R3156 a_10219_989.n2 a_10219_989.t8 370.613
R3157 a_10219_989.n7 a_10219_989.t13 255.965
R3158 a_10219_989.n12 a_10219_989.n11 252.498
R3159 a_10219_989.n7 a_10219_989.n6 227.006
R3160 a_10219_989.n16 a_10219_989.n15 161.352
R3161 a_10219_989.n14 a_10219_989.n13 151.34
R3162 a_10219_989.n2 a_10219_989.n1 128.028
R3163 a_10219_989.n4 a_10219_989.n3 126.97
R3164 a_10219_989.n14 a_10219_989.n0 95.095
R3165 a_10219_989.n17 a_10219_989.n16 95.094
R3166 a_10219_989.n13 a_10219_989.n12 83.576
R3167 a_10219_989.n16 a_10219_989.n14 66.258
R3168 a_10219_989.n11 a_10219_989.n10 30
R3169 a_10219_989.n13 a_10219_989.n5 27.875
R3170 a_10219_989.n9 a_10219_989.n8 24.383
R3171 a_10219_989.n11 a_10219_989.n9 23.684
R3172 a_10219_989.n0 a_10219_989.t3 14.282
R3173 a_10219_989.n0 a_10219_989.t4 14.282
R3174 a_10219_989.n15 a_10219_989.t6 14.282
R3175 a_10219_989.n15 a_10219_989.t5 14.282
R3176 a_10219_989.n17 a_10219_989.t0 14.282
R3177 a_10219_989.t1 a_10219_989.n17 14.282
R3178 a_10219_989.n12 a_10219_989.n7 13.335
R3179 a_10219_989.n5 a_10219_989.n2 9.501
R3180 a_10219_989.n5 a_10219_989.n4 4.65
R3181 a_6371_989.n0 a_6371_989.t10 512.525
R3182 a_6371_989.n2 a_6371_989.t12 454.685
R3183 a_6371_989.n2 a_6371_989.t8 428.979
R3184 a_6371_989.n0 a_6371_989.t7 371.139
R3185 a_6371_989.n1 a_6371_989.t9 361.392
R3186 a_6371_989.n3 a_6371_989.t11 311.683
R3187 a_6371_989.n9 a_6371_989.n8 308.216
R3188 a_6371_989.n1 a_6371_989.n0 235.554
R3189 a_6371_989.n13 a_6371_989.n9 179.199
R3190 a_6371_989.n3 a_6371_989.n2 171.288
R3191 a_6371_989.n12 a_6371_989.n11 161.352
R3192 a_6371_989.n12 a_6371_989.n10 95.095
R3193 a_6371_989.n14 a_6371_989.n13 95.094
R3194 a_6371_989.n13 a_6371_989.n12 66.258
R3195 a_6371_989.n8 a_6371_989.n7 30
R3196 a_6371_989.n6 a_6371_989.n5 24.383
R3197 a_6371_989.n8 a_6371_989.n6 23.684
R3198 a_6371_989.n10 a_6371_989.t5 14.282
R3199 a_6371_989.n10 a_6371_989.t6 14.282
R3200 a_6371_989.n11 a_6371_989.t0 14.282
R3201 a_6371_989.n11 a_6371_989.t4 14.282
R3202 a_6371_989.t3 a_6371_989.n14 14.282
R3203 a_6371_989.n14 a_6371_989.t2 14.282
R3204 a_6371_989.n4 a_6371_989.n1 13.038
R3205 a_6371_989.n4 a_6371_989.n3 8.685
R3206 a_6371_989.n9 a_6371_989.n4 4.65
R3207 a_4901_103.n5 a_4901_103.n4 66.708
R3208 a_4901_103.n2 a_4901_103.n0 32.662
R3209 a_4901_103.n5 a_4901_103.n3 19.496
R3210 a_4901_103.t0 a_4901_103.n5 13.756
R3211 a_4901_103.t0 a_4901_103.n2 3.034
R3212 a_4901_103.n2 a_4901_103.n1 0.443
R3213 a_5182_210.n12 a_5182_210.n10 171.558
R3214 a_5182_210.n7 a_5182_210.n6 117.622
R3215 a_5182_210.n5 a_5182_210.n4 92.5
R3216 a_5182_210.n9 a_5182_210.n8 92.5
R3217 a_5182_210.n10 a_5182_210.t1 75.764
R3218 a_5182_210.n5 a_5182_210.n3 65.02
R3219 a_5182_210.n13 a_5182_210.n0 49.6
R3220 a_5182_210.n7 a_5182_210.n5 36.517
R3221 a_5182_210.n3 a_5182_210.n2 35.865
R3222 a_5182_210.n12 a_5182_210.n11 27.2
R3223 a_5182_210.n13 a_5182_210.n12 22.4
R3224 a_5182_210.n9 a_5182_210.n7 19.952
R3225 a_5182_210.t1 a_5182_210.n1 7.04
R3226 a_5182_210.n10 a_5182_210.n9 1.505
R3227 a_6825_103.n5 a_6825_103.n4 66.708
R3228 a_6825_103.n2 a_6825_103.n0 32.662
R3229 a_6825_103.n5 a_6825_103.n3 19.496
R3230 a_6825_103.t0 a_6825_103.n5 13.756
R3231 a_6825_103.t0 a_6825_103.n2 3.034
R3232 a_6825_103.n2 a_6825_103.n1 0.443
R3233 a_7106_210.n8 a_7106_210.n6 185.173
R3234 a_7106_210.t0 a_7106_210.n8 75.765
R3235 a_7106_210.n3 a_7106_210.n1 74.827
R3236 a_7106_210.n3 a_7106_210.n2 27.476
R3237 a_7106_210.n6 a_7106_210.n5 22.349
R3238 a_7106_210.t0 a_7106_210.n10 20.241
R3239 a_7106_210.t0 a_7106_210.n3 13.984
R3240 a_7106_210.n10 a_7106_210.n9 13.494
R3241 a_7106_210.n6 a_7106_210.n4 8.443
R3242 a_7106_210.t0 a_7106_210.n0 8.137
R3243 a_7106_210.n8 a_7106_210.n7 1.505
R3244 a_1053_103.n5 a_1053_103.n4 66.708
R3245 a_1053_103.n2 a_1053_103.n0 32.662
R3246 a_1053_103.n5 a_1053_103.n3 19.496
R3247 a_1053_103.t0 a_1053_103.n5 13.756
R3248 a_1053_103.t0 a_1053_103.n2 3.034
R3249 a_1053_103.n2 a_1053_103.n1 0.443
R3250 a_1334_210.n8 a_1334_210.n6 185.173
R3251 a_1334_210.t0 a_1334_210.n8 75.765
R3252 a_1334_210.n3 a_1334_210.n1 74.827
R3253 a_1334_210.n3 a_1334_210.n2 27.476
R3254 a_1334_210.n6 a_1334_210.n5 22.349
R3255 a_1334_210.t0 a_1334_210.n10 20.241
R3256 a_1334_210.t0 a_1334_210.n3 13.984
R3257 a_1334_210.n10 a_1334_210.n9 13.494
R3258 a_1334_210.n6 a_1334_210.n4 8.443
R3259 a_1334_210.t0 a_1334_210.n0 8.137
R3260 a_1334_210.n8 a_1334_210.n7 1.505
R3261 a_15991_989.n3 a_15991_989.t15 512.525
R3262 a_15991_989.n1 a_15991_989.t13 477.179
R3263 a_15991_989.n6 a_15991_989.t14 454.685
R3264 a_15991_989.n2 a_15991_989.t9 440.954
R3265 a_15991_989.n6 a_15991_989.t11 428.979
R3266 a_15991_989.n1 a_15991_989.t10 406.485
R3267 a_15991_989.n5 a_15991_989.t12 378.636
R3268 a_15991_989.n3 a_15991_989.t8 371.139
R3269 a_15991_989.n7 a_15991_989.t7 255.965
R3270 a_15991_989.n12 a_15991_989.n11 252.498
R3271 a_15991_989.n7 a_15991_989.n6 227.006
R3272 a_15991_989.n16 a_15991_989.n15 161.352
R3273 a_15991_989.n14 a_15991_989.n13 151.34
R3274 a_15991_989.n14 a_15991_989.n0 95.095
R3275 a_15991_989.n17 a_15991_989.n16 95.094
R3276 a_15991_989.n13 a_15991_989.n12 83.576
R3277 a_15991_989.n4 a_15991_989.n3 77.972
R3278 a_15991_989.n16 a_15991_989.n14 66.258
R3279 a_15991_989.n5 a_15991_989.n4 55.891
R3280 a_15991_989.n11 a_15991_989.n10 30
R3281 a_15991_989.n9 a_15991_989.n8 24.383
R3282 a_15991_989.n11 a_15991_989.n9 23.684
R3283 a_15991_989.n2 a_15991_989.n1 21.4
R3284 a_15991_989.n0 a_15991_989.t6 14.282
R3285 a_15991_989.n0 a_15991_989.t5 14.282
R3286 a_15991_989.n15 a_15991_989.t2 14.282
R3287 a_15991_989.n15 a_15991_989.t3 14.282
R3288 a_15991_989.n17 a_15991_989.t0 14.282
R3289 a_15991_989.t1 a_15991_989.n17 14.282
R3290 a_15991_989.n12 a_15991_989.n7 13.335
R3291 a_15991_989.n13 a_15991_989.n5 10.343
R3292 a_15991_989.n4 a_15991_989.n2 6.833
R3293 a_15764_210.n9 a_15764_210.n7 171.558
R3294 a_15764_210.t0 a_15764_210.n9 75.765
R3295 a_15764_210.n3 a_15764_210.n1 74.827
R3296 a_15764_210.n3 a_15764_210.n2 27.476
R3297 a_15764_210.n7 a_15764_210.n6 27.2
R3298 a_15764_210.n5 a_15764_210.n4 23.498
R3299 a_15764_210.n7 a_15764_210.n5 22.4
R3300 a_15764_210.t0 a_15764_210.n11 20.241
R3301 a_15764_210.t0 a_15764_210.n3 13.984
R3302 a_15764_210.n11 a_15764_210.n10 13.494
R3303 a_15764_210.t0 a_15764_210.n0 8.137
R3304 a_15764_210.n9 a_15764_210.n8 1.505
R3305 a_2977_103.n5 a_2977_103.n4 66.708
R3306 a_2977_103.n2 a_2977_103.n0 32.662
R3307 a_2977_103.n5 a_2977_103.n3 19.496
R3308 a_2977_103.t0 a_2977_103.n5 13.756
R3309 a_2977_103.t0 a_2977_103.n2 3.034
R3310 a_2977_103.n2 a_2977_103.n1 0.443
R3311 a_3258_210.n8 a_3258_210.n6 185.173
R3312 a_3258_210.t0 a_3258_210.n8 75.765
R3313 a_3258_210.n3 a_3258_210.n1 74.827
R3314 a_3258_210.n3 a_3258_210.n2 27.476
R3315 a_3258_210.n6 a_3258_210.n5 22.349
R3316 a_3258_210.t0 a_3258_210.n10 20.241
R3317 a_3258_210.t0 a_3258_210.n3 13.984
R3318 a_3258_210.n10 a_3258_210.n9 13.494
R3319 a_3258_210.n6 a_3258_210.n4 8.443
R3320 a_3258_210.t0 a_3258_210.n0 8.137
R3321 a_3258_210.n8 a_3258_210.n7 1.505
R3322 a_6049_1050.n2 a_6049_1050.t12 512.525
R3323 a_6049_1050.n0 a_6049_1050.t10 512.525
R3324 a_6049_1050.n2 a_6049_1050.t7 371.139
R3325 a_6049_1050.n0 a_6049_1050.t11 371.139
R3326 a_6049_1050.n3 a_6049_1050.t8 306.051
R3327 a_6049_1050.n1 a_6049_1050.t9 306.051
R3328 a_6049_1050.n3 a_6049_1050.n2 290.895
R3329 a_6049_1050.n1 a_6049_1050.n0 290.895
R3330 a_6049_1050.n9 a_6049_1050.n8 252.875
R3331 a_6049_1050.n13 a_6049_1050.n9 234.54
R3332 a_6049_1050.n12 a_6049_1050.n11 161.352
R3333 a_6049_1050.n12 a_6049_1050.n10 95.095
R3334 a_6049_1050.n14 a_6049_1050.n13 95.094
R3335 a_6049_1050.n13 a_6049_1050.n12 66.258
R3336 a_6049_1050.n8 a_6049_1050.n7 30
R3337 a_6049_1050.n6 a_6049_1050.n5 24.383
R3338 a_6049_1050.n8 a_6049_1050.n6 23.684
R3339 a_6049_1050.n10 a_6049_1050.t6 14.282
R3340 a_6049_1050.n10 a_6049_1050.t5 14.282
R3341 a_6049_1050.n11 a_6049_1050.t1 14.282
R3342 a_6049_1050.n11 a_6049_1050.t0 14.282
R3343 a_6049_1050.t4 a_6049_1050.n14 14.282
R3344 a_6049_1050.n14 a_6049_1050.t3 14.282
R3345 a_6049_1050.n4 a_6049_1050.n1 8.141
R3346 a_6049_1050.n9 a_6049_1050.n4 5.965
R3347 a_6049_1050.n4 a_6049_1050.n3 4.65
R3348 a_13840_210.n10 a_13840_210.n8 171.558
R3349 a_13840_210.n8 a_13840_210.t1 75.764
R3350 a_13840_210.n3 a_13840_210.n2 27.476
R3351 a_13840_210.n10 a_13840_210.n9 27.2
R3352 a_13840_210.n11 a_13840_210.n0 23.498
R3353 a_13840_210.n11 a_13840_210.n10 22.4
R3354 a_13840_210.t1 a_13840_210.n5 20.241
R3355 a_13840_210.n7 a_13840_210.n6 19.952
R3356 a_13840_210.t1 a_13840_210.n3 13.984
R3357 a_13840_210.n5 a_13840_210.n4 13.494
R3358 a_13840_210.t1 a_13840_210.n1 7.04
R3359 a_13840_210.n8 a_13840_210.n7 1.505
R3360 a_7973_1050.n2 a_7973_1050.t7 512.525
R3361 a_7973_1050.n2 a_7973_1050.t8 371.139
R3362 a_7973_1050.n3 a_7973_1050.t9 305.674
R3363 a_7973_1050.n3 a_7973_1050.n2 291.272
R3364 a_7973_1050.n8 a_7973_1050.n7 252.498
R3365 a_7973_1050.n9 a_7973_1050.n8 234.917
R3366 a_7973_1050.n11 a_7973_1050.n10 161.352
R3367 a_7973_1050.n9 a_7973_1050.n1 95.095
R3368 a_7973_1050.n10 a_7973_1050.n0 95.095
R3369 a_7973_1050.n10 a_7973_1050.n9 66.258
R3370 a_7973_1050.n7 a_7973_1050.n6 30
R3371 a_7973_1050.n5 a_7973_1050.n4 24.383
R3372 a_7973_1050.n7 a_7973_1050.n5 23.684
R3373 a_7973_1050.n1 a_7973_1050.t5 14.282
R3374 a_7973_1050.n1 a_7973_1050.t6 14.282
R3375 a_7973_1050.n0 a_7973_1050.t3 14.282
R3376 a_7973_1050.n0 a_7973_1050.t2 14.282
R3377 a_7973_1050.t1 a_7973_1050.n11 14.282
R3378 a_7973_1050.n11 a_7973_1050.t0 14.282
R3379 a_7973_1050.n8 a_7973_1050.n3 10.615
R3380 a_17533_1051.n2 a_17533_1051.t0 179.895
R3381 a_17533_1051.n5 a_17533_1051.n4 157.021
R3382 a_17533_1051.n4 a_17533_1051.n0 124.955
R3383 a_17533_1051.n3 a_17533_1051.n2 106.183
R3384 a_17533_1051.n2 a_17533_1051.n1 99.355
R3385 a_17533_1051.n4 a_17533_1051.n3 82.65
R3386 a_17533_1051.n3 a_17533_1051.t2 73.712
R3387 a_17533_1051.n0 a_17533_1051.t6 14.282
R3388 a_17533_1051.n0 a_17533_1051.t7 14.282
R3389 a_17533_1051.n1 a_17533_1051.t1 14.282
R3390 a_17533_1051.n1 a_17533_1051.t3 14.282
R3391 a_17533_1051.n5 a_17533_1051.t4 14.282
R3392 a_17533_1051.t5 a_17533_1051.n5 14.282
R3393 a_4125_1050.n2 a_4125_1050.t8 512.525
R3394 a_4125_1050.n2 a_4125_1050.t9 371.139
R3395 a_4125_1050.n3 a_4125_1050.t7 361.392
R3396 a_4125_1050.n5 a_4125_1050.n4 329.955
R3397 a_4125_1050.n3 a_4125_1050.n2 235.554
R3398 a_4125_1050.n6 a_4125_1050.n5 179.199
R3399 a_4125_1050.n8 a_4125_1050.n7 161.352
R3400 a_4125_1050.n6 a_4125_1050.n1 95.095
R3401 a_4125_1050.n7 a_4125_1050.n0 95.095
R3402 a_4125_1050.n7 a_4125_1050.n6 66.258
R3403 a_4125_1050.n1 a_4125_1050.t6 14.282
R3404 a_4125_1050.n1 a_4125_1050.t1 14.282
R3405 a_4125_1050.n0 a_4125_1050.t4 14.282
R3406 a_4125_1050.n0 a_4125_1050.t5 14.282
R3407 a_4125_1050.n8 a_4125_1050.t2 14.282
R3408 a_4125_1050.t3 a_4125_1050.n8 14.282
R3409 a_4125_1050.n5 a_4125_1050.n3 10.615
R3410 a_4447_989.n3 a_4447_989.t10 512.525
R3411 a_4447_989.n2 a_4447_989.t9 512.525
R3412 a_4447_989.n7 a_4447_989.t7 454.685
R3413 a_4447_989.n7 a_4447_989.t13 428.979
R3414 a_4447_989.n3 a_4447_989.t14 371.139
R3415 a_4447_989.n2 a_4447_989.t15 371.139
R3416 a_4447_989.n4 a_4447_989.n3 343.521
R3417 a_4447_989.n13 a_4447_989.n12 295.88
R3418 a_4447_989.n8 a_4447_989.t12 272.577
R3419 a_4447_989.n6 a_4447_989.n2 259.945
R3420 a_4447_989.n14 a_4447_989.n13 207.058
R3421 a_4447_989.n8 a_4447_989.n7 199.147
R3422 a_4447_989.n4 a_4447_989.t8 172.106
R3423 a_4447_989.n5 a_4447_989.t11 165.68
R3424 a_4447_989.n16 a_4447_989.n15 161.352
R3425 a_4447_989.n14 a_4447_989.n1 95.095
R3426 a_4447_989.n15 a_4447_989.n0 95.095
R3427 a_4447_989.n6 a_4447_989.n5 83.576
R3428 a_4447_989.n15 a_4447_989.n14 66.258
R3429 a_4447_989.n9 a_4447_989.n6 51.943
R3430 a_4447_989.n12 a_4447_989.n11 22.578
R3431 a_4447_989.n1 a_4447_989.t6 14.282
R3432 a_4447_989.n1 a_4447_989.t5 14.282
R3433 a_4447_989.n0 a_4447_989.t3 14.282
R3434 a_4447_989.n0 a_4447_989.t2 14.282
R3435 a_4447_989.t1 a_4447_989.n16 14.282
R3436 a_4447_989.n16 a_4447_989.t0 14.282
R3437 a_4447_989.n5 a_4447_989.n4 10.343
R3438 a_4447_989.n9 a_4447_989.n8 8.685
R3439 a_4447_989.n12 a_4447_989.n10 8.58
R3440 a_4447_989.n13 a_4447_989.n9 4.65
R3441 a_18760_101.n3 a_18760_101.n1 42.788
R3442 a_18760_101.t0 a_18760_101.n0 8.137
R3443 a_18760_101.n3 a_18760_101.n2 4.665
R3444 a_18760_101.t0 a_18760_101.n3 0.06
R3445 a_18094_101.n2 a_18094_101.n0 42.761
R3446 a_18094_101.n2 a_18094_101.n1 2.167
R3447 a_18094_101.t0 a_18094_101.n2 0.099
R3448 a_18197_1051.n2 a_18197_1051.t6 179.895
R3449 a_18197_1051.n4 a_18197_1051.n0 165.613
R3450 a_18197_1051.n5 a_18197_1051.n4 142.653
R3451 a_18197_1051.n3 a_18197_1051.n2 106.183
R3452 a_18197_1051.n2 a_18197_1051.n1 99.355
R3453 a_18197_1051.n4 a_18197_1051.n3 82.665
R3454 a_18197_1051.n3 a_18197_1051.t2 73.712
R3455 a_18197_1051.n1 a_18197_1051.t7 14.282
R3456 a_18197_1051.n1 a_18197_1051.t3 14.282
R3457 a_18197_1051.n0 a_18197_1051.t4 14.282
R3458 a_18197_1051.n0 a_18197_1051.t5 14.282
R3459 a_18197_1051.n5 a_18197_1051.t0 14.282
R3460 a_18197_1051.t1 a_18197_1051.n5 14.282
R3461 a_5863_103.t0 a_5863_103.n7 59.616
R3462 a_5863_103.n4 a_5863_103.n2 54.496
R3463 a_5863_103.n4 a_5863_103.n3 54.496
R3464 a_5863_103.n1 a_5863_103.n0 24.679
R3465 a_5863_103.n6 a_5863_103.n4 7.859
R3466 a_5863_103.t0 a_5863_103.n1 7.505
R3467 a_5863_103.t0 a_5863_103.n6 3.034
R3468 a_5863_103.n6 a_5863_103.n5 0.443
R3469 a_6144_210.n8 a_6144_210.n6 185.173
R3470 a_6144_210.t0 a_6144_210.n8 75.765
R3471 a_6144_210.n3 a_6144_210.n1 74.827
R3472 a_6144_210.n3 a_6144_210.n2 27.476
R3473 a_6144_210.n6 a_6144_210.n5 22.349
R3474 a_6144_210.t0 a_6144_210.n10 20.241
R3475 a_6144_210.t0 a_6144_210.n3 13.984
R3476 a_6144_210.n10 a_6144_210.n9 13.494
R3477 a_6144_210.n6 a_6144_210.n4 8.443
R3478 a_6144_210.t0 a_6144_210.n0 8.137
R3479 a_6144_210.n8 a_6144_210.n7 1.505
R3480 D.n5 D.t7 512.525
R3481 D.n2 D.t6 512.525
R3482 D.n0 D.t8 512.525
R3483 D.n6 D.t4 417.109
R3484 D.n3 D.t1 417.109
R3485 D.n1 D.t0 417.109
R3486 D.n5 D.t3 371.139
R3487 D.n2 D.t2 371.139
R3488 D.n0 D.t5 371.139
R3489 D.n6 D.n5 179.837
R3490 D.n3 D.n2 179.837
R3491 D.n1 D.n0 179.837
R3492 D.n4 D.n1 25.825
R3493 D.n7 D.n4 21.175
R3494 D.n4 D.n3 4.65
R3495 D.n7 D.n6 4.65
R3496 D.n7 D 0.046
R3497 a_11635_103.n5 a_11635_103.n4 66.708
R3498 a_11635_103.n2 a_11635_103.n0 32.662
R3499 a_11635_103.n5 a_11635_103.n3 19.496
R3500 a_11635_103.t0 a_11635_103.n5 13.756
R3501 a_11635_103.t0 a_11635_103.n2 3.034
R3502 a_11635_103.n2 a_11635_103.n1 0.443
R3503 a_16726_210.n10 a_16726_210.n8 171.558
R3504 a_16726_210.n8 a_16726_210.t1 75.764
R3505 a_16726_210.n3 a_16726_210.n2 27.476
R3506 a_16726_210.n10 a_16726_210.n9 27.2
R3507 a_16726_210.n11 a_16726_210.n0 23.498
R3508 a_16726_210.n11 a_16726_210.n10 22.4
R3509 a_16726_210.t1 a_16726_210.n5 20.241
R3510 a_16726_210.n7 a_16726_210.n6 19.952
R3511 a_16726_210.t1 a_16726_210.n3 13.984
R3512 a_16726_210.n5 a_16726_210.n4 13.494
R3513 a_16726_210.t1 a_16726_210.n1 7.04
R3514 a_16726_210.n8 a_16726_210.n7 1.505
R3515 a_7787_103.n5 a_7787_103.n4 66.708
R3516 a_7787_103.n2 a_7787_103.n0 32.662
R3517 a_7787_103.n5 a_7787_103.n3 19.496
R3518 a_7787_103.t0 a_7787_103.n5 13.756
R3519 a_7787_103.t0 a_7787_103.n2 3.034
R3520 a_7787_103.n2 a_7787_103.n1 0.443
R3521 a_8068_210.n10 a_8068_210.n8 171.558
R3522 a_8068_210.n8 a_8068_210.t1 75.764
R3523 a_8068_210.n11 a_8068_210.n0 49.6
R3524 a_8068_210.n3 a_8068_210.n2 27.476
R3525 a_8068_210.n10 a_8068_210.n9 27.2
R3526 a_8068_210.n11 a_8068_210.n10 22.4
R3527 a_8068_210.t1 a_8068_210.n5 20.241
R3528 a_8068_210.n7 a_8068_210.n6 19.952
R3529 a_8068_210.t1 a_8068_210.n3 13.984
R3530 a_8068_210.n5 a_8068_210.n4 13.494
R3531 a_8068_210.t1 a_8068_210.n1 7.04
R3532 a_8068_210.n8 a_8068_210.n7 1.505
R3533 a_9711_103.n5 a_9711_103.n4 66.708
R3534 a_9711_103.n2 a_9711_103.n0 32.662
R3535 a_9711_103.n5 a_9711_103.n3 19.496
R3536 a_9711_103.t0 a_9711_103.n5 13.756
R3537 a_9711_103.t0 a_9711_103.n2 3.034
R3538 a_9711_103.n2 a_9711_103.n1 0.443
R3539 a_17708_209.n1 a_17708_209.t7 512.525
R3540 a_17708_209.n1 a_17708_209.t9 371.139
R3541 a_17708_209.n2 a_17708_209.t8 338.57
R3542 a_17708_209.n13 a_17708_209.n12 227.387
R3543 a_17708_209.n2 a_17708_209.n1 191.629
R3544 a_17708_209.n15 a_17708_209.n14 165.613
R3545 a_17708_209.n14 a_17708_209.n13 132.893
R3546 a_17708_209.n12 a_17708_209.n11 127.909
R3547 a_17708_209.n10 a_17708_209.n5 126.225
R3548 a_17708_209.n10 a_17708_209.n9 112.771
R3549 a_17708_209.n14 a_17708_209.n0 99.355
R3550 a_17708_209.n9 a_17708_209.n8 30
R3551 a_17708_209.n7 a_17708_209.n6 24.383
R3552 a_17708_209.n9 a_17708_209.n7 23.684
R3553 a_17708_209.n5 a_17708_209.n4 22.578
R3554 a_17708_209.n0 a_17708_209.t3 14.282
R3555 a_17708_209.n0 a_17708_209.t4 14.282
R3556 a_17708_209.t1 a_17708_209.n15 14.282
R3557 a_17708_209.n15 a_17708_209.t0 14.282
R3558 a_17708_209.n13 a_17708_209.n2 10.343
R3559 a_17708_209.n5 a_17708_209.n3 8.58
R3560 a_17708_209.n12 a_17708_209.n10 7.053
R3561 Q.n2 Q.n1 349.908
R3562 Q.n2 Q.n0 215.564
R3563 Q.n0 Q.t1 14.282
R3564 Q.n0 Q.t0 14.282
R3565 Q.n3 Q.n2 4.65
R3566 Q.n3 Q 0.046
R3567 a_372_210.n9 a_372_210.n7 171.558
R3568 a_372_210.t0 a_372_210.n9 75.765
R3569 a_372_210.n3 a_372_210.n1 74.827
R3570 a_372_210.n3 a_372_210.n2 27.476
R3571 a_372_210.n7 a_372_210.n6 27.2
R3572 a_372_210.n5 a_372_210.n4 23.498
R3573 a_372_210.n7 a_372_210.n5 22.4
R3574 a_372_210.t0 a_372_210.n11 20.241
R3575 a_372_210.t0 a_372_210.n3 13.984
R3576 a_372_210.n11 a_372_210.n10 13.494
R3577 a_372_210.t0 a_372_210.n0 8.137
R3578 a_372_210.n9 a_372_210.n8 1.505
R3579 a_8749_103.n5 a_8749_103.n4 66.708
R3580 a_8749_103.n2 a_8749_103.n0 25.439
R3581 a_8749_103.n5 a_8749_103.n3 19.496
R3582 a_8749_103.t0 a_8749_103.n5 13.756
R3583 a_8749_103.n2 a_8749_103.n1 2.455
R3584 a_8749_103.t0 a_8749_103.n2 0.246
R3585 a_12597_103.n5 a_12597_103.n4 66.708
R3586 a_12597_103.n2 a_12597_103.n0 32.662
R3587 a_12597_103.n5 a_12597_103.n3 19.496
R3588 a_12597_103.t0 a_12597_103.n5 13.756
R3589 a_12597_103.t0 a_12597_103.n2 3.034
R3590 a_12597_103.n2 a_12597_103.n1 0.443
R3591 a_14521_103.n5 a_14521_103.n4 66.708
R3592 a_14521_103.n2 a_14521_103.n0 25.439
R3593 a_14521_103.n5 a_14521_103.n3 19.496
R3594 a_14521_103.t0 a_14521_103.n5 13.756
R3595 a_14521_103.n2 a_14521_103.n1 2.455
R3596 a_14521_103.t0 a_14521_103.n2 0.246
R3597 a_10673_103.t0 a_10673_103.n7 59.616
R3598 a_10673_103.n4 a_10673_103.n2 54.496
R3599 a_10673_103.n4 a_10673_103.n3 54.496
R3600 a_10673_103.n1 a_10673_103.n0 24.679
R3601 a_10673_103.n6 a_10673_103.n4 7.859
R3602 a_10673_103.t0 a_10673_103.n1 7.505
R3603 a_10673_103.t0 a_10673_103.n6 3.034
R3604 a_10673_103.n6 a_10673_103.n5 0.443
R3605 a_91_103.n5 a_91_103.n4 66.708
R3606 a_91_103.n2 a_91_103.n0 25.439
R3607 a_91_103.n5 a_91_103.n3 19.496
R3608 a_91_103.t0 a_91_103.n5 13.756
R3609 a_91_103.n2 a_91_103.n1 2.455
R3610 a_91_103.t0 a_91_103.n2 0.246
R3611 a_11916_210.n8 a_11916_210.n6 185.173
R3612 a_11916_210.t0 a_11916_210.n8 75.765
R3613 a_11916_210.n3 a_11916_210.n1 74.827
R3614 a_11916_210.n3 a_11916_210.n2 27.476
R3615 a_11916_210.n6 a_11916_210.n5 22.349
R3616 a_11916_210.t0 a_11916_210.n10 20.241
R3617 a_11916_210.t0 a_11916_210.n3 13.984
R3618 a_11916_210.n10 a_11916_210.n9 13.494
R3619 a_11916_210.n6 a_11916_210.n4 8.443
R3620 a_11916_210.t0 a_11916_210.n0 8.137
R3621 a_11916_210.n8 a_11916_210.n7 1.505
R3622 a_9992_210.n8 a_9992_210.n6 185.173
R3623 a_9992_210.t0 a_9992_210.n8 75.765
R3624 a_9992_210.n3 a_9992_210.n1 74.827
R3625 a_9992_210.n3 a_9992_210.n2 27.476
R3626 a_9992_210.n6 a_9992_210.n5 22.349
R3627 a_9992_210.t0 a_9992_210.n10 20.241
R3628 a_9992_210.t0 a_9992_210.n3 13.984
R3629 a_9992_210.n10 a_9992_210.n9 13.494
R3630 a_9992_210.n6 a_9992_210.n4 8.443
R3631 a_9992_210.t0 a_9992_210.n0 8.137
R3632 a_9992_210.n8 a_9992_210.n7 1.505
R3633 a_17428_101.n3 a_17428_101.n2 62.817
R3634 a_17428_101.n11 a_17428_101.n10 46.054
R3635 a_17428_101.n7 a_17428_101.n6 38.626
R3636 a_17428_101.n6 a_17428_101.n5 35.955
R3637 a_17428_101.n12 a_17428_101.n11 27.923
R3638 a_17428_101.n3 a_17428_101.n1 26.202
R3639 a_17428_101.t0 a_17428_101.n3 19.737
R3640 a_17428_101.t0 a_17428_101.n4 7.273
R3641 a_17428_101.n9 a_17428_101.n8 6.883
R3642 a_17428_101.t0 a_17428_101.n0 6.109
R3643 a_17428_101.t1 a_17428_101.n7 4.864
R3644 a_17428_101.t0 a_17428_101.n13 2.074
R3645 a_17428_101.t1 a_17428_101.n9 1.179
R3646 a_17428_101.t1 a_17428_101.n12 0.958
R3647 a_17428_101.n13 a_17428_101.t1 0.937
R3648 a_13559_103.t0 a_13559_103.n7 59.616
R3649 a_13559_103.n4 a_13559_103.n2 54.496
R3650 a_13559_103.n4 a_13559_103.n3 54.496
R3651 a_13559_103.n1 a_13559_103.n0 24.679
R3652 a_13559_103.t0 a_13559_103.n1 7.505
R3653 a_13559_103.n6 a_13559_103.n5 2.455
R3654 a_13559_103.n6 a_13559_103.n4 0.636
R3655 a_13559_103.t0 a_13559_103.n6 0.246
R3656 a_15483_103.n5 a_15483_103.n4 66.708
R3657 a_15483_103.n2 a_15483_103.n0 25.439
R3658 a_15483_103.n5 a_15483_103.n3 19.496
R3659 a_15483_103.t0 a_15483_103.n5 13.756
R3660 a_15483_103.n2 a_15483_103.n1 2.455
R3661 a_15483_103.t0 a_15483_103.n2 0.246
R3662 a_10954_210.n10 a_10954_210.n8 171.558
R3663 a_10954_210.n8 a_10954_210.t1 75.764
R3664 a_10954_210.n11 a_10954_210.n0 49.6
R3665 a_10954_210.n3 a_10954_210.n2 27.476
R3666 a_10954_210.n10 a_10954_210.n9 27.2
R3667 a_10954_210.n11 a_10954_210.n10 22.4
R3668 a_10954_210.t1 a_10954_210.n5 20.241
R3669 a_10954_210.n7 a_10954_210.n6 19.952
R3670 a_10954_210.t1 a_10954_210.n3 13.984
R3671 a_10954_210.n5 a_10954_210.n4 13.494
R3672 a_10954_210.t1 a_10954_210.n1 7.04
R3673 a_10954_210.n8 a_10954_210.n7 1.505
R3674 a_16445_103.t0 a_16445_103.n7 59.616
R3675 a_16445_103.n4 a_16445_103.n2 54.496
R3676 a_16445_103.n4 a_16445_103.n3 54.496
R3677 a_16445_103.n1 a_16445_103.n0 24.679
R3678 a_16445_103.t0 a_16445_103.n1 7.505
R3679 a_16445_103.n6 a_16445_103.n5 2.455
R3680 a_16445_103.n6 a_16445_103.n4 0.636
R3681 a_16445_103.t0 a_16445_103.n6 0.246
R3682 a_12878_210.n10 a_12878_210.n8 171.558
R3683 a_12878_210.n8 a_12878_210.t1 75.764
R3684 a_12878_210.n11 a_12878_210.n0 49.6
R3685 a_12878_210.n3 a_12878_210.n2 27.476
R3686 a_12878_210.n10 a_12878_210.n9 27.2
R3687 a_12878_210.n11 a_12878_210.n10 22.4
R3688 a_12878_210.t1 a_12878_210.n5 20.241
R3689 a_12878_210.n7 a_12878_210.n6 19.952
R3690 a_12878_210.t1 a_12878_210.n3 13.984
R3691 a_12878_210.n5 a_12878_210.n4 13.494
R3692 a_12878_210.t1 a_12878_210.n1 7.04
R3693 a_12878_210.n8 a_12878_210.n7 1.505
R3694 a_2296_210.n10 a_2296_210.n8 171.558
R3695 a_2296_210.n8 a_2296_210.t1 75.764
R3696 a_2296_210.n3 a_2296_210.n2 27.476
R3697 a_2296_210.n10 a_2296_210.n9 27.2
R3698 a_2296_210.n11 a_2296_210.n0 23.498
R3699 a_2296_210.n11 a_2296_210.n10 22.4
R3700 a_2296_210.t1 a_2296_210.n5 20.241
R3701 a_2296_210.n7 a_2296_210.n6 19.952
R3702 a_2296_210.t1 a_2296_210.n3 13.984
R3703 a_2296_210.n5 a_2296_210.n4 13.494
R3704 a_2296_210.t1 a_2296_210.n1 7.04
R3705 a_2296_210.n8 a_2296_210.n7 1.505
R3706 a_4220_210.n8 a_4220_210.n6 185.173
R3707 a_4220_210.t0 a_4220_210.n8 75.765
R3708 a_4220_210.n3 a_4220_210.n1 74.827
R3709 a_4220_210.n3 a_4220_210.n2 27.476
R3710 a_4220_210.n6 a_4220_210.n5 22.349
R3711 a_4220_210.t0 a_4220_210.n10 20.241
R3712 a_4220_210.t0 a_4220_210.n3 13.984
R3713 a_4220_210.n10 a_4220_210.n9 13.494
R3714 a_4220_210.n6 a_4220_210.n4 8.443
R3715 a_4220_210.t0 a_4220_210.n0 8.137
R3716 a_4220_210.n8 a_4220_210.n7 1.505
R3717 a_2015_103.t0 a_2015_103.n7 59.616
R3718 a_2015_103.n4 a_2015_103.n2 54.496
R3719 a_2015_103.n4 a_2015_103.n3 54.496
R3720 a_2015_103.n1 a_2015_103.n0 24.679
R3721 a_2015_103.t0 a_2015_103.n1 7.505
R3722 a_2015_103.n6 a_2015_103.n5 2.455
R3723 a_2015_103.n6 a_2015_103.n4 0.636
R3724 a_2015_103.t0 a_2015_103.n6 0.246
C11 SN GND 7.80fF
C12 RN GND 8.38fF
C13 VDD GND 32.50fF
C14 a_2015_103.n0 GND 0.08fF
C15 a_2015_103.n1 GND 0.07fF
C16 a_2015_103.n2 GND 0.04fF
C17 a_2015_103.n3 GND 0.06fF
C18 a_2015_103.n4 GND 0.03fF
C19 a_2015_103.n5 GND 0.04fF
C20 a_2015_103.n7 GND 0.08fF
C21 a_4220_210.n0 GND 0.07fF
C22 a_4220_210.n1 GND 0.09fF
C23 a_4220_210.n2 GND 0.12fF
C24 a_4220_210.n3 GND 0.08fF
C25 a_4220_210.n4 GND 0.02fF
C26 a_4220_210.n5 GND 0.03fF
C27 a_4220_210.n6 GND 0.05fF
C28 a_4220_210.n7 GND 0.02fF
C29 a_4220_210.n8 GND 0.14fF
C30 a_4220_210.n9 GND 0.08fF
C31 a_4220_210.n10 GND 0.02fF
C32 a_4220_210.t0 GND 0.31fF
C33 a_2296_210.n0 GND 0.02fF
C34 a_2296_210.n1 GND 0.09fF
C35 a_2296_210.n2 GND 0.12fF
C36 a_2296_210.n3 GND 0.08fF
C37 a_2296_210.n4 GND 0.08fF
C38 a_2296_210.n5 GND 0.02fF
C39 a_2296_210.t1 GND 0.29fF
C40 a_2296_210.n6 GND 0.09fF
C41 a_2296_210.n7 GND 0.02fF
C42 a_2296_210.n8 GND 0.13fF
C43 a_2296_210.n9 GND 0.02fF
C44 a_2296_210.n10 GND 0.03fF
C45 a_2296_210.n11 GND 0.03fF
C46 a_12878_210.n0 GND 0.02fF
C47 a_12878_210.n1 GND 0.09fF
C48 a_12878_210.n2 GND 0.12fF
C49 a_12878_210.n3 GND 0.08fF
C50 a_12878_210.n4 GND 0.08fF
C51 a_12878_210.n5 GND 0.02fF
C52 a_12878_210.t1 GND 0.29fF
C53 a_12878_210.n6 GND 0.09fF
C54 a_12878_210.n7 GND 0.02fF
C55 a_12878_210.n8 GND 0.13fF
C56 a_12878_210.n9 GND 0.02fF
C57 a_12878_210.n10 GND 0.03fF
C58 a_12878_210.n11 GND 0.02fF
C59 a_16445_103.n0 GND 0.08fF
C60 a_16445_103.n1 GND 0.07fF
C61 a_16445_103.n2 GND 0.04fF
C62 a_16445_103.n3 GND 0.06fF
C63 a_16445_103.n4 GND 0.03fF
C64 a_16445_103.n5 GND 0.04fF
C65 a_16445_103.n7 GND 0.08fF
C66 a_10954_210.n0 GND 0.02fF
C67 a_10954_210.n1 GND 0.09fF
C68 a_10954_210.n2 GND 0.12fF
C69 a_10954_210.n3 GND 0.08fF
C70 a_10954_210.n4 GND 0.08fF
C71 a_10954_210.n5 GND 0.02fF
C72 a_10954_210.t1 GND 0.29fF
C73 a_10954_210.n6 GND 0.09fF
C74 a_10954_210.n7 GND 0.02fF
C75 a_10954_210.n8 GND 0.13fF
C76 a_10954_210.n9 GND 0.02fF
C77 a_10954_210.n10 GND 0.03fF
C78 a_10954_210.n11 GND 0.02fF
C79 a_15483_103.n0 GND 0.11fF
C80 a_15483_103.n1 GND 0.04fF
C81 a_15483_103.n2 GND 0.03fF
C82 a_15483_103.n3 GND 0.07fF
C83 a_15483_103.n4 GND 0.08fF
C84 a_15483_103.n5 GND 0.03fF
C85 a_13559_103.n0 GND 0.08fF
C86 a_13559_103.n1 GND 0.07fF
C87 a_13559_103.n2 GND 0.04fF
C88 a_13559_103.n3 GND 0.06fF
C89 a_13559_103.n4 GND 0.03fF
C90 a_13559_103.n5 GND 0.04fF
C91 a_13559_103.n7 GND 0.08fF
C92 a_17428_101.n0 GND 0.02fF
C93 a_17428_101.n1 GND 0.09fF
C94 a_17428_101.n2 GND 0.07fF
C95 a_17428_101.n3 GND 0.03fF
C96 a_17428_101.n4 GND 0.01fF
C97 a_17428_101.n5 GND 0.03fF
C98 a_17428_101.n6 GND 0.04fF
C99 a_17428_101.n7 GND 0.02fF
C100 a_17428_101.n8 GND 0.04fF
C101 a_17428_101.n9 GND 0.08fF
C102 a_17428_101.n10 GND 0.04fF
C103 a_17428_101.n11 GND 0.12fF
C104 a_17428_101.n12 GND 0.14fF
C105 a_17428_101.t1 GND 0.16fF
C106 a_17428_101.n13 GND 0.01fF
C107 a_9992_210.n0 GND 0.07fF
C108 a_9992_210.n1 GND 0.09fF
C109 a_9992_210.n2 GND 0.12fF
C110 a_9992_210.n3 GND 0.08fF
C111 a_9992_210.n4 GND 0.02fF
C112 a_9992_210.n5 GND 0.03fF
C113 a_9992_210.n6 GND 0.05fF
C114 a_9992_210.n7 GND 0.02fF
C115 a_9992_210.n8 GND 0.14fF
C116 a_9992_210.n9 GND 0.08fF
C117 a_9992_210.n10 GND 0.02fF
C118 a_9992_210.t0 GND 0.31fF
C119 a_11916_210.n0 GND 0.07fF
C120 a_11916_210.n1 GND 0.09fF
C121 a_11916_210.n2 GND 0.12fF
C122 a_11916_210.n3 GND 0.08fF
C123 a_11916_210.n4 GND 0.02fF
C124 a_11916_210.n5 GND 0.03fF
C125 a_11916_210.n6 GND 0.05fF
C126 a_11916_210.n7 GND 0.02fF
C127 a_11916_210.n8 GND 0.14fF
C128 a_11916_210.n9 GND 0.08fF
C129 a_11916_210.n10 GND 0.02fF
C130 a_11916_210.t0 GND 0.31fF
C131 a_91_103.n0 GND 0.10fF
C132 a_91_103.n1 GND 0.03fF
C133 a_91_103.n2 GND 0.03fF
C134 a_91_103.n3 GND 0.07fF
C135 a_91_103.n4 GND 0.08fF
C136 a_91_103.n5 GND 0.03fF
C137 a_10673_103.n0 GND 0.08fF
C138 a_10673_103.n1 GND 0.07fF
C139 a_10673_103.n2 GND 0.04fF
C140 a_10673_103.n3 GND 0.06fF
C141 a_10673_103.n4 GND 0.11fF
C142 a_10673_103.n5 GND 0.04fF
C143 a_10673_103.n7 GND 0.08fF
C144 a_14521_103.n0 GND 0.11fF
C145 a_14521_103.n1 GND 0.04fF
C146 a_14521_103.n2 GND 0.03fF
C147 a_14521_103.n3 GND 0.07fF
C148 a_14521_103.n4 GND 0.08fF
C149 a_14521_103.n5 GND 0.03fF
C150 a_12597_103.n0 GND 0.13fF
C151 a_12597_103.n1 GND 0.04fF
C152 a_12597_103.n2 GND 0.09fF
C153 a_12597_103.n3 GND 0.07fF
C154 a_12597_103.n4 GND 0.08fF
C155 a_12597_103.n5 GND 0.03fF
C156 a_8749_103.n0 GND 0.11fF
C157 a_8749_103.n1 GND 0.04fF
C158 a_8749_103.n2 GND 0.03fF
C159 a_8749_103.n3 GND 0.07fF
C160 a_8749_103.n4 GND 0.08fF
C161 a_8749_103.n5 GND 0.03fF
C162 a_372_210.n0 GND 0.07fF
C163 a_372_210.n1 GND 0.09fF
C164 a_372_210.n2 GND 0.12fF
C165 a_372_210.n3 GND 0.08fF
C166 a_372_210.n4 GND 0.02fF
C167 a_372_210.n5 GND 0.03fF
C168 a_372_210.n6 GND 0.02fF
C169 a_372_210.n7 GND 0.03fF
C170 a_372_210.n8 GND 0.02fF
C171 a_372_210.n9 GND 0.13fF
C172 a_372_210.n10 GND 0.08fF
C173 a_372_210.n11 GND 0.02fF
C174 a_372_210.t0 GND 0.31fF
C175 Q.n0 GND 0.58fF
C176 Q.n1 GND 0.36fF
C177 Q.n2 GND 0.66fF
C178 Q.n3 GND 0.01fF
C179 a_17708_209.n0 GND 0.26fF
C180 a_17708_209.n1 GND 0.24fF
C181 a_17708_209.n2 GND 0.47fF
C182 a_17708_209.n3 GND 0.03fF
C183 a_17708_209.n4 GND 0.04fF
C184 a_17708_209.n5 GND 0.05fF
C185 a_17708_209.n6 GND 0.03fF
C186 a_17708_209.n7 GND 0.04fF
C187 a_17708_209.n8 GND 0.03fF
C188 a_17708_209.n9 GND 0.04fF
C189 a_17708_209.n10 GND 0.95fF
C190 a_17708_209.n11 GND 0.12fF
C191 a_17708_209.n12 GND 0.34fF
C192 a_17708_209.n13 GND 0.43fF
C193 a_17708_209.n14 GND 0.41fF
C194 a_17708_209.n15 GND 0.34fF
C195 a_9711_103.n0 GND 0.13fF
C196 a_9711_103.n1 GND 0.04fF
C197 a_9711_103.n2 GND 0.09fF
C198 a_9711_103.n3 GND 0.07fF
C199 a_9711_103.n4 GND 0.08fF
C200 a_9711_103.n5 GND 0.03fF
C201 a_8068_210.n0 GND 0.02fF
C202 a_8068_210.n1 GND 0.09fF
C203 a_8068_210.n2 GND 0.12fF
C204 a_8068_210.n3 GND 0.08fF
C205 a_8068_210.n4 GND 0.08fF
C206 a_8068_210.n5 GND 0.02fF
C207 a_8068_210.t1 GND 0.29fF
C208 a_8068_210.n6 GND 0.09fF
C209 a_8068_210.n7 GND 0.02fF
C210 a_8068_210.n8 GND 0.13fF
C211 a_8068_210.n9 GND 0.02fF
C212 a_8068_210.n10 GND 0.03fF
C213 a_8068_210.n11 GND 0.02fF
C214 a_7787_103.n0 GND 0.13fF
C215 a_7787_103.n1 GND 0.04fF
C216 a_7787_103.n2 GND 0.09fF
C217 a_7787_103.n3 GND 0.07fF
C218 a_7787_103.n4 GND 0.08fF
C219 a_7787_103.n5 GND 0.03fF
C220 a_16726_210.n0 GND 0.02fF
C221 a_16726_210.n1 GND 0.09fF
C222 a_16726_210.n2 GND 0.12fF
C223 a_16726_210.n3 GND 0.08fF
C224 a_16726_210.n4 GND 0.08fF
C225 a_16726_210.n5 GND 0.02fF
C226 a_16726_210.t1 GND 0.29fF
C227 a_16726_210.n6 GND 0.09fF
C228 a_16726_210.n7 GND 0.02fF
C229 a_16726_210.n8 GND 0.13fF
C230 a_16726_210.n9 GND 0.02fF
C231 a_16726_210.n10 GND 0.03fF
C232 a_16726_210.n11 GND 0.03fF
C233 a_11635_103.n0 GND 0.13fF
C234 a_11635_103.n1 GND 0.04fF
C235 a_11635_103.n2 GND 0.09fF
C236 a_11635_103.n3 GND 0.07fF
C237 a_11635_103.n4 GND 0.08fF
C238 a_11635_103.n5 GND 0.03fF
C239 a_6144_210.n0 GND 0.07fF
C240 a_6144_210.n1 GND 0.09fF
C241 a_6144_210.n2 GND 0.12fF
C242 a_6144_210.n3 GND 0.08fF
C243 a_6144_210.n4 GND 0.02fF
C244 a_6144_210.n5 GND 0.03fF
C245 a_6144_210.n6 GND 0.05fF
C246 a_6144_210.n7 GND 0.02fF
C247 a_6144_210.n8 GND 0.14fF
C248 a_6144_210.n9 GND 0.08fF
C249 a_6144_210.n10 GND 0.02fF
C250 a_6144_210.t0 GND 0.31fF
C251 a_5863_103.n0 GND 0.08fF
C252 a_5863_103.n1 GND 0.07fF
C253 a_5863_103.n2 GND 0.04fF
C254 a_5863_103.n3 GND 0.06fF
C255 a_5863_103.n4 GND 0.11fF
C256 a_5863_103.n5 GND 0.04fF
C257 a_5863_103.n7 GND 0.08fF
C258 a_18197_1051.n0 GND 0.37fF
C259 a_18197_1051.n1 GND 0.29fF
C260 a_18197_1051.n2 GND 0.46fF
C261 a_18197_1051.n3 GND 0.27fF
C262 a_18197_1051.n4 GND 0.71fF
C263 a_18197_1051.n5 GND 0.28fF
C264 a_18094_101.n0 GND 0.13fF
C265 a_18094_101.n1 GND 0.16fF
C266 a_18094_101.n2 GND 0.15fF
C267 a_18760_101.n0 GND 0.06fF
C268 a_18760_101.n1 GND 0.13fF
C269 a_18760_101.n2 GND 0.04fF
C270 a_18760_101.n3 GND 0.19fF
C271 a_4447_989.n0 GND 0.88fF
C272 a_4447_989.n1 GND 0.88fF
C273 a_4447_989.n2 GND 0.81fF
C274 a_4447_989.n3 GND 0.99fF
C275 a_4447_989.n4 GND 1.37fF
C276 a_4447_989.t11 GND 0.97fF
C277 a_4447_989.n5 GND 0.82fF
C278 a_4447_989.n6 GND 11.47fF
C279 a_4447_989.n7 GND 0.80fF
C280 a_4447_989.t12 GND 1.15fF
C281 a_4447_989.n8 GND 1.40fF
C282 a_4447_989.n9 GND 14.41fF
C283 a_4447_989.n10 GND 0.10fF
C284 a_4447_989.n11 GND 0.12fF
C285 a_4447_989.n12 GND 0.49fF
C286 a_4447_989.n13 GND 1.20fF
C287 a_4447_989.n14 GND 1.08fF
C288 a_4447_989.n15 GND 1.06fF
C289 a_4447_989.n16 GND 1.12fF
C290 a_4125_1050.n0 GND 0.38fF
C291 a_4125_1050.n1 GND 0.38fF
C292 a_4125_1050.n2 GND 0.32fF
C293 a_4125_1050.n3 GND 0.64fF
C294 a_4125_1050.n4 GND 0.33fF
C295 a_4125_1050.n5 GND 0.70fF
C296 a_4125_1050.n6 GND 0.44fF
C297 a_4125_1050.n7 GND 0.46fF
C298 a_4125_1050.n8 GND 0.49fF
C299 a_17533_1051.n0 GND 0.36fF
C300 a_17533_1051.n1 GND 0.32fF
C301 a_17533_1051.n2 GND 0.52fF
C302 a_17533_1051.n3 GND 0.30fF
C303 a_17533_1051.n4 GND 0.80fF
C304 a_17533_1051.n5 GND 0.43fF
C305 a_7973_1050.n0 GND 0.40fF
C306 a_7973_1050.n1 GND 0.40fF
C307 a_7973_1050.n2 GND 0.38fF
C308 a_7973_1050.n3 GND 0.65fF
C309 a_7973_1050.n4 GND 0.04fF
C310 a_7973_1050.n5 GND 0.05fF
C311 a_7973_1050.n6 GND 0.03fF
C312 a_7973_1050.n7 GND 0.17fF
C313 a_7973_1050.n8 GND 0.70fF
C314 a_7973_1050.n9 GND 0.52fF
C315 a_7973_1050.n10 GND 0.48fF
C316 a_7973_1050.n11 GND 0.50fF
C317 a_13840_210.n0 GND 0.02fF
C318 a_13840_210.n1 GND 0.09fF
C319 a_13840_210.n2 GND 0.12fF
C320 a_13840_210.n3 GND 0.08fF
C321 a_13840_210.n4 GND 0.08fF
C322 a_13840_210.n5 GND 0.02fF
C323 a_13840_210.t1 GND 0.29fF
C324 a_13840_210.n6 GND 0.09fF
C325 a_13840_210.n7 GND 0.02fF
C326 a_13840_210.n8 GND 0.13fF
C327 a_13840_210.n9 GND 0.02fF
C328 a_13840_210.n10 GND 0.03fF
C329 a_13840_210.n11 GND 0.03fF
C330 a_6049_1050.n0 GND 0.48fF
C331 a_6049_1050.n1 GND 0.83fF
C332 a_6049_1050.n2 GND 0.48fF
C333 a_6049_1050.n3 GND 0.60fF
C334 a_6049_1050.n4 GND 1.20fF
C335 a_6049_1050.n5 GND 0.05fF
C336 a_6049_1050.n6 GND 0.07fF
C337 a_6049_1050.n7 GND 0.04fF
C338 a_6049_1050.n8 GND 0.22fF
C339 a_6049_1050.n9 GND 0.72fF
C340 a_6049_1050.n10 GND 0.50fF
C341 a_6049_1050.n11 GND 0.64fF
C342 a_6049_1050.n12 GND 0.61fF
C343 a_6049_1050.n13 GND 0.66fF
C344 a_6049_1050.n14 GND 0.50fF
C345 a_3258_210.n0 GND 0.07fF
C346 a_3258_210.n1 GND 0.09fF
C347 a_3258_210.n2 GND 0.12fF
C348 a_3258_210.n3 GND 0.08fF
C349 a_3258_210.n4 GND 0.02fF
C350 a_3258_210.n5 GND 0.03fF
C351 a_3258_210.n6 GND 0.05fF
C352 a_3258_210.n7 GND 0.02fF
C353 a_3258_210.n8 GND 0.14fF
C354 a_3258_210.n9 GND 0.08fF
C355 a_3258_210.n10 GND 0.02fF
C356 a_3258_210.t0 GND 0.31fF
C357 a_2977_103.n0 GND 0.13fF
C358 a_2977_103.n1 GND 0.04fF
C359 a_2977_103.n2 GND 0.09fF
C360 a_2977_103.n3 GND 0.07fF
C361 a_2977_103.n4 GND 0.08fF
C362 a_2977_103.n5 GND 0.03fF
C363 a_15764_210.n0 GND 0.07fF
C364 a_15764_210.n1 GND 0.09fF
C365 a_15764_210.n2 GND 0.12fF
C366 a_15764_210.n3 GND 0.08fF
C367 a_15764_210.n4 GND 0.02fF
C368 a_15764_210.n5 GND 0.03fF
C369 a_15764_210.n6 GND 0.02fF
C370 a_15764_210.n7 GND 0.03fF
C371 a_15764_210.n8 GND 0.02fF
C372 a_15764_210.n9 GND 0.13fF
C373 a_15764_210.n10 GND 0.08fF
C374 a_15764_210.n11 GND 0.02fF
C375 a_15764_210.t0 GND 0.31fF
C376 a_15991_989.n0 GND 0.40fF
C377 a_15991_989.n1 GND 0.26fF
C378 a_15991_989.n2 GND 0.80fF
C379 a_15991_989.n3 GND 0.25fF
C380 a_15991_989.n4 GND 0.52fF
C381 a_15991_989.n5 GND 0.53fF
C382 a_15991_989.n6 GND 0.40fF
C383 a_15991_989.t7 GND 0.50fF
C384 a_15991_989.n7 GND 0.91fF
C385 a_15991_989.n8 GND 0.04fF
C386 a_15991_989.n9 GND 0.06fF
C387 a_15991_989.n10 GND 0.04fF
C388 a_15991_989.n11 GND 0.17fF
C389 a_15991_989.n12 GND 0.86fF
C390 a_15991_989.n13 GND 0.42fF
C391 a_15991_989.n14 GND 0.43fF
C392 a_15991_989.n15 GND 0.51fF
C393 a_15991_989.n16 GND 0.49fF
C394 a_15991_989.n17 GND 0.40fF
C395 a_1334_210.n0 GND 0.07fF
C396 a_1334_210.n1 GND 0.09fF
C397 a_1334_210.n2 GND 0.12fF
C398 a_1334_210.n3 GND 0.08fF
C399 a_1334_210.n4 GND 0.02fF
C400 a_1334_210.n5 GND 0.03fF
C401 a_1334_210.n6 GND 0.05fF
C402 a_1334_210.n7 GND 0.02fF
C403 a_1334_210.n8 GND 0.14fF
C404 a_1334_210.n9 GND 0.08fF
C405 a_1334_210.n10 GND 0.02fF
C406 a_1334_210.t0 GND 0.31fF
C407 a_1053_103.n0 GND 0.13fF
C408 a_1053_103.n1 GND 0.04fF
C409 a_1053_103.n2 GND 0.09fF
C410 a_1053_103.n3 GND 0.07fF
C411 a_1053_103.n4 GND 0.08fF
C412 a_1053_103.n5 GND 0.03fF
C413 a_7106_210.n0 GND 0.07fF
C414 a_7106_210.n1 GND 0.09fF
C415 a_7106_210.n2 GND 0.12fF
C416 a_7106_210.n3 GND 0.08fF
C417 a_7106_210.n4 GND 0.02fF
C418 a_7106_210.n5 GND 0.03fF
C419 a_7106_210.n6 GND 0.05fF
C420 a_7106_210.n7 GND 0.02fF
C421 a_7106_210.n8 GND 0.14fF
C422 a_7106_210.n9 GND 0.08fF
C423 a_7106_210.n10 GND 0.02fF
C424 a_7106_210.t0 GND 0.31fF
C425 a_6825_103.n0 GND 0.13fF
C426 a_6825_103.n1 GND 0.04fF
C427 a_6825_103.n2 GND 0.09fF
C428 a_6825_103.n3 GND 0.07fF
C429 a_6825_103.n4 GND 0.08fF
C430 a_6825_103.n5 GND 0.03fF
C431 a_5182_210.n0 GND 0.02fF
C432 a_5182_210.n1 GND 0.09fF
C433 a_5182_210.t1 GND 0.23fF
C434 a_5182_210.n2 GND 0.10fF
C435 a_5182_210.n3 GND 0.07fF
C436 a_5182_210.n4 GND 0.04fF
C437 a_5182_210.n5 GND 0.08fF
C438 a_5182_210.n6 GND 0.09fF
C439 a_5182_210.n7 GND 0.04fF
C440 a_5182_210.n8 GND 0.02fF
C441 a_5182_210.n9 GND 0.01fF
C442 a_5182_210.n10 GND 0.13fF
C443 a_5182_210.n11 GND 0.02fF
C444 a_5182_210.n12 GND 0.03fF
C445 a_5182_210.n13 GND 0.02fF
C446 a_4901_103.n0 GND 0.13fF
C447 a_4901_103.n1 GND 0.04fF
C448 a_4901_103.n2 GND 0.09fF
C449 a_4901_103.n3 GND 0.07fF
C450 a_4901_103.n4 GND 0.08fF
C451 a_4901_103.n5 GND 0.03fF
C452 a_6371_989.n0 GND 0.59fF
C453 a_6371_989.n1 GND 1.98fF
C454 a_6371_989.n2 GND 0.60fF
C455 a_6371_989.t11 GND 0.96fF
C456 a_6371_989.n3 GND 1.15fF
C457 a_6371_989.n4 GND 3.61fF
C458 a_6371_989.n5 GND 0.07fF
C459 a_6371_989.n6 GND 0.10fF
C460 a_6371_989.n7 GND 0.06fF
C461 a_6371_989.n8 GND 0.41fF
C462 a_6371_989.n9 GND 0.94fF
C463 a_6371_989.n10 GND 0.71fF
C464 a_6371_989.n11 GND 0.90fF
C465 a_6371_989.n12 GND 0.85fF
C466 a_6371_989.n13 GND 0.81fF
C467 a_6371_989.n14 GND 0.71fF
C468 a_10219_989.n0 GND 0.77fF
C469 a_10219_989.n1 GND 0.58fF
C470 a_10219_989.t8 GND 1.14fF
C471 a_10219_989.n2 GND 1.41fF
C472 a_10219_989.n3 GND 0.55fF
C473 a_10219_989.t12 GND 1.14fF
C474 a_10219_989.n4 GND 0.77fF
C475 a_10219_989.n5 GND 7.58fF
C476 a_10219_989.n6 GND 0.76fF
C477 a_10219_989.t13 GND 0.96fF
C478 a_10219_989.n7 GND 1.73fF
C479 a_10219_989.n8 GND 0.08fF
C480 a_10219_989.n9 GND 0.11fF
C481 a_10219_989.n10 GND 0.07fF
C482 a_10219_989.n11 GND 0.33fF
C483 a_10219_989.n12 GND 1.64fF
C484 a_10219_989.n13 GND 4.82fF
C485 a_10219_989.n14 GND 0.82fF
C486 a_10219_989.n15 GND 0.98fF
C487 a_10219_989.n16 GND 0.93fF
C488 a_10219_989.n17 GND 0.77fF
C489 SN.n0 GND 0.85fF
C490 SN.t10 GND 0.78fF
C491 SN.n1 GND 2.33fF
C492 SN.n2 GND 0.84fF
C493 SN.t12 GND 0.78fF
C494 SN.n3 GND 0.78fF
C495 SN.n4 GND 5.12fF
C496 SN.n5 GND 0.85fF
C497 SN.t9 GND 0.78fF
C498 SN.n6 GND 0.77fF
C499 SN.n7 GND 4.43fF
C500 SN.n8 GND 0.84fF
C501 SN.t3 GND 0.78fF
C502 SN.n9 GND 0.78fF
C503 SN.n10 GND 4.43fF
C504 SN.n11 GND 0.85fF
C505 SN.t1 GND 0.78fF
C506 SN.n12 GND 0.77fF
C507 SN.n13 GND 4.43fF
C508 SN.t17 GND 0.78fF
C509 SN.n14 GND 0.84fF
C510 SN.n15 GND 0.78fF
C511 SN.n16 GND 2.23fF
C512 a_2201_1050.n0 GND 0.36fF
C513 a_2201_1050.n1 GND 0.36fF
C514 a_2201_1050.n2 GND 0.35fF
C515 a_2201_1050.n3 GND 0.59fF
C516 a_2201_1050.n4 GND 0.04fF
C517 a_2201_1050.n5 GND 0.05fF
C518 a_2201_1050.n6 GND 0.03fF
C519 a_2201_1050.n7 GND 0.15fF
C520 a_2201_1050.n8 GND 0.64fF
C521 a_2201_1050.n9 GND 0.47fF
C522 a_2201_1050.n10 GND 0.43fF
C523 a_2201_1050.n11 GND 0.46fF
C524 a_277_1050.n0 GND 0.37fF
C525 a_277_1050.n1 GND 0.63fF
C526 a_277_1050.n2 GND 0.37fF
C527 a_277_1050.n3 GND 0.46fF
C528 a_277_1050.n4 GND 0.91fF
C529 a_277_1050.n5 GND 0.04fF
C530 a_277_1050.n6 GND 0.05fF
C531 a_277_1050.n7 GND 0.03fF
C532 a_277_1050.n8 GND 0.16fF
C533 a_277_1050.n9 GND 0.55fF
C534 a_277_1050.n10 GND 0.38fF
C535 a_277_1050.n11 GND 0.49fF
C536 a_277_1050.n12 GND 0.46fF
C537 a_277_1050.n13 GND 0.50fF
C538 a_277_1050.n14 GND 0.38fF
C539 a_13745_1050.n0 GND 0.40fF
C540 a_13745_1050.n1 GND 0.40fF
C541 a_13745_1050.n2 GND 0.38fF
C542 a_13745_1050.n3 GND 0.65fF
C543 a_13745_1050.n4 GND 0.04fF
C544 a_13745_1050.n5 GND 0.05fF
C545 a_13745_1050.n6 GND 0.03fF
C546 a_13745_1050.n7 GND 0.17fF
C547 a_13745_1050.n8 GND 0.70fF
C548 a_13745_1050.n9 GND 0.52fF
C549 a_13745_1050.n10 GND 0.48fF
C550 a_13745_1050.n11 GND 0.50fF
C551 a_7333_989.n0 GND 0.53fF
C552 a_7333_989.t15 GND 0.97fF
C553 a_7333_989.n1 GND 1.49fF
C554 a_7333_989.n2 GND 0.53fF
C555 a_7333_989.t13 GND 0.97fF
C556 a_7333_989.n3 GND 0.73fF
C557 a_7333_989.n4 GND 0.53fF
C558 a_7333_989.t12 GND 0.97fF
C559 a_7333_989.n5 GND 1.04fF
C560 a_7333_989.n6 GND 1.92fF
C561 a_7333_989.n7 GND 2.63fF
C562 a_7333_989.n8 GND 0.64fF
C563 a_7333_989.n9 GND 0.95fF
C564 a_7333_989.n10 GND 0.69fF
C565 a_7333_989.n11 GND 0.87fF
C566 a_7333_989.n12 GND 0.83fF
C567 a_7333_989.n13 GND 0.73fF
C568 a_7333_989.n14 GND 0.69fF
C569 a_9030_210.n0 GND 0.04fF
C570 a_9030_210.n1 GND 0.10fF
C571 a_9030_210.n2 GND 0.08fF
C572 a_9030_210.n3 GND 0.07fF
C573 a_9030_210.n4 GND 0.07fF
C574 a_9030_210.n5 GND 0.02fF
C575 a_9030_210.n6 GND 0.03fF
C576 a_9030_210.n7 GND 0.02fF
C577 a_9030_210.n8 GND 0.03fF
C578 a_9030_210.n9 GND 0.04fF
C579 a_9030_210.n10 GND 0.01fF
C580 a_9030_210.n11 GND 0.13fF
C581 a_9030_210.n12 GND 0.09fF
C582 a_9030_210.n13 GND 0.02fF
C583 a_9030_210.t0 GND 0.25fF
C584 a_11821_1050.n0 GND 0.48fF
C585 a_11821_1050.n1 GND 0.83fF
C586 a_11821_1050.n2 GND 0.48fF
C587 a_11821_1050.n3 GND 0.60fF
C588 a_11821_1050.n4 GND 1.20fF
C589 a_11821_1050.n5 GND 0.05fF
C590 a_11821_1050.n6 GND 0.07fF
C591 a_11821_1050.n7 GND 0.04fF
C592 a_11821_1050.n8 GND 0.22fF
C593 a_11821_1050.n9 GND 0.72fF
C594 a_11821_1050.n10 GND 0.50fF
C595 a_11821_1050.n11 GND 0.64fF
C596 a_11821_1050.n12 GND 0.61fF
C597 a_11821_1050.n13 GND 0.66fF
C598 a_11821_1050.n14 GND 0.50fF
C599 a_12143_989.n0 GND 0.70fF
C600 a_12143_989.n1 GND 0.58fF
C601 a_12143_989.n2 GND 1.96fF
C602 a_12143_989.n3 GND 0.59fF
C603 a_12143_989.t11 GND 0.95fF
C604 a_12143_989.n4 GND 1.13fF
C605 a_12143_989.n5 GND 3.56fF
C606 a_12143_989.n6 GND 0.07fF
C607 a_12143_989.n7 GND 0.10fF
C608 a_12143_989.n8 GND 0.06fF
C609 a_12143_989.n9 GND 0.40fF
C610 a_12143_989.n10 GND 0.93fF
C611 a_12143_989.n11 GND 0.80fF
C612 a_12143_989.n12 GND 0.89fF
C613 a_12143_989.n13 GND 0.84fF
C614 a_12143_989.n14 GND 0.70fF
C615 a_1561_989.n0 GND 0.49fF
C616 a_1561_989.t14 GND 0.89fF
C617 a_1561_989.n1 GND 1.37fF
C618 a_1561_989.n2 GND 0.49fF
C619 a_1561_989.t11 GND 0.89fF
C620 a_1561_989.n3 GND 0.67fF
C621 a_1561_989.n4 GND 0.49fF
C622 a_1561_989.t13 GND 0.89fF
C623 a_1561_989.n5 GND 0.96fF
C624 a_1561_989.n6 GND 1.76fF
C625 a_1561_989.n7 GND 2.42fF
C626 a_1561_989.n8 GND 0.06fF
C627 a_1561_989.n9 GND 0.09fF
C628 a_1561_989.n10 GND 0.05fF
C629 a_1561_989.n11 GND 0.41fF
C630 a_1561_989.n12 GND 0.84fF
C631 a_1561_989.n13 GND 0.63fF
C632 a_1561_989.n14 GND 0.80fF
C633 a_1561_989.n15 GND 0.76fF
C634 a_1561_989.n16 GND 0.67fF
C635 a_1561_989.n17 GND 0.63fF
C636 a_3939_103.n0 GND 0.13fF
C637 a_3939_103.n1 GND 0.04fF
C638 a_3939_103.n2 GND 0.09fF
C639 a_3939_103.n3 GND 0.07fF
C640 a_3939_103.n4 GND 0.08fF
C641 a_3939_103.n5 GND 0.03fF
C642 a_9897_1050.n0 GND 0.40fF
C643 a_9897_1050.n1 GND 0.33fF
C644 a_9897_1050.n2 GND 0.67fF
C645 a_9897_1050.n3 GND 0.35fF
C646 a_9897_1050.n4 GND 0.73fF
C647 a_9897_1050.n5 GND 0.46fF
C648 a_9897_1050.n6 GND 0.51fF
C649 a_9897_1050.n7 GND 0.48fF
C650 a_9897_1050.n8 GND 0.40fF
C651 a_599_989.n0 GND 0.53fF
C652 a_599_989.n1 GND 0.44fF
C653 a_599_989.n2 GND 1.48fF
C654 a_599_989.n3 GND 0.45fF
C655 a_599_989.t10 GND 0.72fF
C656 a_599_989.n4 GND 0.86fF
C657 a_599_989.n5 GND 2.70fF
C658 a_599_989.n6 GND 0.46fF
C659 a_599_989.n7 GND 0.73fF
C660 a_599_989.n8 GND 0.61fF
C661 a_599_989.n9 GND 0.68fF
C662 a_599_989.n10 GND 0.64fF
C663 a_599_989.n11 GND 0.53fF
C664 VDD.n1 GND 0.03fF
C665 VDD.n2 GND 0.11fF
C666 VDD.n3 GND 0.03fF
C667 VDD.n4 GND 0.02fF
C668 VDD.n5 GND 0.06fF
C669 VDD.n6 GND 0.02fF
C670 VDD.n7 GND 0.02fF
C671 VDD.n8 GND 0.02fF
C672 VDD.n9 GND 0.02fF
C673 VDD.n10 GND 0.02fF
C674 VDD.n11 GND 0.02fF
C675 VDD.n12 GND 0.02fF
C676 VDD.n13 GND 0.02fF
C677 VDD.n14 GND 0.04fF
C678 VDD.n15 GND 0.01fF
C679 VDD.n20 GND 0.48fF
C680 VDD.n21 GND 0.29fF
C681 VDD.n22 GND 0.02fF
C682 VDD.n23 GND 0.03fF
C683 VDD.n24 GND 0.07fF
C684 VDD.n25 GND 0.21fF
C685 VDD.n26 GND 0.01fF
C686 VDD.n27 GND 0.01fF
C687 VDD.n28 GND 0.07fF
C688 VDD.n29 GND 0.18fF
C689 VDD.n30 GND 0.01fF
C690 VDD.n31 GND 0.03fF
C691 VDD.n32 GND 0.03fF
C692 VDD.n33 GND 0.21fF
C693 VDD.n34 GND 0.01fF
C694 VDD.n35 GND 0.07fF
C695 VDD.n36 GND 0.01fF
C696 VDD.n37 GND 0.03fF
C697 VDD.n38 GND 0.29fF
C698 VDD.n39 GND 0.01fF
C699 VDD.n40 GND 0.02fF
C700 VDD.n41 GND 0.04fF
C701 VDD.n42 GND 0.06fF
C702 VDD.n43 GND 0.02fF
C703 VDD.n44 GND 0.02fF
C704 VDD.n45 GND 0.02fF
C705 VDD.n46 GND 0.02fF
C706 VDD.n47 GND 0.02fF
C707 VDD.n48 GND 0.02fF
C708 VDD.n49 GND 0.02fF
C709 VDD.n50 GND 0.02fF
C710 VDD.n51 GND 0.02fF
C711 VDD.n52 GND 0.02fF
C712 VDD.n53 GND 0.02fF
C713 VDD.n54 GND 0.03fF
C714 VDD.n55 GND 0.02fF
C715 VDD.n56 GND 0.19fF
C716 VDD.n57 GND 0.02fF
C717 VDD.n58 GND 0.02fF
C718 VDD.n60 GND 0.02fF
C719 VDD.n64 GND 0.29fF
C720 VDD.n65 GND 0.29fF
C721 VDD.n66 GND 0.01fF
C722 VDD.n67 GND 0.02fF
C723 VDD.n68 GND 0.04fF
C724 VDD.n69 GND 0.26fF
C725 VDD.n70 GND 0.01fF
C726 VDD.n71 GND 0.02fF
C727 VDD.n72 GND 0.02fF
C728 VDD.n73 GND 0.18fF
C729 VDD.n74 GND 0.01fF
C730 VDD.n75 GND 0.02fF
C731 VDD.n76 GND 0.02fF
C732 VDD.n77 GND 0.01fF
C733 VDD.n78 GND 0.03fF
C734 VDD.n79 GND 0.03fF
C735 VDD.n80 GND 0.15fF
C736 VDD.n81 GND 0.01fF
C737 VDD.n82 GND 0.03fF
C738 VDD.n83 GND 0.03fF
C739 VDD.n84 GND 0.17fF
C740 VDD.n85 GND 0.01fF
C741 VDD.n86 GND 0.02fF
C742 VDD.n87 GND 0.02fF
C743 VDD.n88 GND 0.26fF
C744 VDD.n89 GND 0.01fF
C745 VDD.n90 GND 0.02fF
C746 VDD.n91 GND 0.02fF
C747 VDD.n92 GND 0.29fF
C748 VDD.n93 GND 0.01fF
C749 VDD.n94 GND 0.02fF
C750 VDD.n95 GND 0.04fF
C751 VDD.n96 GND 0.23fF
C752 VDD.n97 GND 0.02fF
C753 VDD.n98 GND 0.02fF
C754 VDD.n99 GND 0.02fF
C755 VDD.n100 GND 0.06fF
C756 VDD.n101 GND 0.02fF
C757 VDD.n102 GND 0.02fF
C758 VDD.n103 GND 0.02fF
C759 VDD.n104 GND 0.02fF
C760 VDD.n105 GND 0.02fF
C761 VDD.n106 GND 0.02fF
C762 VDD.n107 GND 0.02fF
C763 VDD.n108 GND 0.02fF
C764 VDD.n109 GND 0.02fF
C765 VDD.n110 GND 0.02fF
C766 VDD.n111 GND 0.03fF
C767 VDD.n112 GND 0.02fF
C768 VDD.n113 GND 0.02fF
C769 VDD.n117 GND 0.29fF
C770 VDD.n118 GND 0.29fF
C771 VDD.n119 GND 0.01fF
C772 VDD.n120 GND 0.02fF
C773 VDD.n121 GND 0.04fF
C774 VDD.n122 GND 0.26fF
C775 VDD.n123 GND 0.01fF
C776 VDD.n124 GND 0.02fF
C777 VDD.n125 GND 0.02fF
C778 VDD.n126 GND 0.17fF
C779 VDD.n127 GND 0.01fF
C780 VDD.n128 GND 0.02fF
C781 VDD.n129 GND 0.02fF
C782 VDD.n130 GND 0.15fF
C783 VDD.n131 GND 0.01fF
C784 VDD.n132 GND 0.03fF
C785 VDD.n133 GND 0.03fF
C786 VDD.n134 GND 0.01fF
C787 VDD.n135 GND 0.03fF
C788 VDD.n136 GND 0.03fF
C789 VDD.n137 GND 0.18fF
C790 VDD.n138 GND 0.01fF
C791 VDD.n139 GND 0.02fF
C792 VDD.n140 GND 0.02fF
C793 VDD.n141 GND 0.26fF
C794 VDD.n142 GND 0.01fF
C795 VDD.n143 GND 0.02fF
C796 VDD.n144 GND 0.02fF
C797 VDD.n145 GND 0.29fF
C798 VDD.n146 GND 0.01fF
C799 VDD.n147 GND 0.02fF
C800 VDD.n148 GND 0.04fF
C801 VDD.n149 GND 0.23fF
C802 VDD.n150 GND 0.02fF
C803 VDD.n151 GND 0.02fF
C804 VDD.n152 GND 0.02fF
C805 VDD.n153 GND 0.06fF
C806 VDD.n154 GND 0.02fF
C807 VDD.n155 GND 0.02fF
C808 VDD.n156 GND 0.02fF
C809 VDD.n157 GND 0.02fF
C810 VDD.n158 GND 0.02fF
C811 VDD.n159 GND 0.02fF
C812 VDD.n160 GND 0.02fF
C813 VDD.n161 GND 0.02fF
C814 VDD.n162 GND 0.02fF
C815 VDD.n163 GND 0.02fF
C816 VDD.n164 GND 0.03fF
C817 VDD.n165 GND 0.02fF
C818 VDD.n166 GND 0.02fF
C819 VDD.n170 GND 0.29fF
C820 VDD.n171 GND 0.29fF
C821 VDD.n172 GND 0.01fF
C822 VDD.n173 GND 0.02fF
C823 VDD.n174 GND 0.04fF
C824 VDD.n175 GND 0.07fF
C825 VDD.n176 GND 0.26fF
C826 VDD.n177 GND 0.01fF
C827 VDD.n178 GND 0.01fF
C828 VDD.n179 GND 0.02fF
C829 VDD.n180 GND 0.18fF
C830 VDD.n181 GND 0.01fF
C831 VDD.n182 GND 0.02fF
C832 VDD.n183 GND 0.02fF
C833 VDD.n184 GND 0.09fF
C834 VDD.n185 GND 0.05fF
C835 VDD.n186 GND 0.01fF
C836 VDD.n187 GND 0.02fF
C837 VDD.n188 GND 0.03fF
C838 VDD.n189 GND 0.15fF
C839 VDD.n190 GND 0.01fF
C840 VDD.n191 GND 0.02fF
C841 VDD.n192 GND 0.03fF
C842 VDD.n193 GND 0.17fF
C843 VDD.n194 GND 0.01fF
C844 VDD.n195 GND 0.02fF
C845 VDD.n196 GND 0.02fF
C846 VDD.n197 GND 0.07fF
C847 VDD.n198 GND 0.26fF
C848 VDD.n199 GND 0.01fF
C849 VDD.n200 GND 0.01fF
C850 VDD.n201 GND 0.02fF
C851 VDD.n202 GND 0.29fF
C852 VDD.n203 GND 0.01fF
C853 VDD.n204 GND 0.02fF
C854 VDD.n205 GND 0.04fF
C855 VDD.n206 GND 0.28fF
C856 VDD.n207 GND 0.02fF
C857 VDD.n208 GND 0.02fF
C858 VDD.n209 GND 0.02fF
C859 VDD.n210 GND 0.06fF
C860 VDD.n211 GND 0.02fF
C861 VDD.n212 GND 0.02fF
C862 VDD.n213 GND 0.02fF
C863 VDD.n214 GND 0.02fF
C864 VDD.n215 GND 0.02fF
C865 VDD.n216 GND 0.02fF
C866 VDD.n217 GND 0.02fF
C867 VDD.n218 GND 0.02fF
C868 VDD.n219 GND 0.02fF
C869 VDD.n220 GND 0.02fF
C870 VDD.n221 GND 0.03fF
C871 VDD.n222 GND 0.02fF
C872 VDD.n223 GND 0.02fF
C873 VDD.n227 GND 0.29fF
C874 VDD.n228 GND 0.29fF
C875 VDD.n229 GND 0.01fF
C876 VDD.n230 GND 0.02fF
C877 VDD.n231 GND 0.04fF
C878 VDD.n232 GND 0.29fF
C879 VDD.n233 GND 0.01fF
C880 VDD.n234 GND 0.02fF
C881 VDD.n235 GND 0.02fF
C882 VDD.n236 GND 0.23fF
C883 VDD.n237 GND 0.01fF
C884 VDD.n238 GND 0.07fF
C885 VDD.n239 GND 0.02fF
C886 VDD.n240 GND 0.18fF
C887 VDD.n241 GND 0.01fF
C888 VDD.n242 GND 0.02fF
C889 VDD.n243 GND 0.02fF
C890 VDD.n244 GND 0.17fF
C891 VDD.n245 GND 0.01fF
C892 VDD.n246 GND 0.09fF
C893 VDD.n247 GND 0.05fF
C894 VDD.n248 GND 0.02fF
C895 VDD.n249 GND 0.02fF
C896 VDD.n250 GND 0.15fF
C897 VDD.n251 GND 0.02fF
C898 VDD.n252 GND 0.02fF
C899 VDD.n253 GND 0.03fF
C900 VDD.n254 GND 0.16fF
C901 VDD.n255 GND 0.02fF
C902 VDD.n256 GND 0.02fF
C903 VDD.n257 GND 0.03fF
C904 VDD.n258 GND 0.09fF
C905 VDD.n259 GND 0.05fF
C906 VDD.n260 GND 0.17fF
C907 VDD.n261 GND 0.01fF
C908 VDD.n262 GND 0.02fF
C909 VDD.n263 GND 0.02fF
C910 VDD.n264 GND 0.18fF
C911 VDD.n265 GND 0.01fF
C912 VDD.n266 GND 0.02fF
C913 VDD.n267 GND 0.02fF
C914 VDD.n268 GND 0.07fF
C915 VDD.n269 GND 0.24fF
C916 VDD.n270 GND 0.01fF
C917 VDD.n271 GND 0.01fF
C918 VDD.n272 GND 0.02fF
C919 VDD.n273 GND 0.29fF
C920 VDD.n274 GND 0.01fF
C921 VDD.n275 GND 0.02fF
C922 VDD.n276 GND 0.02fF
C923 VDD.n277 GND 0.29fF
C924 VDD.n278 GND 0.01fF
C925 VDD.n279 GND 0.02fF
C926 VDD.n280 GND 0.04fF
C927 VDD.n281 GND 0.33fF
C928 VDD.n282 GND 0.02fF
C929 VDD.n283 GND 0.02fF
C930 VDD.n284 GND 0.02fF
C931 VDD.n285 GND 0.06fF
C932 VDD.n286 GND 0.02fF
C933 VDD.n287 GND 0.02fF
C934 VDD.n288 GND 0.02fF
C935 VDD.n289 GND 0.02fF
C936 VDD.n290 GND 0.02fF
C937 VDD.n291 GND 0.02fF
C938 VDD.n292 GND 0.02fF
C939 VDD.n293 GND 0.02fF
C940 VDD.n294 GND 0.02fF
C941 VDD.n295 GND 0.02fF
C942 VDD.n296 GND 0.03fF
C943 VDD.n297 GND 0.02fF
C944 VDD.n298 GND 0.02fF
C945 VDD.n302 GND 0.29fF
C946 VDD.n303 GND 0.29fF
C947 VDD.n304 GND 0.01fF
C948 VDD.n305 GND 0.02fF
C949 VDD.n306 GND 0.04fF
C950 VDD.n307 GND 0.29fF
C951 VDD.n308 GND 0.01fF
C952 VDD.n309 GND 0.02fF
C953 VDD.n310 GND 0.02fF
C954 VDD.n311 GND 0.23fF
C955 VDD.n312 GND 0.01fF
C956 VDD.n313 GND 0.07fF
C957 VDD.n314 GND 0.02fF
C958 VDD.n315 GND 0.18fF
C959 VDD.n316 GND 0.01fF
C960 VDD.n317 GND 0.02fF
C961 VDD.n318 GND 0.02fF
C962 VDD.n319 GND 0.17fF
C963 VDD.n320 GND 0.01fF
C964 VDD.n321 GND 0.09fF
C965 VDD.n322 GND 0.05fF
C966 VDD.n323 GND 0.02fF
C967 VDD.n324 GND 0.02fF
C968 VDD.n325 GND 0.15fF
C969 VDD.n326 GND 0.02fF
C970 VDD.n327 GND 0.02fF
C971 VDD.n328 GND 0.03fF
C972 VDD.n329 GND 0.16fF
C973 VDD.n330 GND 0.02fF
C974 VDD.n331 GND 0.02fF
C975 VDD.n332 GND 0.03fF
C976 VDD.n333 GND 0.09fF
C977 VDD.n334 GND 0.05fF
C978 VDD.n335 GND 0.17fF
C979 VDD.n336 GND 0.01fF
C980 VDD.n337 GND 0.02fF
C981 VDD.n338 GND 0.02fF
C982 VDD.n339 GND 0.18fF
C983 VDD.n340 GND 0.01fF
C984 VDD.n341 GND 0.02fF
C985 VDD.n342 GND 0.02fF
C986 VDD.n343 GND 0.07fF
C987 VDD.n344 GND 0.24fF
C988 VDD.n345 GND 0.01fF
C989 VDD.n346 GND 0.01fF
C990 VDD.n347 GND 0.02fF
C991 VDD.n348 GND 0.29fF
C992 VDD.n349 GND 0.01fF
C993 VDD.n350 GND 0.02fF
C994 VDD.n351 GND 0.02fF
C995 VDD.n352 GND 0.29fF
C996 VDD.n353 GND 0.01fF
C997 VDD.n354 GND 0.02fF
C998 VDD.n355 GND 0.04fF
C999 VDD.n356 GND 0.33fF
C1000 VDD.n357 GND 0.02fF
C1001 VDD.n358 GND 0.02fF
C1002 VDD.n359 GND 0.02fF
C1003 VDD.n360 GND 0.06fF
C1004 VDD.n361 GND 0.02fF
C1005 VDD.n362 GND 0.02fF
C1006 VDD.n363 GND 0.02fF
C1007 VDD.n364 GND 0.02fF
C1008 VDD.n365 GND 0.02fF
C1009 VDD.n366 GND 0.02fF
C1010 VDD.n367 GND 0.02fF
C1011 VDD.n368 GND 0.02fF
C1012 VDD.n369 GND 0.02fF
C1013 VDD.n370 GND 0.02fF
C1014 VDD.n371 GND 0.03fF
C1015 VDD.n372 GND 0.02fF
C1016 VDD.n373 GND 0.02fF
C1017 VDD.n377 GND 0.29fF
C1018 VDD.n378 GND 0.29fF
C1019 VDD.n379 GND 0.01fF
C1020 VDD.n380 GND 0.02fF
C1021 VDD.n381 GND 0.04fF
C1022 VDD.n382 GND 0.29fF
C1023 VDD.n383 GND 0.01fF
C1024 VDD.n384 GND 0.02fF
C1025 VDD.n385 GND 0.02fF
C1026 VDD.n386 GND 0.23fF
C1027 VDD.n387 GND 0.01fF
C1028 VDD.n388 GND 0.07fF
C1029 VDD.n389 GND 0.02fF
C1030 VDD.n390 GND 0.18fF
C1031 VDD.n391 GND 0.01fF
C1032 VDD.n392 GND 0.02fF
C1033 VDD.n393 GND 0.02fF
C1034 VDD.n394 GND 0.17fF
C1035 VDD.n395 GND 0.01fF
C1036 VDD.n396 GND 0.09fF
C1037 VDD.n397 GND 0.05fF
C1038 VDD.n398 GND 0.02fF
C1039 VDD.n399 GND 0.02fF
C1040 VDD.n400 GND 0.15fF
C1041 VDD.n401 GND 0.02fF
C1042 VDD.n402 GND 0.02fF
C1043 VDD.n403 GND 0.03fF
C1044 VDD.n404 GND 0.16fF
C1045 VDD.n405 GND 0.02fF
C1046 VDD.n406 GND 0.02fF
C1047 VDD.n407 GND 0.03fF
C1048 VDD.n408 GND 0.09fF
C1049 VDD.n409 GND 0.05fF
C1050 VDD.n410 GND 0.17fF
C1051 VDD.n411 GND 0.01fF
C1052 VDD.n412 GND 0.02fF
C1053 VDD.n413 GND 0.02fF
C1054 VDD.n414 GND 0.18fF
C1055 VDD.n415 GND 0.01fF
C1056 VDD.n416 GND 0.02fF
C1057 VDD.n417 GND 0.02fF
C1058 VDD.n418 GND 0.07fF
C1059 VDD.n419 GND 0.24fF
C1060 VDD.n420 GND 0.01fF
C1061 VDD.n421 GND 0.01fF
C1062 VDD.n422 GND 0.02fF
C1063 VDD.n423 GND 0.29fF
C1064 VDD.n424 GND 0.01fF
C1065 VDD.n425 GND 0.02fF
C1066 VDD.n426 GND 0.02fF
C1067 VDD.n427 GND 0.29fF
C1068 VDD.n428 GND 0.01fF
C1069 VDD.n429 GND 0.02fF
C1070 VDD.n430 GND 0.04fF
C1071 VDD.n431 GND 0.33fF
C1072 VDD.n432 GND 0.02fF
C1073 VDD.n433 GND 0.02fF
C1074 VDD.n434 GND 0.02fF
C1075 VDD.n435 GND 0.06fF
C1076 VDD.n436 GND 0.02fF
C1077 VDD.n437 GND 0.02fF
C1078 VDD.n438 GND 0.02fF
C1079 VDD.n439 GND 0.02fF
C1080 VDD.n440 GND 0.02fF
C1081 VDD.n441 GND 0.02fF
C1082 VDD.n442 GND 0.02fF
C1083 VDD.n443 GND 0.02fF
C1084 VDD.n444 GND 0.02fF
C1085 VDD.n445 GND 0.02fF
C1086 VDD.n446 GND 0.03fF
C1087 VDD.n447 GND 0.02fF
C1088 VDD.n448 GND 0.02fF
C1089 VDD.n452 GND 0.29fF
C1090 VDD.n453 GND 0.29fF
C1091 VDD.n454 GND 0.01fF
C1092 VDD.n455 GND 0.02fF
C1093 VDD.n456 GND 0.04fF
C1094 VDD.n457 GND 0.29fF
C1095 VDD.n458 GND 0.01fF
C1096 VDD.n459 GND 0.02fF
C1097 VDD.n460 GND 0.02fF
C1098 VDD.n461 GND 0.23fF
C1099 VDD.n462 GND 0.01fF
C1100 VDD.n463 GND 0.07fF
C1101 VDD.n464 GND 0.02fF
C1102 VDD.n465 GND 0.18fF
C1103 VDD.n466 GND 0.01fF
C1104 VDD.n467 GND 0.02fF
C1105 VDD.n468 GND 0.02fF
C1106 VDD.n469 GND 0.17fF
C1107 VDD.n470 GND 0.01fF
C1108 VDD.n471 GND 0.09fF
C1109 VDD.n472 GND 0.05fF
C1110 VDD.n473 GND 0.02fF
C1111 VDD.n474 GND 0.02fF
C1112 VDD.n475 GND 0.15fF
C1113 VDD.n476 GND 0.02fF
C1114 VDD.n477 GND 0.02fF
C1115 VDD.n478 GND 0.03fF
C1116 VDD.n479 GND 0.16fF
C1117 VDD.n480 GND 0.02fF
C1118 VDD.n481 GND 0.02fF
C1119 VDD.n482 GND 0.03fF
C1120 VDD.n483 GND 0.09fF
C1121 VDD.n484 GND 0.05fF
C1122 VDD.n485 GND 0.17fF
C1123 VDD.n486 GND 0.01fF
C1124 VDD.n487 GND 0.02fF
C1125 VDD.n488 GND 0.02fF
C1126 VDD.n489 GND 0.18fF
C1127 VDD.n490 GND 0.01fF
C1128 VDD.n491 GND 0.02fF
C1129 VDD.n492 GND 0.02fF
C1130 VDD.n493 GND 0.07fF
C1131 VDD.n494 GND 0.24fF
C1132 VDD.n495 GND 0.01fF
C1133 VDD.n496 GND 0.01fF
C1134 VDD.n497 GND 0.02fF
C1135 VDD.n498 GND 0.29fF
C1136 VDD.n499 GND 0.01fF
C1137 VDD.n500 GND 0.02fF
C1138 VDD.n501 GND 0.02fF
C1139 VDD.n502 GND 0.29fF
C1140 VDD.n503 GND 0.01fF
C1141 VDD.n504 GND 0.02fF
C1142 VDD.n505 GND 0.04fF
C1143 VDD.n506 GND 0.33fF
C1144 VDD.n507 GND 0.02fF
C1145 VDD.n508 GND 0.02fF
C1146 VDD.n509 GND 0.02fF
C1147 VDD.n510 GND 0.06fF
C1148 VDD.n511 GND 0.02fF
C1149 VDD.n512 GND 0.02fF
C1150 VDD.n513 GND 0.02fF
C1151 VDD.n514 GND 0.02fF
C1152 VDD.n515 GND 0.02fF
C1153 VDD.n516 GND 0.02fF
C1154 VDD.n517 GND 0.02fF
C1155 VDD.n518 GND 0.02fF
C1156 VDD.n519 GND 0.02fF
C1157 VDD.n520 GND 0.02fF
C1158 VDD.n521 GND 0.03fF
C1159 VDD.n522 GND 0.02fF
C1160 VDD.n523 GND 0.02fF
C1161 VDD.n527 GND 0.29fF
C1162 VDD.n528 GND 0.29fF
C1163 VDD.n529 GND 0.01fF
C1164 VDD.n530 GND 0.02fF
C1165 VDD.n531 GND 0.04fF
C1166 VDD.n532 GND 0.29fF
C1167 VDD.n533 GND 0.01fF
C1168 VDD.n534 GND 0.02fF
C1169 VDD.n535 GND 0.02fF
C1170 VDD.n536 GND 0.23fF
C1171 VDD.n537 GND 0.01fF
C1172 VDD.n538 GND 0.07fF
C1173 VDD.n539 GND 0.02fF
C1174 VDD.n540 GND 0.18fF
C1175 VDD.n541 GND 0.01fF
C1176 VDD.n542 GND 0.02fF
C1177 VDD.n543 GND 0.02fF
C1178 VDD.n544 GND 0.17fF
C1179 VDD.n545 GND 0.01fF
C1180 VDD.n546 GND 0.09fF
C1181 VDD.n547 GND 0.05fF
C1182 VDD.n548 GND 0.02fF
C1183 VDD.n549 GND 0.02fF
C1184 VDD.n550 GND 0.15fF
C1185 VDD.n551 GND 0.02fF
C1186 VDD.n552 GND 0.02fF
C1187 VDD.n553 GND 0.03fF
C1188 VDD.n554 GND 0.16fF
C1189 VDD.n555 GND 0.02fF
C1190 VDD.n556 GND 0.02fF
C1191 VDD.n557 GND 0.03fF
C1192 VDD.n558 GND 0.09fF
C1193 VDD.n559 GND 0.05fF
C1194 VDD.n560 GND 0.17fF
C1195 VDD.n561 GND 0.01fF
C1196 VDD.n562 GND 0.02fF
C1197 VDD.n563 GND 0.02fF
C1198 VDD.n564 GND 0.18fF
C1199 VDD.n565 GND 0.01fF
C1200 VDD.n566 GND 0.02fF
C1201 VDD.n567 GND 0.02fF
C1202 VDD.n568 GND 0.07fF
C1203 VDD.n569 GND 0.24fF
C1204 VDD.n570 GND 0.01fF
C1205 VDD.n571 GND 0.01fF
C1206 VDD.n572 GND 0.02fF
C1207 VDD.n573 GND 0.29fF
C1208 VDD.n574 GND 0.01fF
C1209 VDD.n575 GND 0.02fF
C1210 VDD.n576 GND 0.02fF
C1211 VDD.n577 GND 0.29fF
C1212 VDD.n578 GND 0.01fF
C1213 VDD.n579 GND 0.02fF
C1214 VDD.n580 GND 0.04fF
C1215 VDD.n581 GND 0.33fF
C1216 VDD.n582 GND 0.02fF
C1217 VDD.n583 GND 0.02fF
C1218 VDD.n584 GND 0.02fF
C1219 VDD.n585 GND 0.06fF
C1220 VDD.n586 GND 0.02fF
C1221 VDD.n587 GND 0.02fF
C1222 VDD.n588 GND 0.02fF
C1223 VDD.n589 GND 0.02fF
C1224 VDD.n590 GND 0.02fF
C1225 VDD.n591 GND 0.02fF
C1226 VDD.n592 GND 0.02fF
C1227 VDD.n593 GND 0.02fF
C1228 VDD.n594 GND 0.02fF
C1229 VDD.n595 GND 0.02fF
C1230 VDD.n596 GND 0.03fF
C1231 VDD.n597 GND 0.02fF
C1232 VDD.n598 GND 0.02fF
C1233 VDD.n602 GND 0.29fF
C1234 VDD.n603 GND 0.29fF
C1235 VDD.n604 GND 0.01fF
C1236 VDD.n605 GND 0.02fF
C1237 VDD.n606 GND 0.04fF
C1238 VDD.n607 GND 0.29fF
C1239 VDD.n608 GND 0.01fF
C1240 VDD.n609 GND 0.02fF
C1241 VDD.n610 GND 0.02fF
C1242 VDD.n611 GND 0.23fF
C1243 VDD.n612 GND 0.01fF
C1244 VDD.n613 GND 0.07fF
C1245 VDD.n614 GND 0.02fF
C1246 VDD.n615 GND 0.18fF
C1247 VDD.n616 GND 0.01fF
C1248 VDD.n617 GND 0.02fF
C1249 VDD.n618 GND 0.02fF
C1250 VDD.n619 GND 0.17fF
C1251 VDD.n620 GND 0.01fF
C1252 VDD.n621 GND 0.09fF
C1253 VDD.n622 GND 0.05fF
C1254 VDD.n623 GND 0.02fF
C1255 VDD.n624 GND 0.02fF
C1256 VDD.n625 GND 0.15fF
C1257 VDD.n626 GND 0.02fF
C1258 VDD.n627 GND 0.02fF
C1259 VDD.n628 GND 0.03fF
C1260 VDD.n629 GND 0.16fF
C1261 VDD.n630 GND 0.02fF
C1262 VDD.n631 GND 0.02fF
C1263 VDD.n632 GND 0.03fF
C1264 VDD.n633 GND 0.09fF
C1265 VDD.n634 GND 0.05fF
C1266 VDD.n635 GND 0.17fF
C1267 VDD.n636 GND 0.01fF
C1268 VDD.n637 GND 0.02fF
C1269 VDD.n638 GND 0.02fF
C1270 VDD.n639 GND 0.18fF
C1271 VDD.n640 GND 0.01fF
C1272 VDD.n641 GND 0.02fF
C1273 VDD.n642 GND 0.02fF
C1274 VDD.n643 GND 0.07fF
C1275 VDD.n644 GND 0.24fF
C1276 VDD.n645 GND 0.01fF
C1277 VDD.n646 GND 0.01fF
C1278 VDD.n647 GND 0.02fF
C1279 VDD.n648 GND 0.29fF
C1280 VDD.n649 GND 0.01fF
C1281 VDD.n650 GND 0.02fF
C1282 VDD.n651 GND 0.02fF
C1283 VDD.n652 GND 0.29fF
C1284 VDD.n653 GND 0.01fF
C1285 VDD.n654 GND 0.02fF
C1286 VDD.n655 GND 0.04fF
C1287 VDD.n656 GND 0.33fF
C1288 VDD.n657 GND 0.02fF
C1289 VDD.n658 GND 0.02fF
C1290 VDD.n659 GND 0.02fF
C1291 VDD.n660 GND 0.06fF
C1292 VDD.n661 GND 0.02fF
C1293 VDD.n662 GND 0.02fF
C1294 VDD.n663 GND 0.02fF
C1295 VDD.n664 GND 0.02fF
C1296 VDD.n665 GND 0.02fF
C1297 VDD.n666 GND 0.02fF
C1298 VDD.n667 GND 0.02fF
C1299 VDD.n668 GND 0.02fF
C1300 VDD.n669 GND 0.02fF
C1301 VDD.n670 GND 0.02fF
C1302 VDD.n671 GND 0.03fF
C1303 VDD.n672 GND 0.02fF
C1304 VDD.n673 GND 0.02fF
C1305 VDD.n677 GND 0.29fF
C1306 VDD.n678 GND 0.29fF
C1307 VDD.n679 GND 0.01fF
C1308 VDD.n680 GND 0.02fF
C1309 VDD.n681 GND 0.04fF
C1310 VDD.n682 GND 0.29fF
C1311 VDD.n683 GND 0.01fF
C1312 VDD.n684 GND 0.02fF
C1313 VDD.n685 GND 0.02fF
C1314 VDD.n686 GND 0.23fF
C1315 VDD.n687 GND 0.01fF
C1316 VDD.n688 GND 0.07fF
C1317 VDD.n689 GND 0.02fF
C1318 VDD.n690 GND 0.18fF
C1319 VDD.n691 GND 0.01fF
C1320 VDD.n692 GND 0.02fF
C1321 VDD.n693 GND 0.02fF
C1322 VDD.n694 GND 0.17fF
C1323 VDD.n695 GND 0.01fF
C1324 VDD.n696 GND 0.09fF
C1325 VDD.n697 GND 0.05fF
C1326 VDD.n698 GND 0.02fF
C1327 VDD.n699 GND 0.02fF
C1328 VDD.n700 GND 0.15fF
C1329 VDD.n701 GND 0.02fF
C1330 VDD.n702 GND 0.02fF
C1331 VDD.n703 GND 0.03fF
C1332 VDD.n704 GND 0.16fF
C1333 VDD.n705 GND 0.02fF
C1334 VDD.n706 GND 0.02fF
C1335 VDD.n707 GND 0.03fF
C1336 VDD.n708 GND 0.09fF
C1337 VDD.n709 GND 0.05fF
C1338 VDD.n710 GND 0.17fF
C1339 VDD.n711 GND 0.01fF
C1340 VDD.n712 GND 0.02fF
C1341 VDD.n713 GND 0.02fF
C1342 VDD.n714 GND 0.18fF
C1343 VDD.n715 GND 0.01fF
C1344 VDD.n716 GND 0.02fF
C1345 VDD.n717 GND 0.02fF
C1346 VDD.n718 GND 0.07fF
C1347 VDD.n719 GND 0.24fF
C1348 VDD.n720 GND 0.01fF
C1349 VDD.n721 GND 0.01fF
C1350 VDD.n722 GND 0.02fF
C1351 VDD.n723 GND 0.29fF
C1352 VDD.n724 GND 0.01fF
C1353 VDD.n725 GND 0.02fF
C1354 VDD.n726 GND 0.02fF
C1355 VDD.n727 GND 0.29fF
C1356 VDD.n728 GND 0.01fF
C1357 VDD.n729 GND 0.02fF
C1358 VDD.n730 GND 0.04fF
C1359 VDD.n731 GND 0.33fF
C1360 VDD.n732 GND 0.02fF
C1361 VDD.n733 GND 0.02fF
C1362 VDD.n734 GND 0.02fF
C1363 VDD.n735 GND 0.06fF
C1364 VDD.n736 GND 0.02fF
C1365 VDD.n737 GND 0.02fF
C1366 VDD.n738 GND 0.02fF
C1367 VDD.n739 GND 0.02fF
C1368 VDD.n740 GND 0.02fF
C1369 VDD.n741 GND 0.02fF
C1370 VDD.n742 GND 0.02fF
C1371 VDD.n743 GND 0.02fF
C1372 VDD.n744 GND 0.02fF
C1373 VDD.n745 GND 0.02fF
C1374 VDD.n746 GND 0.03fF
C1375 VDD.n747 GND 0.02fF
C1376 VDD.n748 GND 0.02fF
C1377 VDD.n752 GND 0.29fF
C1378 VDD.n753 GND 0.29fF
C1379 VDD.n754 GND 0.01fF
C1380 VDD.n755 GND 0.02fF
C1381 VDD.n756 GND 0.04fF
C1382 VDD.n757 GND 0.29fF
C1383 VDD.n758 GND 0.01fF
C1384 VDD.n759 GND 0.02fF
C1385 VDD.n760 GND 0.02fF
C1386 VDD.n761 GND 0.23fF
C1387 VDD.n762 GND 0.01fF
C1388 VDD.n763 GND 0.07fF
C1389 VDD.n764 GND 0.02fF
C1390 VDD.n765 GND 0.18fF
C1391 VDD.n766 GND 0.01fF
C1392 VDD.n767 GND 0.02fF
C1393 VDD.n768 GND 0.02fF
C1394 VDD.n769 GND 0.17fF
C1395 VDD.n770 GND 0.01fF
C1396 VDD.n771 GND 0.09fF
C1397 VDD.n772 GND 0.05fF
C1398 VDD.n773 GND 0.02fF
C1399 VDD.n774 GND 0.02fF
C1400 VDD.n775 GND 0.15fF
C1401 VDD.n776 GND 0.02fF
C1402 VDD.n777 GND 0.02fF
C1403 VDD.n778 GND 0.03fF
C1404 VDD.n779 GND 0.16fF
C1405 VDD.n780 GND 0.02fF
C1406 VDD.n781 GND 0.02fF
C1407 VDD.n782 GND 0.03fF
C1408 VDD.n783 GND 0.09fF
C1409 VDD.n784 GND 0.05fF
C1410 VDD.n785 GND 0.17fF
C1411 VDD.n786 GND 0.01fF
C1412 VDD.n787 GND 0.02fF
C1413 VDD.n788 GND 0.02fF
C1414 VDD.n789 GND 0.18fF
C1415 VDD.n790 GND 0.01fF
C1416 VDD.n791 GND 0.02fF
C1417 VDD.n792 GND 0.02fF
C1418 VDD.n793 GND 0.19fF
C1419 VDD.n794 GND 0.02fF
C1420 VDD.n795 GND 0.02fF
C1421 VDD.n796 GND 0.06fF
C1422 VDD.n797 GND 0.02fF
C1423 VDD.n798 GND 0.02fF
C1424 VDD.n799 GND 0.02fF
C1425 VDD.n800 GND 0.02fF
C1426 VDD.n801 GND 0.02fF
C1427 VDD.n802 GND 0.02fF
C1428 VDD.n803 GND 0.02fF
C1429 VDD.n804 GND 0.02fF
C1430 VDD.n805 GND 0.03fF
C1431 VDD.n806 GND 0.04fF
C1432 VDD.n807 GND 0.02fF
C1433 VDD.n811 GND 0.48fF
C1434 VDD.n812 GND 0.29fF
C1435 VDD.n813 GND 0.02fF
C1436 VDD.n814 GND 0.03fF
C1437 VDD.n815 GND 0.03fF
C1438 VDD.n816 GND 0.29fF
C1439 VDD.n817 GND 0.01fF
C1440 VDD.n818 GND 0.02fF
C1441 VDD.n819 GND 0.02fF
C1442 VDD.n820 GND 0.07fF
C1443 VDD.n821 GND 0.24fF
C1444 VDD.n822 GND 0.01fF
C1445 VDD.n823 GND 0.01fF
C1446 VDD.n824 GND 0.02fF
C1447 VDD.n825 GND 0.18fF
C1448 VDD.n826 GND 0.01fF
C1449 VDD.n827 GND 0.02fF
C1450 VDD.n828 GND 0.02fF
C1451 VDD.n829 GND 0.09fF
C1452 VDD.n830 GND 0.05fF
C1453 VDD.n831 GND 0.17fF
C1454 VDD.n832 GND 0.01fF
C1455 VDD.n833 GND 0.02fF
C1456 VDD.n834 GND 0.02fF
C1457 VDD.n835 GND 0.16fF
C1458 VDD.n836 GND 0.02fF
C1459 VDD.n837 GND 0.02fF
C1460 VDD.n838 GND 0.03fF
C1461 VDD.n839 GND 0.15fF
C1462 VDD.n840 GND 0.02fF
C1463 VDD.n841 GND 0.02fF
C1464 VDD.n842 GND 0.03fF
C1465 VDD.n843 GND 0.17fF
C1466 VDD.n844 GND 0.01fF
C1467 VDD.n845 GND 0.09fF
C1468 VDD.n846 GND 0.05fF
C1469 VDD.n847 GND 0.02fF
C1470 VDD.n848 GND 0.02fF
C1471 VDD.n849 GND 0.18fF
C1472 VDD.n850 GND 0.01fF
C1473 VDD.n851 GND 0.02fF
C1474 VDD.n852 GND 0.02fF
C1475 VDD.n853 GND 0.23fF
C1476 VDD.n854 GND 0.01fF
C1477 VDD.n855 GND 0.07fF
C1478 VDD.n856 GND 0.02fF
C1479 VDD.n857 GND 0.29fF
C1480 VDD.n858 GND 0.01fF
C1481 VDD.n859 GND 0.02fF
C1482 VDD.n860 GND 0.02fF
C1483 VDD.n861 GND 0.29fF
C1484 VDD.n862 GND 0.01fF
C1485 VDD.n863 GND 0.02fF
C1486 VDD.n864 GND 0.04fF
C1487 VDD.n865 GND 0.06fF
C1488 VDD.n866 GND 0.02fF
C1489 VDD.n867 GND 0.02fF
C1490 VDD.n868 GND 0.02fF
C1491 VDD.n869 GND 0.02fF
C1492 VDD.n870 GND 0.02fF
C1493 VDD.n871 GND 0.02fF
C1494 VDD.n872 GND 0.02fF
C1495 VDD.n873 GND 0.02fF
C1496 VDD.n874 GND 0.02fF
C1497 VDD.n875 GND 0.02fF
C1498 VDD.n876 GND 0.02fF
C1499 VDD.n877 GND 0.03fF
C1500 VDD.n878 GND 0.02fF
C1501 VDD.n881 GND 0.02fF
C1502 VDD.n883 GND 0.02fF
C1503 VDD.n884 GND 0.33fF
C1504 VDD.n885 GND 0.02fF
C1505 VDD.n887 GND 0.29fF
C1506 VDD.n888 GND 0.29fF
C1507 VDD.n889 GND 0.01fF
C1508 VDD.n890 GND 0.02fF
C1509 VDD.n891 GND 0.04fF
C1510 VDD.n892 GND 0.29fF
C1511 VDD.n893 GND 0.01fF
C1512 VDD.n894 GND 0.02fF
C1513 VDD.n895 GND 0.02fF
C1514 VDD.n896 GND 0.07fF
C1515 VDD.n897 GND 0.24fF
C1516 VDD.n898 GND 0.01fF
C1517 VDD.n899 GND 0.01fF
C1518 VDD.n900 GND 0.02fF
C1519 VDD.n901 GND 0.18fF
C1520 VDD.n902 GND 0.01fF
C1521 VDD.n903 GND 0.02fF
C1522 VDD.n904 GND 0.02fF
C1523 VDD.n905 GND 0.09fF
C1524 VDD.n906 GND 0.05fF
C1525 VDD.n907 GND 0.17fF
C1526 VDD.n908 GND 0.01fF
C1527 VDD.n909 GND 0.02fF
C1528 VDD.n910 GND 0.02fF
C1529 VDD.n911 GND 0.16fF
C1530 VDD.n912 GND 0.02fF
C1531 VDD.n913 GND 0.02fF
C1532 VDD.n914 GND 0.03fF
C1533 VDD.n915 GND 0.15fF
C1534 VDD.n916 GND 0.02fF
C1535 VDD.n917 GND 0.02fF
C1536 VDD.n918 GND 0.03fF
C1537 VDD.n919 GND 0.17fF
C1538 VDD.n920 GND 0.01fF
C1539 VDD.n921 GND 0.09fF
C1540 VDD.n922 GND 0.05fF
C1541 VDD.n923 GND 0.02fF
C1542 VDD.n924 GND 0.02fF
C1543 VDD.n925 GND 0.18fF
C1544 VDD.n926 GND 0.01fF
C1545 VDD.n927 GND 0.02fF
C1546 VDD.n928 GND 0.02fF
C1547 VDD.n929 GND 0.23fF
C1548 VDD.n930 GND 0.01fF
C1549 VDD.n931 GND 0.07fF
C1550 VDD.n932 GND 0.02fF
C1551 VDD.n933 GND 0.29fF
C1552 VDD.n934 GND 0.01fF
C1553 VDD.n935 GND 0.02fF
C1554 VDD.n936 GND 0.02fF
C1555 VDD.n937 GND 0.29fF
C1556 VDD.n938 GND 0.01fF
C1557 VDD.n939 GND 0.02fF
C1558 VDD.n940 GND 0.04fF
C1559 VDD.n941 GND 0.33fF
C1560 VDD.n942 GND 0.02fF
C1561 VDD.n943 GND 0.02fF
C1562 VDD.n944 GND 0.02fF
C1563 VDD.n945 GND 0.06fF
C1564 VDD.n946 GND 0.02fF
C1565 VDD.n947 GND 0.02fF
C1566 VDD.n948 GND 0.02fF
C1567 VDD.n949 GND 0.02fF
C1568 VDD.n950 GND 0.02fF
C1569 VDD.n951 GND 0.02fF
C1570 VDD.n952 GND 0.02fF
C1571 VDD.n953 GND 0.02fF
C1572 VDD.n954 GND 0.02fF
C1573 VDD.n955 GND 0.02fF
C1574 VDD.n956 GND 0.03fF
C1575 VDD.n957 GND 0.02fF
C1576 VDD.n958 GND 0.02fF
C1577 VDD.n962 GND 0.29fF
C1578 VDD.n963 GND 0.29fF
C1579 VDD.n964 GND 0.01fF
C1580 VDD.n965 GND 0.02fF
C1581 VDD.n966 GND 0.04fF
C1582 VDD.n967 GND 0.29fF
C1583 VDD.n968 GND 0.01fF
C1584 VDD.n969 GND 0.02fF
C1585 VDD.n970 GND 0.02fF
C1586 VDD.n971 GND 0.07fF
C1587 VDD.n972 GND 0.24fF
C1588 VDD.n973 GND 0.01fF
C1589 VDD.n974 GND 0.01fF
C1590 VDD.n975 GND 0.02fF
C1591 VDD.n976 GND 0.18fF
C1592 VDD.n977 GND 0.01fF
C1593 VDD.n978 GND 0.02fF
C1594 VDD.n979 GND 0.02fF
C1595 VDD.n980 GND 0.09fF
C1596 VDD.n981 GND 0.05fF
C1597 VDD.n982 GND 0.17fF
C1598 VDD.n983 GND 0.01fF
C1599 VDD.n984 GND 0.02fF
C1600 VDD.n985 GND 0.02fF
C1601 VDD.n986 GND 0.16fF
C1602 VDD.n987 GND 0.02fF
C1603 VDD.n988 GND 0.02fF
C1604 VDD.n989 GND 0.03fF
C1605 VDD.n990 GND 0.15fF
C1606 VDD.n991 GND 0.02fF
C1607 VDD.n992 GND 0.02fF
C1608 VDD.n993 GND 0.03fF
C1609 VDD.n994 GND 0.17fF
C1610 VDD.n995 GND 0.01fF
C1611 VDD.n996 GND 0.09fF
C1612 VDD.n997 GND 0.05fF
C1613 VDD.n998 GND 0.02fF
C1614 VDD.n999 GND 0.02fF
C1615 VDD.n1000 GND 0.18fF
C1616 VDD.n1001 GND 0.01fF
C1617 VDD.n1002 GND 0.02fF
C1618 VDD.n1003 GND 0.02fF
C1619 VDD.n1004 GND 0.23fF
C1620 VDD.n1005 GND 0.01fF
C1621 VDD.n1006 GND 0.07fF
C1622 VDD.n1007 GND 0.02fF
C1623 VDD.n1008 GND 0.29fF
C1624 VDD.n1009 GND 0.01fF
C1625 VDD.n1010 GND 0.02fF
C1626 VDD.n1011 GND 0.02fF
C1627 VDD.n1012 GND 0.29fF
C1628 VDD.n1013 GND 0.01fF
C1629 VDD.n1014 GND 0.02fF
C1630 VDD.n1015 GND 0.04fF
C1631 VDD.n1016 GND 0.33fF
C1632 VDD.n1017 GND 0.02fF
C1633 VDD.n1018 GND 0.02fF
C1634 VDD.n1019 GND 0.02fF
C1635 VDD.n1020 GND 0.06fF
C1636 VDD.n1021 GND 0.02fF
C1637 VDD.n1022 GND 0.02fF
C1638 VDD.n1023 GND 0.02fF
C1639 VDD.n1024 GND 0.02fF
C1640 VDD.n1025 GND 0.02fF
C1641 VDD.n1026 GND 0.02fF
C1642 VDD.n1027 GND 0.02fF
C1643 VDD.n1028 GND 0.02fF
C1644 VDD.n1029 GND 0.02fF
C1645 VDD.n1030 GND 0.02fF
C1646 VDD.n1031 GND 0.03fF
C1647 VDD.n1032 GND 0.02fF
C1648 VDD.n1033 GND 0.02fF
C1649 VDD.n1037 GND 0.29fF
C1650 VDD.n1038 GND 0.29fF
C1651 VDD.n1039 GND 0.01fF
C1652 VDD.n1040 GND 0.02fF
C1653 VDD.n1041 GND 0.04fF
C1654 VDD.n1042 GND 0.29fF
C1655 VDD.n1043 GND 0.01fF
C1656 VDD.n1044 GND 0.02fF
C1657 VDD.n1045 GND 0.02fF
C1658 VDD.n1046 GND 0.07fF
C1659 VDD.n1047 GND 0.24fF
C1660 VDD.n1048 GND 0.01fF
C1661 VDD.n1049 GND 0.01fF
C1662 VDD.n1050 GND 0.02fF
C1663 VDD.n1051 GND 0.18fF
C1664 VDD.n1052 GND 0.01fF
C1665 VDD.n1053 GND 0.02fF
C1666 VDD.n1054 GND 0.02fF
C1667 VDD.n1055 GND 0.09fF
C1668 VDD.n1056 GND 0.05fF
C1669 VDD.n1057 GND 0.17fF
C1670 VDD.n1058 GND 0.01fF
C1671 VDD.n1059 GND 0.02fF
C1672 VDD.n1060 GND 0.02fF
C1673 VDD.n1061 GND 0.16fF
C1674 VDD.n1062 GND 0.02fF
C1675 VDD.n1063 GND 0.02fF
C1676 VDD.n1064 GND 0.03fF
C1677 VDD.n1065 GND 0.15fF
C1678 VDD.n1066 GND 0.02fF
C1679 VDD.n1067 GND 0.02fF
C1680 VDD.n1068 GND 0.03fF
C1681 VDD.n1069 GND 0.17fF
C1682 VDD.n1070 GND 0.01fF
C1683 VDD.n1071 GND 0.09fF
C1684 VDD.n1072 GND 0.05fF
C1685 VDD.n1073 GND 0.02fF
C1686 VDD.n1074 GND 0.02fF
C1687 VDD.n1075 GND 0.18fF
C1688 VDD.n1076 GND 0.01fF
C1689 VDD.n1077 GND 0.02fF
C1690 VDD.n1078 GND 0.02fF
C1691 VDD.n1079 GND 0.23fF
C1692 VDD.n1080 GND 0.01fF
C1693 VDD.n1081 GND 0.07fF
C1694 VDD.n1082 GND 0.02fF
C1695 VDD.n1083 GND 0.29fF
C1696 VDD.n1084 GND 0.01fF
C1697 VDD.n1085 GND 0.02fF
C1698 VDD.n1086 GND 0.02fF
C1699 VDD.n1087 GND 0.29fF
C1700 VDD.n1088 GND 0.01fF
C1701 VDD.n1089 GND 0.02fF
C1702 VDD.n1090 GND 0.04fF
C1703 VDD.n1091 GND 0.33fF
C1704 VDD.n1092 GND 0.02fF
C1705 VDD.n1093 GND 0.02fF
C1706 VDD.n1094 GND 0.02fF
C1707 VDD.n1095 GND 0.06fF
C1708 VDD.n1096 GND 0.02fF
C1709 VDD.n1097 GND 0.02fF
C1710 VDD.n1098 GND 0.02fF
C1711 VDD.n1099 GND 0.02fF
C1712 VDD.n1100 GND 0.02fF
C1713 VDD.n1101 GND 0.02fF
C1714 VDD.n1102 GND 0.02fF
C1715 VDD.n1103 GND 0.02fF
C1716 VDD.n1104 GND 0.02fF
C1717 VDD.n1105 GND 0.02fF
C1718 VDD.n1106 GND 0.03fF
C1719 VDD.n1107 GND 0.02fF
C1720 VDD.n1108 GND 0.02fF
C1721 VDD.n1112 GND 0.29fF
C1722 VDD.n1113 GND 0.29fF
C1723 VDD.n1114 GND 0.01fF
C1724 VDD.n1115 GND 0.02fF
C1725 VDD.n1116 GND 0.04fF
C1726 VDD.n1117 GND 0.29fF
C1727 VDD.n1118 GND 0.01fF
C1728 VDD.n1119 GND 0.02fF
C1729 VDD.n1120 GND 0.02fF
C1730 VDD.n1121 GND 0.07fF
C1731 VDD.n1122 GND 0.24fF
C1732 VDD.n1123 GND 0.01fF
C1733 VDD.n1124 GND 0.01fF
C1734 VDD.n1125 GND 0.02fF
C1735 VDD.n1126 GND 0.18fF
C1736 VDD.n1127 GND 0.01fF
C1737 VDD.n1128 GND 0.02fF
C1738 VDD.n1129 GND 0.02fF
C1739 VDD.n1130 GND 0.09fF
C1740 VDD.n1131 GND 0.05fF
C1741 VDD.n1132 GND 0.17fF
C1742 VDD.n1133 GND 0.01fF
C1743 VDD.n1134 GND 0.02fF
C1744 VDD.n1135 GND 0.02fF
C1745 VDD.n1136 GND 0.16fF
C1746 VDD.n1137 GND 0.02fF
C1747 VDD.n1138 GND 0.02fF
C1748 VDD.n1139 GND 0.03fF
C1749 VDD.n1140 GND 0.15fF
C1750 VDD.n1141 GND 0.02fF
C1751 VDD.n1142 GND 0.02fF
C1752 VDD.n1143 GND 0.03fF
C1753 VDD.n1144 GND 0.17fF
C1754 VDD.n1145 GND 0.01fF
C1755 VDD.n1146 GND 0.09fF
C1756 VDD.n1147 GND 0.05fF
C1757 VDD.n1148 GND 0.02fF
C1758 VDD.n1149 GND 0.02fF
C1759 VDD.n1150 GND 0.18fF
C1760 VDD.n1151 GND 0.01fF
C1761 VDD.n1152 GND 0.02fF
C1762 VDD.n1153 GND 0.02fF
C1763 VDD.n1154 GND 0.23fF
C1764 VDD.n1155 GND 0.01fF
C1765 VDD.n1156 GND 0.07fF
C1766 VDD.n1157 GND 0.02fF
C1767 VDD.n1158 GND 0.29fF
C1768 VDD.n1159 GND 0.01fF
C1769 VDD.n1160 GND 0.02fF
C1770 VDD.n1161 GND 0.02fF
C1771 VDD.n1162 GND 0.29fF
C1772 VDD.n1163 GND 0.01fF
C1773 VDD.n1164 GND 0.02fF
C1774 VDD.n1165 GND 0.04fF
C1775 VDD.n1166 GND 0.33fF
C1776 VDD.n1167 GND 0.02fF
C1777 VDD.n1168 GND 0.02fF
C1778 VDD.n1169 GND 0.02fF
C1779 VDD.n1170 GND 0.06fF
C1780 VDD.n1171 GND 0.02fF
C1781 VDD.n1172 GND 0.02fF
C1782 VDD.n1173 GND 0.02fF
C1783 VDD.n1174 GND 0.02fF
C1784 VDD.n1175 GND 0.02fF
C1785 VDD.n1176 GND 0.02fF
C1786 VDD.n1177 GND 0.02fF
C1787 VDD.n1178 GND 0.02fF
C1788 VDD.n1179 GND 0.02fF
C1789 VDD.n1180 GND 0.02fF
C1790 VDD.n1181 GND 0.03fF
C1791 VDD.n1182 GND 0.02fF
C1792 VDD.n1183 GND 0.02fF
C1793 VDD.n1187 GND 0.29fF
C1794 VDD.n1188 GND 0.29fF
C1795 VDD.n1189 GND 0.01fF
C1796 VDD.n1190 GND 0.02fF
C1797 VDD.n1191 GND 0.04fF
C1798 VDD.n1192 GND 0.29fF
C1799 VDD.n1193 GND 0.01fF
C1800 VDD.n1194 GND 0.02fF
C1801 VDD.n1195 GND 0.02fF
C1802 VDD.n1196 GND 0.07fF
C1803 VDD.n1197 GND 0.24fF
C1804 VDD.n1198 GND 0.01fF
C1805 VDD.n1199 GND 0.01fF
C1806 VDD.n1200 GND 0.02fF
C1807 VDD.n1201 GND 0.18fF
C1808 VDD.n1202 GND 0.01fF
C1809 VDD.n1203 GND 0.02fF
C1810 VDD.n1204 GND 0.02fF
C1811 VDD.n1205 GND 0.09fF
C1812 VDD.n1206 GND 0.05fF
C1813 VDD.n1207 GND 0.17fF
C1814 VDD.n1208 GND 0.01fF
C1815 VDD.n1209 GND 0.02fF
C1816 VDD.n1210 GND 0.02fF
C1817 VDD.n1211 GND 0.16fF
C1818 VDD.n1212 GND 0.02fF
C1819 VDD.n1213 GND 0.02fF
C1820 VDD.n1214 GND 0.03fF
C1821 VDD.n1215 GND 0.15fF
C1822 VDD.n1216 GND 0.02fF
C1823 VDD.n1217 GND 0.02fF
C1824 VDD.n1218 GND 0.03fF
C1825 VDD.n1219 GND 0.17fF
C1826 VDD.n1220 GND 0.01fF
C1827 VDD.n1221 GND 0.09fF
C1828 VDD.n1222 GND 0.05fF
C1829 VDD.n1223 GND 0.02fF
C1830 VDD.n1224 GND 0.02fF
C1831 VDD.n1225 GND 0.18fF
C1832 VDD.n1226 GND 0.01fF
C1833 VDD.n1227 GND 0.02fF
C1834 VDD.n1228 GND 0.02fF
C1835 VDD.n1229 GND 0.23fF
C1836 VDD.n1230 GND 0.01fF
C1837 VDD.n1231 GND 0.07fF
C1838 VDD.n1232 GND 0.02fF
C1839 VDD.n1233 GND 0.29fF
C1840 VDD.n1234 GND 0.01fF
C1841 VDD.n1235 GND 0.02fF
C1842 VDD.n1236 GND 0.02fF
C1843 VDD.n1237 GND 0.29fF
C1844 VDD.n1238 GND 0.01fF
C1845 VDD.n1239 GND 0.02fF
C1846 VDD.n1240 GND 0.04fF
C1847 VDD.n1241 GND 0.33fF
C1848 VDD.n1242 GND 0.02fF
C1849 VDD.n1243 GND 0.02fF
C1850 VDD.n1244 GND 0.02fF
C1851 VDD.n1245 GND 0.06fF
C1852 VDD.n1246 GND 0.02fF
C1853 VDD.n1247 GND 0.02fF
C1854 VDD.n1248 GND 0.02fF
C1855 VDD.n1249 GND 0.02fF
C1856 VDD.n1250 GND 0.02fF
C1857 VDD.n1251 GND 0.02fF
C1858 VDD.n1252 GND 0.02fF
C1859 VDD.n1253 GND 0.02fF
C1860 VDD.n1254 GND 0.02fF
C1861 VDD.n1255 GND 0.02fF
C1862 VDD.n1256 GND 0.03fF
C1863 VDD.n1257 GND 0.02fF
C1864 VDD.n1258 GND 0.02fF
C1865 VDD.n1262 GND 0.29fF
C1866 VDD.n1263 GND 0.29fF
C1867 VDD.n1264 GND 0.01fF
C1868 VDD.n1265 GND 0.02fF
C1869 VDD.n1266 GND 0.04fF
C1870 VDD.n1267 GND 0.29fF
C1871 VDD.n1268 GND 0.01fF
C1872 VDD.n1269 GND 0.02fF
C1873 VDD.n1270 GND 0.02fF
C1874 VDD.n1271 GND 0.07fF
C1875 VDD.n1272 GND 0.24fF
C1876 VDD.n1273 GND 0.01fF
C1877 VDD.n1274 GND 0.01fF
C1878 VDD.n1275 GND 0.02fF
C1879 VDD.n1276 GND 0.18fF
C1880 VDD.n1277 GND 0.01fF
C1881 VDD.n1278 GND 0.02fF
C1882 VDD.n1279 GND 0.02fF
C1883 VDD.n1280 GND 0.09fF
C1884 VDD.n1281 GND 0.05fF
C1885 VDD.n1282 GND 0.17fF
C1886 VDD.n1283 GND 0.01fF
C1887 VDD.n1284 GND 0.02fF
C1888 VDD.n1285 GND 0.02fF
C1889 VDD.n1286 GND 0.16fF
C1890 VDD.n1287 GND 0.02fF
C1891 VDD.n1288 GND 0.02fF
C1892 VDD.n1289 GND 0.03fF
C1893 VDD.n1290 GND 0.15fF
C1894 VDD.n1291 GND 0.02fF
C1895 VDD.n1292 GND 0.02fF
C1896 VDD.n1293 GND 0.03fF
C1897 VDD.n1294 GND 0.17fF
C1898 VDD.n1295 GND 0.01fF
C1899 VDD.n1296 GND 0.09fF
C1900 VDD.n1297 GND 0.05fF
C1901 VDD.n1298 GND 0.02fF
C1902 VDD.n1299 GND 0.02fF
C1903 VDD.n1300 GND 0.18fF
C1904 VDD.n1301 GND 0.01fF
C1905 VDD.n1302 GND 0.02fF
C1906 VDD.n1303 GND 0.02fF
C1907 VDD.n1304 GND 0.23fF
C1908 VDD.n1305 GND 0.01fF
C1909 VDD.n1306 GND 0.07fF
C1910 VDD.n1307 GND 0.02fF
C1911 VDD.n1308 GND 0.29fF
C1912 VDD.n1309 GND 0.01fF
C1913 VDD.n1310 GND 0.02fF
C1914 VDD.n1311 GND 0.02fF
C1915 VDD.n1312 GND 0.29fF
C1916 VDD.n1313 GND 0.01fF
C1917 VDD.n1314 GND 0.02fF
C1918 VDD.n1315 GND 0.04fF
C1919 VDD.n1316 GND 0.33fF
C1920 VDD.n1317 GND 0.02fF
C1921 VDD.n1318 GND 0.02fF
C1922 VDD.n1319 GND 0.02fF
C1923 VDD.n1320 GND 0.06fF
C1924 VDD.n1321 GND 0.02fF
C1925 VDD.n1322 GND 0.02fF
C1926 VDD.n1323 GND 0.02fF
C1927 VDD.n1324 GND 0.02fF
C1928 VDD.n1325 GND 0.02fF
C1929 VDD.n1326 GND 0.02fF
C1930 VDD.n1327 GND 0.02fF
C1931 VDD.n1328 GND 0.02fF
C1932 VDD.n1329 GND 0.02fF
C1933 VDD.n1330 GND 0.02fF
C1934 VDD.n1331 GND 0.03fF
C1935 VDD.n1332 GND 0.02fF
C1936 VDD.n1333 GND 0.02fF
C1937 VDD.n1337 GND 0.29fF
C1938 VDD.n1338 GND 0.29fF
C1939 VDD.n1339 GND 0.01fF
C1940 VDD.n1340 GND 0.02fF
C1941 VDD.n1341 GND 0.04fF
C1942 VDD.n1342 GND 0.29fF
C1943 VDD.n1343 GND 0.01fF
C1944 VDD.n1344 GND 0.02fF
C1945 VDD.n1345 GND 0.02fF
C1946 VDD.n1346 GND 0.07fF
C1947 VDD.n1347 GND 0.24fF
C1948 VDD.n1348 GND 0.01fF
C1949 VDD.n1349 GND 0.01fF
C1950 VDD.n1350 GND 0.02fF
C1951 VDD.n1351 GND 0.18fF
C1952 VDD.n1352 GND 0.01fF
C1953 VDD.n1353 GND 0.02fF
C1954 VDD.n1354 GND 0.02fF
C1955 VDD.n1355 GND 0.09fF
C1956 VDD.n1356 GND 0.05fF
C1957 VDD.n1357 GND 0.17fF
C1958 VDD.n1358 GND 0.01fF
C1959 VDD.n1359 GND 0.02fF
C1960 VDD.n1360 GND 0.02fF
C1961 VDD.n1361 GND 0.16fF
C1962 VDD.n1362 GND 0.02fF
C1963 VDD.n1363 GND 0.02fF
C1964 VDD.n1364 GND 0.03fF
C1965 VDD.n1365 GND 0.15fF
C1966 VDD.n1366 GND 0.02fF
C1967 VDD.n1367 GND 0.02fF
C1968 VDD.n1368 GND 0.03fF
C1969 VDD.n1369 GND 0.17fF
C1970 VDD.n1370 GND 0.01fF
C1971 VDD.n1371 GND 0.09fF
C1972 VDD.n1372 GND 0.05fF
C1973 VDD.n1373 GND 0.02fF
C1974 VDD.n1374 GND 0.02fF
C1975 VDD.n1375 GND 0.18fF
C1976 VDD.n1376 GND 0.01fF
C1977 VDD.n1377 GND 0.02fF
C1978 VDD.n1378 GND 0.02fF
C1979 VDD.n1379 GND 0.23fF
C1980 VDD.n1380 GND 0.01fF
C1981 VDD.n1381 GND 0.07fF
C1982 VDD.n1382 GND 0.02fF
C1983 VDD.n1383 GND 0.29fF
C1984 VDD.n1384 GND 0.01fF
C1985 VDD.n1385 GND 0.02fF
C1986 VDD.n1386 GND 0.02fF
C1987 VDD.n1387 GND 0.29fF
C1988 VDD.n1388 GND 0.01fF
C1989 VDD.n1389 GND 0.02fF
C1990 VDD.n1390 GND 0.04fF
C1991 VDD.n1391 GND 0.33fF
C1992 VDD.n1392 GND 0.02fF
C1993 VDD.n1393 GND 0.02fF
C1994 VDD.n1394 GND 0.02fF
C1995 VDD.n1395 GND 0.06fF
C1996 VDD.n1396 GND 0.02fF
C1997 VDD.n1397 GND 0.02fF
C1998 VDD.n1398 GND 0.02fF
C1999 VDD.n1399 GND 0.02fF
C2000 VDD.n1400 GND 0.02fF
C2001 VDD.n1401 GND 0.02fF
C2002 VDD.n1402 GND 0.02fF
C2003 VDD.n1403 GND 0.02fF
C2004 VDD.n1404 GND 0.02fF
C2005 VDD.n1405 GND 0.02fF
C2006 VDD.n1406 GND 0.03fF
C2007 VDD.n1407 GND 0.02fF
C2008 VDD.n1408 GND 0.02fF
C2009 VDD.n1412 GND 0.29fF
C2010 VDD.n1413 GND 0.29fF
C2011 VDD.n1414 GND 0.01fF
C2012 VDD.n1415 GND 0.02fF
C2013 VDD.n1416 GND 0.04fF
C2014 VDD.n1417 GND 0.29fF
C2015 VDD.n1418 GND 0.01fF
C2016 VDD.n1419 GND 0.02fF
C2017 VDD.n1420 GND 0.02fF
C2018 VDD.n1421 GND 0.07fF
C2019 VDD.n1422 GND 0.24fF
C2020 VDD.n1423 GND 0.01fF
C2021 VDD.n1424 GND 0.01fF
C2022 VDD.n1425 GND 0.02fF
C2023 VDD.n1426 GND 0.18fF
C2024 VDD.n1427 GND 0.01fF
C2025 VDD.n1428 GND 0.02fF
C2026 VDD.n1429 GND 0.02fF
C2027 VDD.n1430 GND 0.09fF
C2028 VDD.n1431 GND 0.05fF
C2029 VDD.n1432 GND 0.17fF
C2030 VDD.n1433 GND 0.01fF
C2031 VDD.n1434 GND 0.02fF
C2032 VDD.n1435 GND 0.02fF
C2033 VDD.n1436 GND 0.16fF
C2034 VDD.n1437 GND 0.02fF
C2035 VDD.n1438 GND 0.02fF
C2036 VDD.n1439 GND 0.03fF
C2037 VDD.n1440 GND 0.15fF
C2038 VDD.n1441 GND 0.02fF
C2039 VDD.n1442 GND 0.02fF
C2040 VDD.n1443 GND 0.03fF
C2041 VDD.n1444 GND 0.17fF
C2042 VDD.n1445 GND 0.01fF
C2043 VDD.n1446 GND 0.09fF
C2044 VDD.n1447 GND 0.05fF
C2045 VDD.n1448 GND 0.02fF
C2046 VDD.n1449 GND 0.02fF
C2047 VDD.n1450 GND 0.18fF
C2048 VDD.n1451 GND 0.01fF
C2049 VDD.n1452 GND 0.02fF
C2050 VDD.n1453 GND 0.02fF
C2051 VDD.n1454 GND 0.23fF
C2052 VDD.n1455 GND 0.01fF
C2053 VDD.n1456 GND 0.07fF
C2054 VDD.n1457 GND 0.02fF
C2055 VDD.n1458 GND 0.29fF
C2056 VDD.n1459 GND 0.01fF
C2057 VDD.n1460 GND 0.02fF
C2058 VDD.n1461 GND 0.02fF
C2059 VDD.n1462 GND 0.29fF
C2060 VDD.n1463 GND 0.01fF
C2061 VDD.n1464 GND 0.02fF
C2062 VDD.n1465 GND 0.04fF
C2063 VDD.n1466 GND 0.33fF
C2064 VDD.n1467 GND 0.02fF
C2065 VDD.n1468 GND 0.02fF
C2066 VDD.n1469 GND 0.02fF
C2067 VDD.n1470 GND 0.06fF
C2068 VDD.n1471 GND 0.02fF
C2069 VDD.n1472 GND 0.02fF
C2070 VDD.n1473 GND 0.02fF
C2071 VDD.n1474 GND 0.02fF
C2072 VDD.n1475 GND 0.02fF
C2073 VDD.n1476 GND 0.02fF
C2074 VDD.n1477 GND 0.02fF
C2075 VDD.n1478 GND 0.02fF
C2076 VDD.n1479 GND 0.02fF
C2077 VDD.n1480 GND 0.02fF
C2078 VDD.n1481 GND 0.03fF
C2079 VDD.n1482 GND 0.02fF
C2080 VDD.n1483 GND 0.02fF
C2081 VDD.n1487 GND 0.29fF
C2082 VDD.n1488 GND 0.29fF
C2083 VDD.n1489 GND 0.01fF
C2084 VDD.n1490 GND 0.02fF
C2085 VDD.n1491 GND 0.04fF
C2086 VDD.n1492 GND 0.29fF
C2087 VDD.n1493 GND 0.01fF
C2088 VDD.n1494 GND 0.02fF
C2089 VDD.n1495 GND 0.02fF
C2090 VDD.n1496 GND 0.07fF
C2091 VDD.n1497 GND 0.24fF
C2092 VDD.n1498 GND 0.01fF
C2093 VDD.n1499 GND 0.01fF
C2094 VDD.n1500 GND 0.02fF
C2095 VDD.n1501 GND 0.18fF
C2096 VDD.n1502 GND 0.01fF
C2097 VDD.n1503 GND 0.02fF
C2098 VDD.n1504 GND 0.02fF
C2099 VDD.n1505 GND 0.09fF
C2100 VDD.n1506 GND 0.05fF
C2101 VDD.n1507 GND 0.17fF
C2102 VDD.n1508 GND 0.01fF
C2103 VDD.n1509 GND 0.02fF
C2104 VDD.n1510 GND 0.02fF
C2105 VDD.n1511 GND 0.16fF
C2106 VDD.n1512 GND 0.02fF
C2107 VDD.n1513 GND 0.02fF
C2108 VDD.n1514 GND 0.03fF
C2109 VDD.n1515 GND 0.15fF
C2110 VDD.n1516 GND 0.02fF
C2111 VDD.n1517 GND 0.02fF
C2112 VDD.n1518 GND 0.03fF
C2113 VDD.n1519 GND 0.17fF
C2114 VDD.n1520 GND 0.01fF
C2115 VDD.n1521 GND 0.09fF
C2116 VDD.n1522 GND 0.05fF
C2117 VDD.n1523 GND 0.02fF
C2118 VDD.n1524 GND 0.02fF
C2119 VDD.n1525 GND 0.18fF
C2120 VDD.n1526 GND 0.01fF
C2121 VDD.n1527 GND 0.02fF
C2122 VDD.n1528 GND 0.02fF
C2123 VDD.n1529 GND 0.23fF
C2124 VDD.n1530 GND 0.01fF
C2125 VDD.n1531 GND 0.07fF
C2126 VDD.n1532 GND 0.02fF
C2127 VDD.n1533 GND 0.29fF
C2128 VDD.n1534 GND 0.01fF
C2129 VDD.n1535 GND 0.02fF
C2130 VDD.n1536 GND 0.02fF
C2131 VDD.n1537 GND 0.29fF
C2132 VDD.n1538 GND 0.01fF
C2133 VDD.n1539 GND 0.02fF
C2134 VDD.n1540 GND 0.04fF
C2135 VDD.n1541 GND 0.33fF
C2136 VDD.n1542 GND 0.02fF
C2137 VDD.n1543 GND 0.02fF
C2138 VDD.n1544 GND 0.02fF
C2139 VDD.n1545 GND 0.06fF
C2140 VDD.n1546 GND 0.02fF
C2141 VDD.n1547 GND 0.02fF
C2142 VDD.n1548 GND 0.02fF
C2143 VDD.n1549 GND 0.02fF
C2144 VDD.n1550 GND 0.02fF
C2145 VDD.n1551 GND 0.02fF
C2146 VDD.n1552 GND 0.02fF
C2147 VDD.n1553 GND 0.02fF
C2148 VDD.n1554 GND 0.02fF
C2149 VDD.n1555 GND 0.02fF
C2150 VDD.n1556 GND 0.03fF
C2151 VDD.n1557 GND 0.02fF
C2152 VDD.n1558 GND 0.02fF
C2153 VDD.n1562 GND 0.29fF
C2154 VDD.n1563 GND 0.29fF
C2155 VDD.n1564 GND 0.01fF
C2156 VDD.n1565 GND 0.02fF
C2157 VDD.n1566 GND 0.04fF
C2158 VDD.n1567 GND 0.29fF
C2159 VDD.n1568 GND 0.01fF
C2160 VDD.n1569 GND 0.02fF
C2161 VDD.n1570 GND 0.02fF
C2162 VDD.n1571 GND 0.07fF
C2163 VDD.n1572 GND 0.24fF
C2164 VDD.n1573 GND 0.01fF
C2165 VDD.n1574 GND 0.01fF
C2166 VDD.n1575 GND 0.02fF
C2167 a_15669_1050.n0 GND 0.38fF
C2168 a_15669_1050.n1 GND 0.38fF
C2169 a_15669_1050.n2 GND 0.48fF
C2170 a_15669_1050.n3 GND 0.45fF
C2171 a_15669_1050.n4 GND 0.43fF
C2172 a_15669_1050.n5 GND 0.31fF
C2173 a_15669_1050.n6 GND 0.63fF
C2174 a_15669_1050.n7 GND 0.68fF
C2175 a_15669_1050.n8 GND 0.08fF
C2176 a_15669_1050.n9 GND 0.21fF
C2177 a_15669_1050.n10 GND 0.04fF
C2178 a_13105_989.n0 GND 0.65fF
C2179 a_13105_989.n1 GND 0.65fF
C2180 a_13105_989.n2 GND 0.82fF
C2181 a_13105_989.n3 GND 0.78fF
C2182 a_13105_989.n4 GN