* SPICE3 file created from INVX1.ext - technology: sky130A

.subckt INVX1 Y A VDD GND
M1000 Y A GND GND nshort w=3u l=0.15u
+  ad=0.1791p pd=1.57u as=1.1408p ps=8.1u
M1001 Y.t2 A.t1 VDD.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 VDD.t0 A.t2 Y.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y A.t0 GND.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
C0 A Y 0.31fF
C1 Y VDD 0.76fF
C2 A VDD 0.12fF
R0 A.n0 A.t2 512.525
R1 A.n0 A.t1 371.139
R2 A.n1 A.t0 210.434
R3 A.n1 A.n0 173.2
R4 A.n2 A.n1 76
R5 A.n2 A 0.046
R6 GND.n9 GND.n1 76.145
R7 GND.n12 GND.n11 76
R8 GND.n9 GND.n8 76
R9 GND.n29 GND.n28 76
R10 GND.n21 GND.n20 76
R11 GND.n17 GND.t0 39.412
R12 GND.n5 GND.n4 35.01
R13 GND.n6 GND.n5 19.735
R14 GND.n26 GND.n25 19.735
R15 GND.n19 GND.n18 19.735
R16 GND.n5 GND.n3 19.017
R17 GND.n17 GND.n16 17.185
R18 GND.n20 GND.n13 13.653
R19 GND.n28 GND.n27 13.653
R20 GND.n8 GND.n7 13.653
R21 GND.n3 GND.n2 7.5
R22 GND.n24 GND.n23 7.5
R23 GND.n18 GND.n17 6.139
R24 GND.n15 GND.n14 4.551
R25 GND.n8 GND.n6 3.935
R26 GND.n20 GND.n19 3.541
R27 GND.t0 GND.n15 2.238
R28 GND.n23 GND.n22 1.935
R29 GND.n1 GND.n0 0.596
R30 GND.n11 GND.n10 0.596
R31 GND.n25 GND.n24 0.358
R32 GND.n12 GND 0.207
R33 GND.n28 GND.n26 0.196
R34 GND.n29 GND.n9 0.157
R35 GND.n29 GND.n21 0.157
R36 GND.n21 GND.n12 0.145
R37 Y.n2 Y.n1 200.754
R38 Y.n2 Y.n0 184.007
R39 Y.n3 Y.n2 76
R40 Y.n0 Y.t1 14.282
R41 Y.n0 Y.t2 14.282
R42 Y.n3 Y 0.046
R43 VDD.n26 VDD.n25 77.792
R44 VDD.n55 VDD.n54 77.792
R45 VDD.n29 VDD.n23 76.145
R46 VDD.n29 VDD.n28 76
R47 VDD.n63 VDD.n62 76
R48 VDD.n59 VDD.n58 76
R49 VDD.n53 VDD.n52 76
R50 VDD.n57 VDD.t1 55.106
R51 VDD.n24 VDD.t0 55.106
R52 VDD.n52 VDD.n49 21.841
R53 VDD.n23 VDD.n20 21.841
R54 VDD.n49 VDD.n31 14.167
R55 VDD.n31 VDD.n30 14.167
R56 VDD.n20 VDD.n19 14.167
R57 VDD.n19 VDD.n17 14.167
R58 VDD.n23 VDD.n22 13.653
R59 VDD.n22 VDD.n21 13.653
R60 VDD.n28 VDD.n27 13.653
R61 VDD.n27 VDD.n26 13.653
R62 VDD.n62 VDD.n61 13.653
R63 VDD.n61 VDD.n60 13.653
R64 VDD.n58 VDD.n56 13.653
R65 VDD.n56 VDD.n55 13.653
R66 VDD.n52 VDD.n51 13.653
R67 VDD.n51 VDD.n50 13.653
R68 VDD.n4 VDD.n2 12.915
R69 VDD.n4 VDD.n3 12.66
R70 VDD.n12 VDD.n11 12.343
R71 VDD.n10 VDD.n9 12.343
R72 VDD.n7 VDD.n6 12.343
R73 VDD.n35 VDD.n34 7.5
R74 VDD.n38 VDD.n37 7.5
R75 VDD.n40 VDD.n39 7.5
R76 VDD.n43 VDD.n42 7.5
R77 VDD.n49 VDD.n48 7.5
R78 VDD.n20 VDD.n16 7.5
R79 VDD.n2 VDD.n1 7.5
R80 VDD.n6 VDD.n5 7.5
R81 VDD.n9 VDD.n8 7.5
R82 VDD.n19 VDD.n18 7.5
R83 VDD.n14 VDD.n0 7.5
R84 VDD.n48 VDD.n47 6.772
R85 VDD.n36 VDD.n33 6.772
R86 VDD.n41 VDD.n38 6.772
R87 VDD.n45 VDD.n43 6.772
R88 VDD.n45 VDD.n44 6.772
R89 VDD.n41 VDD.n40 6.772
R90 VDD.n36 VDD.n35 6.772
R91 VDD.n47 VDD.n32 6.772
R92 VDD.n16 VDD.n15 6.458
R93 VDD.n28 VDD.n24 1.967
R94 VDD.n58 VDD.n57 1.967
R95 VDD.n14 VDD.n7 1.329
R96 VDD.n14 VDD.n10 1.329
R97 VDD.n14 VDD.n12 1.329
R98 VDD.n14 VDD.n13 1.329
R99 VDD.n15 VDD.n14 0.696
R100 VDD.n14 VDD.n4 0.696
R101 VDD.n46 VDD.n45 0.365
R102 VDD.n46 VDD.n41 0.365
R103 VDD.n46 VDD.n36 0.365
R104 VDD.n47 VDD.n46 0.365
R105 VDD.n53 VDD 0.207
R106 VDD.n63 VDD.n29 0.157
R107 VDD.n63 VDD.n59 0.157
R108 VDD.n59 VDD.n53 0.145
C3 VDD GND 2.55fF
C4 VDD.n0 GND 0.10fF
C5 VDD.n1 GND 0.02fF
C6 VDD.n2 GND 0.02fF
C7 VDD.n3 GND 0.04fF
C8 VDD.n4 GND 0.01fF
C9 VDD.n5 GND 0.02fF
C10 VDD.n6 GND 0.02fF
C11 VDD.n8 GND 0.02fF
C12 VDD.n9 GND 0.02fF
C13 VDD.n11 GND 0.02fF
C14 VDD.n14 GND 0.39fF
C15 VDD.n16 GND 0.03fF
C16 VDD.n17 GND 0.02fF
C17 VDD.n18 GND 0.02fF
C18 VDD.n19 GND 0.02fF
C19 VDD.n20 GND 0.03fF
C20 VDD.n21 GND 0.23fF
C21 VDD.n22 GND 0.02fF
C22 VDD.n23 GND 0.03fF
C23 VDD.n24 GND 0.05fF
C24 VDD.n25 GND 0.13fF
C25 VDD.n26 GND 0.17fF
C26 VDD.n27 GND 0.01fF
C27 VDD.n28 GND 0.01fF
C28 VDD.n29 GND 0.06fF
C29 VDD.n30 GND 0.02fF
C30 VDD.n31 GND 0.02fF
C31 VDD.n32 GND 0.02fF
C32 VDD.n33 GND 0.02fF
C33 VDD.n34 GND 0.02fF
C34 VDD.n35 GND 0.02fF
C35 VDD.n37 GND 0.02fF
C36 VDD.n38 GND 0.02fF
C37 VDD.n39 GND 0.02fF
C38 VDD.n40 GND 0.02fF
C39 VDD.n42 GND 0.03fF
C40 VDD.n43 GND 0.02fF
C41 VDD.n44 GND 0.10fF
C42 VDD.n46 GND 0.39fF
C43 VDD.n48 GND 0.03fF
C44 VDD.n49 GND 0.03fF
C45 VDD.n50 GND 0.23fF
C46 VDD.n51 GND 0.02fF
C47 VDD.n52 GND 0.03fF
C48 VDD.n53 GND 0.02fF
C49 VDD.n54 GND 0.13fF
C50 VDD.n55 GND 0.17fF
C51 VDD.n56 GND 0.01fF
C52 VDD.n57 GND 0.05fF
C53 VDD.n58 GND 0.01fF
C54 VDD.n59 GND 0.02fF
C55 VDD.n60 GND 0.14fF
C56 VDD.n61 GND 0.01fF
C57 VDD.n62 GND 0.02fF
C58 VDD.n63 GND 0.02fF
C59 Y.n0 GND 0.79fF
C60 Y.n1 GND 0.37fF
C61 Y.n2 GND 0.49fF
C62 Y.n3 GND 0.01fF
.ends
