* SPICE3 file created from TMRDFFQX1.ext - technology: sky130A

.subckt TMRDFFQX1 D CLK Q VDD GND
X0 GND a_3303_411.t6 a_14320_101.t0 GND sky130_fd_pr__nfet_01v8 ad=4.9019p pd=4.107u as=0p ps=0u w=0u l=0u
X1 VDD.t137 a_8731_187.t5 a_8861_1050.t4 PF;*V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X2 a_3177_1050.t3 a_277_1050.t7 VDD.t92 �aI*V sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X3 VDD.t59 a_1845_1050.t5 a_147_187.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X4 a_11887_411.t1 a_11761_1050.t5 VDD.t139 VDD.t138 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X5 VDD.t147 D.t0 a_9183_989.t1 |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X6 VDD.t150 D.t1 a_4891_989.t1 |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X7 VDD.t7 a_7469_1050.t5 a_7595_411.t1 |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X8 GND a_8731_187.t8 a_8675_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X9 VDD.t112 CLK.t0 a_277_1050.t4  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X10 GND a_7469_1050.t6 a_8030_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X11 a_13757_1051.t3 a_7595_411.t6 a_13268_209.t5 VDD.t115 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X12 a_3177_1050.t1 a_3303_411.t7 VDD.t21  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X13 VDD.t110 CLK.t1 a_147_187.t4 VDD.t109 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X14 a_11887_411.t4 a_8731_187.t7 VDD.t135  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X15 VDD.t28 a_11887_411.t5 a_11761_1050.t0 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X16 GND a_1845_1050.t6 a_2406_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X17 VDD.t108 CLK.t2 a_4439_187.t3  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X18 a_9183_989.t0 D.t2 VDD.t145 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X19 GND a_8861_1050.t8 a_9658_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X20 a_3303_411.t4 a_3177_1050.t5 VDD.t167  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X21 VDD.t40 a_599_989.t5 a_277_1050.t1 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X22 VDD.t156 a_277_1050.t9 a_599_989.t4  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X23 a_8731_187.t4 a_10429_1050.t5 VDD.t114 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X24 a_4569_1050.t3 a_4891_989.t6 VDD.t73  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X25 a_13757_1051.t5 a_3303_411.t8 a_13268_209.t2 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X26 VDD.t94 a_9183_989.t5 a_10429_1050.t1  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X27 VDD.t175 a_147_187.t6 a_3303_411.t1 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X28 a_7595_411.t0 a_7469_1050.t7 VDD.t5  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X29 Q.t1 a_13268_209.t7 VDD.t48 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X30 VDD.t32 a_4569_1050.t7 a_7469_1050.t0  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X31 a_4439_187.t2 CLK.t3 VDD.t106 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X32 a_1845_1050.t1 a_147_187.t7 VDD.t56  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X33 a_8861_1050.t1 a_9183_989.t6 VDD.t84 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X34 VDD.t34 a_4439_187.t5 a_4569_1050.t6  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X35 GND a_147_187.t10 a_91_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X36 a_6137_1050.t0 a_4439_187.t6 VDD.t3 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X37 a_9183_989.t4 a_8861_1050.t7 VDD.t125  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X38 GND a_8861_1050.t10 a_11656_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X39 a_13093_1051.t7 a_3303_411.t9 a_13757_1051.t7 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X40 a_11761_1050.t1 a_11887_411.t6 VDD.t77  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X41 a_3303_411.t0 a_147_187.t8 VDD.t165 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X42 VDD.t143 a_7595_411.t8 a_13093_1051.t5  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X43 VDD.t160 D.t4 a_599_989.t1 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X44 GND a_10429_1050.t6 a_10990_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X45 GND a_4439_187.t8 a_4383_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X46 a_13757_1051.t0 a_11887_411.t7 a_13093_1051.t3  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X47 a_8731_187.t3 CLK.t4 VDD.t104 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X48 VDD.t133 a_8731_187.t10 a_10429_1050.t3  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X49 a_277_1050.t0 a_147_187.t9 VDD.t23 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X50 a_4439_187.t1 a_6137_1050.t6 VDD.t81  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X51 VDD.t11 a_7595_411.t9 a_7469_1050.t3 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X52 VDD.t102 CLK.t5 a_4569_1050.t1  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X53 VDD.t158 a_599_989.t7 a_1845_1050.t3 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X54 a_11761_1050.t3 a_8861_1050.t9 VDD.t123  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X55 GND a_599_989.t8 a_1740_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X56 Q a_13268_209.t8 GND.t0 GND sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=0p ps=0u w=0u l=0u
X57 GND a_4569_1050.t8 a_5366_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X58 VDD.t65 a_11887_411.t8 a_13093_1051.t1 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X59 GND a_11887_411.t9 a_13654_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X60 a_4891_989.t0 D.t5 VDD.t15  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X61 a_13757_1051.t6 a_3303_411.t11 a_13093_1051.t6 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X62 GND a_11887_411.t10 a_12988_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X63 a_277_1050.t3 CLK.t8 VDD.t100  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X64 VDD.t71 a_4891_989.t8 a_4569_1050.t2 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X65 VDD.t25 a_277_1050.t10 a_3177_1050.t2  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X66 a_147_187.t3 CLK.t9 VDD.t96 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X67 VDD.t173 a_11761_1050.t6 a_11887_411.t0  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X68 GND a_3177_1050.t6 a_3738_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X69 GND a_4569_1050.t11 a_7364_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X70 a_4891_989.t3 a_4569_1050.t9 VDD.t17 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X71 GND a_9183_989.t8 a_10324_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X72 a_7595_411.t3 a_4439_187.t10 VDD.t152  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X73 a_277_1050.t6 a_599_989.t9 VDD.t171 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X74 a_599_989.t3 a_277_1050.t11 VDD.t52  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X75 a_8861_1050.t5 a_8731_187.t11 VDD.t131 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X76 a_13268_209.t3 a_3303_411.t12 a_13757_1051.t4  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X77 VDD.t63 CLK.t12 a_8731_187.t1 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X78 a_10429_1050.t0 a_9183_989.t7 VDD.t79  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X79 a_7469_1050.t1 a_4569_1050.t10 VDD.t42 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X80 a_147_187.t0 a_1845_1050.t7 VDD.t154  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X81 VDD.t75 a_3303_411.t13 a_3177_1050.t4 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X82 VDD.t129 a_8731_187.t12 a_11887_411.t3  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X83 VDD.t90 CLK.t14 a_8861_1050.t3 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X84 GND a_277_1050.t12 a_1074_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X85 a_4569_1050.t5 a_4439_187.t11 VDD.t162  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X86 VDD.t69 a_4891_989.t9 a_6137_1050.t4 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X87 VDD.t121 a_8861_1050.t11 a_11761_1050.t2  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X88 VDD.t61 a_3177_1050.t7 a_3303_411.t3 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X89 a_13093_1051.t4 a_7595_411.t11 VDD.t141  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X90 a_599_989.t0 D.t7 VDD.t9 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X91 VDD.t37 a_10429_1050.t7 a_8731_187.t0  |�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X92 a_13268_209.t6 a_7595_411.t12 a_13757_1051.t2 �{�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X93 a_10429_1050.t2 a_8731_187.t13 VDD.t127 0|�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X94 GND a_11761_1050.t7 a_12322_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X95 VDD.t54 a_13268_209.t9 Q.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X96 a_7469_1050.t2 a_7595_411.t13 VDD.t19 0|�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X97 VDD.t1 a_9183_989.t10 a_8861_1050.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X98 a_4569_1050.t0 CLK.t16 VDD.t88 0|�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X99 VDD.t13 a_4439_187.t12 a_6137_1050.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X100 VDD.t119 a_8861_1050.t12 a_9183_989.t3 0|�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X101 a_1845_1050.t4 a_599_989.t10 VDD.t169  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X102 a_8861_1050.t2 CLK.t17 VDD.t86 0|�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X103 GND a_6137_1050.t5 a_6698_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X104 a_13093_1051.t0 a_11887_411.t12 VDD.t46  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X105 GND a_277_1050.t8 a_3072_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X106 VDD.t44 a_147_187.t11 a_1845_1050.t0 0|�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X107 a_6137_1050.t3 a_4891_989.t10 VDD.t67  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X108 VDD.t117 a_4569_1050.t12 a_4891_989.t4 0|�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X109 a_13093_1051.t2 a_11887_411.t13 a_13757_1051.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X110 VDD.t98 a_4439_187.t13 a_7595_411.t2 0|�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X111 GND a_4891_989.t5 a_6032_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X112 VDD.t50 a_147_187.t13 a_277_1050.t2  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X113 VDD.t30 a_6137_1050.t7 a_4439_187.t0 0|�� sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
C0 VDD CLK 7.71fF
C1 VDD D 0.97fF
C2 CLK D 0.45fF
C3 VDD Q 1.05fF
R0 a_8731_187.n7 a_8731_187.t5 512.525
R1 a_8731_187.n5 a_8731_187.t10 472.359
R2 a_8731_187.n3 a_8731_187.t12 472.359
R3 a_8731_187.n8 a_8731_187.t8 417.109
R4 a_8731_187.n5 a_8731_187.t13 384.527
R5 a_8731_187.n3 a_8731_187.t7 384.527
R6 a_8731_187.n7 a_8731_187.t11 371.139
R7 a_8731_187.n6 a_8731_187.t6 370.613
R8 a_8731_187.n4 a_8731_187.t9 370.613
R9 a_8731_187.n13 a_8731_187.n11 367.82
R10 a_8731_187.n8 a_8731_187.n7 179.837
R11 a_8731_187.n2 a_8731_187.n1 157.964
R12 a_8731_187.n6 a_8731_187.n5 127.096
R13 a_8731_187.n4 a_8731_187.n3 127.096
R14 a_8731_187.n11 a_8731_187.n2 104.282
R15 a_8731_187.n2 a_8731_187.n0 91.706
R16 a_8731_187.n13 a_8731_187.n12 15.218
R17 a_8731_187.n0 a_8731_187.t1 14.282
R18 a_8731_187.n0 a_8731_187.t3 14.282
R19 a_8731_187.n1 a_8731_187.t0 14.282
R20 a_8731_187.n1 a_8731_187.t4 14.282
R21 a_8731_187.n14 a_8731_187.n13 12.014
R22 a_8731_187.n9 a_8731_187.n8 11.134
R23 a_8731_187.n10 a_8731_187.n4 8.957
R24 a_8731_187.n9 a_8731_187.n6 4.65
R25 a_8731_187.n11 a_8731_187.n10 4.65
R26 a_8731_187.n10 a_8731_187.n9 2.947
R27 a_8861_1050.n7 a_8861_1050.t12 480.392
R28 a_8861_1050.n5 a_8861_1050.t11 480.392
R29 a_8861_1050.n7 a_8861_1050.t7 403.272
R30 a_8861_1050.n5 a_8861_1050.t9 403.272
R31 a_8861_1050.n8 a_8861_1050.t8 385.063
R32 a_8861_1050.n6 a_8861_1050.t10 385.063
R33 a_8861_1050.n12 a_8861_1050.n10 342.597
R34 a_8861_1050.n3 a_8861_1050.n2 161.352
R35 a_8861_1050.n10 a_8861_1050.n4 151.34
R36 a_8861_1050.n8 a_8861_1050.n7 143.429
R37 a_8861_1050.n6 a_8861_1050.n5 143.429
R38 a_8861_1050.n4 a_8861_1050.n0 95.095
R39 a_8861_1050.n3 a_8861_1050.n1 95.095
R40 a_8861_1050.n4 a_8861_1050.n3 66.258
R41 a_8861_1050.n12 a_8861_1050.n11 15.218
R42 a_8861_1050.n0 a_8861_1050.t0 14.282
R43 a_8861_1050.n0 a_8861_1050.t1 14.282
R44 a_8861_1050.n1 a_8861_1050.t3 14.282
R45 a_8861_1050.n1 a_8861_1050.t2 14.282
R46 a_8861_1050.n2 a_8861_1050.t4 14.282
R47 a_8861_1050.n2 a_8861_1050.t5 14.282
R48 a_8861_1050.n13 a_8861_1050.n12 12.014
R49 a_8861_1050.n9 a_8861_1050.n6 11.95
R50 a_8861_1050.n10 a_8861_1050.n9 5.965
R51 a_8861_1050.n9 a_8861_1050.n8 4.65
R52 VDD.n754 VDD.n743 144.705
R53 VDD.n811 VDD.n804 144.705
R54 VDD.n868 VDD.n861 144.705
R55 VDD.n925 VDD.n918 144.705
R56 VDD.n982 VDD.n975 144.705
R57 VDD.n1039 VDD.n1032 144.705
R58 VDD.n1114 VDD.n1107 144.705
R59 VDD.n1171 VDD.n1164 144.705
R60 VDD.n1228 VDD.n1221 144.705
R61 VDD.n646 VDD.n639 144.705
R62 VDD.n1285 VDD.n1278 144.705
R63 VDD.n589 VDD.n582 144.705
R64 VDD.n514 VDD.n507 144.705
R65 VDD.n457 VDD.n450 144.705
R66 VDD.n400 VDD.n393 144.705
R67 VDD.n343 VDD.n336 144.705
R68 VDD.n286 VDD.n279 144.705
R69 VDD.n229 VDD.n222 144.705
R70 VDD.n172 VDD.n165 144.705
R71 VDD.n119 VDD.n112 144.705
R72 VDD.n66 VDD.n55 144.705
R73 VDD.n720 VDD.t40 143.754
R74 VDD.n1081 VDD.t71 143.754
R75 VDD.n523 VDD.t1 143.754
R76 VDD.n779 VDD.t160 143.754
R77 VDD.n836 VDD.t44 143.754
R78 VDD.n893 VDD.t110 143.754
R79 VDD.n950 VDD.t75 143.754
R80 VDD.n1007 VDD.t175 143.754
R81 VDD.n1139 VDD.t150 143.754
R82 VDD.n1196 VDD.t13 143.754
R83 VDD.n1253 VDD.t108 143.754
R84 VDD.n649 VDD.t11 143.754
R85 VDD.n592 VDD.t98 143.754
R86 VDD.n460 VDD.t147 143.754
R87 VDD.n403 VDD.t133 143.754
R88 VDD.n346 VDD.t63 143.754
R89 VDD.n289 VDD.t28 143.754
R90 VDD.n232 VDD.t129 143.754
R91 VDD.n197 VDD.t46 135.539
R92 VDD.n175 VDD.t143 135.539
R93 VDD.n685 VDD.t23 135.17
R94 VDD.n757 VDD.t52 135.17
R95 VDD.n814 VDD.t169 135.17
R96 VDD.n871 VDD.t154 135.17
R97 VDD.n928 VDD.t92 135.17
R98 VDD.n985 VDD.t167 135.17
R99 VDD.n1046 VDD.t162 135.17
R100 VDD.n1117 VDD.t17 135.17
R101 VDD.n1174 VDD.t67 135.17
R102 VDD.n1231 VDD.t81 135.17
R103 VDD.n1288 VDD.t42 135.17
R104 VDD.n614 VDD.t5 135.17
R105 VDD.n553 VDD.t131 135.17
R106 VDD.n482 VDD.t125 135.17
R107 VDD.n425 VDD.t79 135.17
R108 VDD.n368 VDD.t114 135.17
R109 VDD.n311 VDD.t123 135.17
R110 VDD.n254 VDD.t139 135.17
R111 VDD.n35 VDD.t48 135.17
R112 VDD.n24 VDD.t54 135.17
R113 VDD.n185 VDD.n184 129.849
R114 VDD.n695 VDD.n694 129.472
R115 VDD.n711 VDD.n710 129.472
R116 VDD.n771 VDD.n770 129.472
R117 VDD.n828 VDD.n827 129.472
R118 VDD.n885 VDD.n884 129.472
R119 VDD.n942 VDD.n941 129.472
R120 VDD.n999 VDD.n998 129.472
R121 VDD.n1056 VDD.n1055 129.472
R122 VDD.n1072 VDD.n1071 129.472
R123 VDD.n1131 VDD.n1130 129.472
R124 VDD.n1188 VDD.n1187 129.472
R125 VDD.n1245 VDD.n1244 129.472
R126 VDD.n1302 VDD.n1301 129.472
R127 VDD.n602 VDD.n601 129.472
R128 VDD.n544 VDD.n543 129.472
R129 VDD.n532 VDD.n531 129.472
R130 VDD.n470 VDD.n469 129.472
R131 VDD.n413 VDD.n412 129.472
R132 VDD.n356 VDD.n355 129.472
R133 VDD.n299 VDD.n298 129.472
R134 VDD.n242 VDD.n241 129.472
R135 VDD.n51 VDD.n50 92.5
R136 VDD.n49 VDD.n48 92.5
R137 VDD.n47 VDD.n46 92.5
R138 VDD.n45 VDD.n44 92.5
R139 VDD.n53 VDD.n52 92.5
R140 VDD.n108 VDD.n107 92.5
R141 VDD.n106 VDD.n105 92.5
R142 VDD.n104 VDD.n103 92.5
R143 VDD.n102 VDD.n101 92.5
R144 VDD.n110 VDD.n109 92.5
R145 VDD.n161 VDD.n160 92.5
R146 VDD.n159 VDD.n158 92.5
R147 VDD.n157 VDD.n156 92.5
R148 VDD.n155 VDD.n154 92.5
R149 VDD.n163 VDD.n162 92.5
R150 VDD.n218 VDD.n217 92.5
R151 VDD.n216 VDD.n215 92.5
R152 VDD.n214 VDD.n213 92.5
R153 VDD.n212 VDD.n211 92.5
R154 VDD.n220 VDD.n219 92.5
R155 VDD.n275 VDD.n274 92.5
R156 VDD.n273 VDD.n272 92.5
R157 VDD.n271 VDD.n270 92.5
R158 VDD.n269 VDD.n268 92.5
R159 VDD.n277 VDD.n276 92.5
R160 VDD.n332 VDD.n331 92.5
R161 VDD.n330 VDD.n329 92.5
R162 VDD.n328 VDD.n327 92.5
R163 VDD.n326 VDD.n325 92.5
R164 VDD.n334 VDD.n333 92.5
R165 VDD.n389 VDD.n388 92.5
R166 VDD.n387 VDD.n386 92.5
R167 VDD.n385 VDD.n384 92.5
R168 VDD.n383 VDD.n382 92.5
R169 VDD.n391 VDD.n390 92.5
R170 VDD.n446 VDD.n445 92.5
R171 VDD.n444 VDD.n443 92.5
R172 VDD.n442 VDD.n441 92.5
R173 VDD.n440 VDD.n439 92.5
R174 VDD.n448 VDD.n447 92.5
R175 VDD.n503 VDD.n502 92.5
R176 VDD.n501 VDD.n500 92.5
R177 VDD.n499 VDD.n498 92.5
R178 VDD.n497 VDD.n496 92.5
R179 VDD.n505 VDD.n504 92.5
R180 VDD.n578 VDD.n577 92.5
R181 VDD.n576 VDD.n575 92.5
R182 VDD.n574 VDD.n573 92.5
R183 VDD.n572 VDD.n571 92.5
R184 VDD.n580 VDD.n579 92.5
R185 VDD.n635 VDD.n634 92.5
R186 VDD.n633 VDD.n632 92.5
R187 VDD.n631 VDD.n630 92.5
R188 VDD.n629 VDD.n628 92.5
R189 VDD.n637 VDD.n636 92.5
R190 VDD.n1274 VDD.n1273 92.5
R191 VDD.n1272 VDD.n1271 92.5
R192 VDD.n1270 VDD.n1269 92.5
R193 VDD.n1268 VDD.n1267 92.5
R194 VDD.n1276 VDD.n1275 92.5
R195 VDD.n1217 VDD.n1216 92.5
R196 VDD.n1215 VDD.n1214 92.5
R197 VDD.n1213 VDD.n1212 92.5
R198 VDD.n1211 VDD.n1210 92.5
R199 VDD.n1219 VDD.n1218 92.5
R200 VDD.n1160 VDD.n1159 92.5
R201 VDD.n1158 VDD.n1157 92.5
R202 VDD.n1156 VDD.n1155 92.5
R203 VDD.n1154 VDD.n1153 92.5
R204 VDD.n1162 VDD.n1161 92.5
R205 VDD.n1103 VDD.n1102 92.5
R206 VDD.n1101 VDD.n1100 92.5
R207 VDD.n1099 VDD.n1098 92.5
R208 VDD.n1097 VDD.n1096 92.5
R209 VDD.n1105 VDD.n1104 92.5
R210 VDD.n1028 VDD.n1027 92.5
R211 VDD.n1026 VDD.n1025 92.5
R212 VDD.n1024 VDD.n1023 92.5
R213 VDD.n1022 VDD.n1021 92.5
R214 VDD.n1030 VDD.n1029 92.5
R215 VDD.n971 VDD.n970 92.5
R216 VDD.n969 VDD.n968 92.5
R217 VDD.n967 VDD.n966 92.5
R218 VDD.n965 VDD.n964 92.5
R219 VDD.n973 VDD.n972 92.5
R220 VDD.n914 VDD.n913 92.5
R221 VDD.n912 VDD.n911 92.5
R222 VDD.n910 VDD.n909 92.5
R223 VDD.n908 VDD.n907 92.5
R224 VDD.n916 VDD.n915 92.5
R225 VDD.n857 VDD.n856 92.5
R226 VDD.n855 VDD.n854 92.5
R227 VDD.n853 VDD.n852 92.5
R228 VDD.n851 VDD.n850 92.5
R229 VDD.n859 VDD.n858 92.5
R230 VDD.n800 VDD.n799 92.5
R231 VDD.n798 VDD.n797 92.5
R232 VDD.n796 VDD.n795 92.5
R233 VDD.n794 VDD.n793 92.5
R234 VDD.n802 VDD.n801 92.5
R235 VDD.n739 VDD.n738 92.5
R236 VDD.n737 VDD.n736 92.5
R237 VDD.n735 VDD.n734 92.5
R238 VDD.n733 VDD.n732 92.5
R239 VDD.n741 VDD.n740 92.5
R240 VDD.n669 VDD.n668 92.5
R241 VDD.n667 VDD.n666 92.5
R242 VDD.n665 VDD.n664 92.5
R243 VDD.n663 VDD.n662 92.5
R244 VDD.n671 VDD.n670 92.5
R245 VDD.n14 VDD.n1 92.5
R246 VDD.n5 VDD.n4 92.5
R247 VDD.n7 VDD.n6 92.5
R248 VDD.n9 VDD.n8 92.5
R249 VDD.n11 VDD.n10 92.5
R250 VDD.n13 VDD.n12 92.5
R251 VDD.n21 VDD.n20 92.059
R252 VDD.n65 VDD.n64 92.059
R253 VDD.n118 VDD.n117 92.059
R254 VDD.n171 VDD.n170 92.059
R255 VDD.n228 VDD.n227 92.059
R256 VDD.n285 VDD.n284 92.059
R257 VDD.n342 VDD.n341 92.059
R258 VDD.n399 VDD.n398 92.059
R259 VDD.n456 VDD.n455 92.059
R260 VDD.n513 VDD.n512 92.059
R261 VDD.n588 VDD.n587 92.059
R262 VDD.n645 VDD.n644 92.059
R263 VDD.n1284 VDD.n1283 92.059
R264 VDD.n1227 VDD.n1226 92.059
R265 VDD.n1170 VDD.n1169 92.059
R266 VDD.n1113 VDD.n1112 92.059
R267 VDD.n1038 VDD.n1037 92.059
R268 VDD.n981 VDD.n980 92.059
R269 VDD.n924 VDD.n923 92.059
R270 VDD.n867 VDD.n866 92.059
R271 VDD.n810 VDD.n809 92.059
R272 VDD.n753 VDD.n752 92.059
R273 VDD.n677 VDD.n676 92.059
R274 VDD.n20 VDD.n16 67.194
R275 VDD.n20 VDD.n17 67.194
R276 VDD.n20 VDD.n18 67.194
R277 VDD.n20 VDD.n19 67.194
R278 VDD.n661 VDD.n660 44.141
R279 VDD.n792 VDD.n791 44.141
R280 VDD.n849 VDD.n848 44.141
R281 VDD.n906 VDD.n905 44.141
R282 VDD.n963 VDD.n962 44.141
R283 VDD.n1020 VDD.n1019 44.141
R284 VDD.n1095 VDD.n1094 44.141
R285 VDD.n1152 VDD.n1151 44.141
R286 VDD.n1209 VDD.n1208 44.141
R287 VDD.n1266 VDD.n1265 44.141
R288 VDD.n627 VDD.n626 44.141
R289 VDD.n570 VDD.n569 44.141
R290 VDD.n495 VDD.n494 44.141
R291 VDD.n438 VDD.n437 44.141
R292 VDD.n381 VDD.n380 44.141
R293 VDD.n324 VDD.n323 44.141
R294 VDD.n267 VDD.n266 44.141
R295 VDD.n210 VDD.n209 44.141
R296 VDD.n153 VDD.n152 44.141
R297 VDD.n100 VDD.n99 44.141
R298 VDD.n5 VDD.n3 44.141
R299 VDD.n791 VDD.n789 44.107
R300 VDD.n848 VDD.n846 44.107
R301 VDD.n905 VDD.n903 44.107
R302 VDD.n962 VDD.n960 44.107
R303 VDD.n1019 VDD.n1017 44.107
R304 VDD.n1094 VDD.n1092 44.107
R305 VDD.n1151 VDD.n1149 44.107
R306 VDD.n1208 VDD.n1206 44.107
R307 VDD.n1265 VDD.n1263 44.107
R308 VDD.n626 VDD.n624 44.107
R309 VDD.n569 VDD.n567 44.107
R310 VDD.n494 VDD.n492 44.107
R311 VDD.n437 VDD.n435 44.107
R312 VDD.n380 VDD.n378 44.107
R313 VDD.n323 VDD.n321 44.107
R314 VDD.n266 VDD.n264 44.107
R315 VDD.n209 VDD.n207 44.107
R316 VDD.n152 VDD.n150 44.107
R317 VDD.n99 VDD.n97 44.107
R318 VDD.n660 VDD.n658 44.107
R319 VDD.n3 VDD.n2 44.107
R320 VDD.n25  43.472
R321 VDD.n33 �{�� 43.472
R322 VDD.n20 VDD.n15 41.052
R323 VDD.n59 VDD.n57 39.742
R324 VDD.n59 VDD.n58 39.742
R325 VDD.n61 VDD.n60 39.742
R326 VDD.n114 VDD.n113 39.742
R327 VDD.n167 VDD.n166 39.742
R328 VDD.n224 VDD.n223 39.742
R329 VDD.n281 VDD.n280 39.742
R330 VDD.n338 VDD.n337 39.742
R331 VDD.n395 VDD.n394 39.742
R332 VDD.n452 VDD.n451 39.742
R333 VDD.n509 VDD.n508 39.742
R334 VDD.n584 VDD.n583 39.742
R335 VDD.n641 VDD.n640 39.742
R336 VDD.n1280 VDD.n1279 39.742
R337 VDD.n1223 VDD.n1222 39.742
R338 VDD.n1166 VDD.n1165 39.742
R339 VDD.n1109 VDD.n1108 39.742
R340 VDD.n1034 VDD.n1033 39.742
R341 VDD.n977 VDD.n976 39.742
R342 VDD.n920 VDD.n919 39.742
R343 VDD.n863 VDD.n862 39.742
R344 VDD.n806 VDD.n805 39.742
R345 VDD.n673 VDD.n672 39.742
R346 VDD.n751 VDD.n748 39.742
R347 VDD.n751 VDD.n750 39.742
R348 VDD.n747 VDD.n746 39.742
R349 VDD.n99 VDD.n98 38
R350 VDD.n152 VDD.n151 38
R351 VDD.n209 VDD.n208 38
R352 VDD.n266 VDD.n265 38
R353 VDD.n323 VDD.n322 38
R354 VDD.n380 VDD.n379 38
R355 VDD.n437 VDD.n436 38
R356 VDD.n494 VDD.n493 38
R357 VDD.n569 VDD.n568 38
R358 VDD.n626 VDD.n625 38
R359 VDD.n1265 VDD.n1264 38
R360 VDD.n1208 VDD.n1207 38
R361 VDD.n1151 VDD.n1150 38
R362 VDD.n1094 VDD.n1093 38
R363 VDD.n1019 VDD.n1018 38
R364 VDD.n962 VDD.n961 38
R365 VDD.n905 VDD.n904 38
R366 VDD.n848 VDD.n847 38
R367 VDD.n791 VDD.n790 38
R368 VDD.n660 VDD.n659 38
R369 VDD.n789 VDD.n788 36.774
R370 VDD.n846 VDD.n845 36.774
R371 VDD.n903 VDD.n902 36.774
R372 VDD.n960 VDD.n959 36.774
R373 VDD.n1017 VDD.n1016 36.774
R374 VDD.n1092 VDD.n1091 36.774
R375 VDD.n1149 VDD.n1148 36.774
R376 VDD.n1206 VDD.n1205 36.774
R377 VDD.n1263 VDD.n1262 36.774
R378 VDD.n624 VDD.n623 36.774
R379 VDD.n567 VDD.n566 36.774
R380 VDD.n492 VDD.n491 36.774
R381 VDD.n435 VDD.n434 36.774
R382 VDD.n378 VDD.n377 36.774
R383 VDD.n321 VDD.n320 36.774
R384 VDD.n264 VDD.n263 36.774
R385 VDD.n207 VDD.n206 36.774
R386 VDD.n150 VDD.n149 36.774
R387 VDD.n97 VDD.n96 36.774
R388 VDD.n57 VDD.n56 36.774
R389 VDD.n750 VDD.n749 36.774
R390 VDD.n525  35.8
R391 VDD.n1075 �+V 35.8
R392 VDD.n714 �{�� 35.8
R393 VDD.n549 �{�� 33.243
R394 VDD.n1051  |�� 33.243
R395 VDD.n690 �;*V 33.243
R396 VDD.n1 VDD.n0 30.923
R397 VDD.n64 VDD.n62 26.38
R398 VDD.n64 VDD.n61 26.38
R399 VDD.n64 VDD.n59 26.38
R400 VDD.n64 VDD.n63 26.38
R401 VDD.n117 VDD.n115 26.38
R402 VDD.n117 VDD.n114 26.38
R403 VDD.n117 VDD.n116 26.38
R404 VDD.n170 VDD.n168 26.38
R405 VDD.n170 VDD.n167 26.38
R406 VDD.n170 VDD.n169 26.38
R407 VDD.n227 VDD.n225 26.38
R408 VDD.n227 VDD.n224 26.38
R409 VDD.n227 VDD.n226 26.38
R410 VDD.n284 VDD.n282 26.38
R411 VDD.n284 VDD.n281 26.38
R412 VDD.n284 VDD.n283 26.38
R413 VDD.n341 VDD.n339 26.38
R414 VDD.n341 VDD.n338 26.38
R415 VDD.n341 VDD.n340 26.38
R416 VDD.n398 VDD.n396 26.38
R417 VDD.n398 VDD.n395 26.38
R418 VDD.n398 VDD.n397 26.38
R419 VDD.n455 VDD.n453 26.38
R420 VDD.n455 VDD.n452 26.38
R421 VDD.n455 VDD.n454 26.38
R422 VDD.n512 VDD.n510 26.38
R423 VDD.n512 VDD.n509 26.38
R424 VDD.n512 VDD.n511 26.38
R425 VDD.n587 VDD.n585 26.38
R426 VDD.n587 VDD.n584 26.38
R427 VDD.n587 VDD.n586 26.38
R428 VDD.n644 VDD.n642 26.38
R429 VDD.n644 VDD.n641 26.38
R430 VDD.n644 VDD.n643 26.38
R431 VDD.n1283 VDD.n1281 26.38
R432 VDD.n1283 VDD.n1280 26.38
R433 VDD.n1283 VDD.n1282 26.38
R434 VDD.n1226 VDD.n1224 26.38
R435 VDD.n1226 VDD.n1223 26.38
R436 VDD.n1226 VDD.n1225 26.38
R437 VDD.n1169 VDD.n1167 26.38
R438 VDD.n1169 VDD.n1166 26.38
R439 VDD.n1169 VDD.n1168 26.38
R440 VDD.n1112 VDD.n1110 26.38
R441 VDD.n1112 VDD.n1109 26.38
R442 VDD.n1112 VDD.n1111 26.38
R443 VDD.n1037 VDD.n1035 26.38
R444 VDD.n1037 VDD.n1034 26.38
R445 VDD.n1037 VDD.n1036 26.38
R446 VDD.n980 VDD.n978 26.38
R447 VDD.n980 VDD.n977 26.38
R448 VDD.n980 VDD.n979 26.38
R449 VDD.n923 VDD.n921 26.38
R450 VDD.n923 VDD.n920 26.38
R451 VDD.n923 VDD.n922 26.38
R452 VDD.n866 VDD.n864 26.38
R453 VDD.n866 VDD.n863 26.38
R454 VDD.n866 VDD.n865 26.38
R455 VDD.n809 VDD.n807 26.38
R456 VDD.n809 VDD.n806 26.38
R457 VDD.n809 VDD.n808 26.38
R458 VDD.n676 VDD.n674 26.38
R459 VDD.n676 VDD.n673 26.38
R460 VDD.n676 VDD.n675 26.38
R461 VDD.n752 VDD.n751 26.38
R462 VDD.n752 VDD.n747 26.38
R463 VDD.n752 VDD.n745 26.38
R464 VDD.n752 VDD.n744 26.38
R465 VDD.n679 VDD.n671 22.915
R466 VDD.n23 VDD.n14 22.915
R467 VDD.n73 VDD.t115 20.457
R468 VDD.n137  |�� 20.457
R469 VDD.n180  |�� 20.457
R470 VDD.n237  |�� 20.457
R471 VDD.n294 `[�*V 20.457
R472 VDD.n351 �{�� 20.457
R473 VDD.n408  |�� 20.457
R474 VDD.n465 |�� 20.457
R475 VDD.n597 0|�� 20.457
R476 VDD.n654 �{�� 20.457
R477 VDD.n1249  |�� 20.457
R478 VDD.n1192  20.457
R479 VDD.n1135 |�� 20.457
R480 VDD.n1003 �{�� 20.457
R481 VDD.n946 �{�� 20.457
R482 VDD.n889 VDD.t109 20.457
R483 VDD.n832 0|�� 20.457
R484 VDD.n775 �{�� 20.457
R485 VDD.n84  |�� 17.9
R486 VDD.n126 �{�� 17.9
R487 VDD.n193  17.9
R488 VDD.n250 VDD.t138 17.9
R489 VDD.n307  |�� 17.9
R490 VDD.n364 �{�� 17.9
R491 VDD.n421  |�� 17.9
R492 VDD.n478  |�� 17.9
R493 VDD.n610  |�� 17.9
R494 VDD.n1293 �{�� 17.9
R495 VDD.n1236  |�� 17.9
R496 VDD.n1179  17.9
R497 VDD.n1122 �{�� 17.9
R498 VDD.n990  |�� 17.9
R499 VDD.n933 �aI*V 17.9
R500 VDD.n876  |�� 17.9
R501 VDD.n819  17.9
R502 VDD.n762  |�� 17.9
R503 VDD.n529 �Xl*V 15.343
R504 VDD.n1069  |�� 15.343
R505 VDD.n708 �{�� 15.343
R506 VDD.n671 VDD.n669 14.864
R507 VDD.n669 VDD.n667 14.864
R508 VDD.n667 VDD.n665 14.864
R509 VDD.n665 VDD.n663 14.864
R510 VDD.n663 VDD.n661 14.864
R511 VDD.n802 VDD.n800 14.864
R512 VDD.n800 VDD.n798 14.864
R513 VDD.n798 VDD.n796 14.864
R514 VDD.n796 VDD.n794 14.864
R515 VDD.n794 VDD.n792 14.864
R516 VDD.n859 VDD.n857 14.864
R517 VDD.n857 VDD.n855 14.864
R518 VDD.n855 VDD.n853 14.864
R519 VDD.n853 VDD.n851 14.864
R520 VDD.n851 VDD.n849 14.864
R521 VDD.n916 VDD.n914 14.864
R522 VDD.n914 VDD.n912 14.864
R523 VDD.n912 VDD.n910 14.864
R524 VDD.n910 VDD.n908 14.864
R525 VDD.n908 VDD.n906 14.864
R526 VDD.n973 VDD.n971 14.864
R527 VDD.n971 VDD.n969 14.864
R528 VDD.n969 VDD.n967 14.864
R529 VDD.n967 VDD.n965 14.864
R530 VDD.n965 VDD.n963 14.864
R531 VDD.n1030 VDD.n1028 14.864
R532 VDD.n1028 VDD.n1026 14.864
R533 VDD.n1026 VDD.n1024 14.864
R534 VDD.n1024 VDD.n1022 14.864
R535 VDD.n1022 VDD.n1020 14.864
R536 VDD.n1105 VDD.n1103 14.864
R537 VDD.n1103 VDD.n1101 14.864
R538 VDD.n1101 VDD.n1099 14.864
R539 VDD.n1099 VDD.n1097 14.864
R540 VDD.n1097 VDD.n1095 14.864
R541 VDD.n1162 VDD.n1160 14.864
R542 VDD.n1160 VDD.n1158 14.864
R543 VDD.n1158 VDD.n1156 14.864
R544 VDD.n1156 VDD.n1154 14.864
R545 VDD.n1154 VDD.n1152 14.864
R546 VDD.n1219 VDD.n1217 14.864
R547 VDD.n1217 VDD.n1215 14.864
R548 VDD.n1215 VDD.n1213 14.864
R549 VDD.n1213 VDD.n1211 14.864
R550 VDD.n1211 VDD.n1209 14.864
R551 VDD.n1276 VDD.n1274 14.864
R552 VDD.n1274 VDD.n1272 14.864
R553 VDD.n1272 VDD.n1270 14.864
R554 VDD.n1270 VDD.n1268 14.864
R555 VDD.n1268 VDD.n1266 14.864
R556 VDD.n637 VDD.n635 14.864
R557 VDD.n635 VDD.n633 14.864
R558 VDD.n633 VDD.n631 14.864
R559 VDD.n631 VDD.n629 14.864
R560 VDD.n629 VDD.n627 14.864
R561 VDD.n580 VDD.n578 14.864
R562 VDD.n578 VDD.n576 14.864
R563 VDD.n576 VDD.n574 14.864
R564 VDD.n574 VDD.n572 14.864
R565 VDD.n572 VDD.n570 14.864
R566 VDD.n505 VDD.n503 14.864
R567 VDD.n503 VDD.n501 14.864
R568 VDD.n501 VDD.n499 14.864
R569 VDD.n499 VDD.n497 14.864
R570 VDD.n497 VDD.n495 14.864
R571 VDD.n448 VDD.n446 14.864
R572 VDD.n446 VDD.n444 14.864
R573 VDD.n444 VDD.n442 14.864
R574 VDD.n442 VDD.n440 14.864
R575 VDD.n440 VDD.n438 14.864
R576 VDD.n391 VDD.n389 14.864
R577 VDD.n389 VDD.n387 14.864
R578 VDD.n387 VDD.n385 14.864
R579 VDD.n385 VDD.n383 14.864
R580 VDD.n383 VDD.n381 14.864
R581 VDD.n334 VDD.n332 14.864
R582 VDD.n332 VDD.n330 14.864
R583 VDD.n330 VDD.n328 14.864
R584 VDD.n328 VDD.n326 14.864
R585 VDD.n326 VDD.n324 14.864
R586 VDD.n277 VDD.n275 14.864
R587 VDD.n275 VDD.n273 14.864
R588 VDD.n273 VDD.n271 14.864
R589 VDD.n271 VDD.n269 14.864
R590 VDD.n269 VDD.n267 14.864
R591 VDD.n220 VDD.n218 14.864
R592 VDD.n218 VDD.n216 14.864
R593 VDD.n216 VDD.n214 14.864
R594 VDD.n214 VDD.n212 14.864
R595 VDD.n212 VDD.n210 14.864
R596 VDD.n163 VDD.n161 14.864
R597 VDD.n161 VDD.n159 14.864
R598 VDD.n159 VDD.n157 14.864
R599 VDD.n157 VDD.n155 14.864
R600 VDD.n155 VDD.n153 14.864
R601 VDD.n110 VDD.n108 14.864
R602 VDD.n108 VDD.n106 14.864
R603 VDD.n106 VDD.n104 14.864
R604 VDD.n104 VDD.n102 14.864
R605 VDD.n102 VDD.n100 14.864
R606 VDD.n53 VDD.n51 14.864
R607 VDD.n51 VDD.n49 14.864
R608 VDD.n49 VDD.n47 14.864
R609 VDD.n47 VDD.n45 14.864
R610 VDD.n45 VDD.n43 14.864
R611 VDD.n43 VDD.n42 14.864
R612 VDD.n741 VDD.n739 14.864
R613 VDD.n739 VDD.n737 14.864
R614 VDD.n737 VDD.n735 14.864
R615 VDD.n735 VDD.n733 14.864
R616 VDD.n733 VDD.n731 14.864
R617 VDD.n731 VDD.n730 14.864
R618 VDD.n14 VDD.n13 14.864
R619 VDD.n13 VDD.n11 14.864
R620 VDD.n11 VDD.n9 14.864
R621 VDD.n9 VDD.n7 14.864
R622 VDD.n7 VDD.n5 14.864
R623 VDD.n67 VDD.n54 14.864
R624 VDD.n120 VDD.n111 14.864
R625 VDD.n173 VDD.n164 14.864
R626 VDD.n230 VDD.n221 14.864
R627 VDD.n287 VDD.n278 14.864
R628 VDD.n344 VDD.n335 14.864
R629 VDD.n401 VDD.n392 14.864
R630 VDD.n458 VDD.n449 14.864
R631 VDD.n515 VDD.n506 14.864
R632 VDD.n590 VDD.n581 14.864
R633 VDD.n647 VDD.n638 14.864
R634 VDD.n1286 VDD.n1277 14.864
R635 VDD.n1229 VDD.n1220 14.864
R636 VDD.n1172 VDD.n1163 14.864
R637 VDD.n1115 VDD.n1106 14.864
R638 VDD.n1040 VDD.n1031 14.864
R639 VDD.n983 VDD.n974 14.864
R640 VDD.n926 VDD.n917 14.864
R641 VDD.n869 VDD.n860 14.864
R642 VDD.n812 VDD.n803 14.864
R643 VDD.n755 VDD.n742 14.864
R644 VDD.n694 VDD.t100 14.282
R645 VDD.n694 VDD.t50 14.282
R646 VDD.n710 VDD.t171 14.282
R647 VDD.n710 VDD.t112 14.282
R648 VDD.n770 VDD.t9 14.282
R649 VDD.n770 VDD.t156 14.282
R650 VDD.n827 VDD.t56 14.282
R651 VDD.n827 VDD.t158 14.282
R652 VDD.n884 VDD.t96 14.282
R653 VDD.n884 VDD.t59 14.282
R654 VDD.n941 VDD.t21 14.282
R655 VDD.n941 VDD.t25 14.282
R656 VDD.n998 VDD.t165 14.282
R657 VDD.n998 VDD.t61 14.282
R658 VDD.n1055 VDD.t88 14.282
R659 VDD.n1055 VDD.t34 14.282
R660 VDD.n1071 VDD.t73 14.282
R661 VDD.n1071 VDD.t102 14.282
R662 VDD.n1130 VDD.t15 14.282
R663 VDD.n1130 VDD.t117 14.282
R664 VDD.n1187 VDD.t3 14.282
R665 VDD.n1187 VDD.t69 14.282
R666 VDD.n1244 VDD.t106 14.282
R667 VDD.n1244 VDD.t30 14.282
R668 VDD.n1301 VDD.t19 14.282
R669 VDD.n1301 VDD.t32 14.282
R670 VDD.n601 VDD.t152 14.282
R671 VDD.n601 VDD.t7 14.282
R672 VDD.n543 VDD.t86 14.282
R673 VDD.n543 VDD.t137 14.282
R674 VDD.n531 VDD.t84 14.282
R675 VDD.n531 VDD.t90 14.282
R676 VDD.n469 VDD.t145 14.282
R677 VDD.n469 VDD.t119 14.282
R678 VDD.n412 VDD.t127 14.282
R679 VDD.n412 VDD.t94 14.282
R680 VDD.n355 VDD.t104 14.282
R681 VDD.n355 VDD.t37 14.282
R682 VDD.n298 VDD.t77 14.282
R683 VDD.n298 VDD.t121 14.282
R684 VDD.n241 VDD.t135 14.282
R685 VDD.n241 VDD.t173 14.282
R686 VDD.n184 VDD.t141 14.282
R687 VDD.n184 VDD.t65 14.282
R688 VDD.n545 PF;*V 12.786
R689 VDD.n1057  |�� 12.786
R690 VDD.n696  12.786
R691 VDD.n187 VDD.n185 9.083
R692 VDD.n244 VDD.n242 9.083
R693 VDD.n301 VDD.n299 9.083
R694 VDD.n358 VDD.n356 9.083
R695 VDD.n415 VDD.n413 9.083
R696 VDD.n472 VDD.n470 9.083
R697 VDD.n604 VDD.n602 9.083
R698 VDD.n1304 VDD.n1302 9.083
R699 VDD.n1247 VDD.n1245 9.083
R700 VDD.n1190 VDD.n1188 9.083
R701 VDD.n1133 VDD.n1131 9.083
R702 VDD.n1001 VDD.n999 9.083
R703 VDD.n944 VDD.n942 9.083
R704 VDD.n887 VDD.n885 9.083
R705 VDD.n830 VDD.n828 9.083
R706 VDD.n773 VDD.n771 9.083
R707 VDD.n23 VDD.n22 8.855
R708 VDD.n22 VDD.n21 8.855
R709 VDD.n27 VDD.n26 8.855
R710 VDD.n26 VDD.n25 8.855
R711 VDD.n31 VDD.n30 8.855
R712 VDD.n30 VDD.n29 8.855
R713 VDD.n36 VDD.n34 8.855
R714 VDD.n34 VDD.n33 8.855
R715 VDD.n40 VDD.n39 8.855
R716 VDD.n39 VDD.n38 8.855
R717 VDD.n67 VDD.n66 8.855
R718 VDD.n66 VDD.n65 8.855
R719 VDD.n71 VDD.n70 8.855
R720 VDD.n70 VDD.n69 8.855
R721 VDD.n75 VDD.n74 8.855
R722 VDD.n74 VDD.n73 8.855
R723 VDD.n78 VDD.n77 8.855
R724 VDD.n77 �{�� 8.855
R725 VDD.n82 VDD.n81 8.855
R726 VDD.n81 VDD.n80 8.855
R727 VDD.n86 VDD.n85 8.855
R728 VDD.n85 VDD.n84 8.855
R729 VDD.n90 VDD.n89 8.855
R730 VDD.n89 VDD.n88 8.855
R731 VDD.n94 VDD.n93 8.855
R732 VDD.n93 VDD.n92 8.855
R733 VDD.n120 VDD.n119 8.855
R734 VDD.n119 VDD.n118 8.855
R735 VDD.n124 VDD.n123 8.855
R736 VDD.n123 VDD.n122 8.855
R737 VDD.n128 VDD.n127 8.855
R738 VDD.n127 VDD.n126 8.855
R739 VDD.n132 VDD.n131 8.855
R740 VDD.n131 VDD.n130 8.855
R741 VDD.n135 VDD.n134 8.855
R742 VDD.n134  8.855
R743 VDD.n139 VDD.n138 8.855
R744 VDD.n138 VDD.n137 8.855
R745 VDD.n143 VDD.n142 8.855
R746 VDD.n142 VDD.n141 8.855
R747 VDD.n147 VDD.n146 8.855
R748 VDD.n146 VDD.n145 8.855
R749 VDD.n173 VDD.n172 8.855
R750 VDD.n172 VDD.n171 8.855
R751 VDD.n178 VDD.n177 8.855
R752 VDD.n177 VDD.n176 8.855
R753 VDD.n182 VDD.n181 8.855
R754 VDD.n181 VDD.n180 8.855
R755 VDD.n187 VDD.n186 8.855
R756 VDD.n186  |�� 8.855
R757 VDD.n191 VDD.n190 8.855
R758 VDD.n190 VDD.n189 8.855
R759 VDD.n195 VDD.n194 8.855
R760 VDD.n194 VDD.n193 8.855
R761 VDD.n200 VDD.n199 8.855
R762 VDD.n199 VDD.n198 8.855
R763 VDD.n204 VDD.n203 8.855
R764 VDD.n203 VDD.n202 8.855
R765 VDD.n230 VDD.n229 8.855
R766 VDD.n229 VDD.n228 8.855
R767 VDD.n235 VDD.n234 8.855
R768 VDD.n234 VDD.n233 8.855
R769 VDD.n239 VDD.n238 8.855
R770 VDD.n238 VDD.n237 8.855
R771 VDD.n244 VDD.n243 8.855
R772 VDD.n243  |�� 8.855
R773 VDD.n248 VDD.n247 8.855
R774 VDD.n247 VDD.n246 8.855
R775 VDD.n252 VDD.n251 8.855
R776 VDD.n251 VDD.n250 8.855
R777 VDD.n257 VDD.n256 8.855
R778 VDD.n256 VDD.n255 8.855
R779 VDD.n261 VDD.n260 8.855
R780 VDD.n260 VDD.n259 8.855
R781 VDD.n287 VDD.n286 8.855
R782 VDD.n286 VDD.n285 8.855
R783 VDD.n292 VDD.n291 8.855
R784 VDD.n291 VDD.n290 8.855
R785 VDD.n296 VDD.n295 8.855
R786 VDD.n295 VDD.n294 8.855
R787 VDD.n301 VDD.n300 8.855
R788 VDD.n300  |�� 8.855
R789 VDD.n305 VDD.n304 8.855
R790 VDD.n304 VDD.n303 8.855
R791 VDD.n309 VDD.n308 8.855
R792 VDD.n308 VDD.n307 8.855
R793 VDD.n314 VDD.n313 8.855
R794 VDD.n313 VDD.n312 8.855
R795 VDD.n318 VDD.n317 8.855
R796 VDD.n317 VDD.n316 8.855
R797 VDD.n344 VDD.n343 8.855
R798 VDD.n343 VDD.n342 8.855
R799 VDD.n349 VDD.n348 8.855
R800 VDD.n348 VDD.n347 8.855
R801 VDD.n353 VDD.n352 8.855
R802 VDD.n352 VDD.n351 8.855
R803 VDD.n358 VDD.n357 8.855
R804 VDD.n357 �{�� 8.855
R805 VDD.n362 VDD.n361 8.855
R806 VDD.n361 VDD.n360 8.855
R807 VDD.n366 VDD.n365 8.855
R808 VDD.n365 VDD.n364 8.855
R809 VDD.n371 VDD.n370 8.855
R810 VDD.n370 VDD.n369 8.855
R811 VDD.n375 VDD.n374 8.855
R812 VDD.n374 VDD.n373 8.855
R813 VDD.n401 VDD.n400 8.855
R814 VDD.n400 VDD.n399 8.855
R815 VDD.n406 VDD.n405 8.855
R816 VDD.n405 VDD.n404 8.855
R817 VDD.n410 VDD.n409 8.855
R818 VDD.n409 VDD.n408 8.855
R819 VDD.n415 VDD.n414 8.855
R820 VDD.n414 0|�� 8.855
R821 VDD.n419 VDD.n418 8.855
R822 VDD.n418 VDD.n417 8.855
R823 VDD.n423 VDD.n422 8.855
R824 VDD.n422 VDD.n421 8.855
R825 VDD.n428 VDD.n427 8.855
R826 VDD.n427 VDD.n426 8.855
R827 VDD.n432 VDD.n431 8.855
R828 VDD.n431 VDD.n430 8.855
R829 VDD.n458 VDD.n457 8.855
R830 VDD.n457 VDD.n456 8.855
R831 VDD.n463 VDD.n462 8.855
R832 VDD.n462 VDD.n461 8.855
R833 VDD.n467 VDD.n466 8.855
R834 VDD.n466 VDD.n465 8.855
R835 VDD.n472 VDD.n471 8.855
R836 VDD.n471 �{�� 8.855
R837 VDD.n476 VDD.n475 8.855
R838 VDD.n475 VDD.n474 8.855
R839 VDD.n480 VDD.n479 8.855
R840 VDD.n479 VDD.n478 8.855
R841 VDD.n485 VDD.n484 8.855
R842 VDD.n484 VDD.n483 8.855
R843 VDD.n489 VDD.n488 8.855
R844 VDD.n488 VDD.n487 8.855
R845 VDD.n515 VDD.n514 8.855
R846 VDD.n514 VDD.n513 8.855
R847 VDD.n519 VDD.n518 8.855
R848 VDD.n518 VDD.n517 8.855
R849 VDD.n523 VDD.n522 8.855
R850 VDD.n522 VDD.n521 8.855
R851 VDD.n527 VDD.n526 8.855
R852 VDD.n526 VDD.n525 8.855
R853 VDD.n533 VDD.n530 8.855
R854 VDD.n530 VDD.n529 8.855
R855 VDD.n537 VDD.n536 8.855
R856 VDD.n536 VDD.n535 8.855
R857 VDD.n541 VDD.n540 8.855
R858 VDD.n540 VDD.n539 8.855
R859 VDD.n547 VDD.n546 8.855
R860 VDD.n546 VDD.n545 8.855
R861 VDD.n551 VDD.n550 8.855
R862 VDD.n550 VDD.n549 8.855
R863 VDD.n556 VDD.n555 8.855
R864 VDD.n555 VDD.n554 8.855
R865 VDD.n560 VDD.n559 8.855
R866 VDD.n559 VDD.n558 8.855
R867 VDD.n564 VDD.n563 8.855
R868 VDD.n563 VDD.n562 8.855
R869 VDD.n590 VDD.n589 8.855
R870 VDD.n589 VDD.n588 8.855
R871 VDD.n595 VDD.n594 8.855
R872 VDD.n594 VDD.n593 8.855
R873 VDD.n599 VDD.n598 8.855
R874 VDD.n598 VDD.n597 8.855
R875 VDD.n604 VDD.n603 8.855
R876 VDD.n603  |�� 8.855
R877 VDD.n608 VDD.n607 8.855
R878 VDD.n607 VDD.n606 8.855
R879 VDD.n612 VDD.n611 8.855
R880 VDD.n611 VDD.n610 8.855
R881 VDD.n617 VDD.n616 8.855
R882 VDD.n616 VDD.n615 8.855
R883 VDD.n621 VDD.n620 8.855
R884 VDD.n620 VDD.n619 8.855
R885 VDD.n647 VDD.n646 8.855
R886 VDD.n646 VDD.n645 8.855
R887 VDD.n652 VDD.n651 8.855
R888 VDD.n651 VDD.n650 8.855
R889 VDD.n656 VDD.n655 8.855
R890 VDD.n655 VDD.n654 8.855
R891 VDD.n1304 VDD.n1303 8.855
R892 VDD.n1303 0|�� 8.855
R893 VDD.n1299 VDD.n1298 8.855
R894 VDD.n1298 VDD.n1297 8.855
R895 VDD.n1295 VDD.n1294 8.855
R896 VDD.n1294 VDD.n1293 8.855
R897 VDD.n1291 VDD.n1290 8.855
R898 VDD.n1290 VDD.n1289 8.855
R899 VDD.n1286 VDD.n1285 8.855
R900 VDD.n1285 VDD.n1284 8.855
R901 VDD.n1260 VDD.n1259 8.855
R902 VDD.n1259 VDD.n1258 8.855
R903 VDD.n1256 VDD.n1255 8.855
R904 VDD.n1255 VDD.n1254 8.855
R905 VDD.n1251 VDD.n1250 8.855
R906 VDD.n1250 VDD.n1249 8.855
R907 VDD.n1247 VDD.n1246 8.855
R908 VDD.n1246 �{�� 8.855
R909 VDD.n1242 VDD.n1241 8.855
R910 VDD.n1241 VDD.n1240 8.855
R911 VDD.n1238 VDD.n1237 8.855
R912 VDD.n1237 VDD.n1236 8.855
R913 VDD.n1234 VDD.n1233 8.855
R914 VDD.n1233 VDD.n1232 8.855
R915 VDD.n1229 VDD.n1228 8.855
R916 VDD.n1228 VDD.n1227 8.855
R917 VDD.n1203 VDD.n1202 8.855
R918 VDD.n1202 VDD.n1201 8.855
R919 VDD.n1199 VDD.n1198 8.855
R920 VDD.n1198 VDD.n1197 8.855
R921 VDD.n1194 VDD.n1193 8.855
R922 VDD.n1193 VDD.n1192 8.855
R923 VDD.n1190 VDD.n1189 8.855
R924 VDD.n1189 �{�� 8.855
R925 VDD.n1185 VDD.n1184 8.855
R926 VDD.n1184 VDD.n1183 8.855
R927 VDD.n1181 VDD.n1180 8.855
R928 VDD.n1180 VDD.n1179 8.855
R929 VDD.n1177 VDD.n1176 8.855
R930 VDD.n1176 VDD.n1175 8.855
R931 VDD.n1172 VDD.n1171 8.855
R932 VDD.n1171 VDD.n1170 8.855
R933 VDD.n1146 VDD.n1145 8.855
R934 VDD.n1145 VDD.n1144 8.855
R935 VDD.n1142 VDD.n1141 8.855
R936 VDD.n1141 VDD.n1140 8.855
R937 VDD.n1137 VDD.n1136 8.855
R938 VDD.n1136 VDD.n1135 8.855
R939 VDD.n1133 VDD.n1132 8.855
R940 VDD.n1132  |�� 8.855
R941 VDD.n1128 VDD.n1127 8.855
R942 VDD.n1127 VDD.n1126 8.855
R943 VDD.n1124 VDD.n1123 8.855
R944 VDD.n1123 VDD.n1122 8.855
R945 VDD.n1120 VDD.n1119 8.855
R946 VDD.n1119 VDD.n1118 8.855
R947 VDD.n1115 VDD.n1114 8.855
R948 VDD.n1114 VDD.n1113 8.855
R949 VDD.n1089 VDD.n1088 8.855
R950 VDD.n1088 VDD.n1087 8.855
R951 VDD.n1085 VDD.n1084 8.855
R952 VDD.n1084 VDD.n1083 8.855
R953 VDD.n1081 VDD.n1080 8.855
R954 VDD.n1080 VDD.n1079 8.855
R955 VDD.n1077 VDD.n1076 8.855
R956 VDD.n1076 VDD.n1075 8.855
R957 VDD.n1073 VDD.n1070 8.855
R958 VDD.n1070 VDD.n1069 8.855
R959 VDD.n1067 VDD.n1066 8.855
R960 VDD.n1066 VDD.n1065 8.855
R961 VDD.n1063 VDD.n1062 8.855
R962 VDD.n1062 VDD.n1061 8.855
R963 VDD.n1059 VDD.n1058 8.855
R964 VDD.n1058 VDD.n1057 8.855
R965 VDD.n1053 VDD.n1052 8.855
R966 VDD.n1052 VDD.n1051 8.855
R967 VDD.n1049 VDD.n1048 8.855
R968 VDD.n1048 VDD.n1047 8.855
R969 VDD.n1044 VDD.n1043 8.855
R970 VDD.n1043 VDD.n1042 8.855
R971 VDD.n1040 VDD.n1039 8.855
R972 VDD.n1039 VDD.n1038 8.855
R973 VDD.n1014 VDD.n1013 8.855
R974 VDD.n1013 VDD.n1012 8.855
R975 VDD.n1010 VDD.n1009 8.855
R976 VDD.n1009 VDD.n1008 8.855
R977 VDD.n1005 VDD.n1004 8.855
R978 VDD.n1004 VDD.n1003 8.855
R979 VDD.n1001 VDD.n1000 8.855
R980 VDD.n1000 �{�� 8.855
R981 VDD.n996 VDD.n995 8.855
R982 VDD.n995 VDD.n994 8.855
R983 VDD.n992 VDD.n991 8.855
R984 VDD.n991 VDD.n990 8.855
R985 VDD.n988 VDD.n987 8.855
R986 VDD.n987 VDD.n986 8.855
R987 VDD.n983 VDD.n982 8.855
R988 VDD.n982 VDD.n981 8.855
R989 VDD.n957 VDD.n956 8.855
R990 VDD.n956 VDD.n955 8.855
R991 VDD.n953 VDD.n952 8.855
R992 VDD.n952 VDD.n951 8.855
R993 VDD.n948 VDD.n947 8.855
R994 VDD.n947 VDD.n946 8.855
R995 VDD.n944 VDD.n943 8.855
R996 VDD.n943  |�� 8.855
R997 VDD.n939 VDD.n938 8.855
R998 VDD.n938 VDD.n937 8.855
R999 VDD.n935 VDD.n934 8.855
R1000 VDD.n934 VDD.n933 8.855
R1001 VDD.n931 VDD.n930 8.855
R1002 VDD.n930 VDD.n929 8.855
R1003 VDD.n926 VDD.n925 8.855
R1004 VDD.n925 VDD.n924 8.855
R1005 VDD.n900 VDD.n899 8.855
R1006 VDD.n899 VDD.n898 8.855
R1007 VDD.n896 VDD.n895 8.855
R1008 VDD.n895 VDD.n894 8.855
R1009 VDD.n891 VDD.n890 8.855
R1010 VDD.n890 VDD.n889 8.855
R1011 VDD.n887 VDD.n886 8.855
R1012 VDD.n886 �{�� 8.855
R1013 VDD.n882 VDD.n881 8.855
R1014 VDD.n881 VDD.n880 8.855
R1015 VDD.n878 VDD.n877 8.855
R1016 VDD.n877 VDD.n876 8.855
R1017 VDD.n874 VDD.n873 8.855
R1018 VDD.n873 VDD.n872 8.855
R1019 VDD.n869 VDD.n868 8.855
R1020 VDD.n868 VDD.n867 8.855
R1021 VDD.n843 VDD.n842 8.855
R1022 VDD.n842 VDD.n841 8.855
R1023 VDD.n839 VDD.n838 8.855
R1024 VDD.n838 VDD.n837 8.855
R1025 VDD.n834 VDD.n833 8.855
R1026 VDD.n833 VDD.n832 8.855
R1027 VDD.n830 VDD.n829 8.855
R1028 VDD.n829  |�� 8.855
R1029 VDD.n825 VDD.n824 8.855
R1030 VDD.n824 VDD.n823 8.855
R1031 VDD.n821 VDD.n820 8.855
R1032 VDD.n820 VDD.n819 8.855
R1033 VDD.n817 VDD.n816 8.855
R1034 VDD.n816 VDD.n815 8.855
R1035 VDD.n812 VDD.n811 8.855
R1036 VDD.n811 VDD.n810 8.855
R1037 VDD.n786 VDD.n785 8.855
R1038 VDD.n785 VDD.n784 8.855
R1039 VDD.n782 VDD.n781 8.855
R1040 VDD.n781 VDD.n780 8.855
R1041 VDD.n777 VDD.n776 8.855
R1042 VDD.n776 VDD.n775 8.855
R1043 VDD.n773 VDD.n772 8.855
R1044 VDD.n772 �{�� 8.855
R1045 VDD.n768 VDD.n767 8.855
R1046 VDD.n767 VDD.n766 8.855
R1047 VDD.n764 VDD.n763 8.855
R1048 VDD.n763 VDD.n762 8.855
R1049 VDD.n760 VDD.n759 8.855
R1050 VDD.n759 VDD.n758 8.855
R1051 VDD.n755 VDD.n754 8.855
R1052 VDD.n754 VDD.n753 8.855
R1053 VDD.n728 VDD.n727 8.855
R1054 VDD.n727 VDD.n726 8.855
R1055 VDD.n724 VDD.n723 8.855
R1056 VDD.n723 VDD.n722 8.855
R1057 VDD.n720 VDD.n719 8.855
R1058 VDD.n719 VDD.n718 8.855
R1059 VDD.n716 VDD.n715 8.855
R1060 VDD.n715 VDD.n714 8.855
R1061 VDD.n712 VDD.n709 8.855
R1062 VDD.n709 VDD.n708 8.855
R1063 VDD.n706 VDD.n705 8.855
R1064 VDD.n705 VDD.n704 8.855
R1065 VDD.n702 VDD.n701 8.855
R1066 VDD.n701 VDD.n700 8.855
R1067 VDD.n698 VDD.n697 8.855
R1068 VDD.n697 VDD.n696 8.855
R1069 VDD.n692 VDD.n691 8.855
R1070 VDD.n691 VDD.n690 8.855
R1071 VDD.n688 VDD.n687 8.855
R1072 VDD.n687 VDD.n686 8.855
R1073 VDD.n683 VDD.n682 8.855
R1074 VDD.n682 VDD.n681 8.855
R1075 VDD.n679 VDD.n678 8.855
R1076 VDD.n678 VDD.n677 8.855
R1077 VDD.n803 VDD.n802 8.051
R1078 VDD.n860 VDD.n859 8.051
R1079 VDD.n917 VDD.n916 8.051
R1080 VDD.n974 VDD.n973 8.051
R1081 VDD.n1031 VDD.n1030 8.051
R1082 VDD.n1106 VDD.n1105 8.051
R1083 VDD.n1163 VDD.n1162 8.051
R1084 VDD.n1220 VDD.n1219 8.051
R1085 VDD.n1277 VDD.n1276 8.051
R1086 VDD.n638 VDD.n637 8.051
R1087 VDD.n581 VDD.n580 8.051
R1088 VDD.n506 VDD.n505 8.051
R1089 VDD.n449 VDD.n448 8.051
R1090 VDD.n392 VDD.n391 8.051
R1091 VDD.n335 VDD.n334 8.051
R1092 VDD.n278 VDD.n277 8.051
R1093 VDD.n221 VDD.n220 8.051
R1094 VDD.n164 VDD.n163 8.051
R1095 VDD.n111 VDD.n110 8.051
R1096 VDD.n54 VDD.n53 8.051
R1097 VDD.n742 VDD.n741 8.051
R1098 VDD.n539 0|�� 7.671
R1099 VDD.n1061 0|�� 7.671
R1100 VDD.n700  |�� 7.671
R1101 VDD.n547 VDD.n544 7.019
R1102 VDD.n1059 VDD.n1056 7.019
R1103 VDD.n698 VDD.n695 7.019
R1104 VDD.n533 VDD.n532 6.606
R1105 VDD.n1073 VDD.n1072 6.606
R1106 VDD.n712 VDD.n711 6.606
R1107 VDD.n535 �{�� 5.114
R1108 VDD.n1065  |�� 5.114
R1109 VDD.n704  |�� 5.114
R1110 VDD.n28 VDD.n23 4.795
R1111 VDD.n28 VDD.n27 4.65
R1112 VDD.n32 VDD.n31 4.65
R1113 VDD.n37 VDD.n36 4.65
R1114 VDD.n41 VDD.n40 4.65
R1115 VDD.n68 VDD.n67 4.65
R1116 VDD.n72 VDD.n71 4.65
R1117 VDD.n76 VDD.n75 4.65
R1118 VDD.n79 VDD.n78 4.65
R1119 VDD.n83 VDD.n82 4.65
R1120 VDD.n87 VDD.n86 4.65
R1121 VDD.n91 VDD.n90 4.65
R1122 VDD.n95 VDD.n94 4.65
R1123 VDD.n121 VDD.n120 4.65
R1124 VDD.n125 VDD.n124 4.65
R1125 VDD.n129 VDD.n128 4.65
R1126 VDD.n133 VDD.n132 4.65
R1127 VDD.n136 VDD.n135 4.65
R1128 VDD.n140 VDD.n139 4.65
R1129 VDD.n144 VDD.n143 4.65
R1130 VDD.n148 VDD.n147 4.65
R1131 VDD.n174 VDD.n173 4.65
R1132 VDD.n179 VDD.n178 4.65
R1133 VDD.n183 VDD.n182 4.65
R1134 VDD.n188 VDD.n187 4.65
R1135 VDD.n192 VDD.n191 4.65
R1136 VDD.n196 VDD.n195 4.65
R1137 VDD.n201 VDD.n200 4.65
R1138 VDD.n205 VDD.n204 4.65
R1139 VDD.n231 VDD.n230 4.65
R1140 VDD.n236 VDD.n235 4.65
R1141 VDD.n240 VDD.n239 4.65
R1142 VDD.n245 VDD.n244 4.65
R1143 VDD.n249 VDD.n248 4.65
R1144 VDD.n253 VDD.n252 4.65
R1145 VDD.n258 VDD.n257 4.65
R1146 VDD.n262 VDD.n261 4.65
R1147 VDD.n288 VDD.n287 4.65
R1148 VDD.n293 VDD.n292 4.65
R1149 VDD.n297 VDD.n296 4.65
R1150 VDD.n302 VDD.n301 4.65
R1151 VDD.n306 VDD.n305 4.65
R1152 VDD.n310 VDD.n309 4.65
R1153 VDD.n315 VDD.n314 4.65
R1154 VDD.n319 VDD.n318 4.65
R1155 VDD.n345 VDD.n344 4.65
R1156 VDD.n350 VDD.n349 4.65
R1157 VDD.n354 VDD.n353 4.65
R1158 VDD.n359 VDD.n358 4.65
R1159 VDD.n363 VDD.n362 4.65
R1160 VDD.n367 VDD.n366 4.65
R1161 VDD.n372 VDD.n371 4.65
R1162 VDD.n376 VDD.n375 4.65
R1163 VDD.n402 VDD.n401 4.65
R1164 VDD.n407 VDD.n406 4.65
R1165 VDD.n411 VDD.n410 4.65
R1166 VDD.n416 VDD.n415 4.65
R1167 VDD.n420 VDD.n419 4.65
R1168 VDD.n424 VDD.n423 4.65
R1169 VDD.n429 VDD.n428 4.65
R1170 VDD.n433 VDD.n432 4.65
R1171 VDD.n459 VDD.n458 4.65
R1172 VDD.n464 VDD.n463 4.65
R1173 VDD.n468 VDD.n467 4.65
R1174 VDD.n473 VDD.n472 4.65
R1175 VDD.n477 VDD.n476 4.65
R1176 VDD.n481 VDD.n480 4.65
R1177 VDD.n486 VDD.n485 4.65
R1178 VDD.n490 VDD.n489 4.65
R1179 VDD.n516 VDD.n515 4.65
R1180 VDD.n520 VDD.n519 4.65
R1181 VDD.n524 VDD.n523 4.65
R1182 VDD.n528 VDD.n527 4.65
R1183 VDD.n534 VDD.n533 4.65
R1184 VDD.n538 VDD.n537 4.65
R1185 VDD.n542 VDD.n541 4.65
R1186 VDD.n548 VDD.n547 4.65
R1187 VDD.n552 VDD.n551 4.65
R1188 VDD.n557 VDD.n556 4.65
R1189 VDD.n561 VDD.n560 4.65
R1190 VDD.n565 VDD.n564 4.65
R1191 VDD.n591 VDD.n590 4.65
R1192 VDD.n596 VDD.n595 4.65
R1193 VDD.n600 VDD.n599 4.65
R1194 VDD.n605 VDD.n604 4.65
R1195 VDD.n609 VDD.n608 4.65
R1196 VDD.n613 VDD.n612 4.65
R1197 VDD.n618 VDD.n617 4.65
R1198 VDD.n622 VDD.n621 4.65
R1199 VDD.n648 VDD.n647 4.65
R1200 VDD.n653 VDD.n652 4.65
R1201 VDD.n657 VDD.n656 4.65
R1202 VDD.n1305 VDD.n1304 4.65
R1203 VDD.n1300 VDD.n1299 4.65
R1204 VDD.n1296 VDD.n1295 4.65
R1205 VDD.n1292 VDD.n1291 4.65
R1206 VDD.n1287 VDD.n1286 4.65
R1207 VDD.n1261 VDD.n1260 4.65
R1208 VDD.n1257 VDD.n1256 4.65
R1209 VDD.n1252 VDD.n1251 4.65
R1210 VDD.n1248 VDD.n1247 4.65
R1211 VDD.n1243 VDD.n1242 4.65
R1212 VDD.n1239 VDD.n1238 4.65
R1213 VDD.n1235 VDD.n1234 4.65
R1214 VDD.n1230 VDD.n1229 4.65
R1215 VDD.n1204 VDD.n1203 4.65
R1216 VDD.n1200 VDD.n1199 4.65
R1217 VDD.n1195 VDD.n1194 4.65
R1218 VDD.n1191 VDD.n1190 4.65
R1219 VDD.n1186 VDD.n1185 4.65
R1220 VDD.n1182 VDD.n1181 4.65
R1221 VDD.n1178 VDD.n1177 4.65
R1222 VDD.n1173 VDD.n1172 4.65
R1223 VDD.n1147 VDD.n1146 4.65
R1224 VDD.n1143 VDD.n1142 4.65
R1225 VDD.n1138 VDD.n1137 4.65
R1226 VDD.n1134 VDD.n1133 4.65
R1227 VDD.n1129 VDD.n1128 4.65
R1228 VDD.n1125 VDD.n1124 4.65
R1229 VDD.n1121 VDD.n1120 4.65
R1230 VDD.n1116 VDD.n1115 4.65
R1231 VDD.n1090 VDD.n1089 4.65
R1232 VDD.n1086 VDD.n1085 4.65
R1233 VDD.n1082 VDD.n1081 4.65
R1234 VDD.n1078 VDD.n1077 4.65
R1235 VDD.n1074 VDD.n1073 4.65
R1236 VDD.n1068 VDD.n1067 4.65
R1237 VDD.n1064 VDD.n1063 4.65
R1238 VDD.n1060 VDD.n1059 4.65
R1239 VDD.n1054 VDD.n1053 4.65
R1240 VDD.n1050 VDD.n1049 4.65
R1241 VDD.n1045 VDD.n1044 4.65
R1242 VDD.n1041 VDD.n1040 4.65
R1243 VDD.n1015 VDD.n1014 4.65
R1244 VDD.n1011 VDD.n1010 4.65
R1245 VDD.n1006 VDD.n1005 4.65
R1246 VDD.n1002 VDD.n1001 4.65
R1247 VDD.n997 VDD.n996 4.65
R1248 VDD.n993 VDD.n992 4.65
R1249 VDD.n989 VDD.n988 4.65
R1250 VDD.n984 VDD.n983 4.65
R1251 VDD.n958 VDD.n957 4.65
R1252 VDD.n954 VDD.n953 4.65
R1253 VDD.n949 VDD.n948 4.65
R1254 VDD.n945 VDD.n944 4.65
R1255 VDD.n940 VDD.n939 4.65
R1256 VDD.n936 VDD.n935 4.65
R1257 VDD.n932 VDD.n931 4.65
R1258 VDD.n927 VDD.n926 4.65
R1259 VDD.n901 VDD.n900 4.65
R1260 VDD.n897 VDD.n896 4.65
R1261 VDD.n892 VDD.n891 4.65
R1262 VDD.n888 VDD.n887 4.65
R1263 VDD.n883 VDD.n882 4.65
R1264 VDD.n879 VDD.n878 4.65
R1265 VDD.n875 VDD.n874 4.65
R1266 VDD.n870 VDD.n869 4.65
R1267 VDD.n844 VDD.n843 4.65
R1268 VDD.n840 VDD.n839 4.65
R1269 VDD.n835 VDD.n834 4.65
R1270 VDD.n831 VDD.n830 4.65
R1271 VDD.n826 VDD.n825 4.65
R1272 VDD.n822 VDD.n821 4.65
R1273 VDD.n818 VDD.n817 4.65
R1274 VDD.n813 VDD.n812 4.65
R1275 VDD.n787 VDD.n786 4.65
R1276 VDD.n783 VDD.n782 4.65
R1277 VDD.n778 VDD.n777 4.65
R1278 VDD.n774 VDD.n773 4.65
R1279 VDD.n769 VDD.n768 4.65
R1280 VDD.n765 VDD.n764 4.65
R1281 VDD.n761 VDD.n760 4.65
R1282 VDD.n756 VDD.n755 4.65
R1283 VDD.n729 VDD.n728 4.65
R1284 VDD.n725 VDD.n724 4.65
R1285 VDD.n721 VDD.n720 4.65
R1286 VDD.n717 VDD.n716 4.65
R1287 VDD.n713 VDD.n712 4.65
R1288 VDD.n707 VDD.n706 4.65
R1289 VDD.n703 VDD.n702 4.65
R1290 VDD.n699 VDD.n698 4.65
R1291 VDD.n693 VDD.n692 4.65
R1292 VDD.n689 VDD.n688 4.65
R1293 VDD.n684 VDD.n683 4.65
R1294 VDD.n680 VDD.n679 4.65
R1295 VDD.n200 VDD.n197 2.89
R1296 VDD.n257 VDD.n254 2.89
R1297 VDD.n314 VDD.n311 2.89
R1298 VDD.n371 VDD.n368 2.89
R1299 VDD.n428 VDD.n425 2.89
R1300 VDD.n485 VDD.n482 2.89
R1301 VDD.n617 VDD.n614 2.89
R1302 VDD.n1291 VDD.n1288 2.89
R1303 VDD.n1234 VDD.n1231 2.89
R1304 VDD.n1177 VDD.n1174 2.89
R1305 VDD.n1120 VDD.n1117 2.89
R1306 VDD.n988 VDD.n985 2.89
R1307 VDD.n931 VDD.n928 2.89
R1308 VDD.n874 VDD.n871 2.89
R1309 VDD.n817 VDD.n814 2.89
R1310 VDD.n760 VDD.n757 2.89
R1311 VDD.n80 �{�� 2.557
R1312 VDD.n130 �{�� 2.557
R1313 VDD.n189 �{�� 2.557
R1314 VDD.n246  |�� 2.557
R1315 VDD.n303  |�� 2.557
R1316 VDD.n360  |�� 2.557
R1317 VDD.n417  |�� 2.557
R1318 VDD.n474 0|�� 2.557
R1319 VDD.n606 |�� 2.557
R1320 VDD.n1297  |�� 2.557
R1321 VDD.n1240 0|�� 2.557
R1322 VDD.n1183 �{�� 2.557
R1323 VDD.n1126 0|�� 2.557
R1324 VDD.n994 �{�� 2.557
R1325 VDD.n937  |�� 2.557
R1326 VDD.n880 ���*V 2.557
R1327 VDD.n823 �{�� 2.557
R1328 VDD.n766  |�� 2.557
R1329 VDD.n178 VDD.n175 2.477
R1330 VDD.n235 VDD.n232 2.477
R1331 VDD.n292 VDD.n289 2.477
R1332 VDD.n349 VDD.n346 2.477
R1333 VDD.n406 VDD.n403 2.477
R1334 VDD.n463 VDD.n460 2.477
R1335 VDD.n595 VDD.n592 2.477
R1336 VDD.n652 VDD.n649 2.477
R1337 VDD.n1256 VDD.n1253 2.477
R1338 VDD.n1199 VDD.n1196 2.477
R1339 VDD.n1142 VDD.n1139 2.477
R1340 VDD.n1010 VDD.n1007 2.477
R1341 VDD.n953 VDD.n950 2.477
R1342 VDD.n896 VDD.n893 2.477
R1343 VDD.n839 VDD.n836 2.477
R1344 VDD.n782 VDD.n779 2.477
R1345 VDD.n27 VDD.n24 2.064
R1346 VDD.n36 VDD.n35 2.064
R1347 VDD.n556 VDD.n553 0.412
R1348 VDD.n1049 VDD.n1046 0.412
R1349 VDD.n688 VDD.n685 0.412
R1350 VDD.n68 VDD.n41 0.29
R1351 VDD.n121 VDD.n95 0.29
R1352 VDD.n174 VDD.n148 0.29
R1353 VDD.n231 VDD.n205 0.29
R1354 VDD.n288 VDD.n262 0.29
R1355 VDD.n345 VDD.n319 0.29
R1356 VDD.n402 VDD.n376 0.29
R1357 VDD.n459 VDD.n433 0.29
R1358 VDD.n516 VDD.n490 0.29
R1359 VDD.n591 VDD.n565 0.29
R1360 VDD.n648 VDD.n622 0.29
R1361 VDD.n1287 VDD.n1261 0.29
R1362 VDD.n1230 VDD.n1204 0.29
R1363 VDD.n1173 VDD.n1147 0.29
R1364 VDD.n1116 VDD.n1090 0.29
R1365 VDD.n1041 VDD.n1015 0.29
R1366 VDD.n984 VDD.n958 0.29
R1367 VDD.n927 VDD.n901 0.29
R1368 VDD.n870 VDD.n844 0.29
R1369 VDD.n813 VDD.n787 0.29
R1370 VDD.n756 VDD.n729 0.29
R1371 VDD.n680 VDD 0.207
R1372 VDD.n542 VDD.n538 0.197
R1373 VDD.n1068 VDD.n1064 0.197
R1374 VDD.n707 VDD.n703 0.197
R1375 VDD.n83 VDD.n79 0.181
R1376 VDD.n136 VDD.n133 0.181
R1377 VDD.n192 VDD.n188 0.181
R1378 VDD.n249 VDD.n245 0.181
R1379 VDD.n306 VDD.n302 0.181
R1380 VDD.n363 VDD.n359 0.181
R1381 VDD.n420 VDD.n416 0.181
R1382 VDD.n477 VDD.n473 0.181
R1383 VDD.n609 VDD.n605 0.181
R1384 VDD.n1305 VDD.n1300 0.181
R1385 VDD.n1248 VDD.n1243 0.181
R1386 VDD.n1191 VDD.n1186 0.181
R1387 VDD.n1134 VDD.n1129 0.181
R1388 VDD.n1002 VDD.n997 0.181
R1389 VDD.n945 VDD.n940 0.181
R1390 VDD.n888 VDD.n883 0.181
R1391 VDD.n831 VDD.n826 0.181
R1392 VDD.n774 VDD.n769 0.181
R1393 VDD.n32 VDD.n28 0.157
R1394 VDD.n37 VDD.n32 0.157
R1395 VDD.n41 VDD.n37 0.145
R1396 VDD.n72 VDD.n68 0.145
R1397 VDD.n76 VDD.n72 0.145
R1398 VDD.n79 VDD.n76 0.145
R1399 VDD.n87 VDD.n83 0.145
R1400 VDD.n91 VDD.n87 0.145
R1401 VDD.n95 VDD.n91 0.145
R1402 VDD.n125 VDD.n121 0.145
R1403 VDD.n129 VDD.n125 0.145
R1404 VDD.n133 VDD.n129 0.145
R1405 VDD.n140 VDD.n136 0.145
R1406 VDD.n144 VDD.n140 0.145
R1407 VDD.n148 VDD.n144 0.145
R1408 VDD.n179 VDD.n174 0.145
R1409 VDD.n183 VDD.n179 0.145
R1410 VDD.n188 VDD.n183 0.145
R1411 VDD.n196 VDD.n192 0.145
R1412 VDD.n201 VDD.n196 0.145
R1413 VDD.n205 VDD.n201 0.145
R1414 VDD.n236 VDD.n231 0.145
R1415 VDD.n240 VDD.n236 0.145
R1416 VDD.n245 VDD.n240 0.145
R1417 VDD.n253 VDD.n249 0.145
R1418 VDD.n258 VDD.n253 0.145
R1419 VDD.n262 VDD.n258 0.145
R1420 VDD.n293 VDD.n288 0.145
R1421 VDD.n297 VDD.n293 0.145
R1422 VDD.n302 VDD.n297 0.145
R1423 VDD.n310 VDD.n306 0.145
R1424 VDD.n315 VDD.n310 0.145
R1425 VDD.n319 VDD.n315 0.145
R1426 VDD.n350 VDD.n345 0.145
R1427 VDD.n354 VDD.n350 0.145
R1428 VDD.n359 VDD.n354 0.145
R1429 VDD.n367 VDD.n363 0.145
R1430 VDD.n372 VDD.n367 0.145
R1431 VDD.n376 VDD.n372 0.145
R1432 VDD.n407 VDD.n402 0.145
R1433 VDD.n411 VDD.n407 0.145
R1434 VDD.n416 VDD.n411 0.145
R1435 VDD.n424 VDD.n420 0.145
R1436 VDD.n429 VDD.n424 0.145
R1437 VDD.n433 VDD.n429 0.145
R1438 VDD.n464 VDD.n459 0.145
R1439 VDD.n468 VDD.n464 0.145
R1440 VDD.n473 VDD.n468 0.145
R1441 VDD.n481 VDD.n477 0.145
R1442 VDD.n486 VDD.n481 0.145
R1443 VDD.n490 VDD.n486 0.145
R1444 VDD.n520 VDD.n516 0.145
R1445 VDD.n524 VDD.n520 0.145
R1446 VDD.n528 VDD.n524 0.145
R1447 VDD.n534 VDD.n528 0.145
R1448 VDD.n538 VDD.n534 0.145
R1449 VDD.n548 VDD.n542 0.145
R1450 VDD.n552 VDD.n548 0.145
R1451 VDD.n557 VDD.n552 0.145
R1452 VDD.n561 VDD.n557 0.145
R1453 VDD.n565 VDD.n561 0.145
R1454 VDD.n596 VDD.n591 0.145
R1455 VDD.n600 VDD.n596 0.145
R1456 VDD.n605 VDD.n600 0.145
R1457 VDD.n613 VDD.n609 0.145
R1458 VDD.n618 VDD.n613 0.145
R1459 VDD.n622 VDD.n618 0.145
R1460 VDD.n653 VDD.n648 0.145
R1461 VDD.n657 VDD.n653 0.145
R1462 VDD.n1300 VDD.n1296 0.145
R1463 VDD.n1296 VDD.n1292 0.145
R1464 VDD.n1292 VDD.n1287 0.145
R1465 VDD.n1261 VDD.n1257 0.145
R1466 VDD.n1257 VDD.n1252 0.145
R1467 VDD.n1252 VDD.n1248 0.145
R1468 VDD.n1243 VDD.n1239 0.145
R1469 VDD.n1239 VDD.n1235 0.145
R1470 VDD.n1235 VDD.n1230 0.145
R1471 VDD.n1204 VDD.n1200 0.145
R1472 VDD.n1200 VDD.n1195 0.145
R1473 VDD.n1195 VDD.n1191 0.145
R1474 VDD.n1186 VDD.n1182 0.145
R1475 VDD.n1182 VDD.n1178 0.145
R1476 VDD.n1178 VDD.n1173 0.145
R1477 VDD.n1147 VDD.n1143 0.145
R1478 VDD.n1143 VDD.n1138 0.145
R1479 VDD.n1138 VDD.n1134 0.145
R1480 VDD.n1129 VDD.n1125 0.145
R1481 VDD.n1125 VDD.n1121 0.145
R1482 VDD.n1121 VDD.n1116 0.145
R1483 VDD.n1090 VDD.n1086 0.145
R1484 VDD.n1086 VDD.n1082 0.145
R1485 VDD.n1082 VDD.n1078 0.145
R1486 VDD.n1078 VDD.n1074 0.145
R1487 VDD.n1074 VDD.n1068 0.145
R1488 VDD.n1064 VDD.n1060 0.145
R1489 VDD.n1060 VDD.n1054 0.145
R1490 VDD.n1054 VDD.n1050 0.145
R1491 VDD.n1050 VDD.n1045 0.145
R1492 VDD.n1045 VDD.n1041 0.145
R1493 VDD.n1015 VDD.n1011 0.145
R1494 VDD.n1011 VDD.n1006 0.145
R1495 VDD.n1006 VDD.n1002 0.145
R1496 VDD.n997 VDD.n993 0.145
R1497 VDD.n993 VDD.n989 0.145
R1498 VDD.n989 VDD.n984 0.145
R1499 VDD.n958 VDD.n954 0.145
R1500 VDD.n954 VDD.n949 0.145
R1501 VDD.n949 VDD.n945 0.145
R1502 VDD.n940 VDD.n936 0.145
R1503 VDD.n936 VDD.n932 0.145
R1504 VDD.n932 VDD.n927 0.145
R1505 VDD.n901 VDD.n897 0.145
R1506 VDD.n897 VDD.n892 0.145
R1507 VDD.n892 VDD.n888 0.145
R1508 VDD.n883 VDD.n879 0.145
R1509 VDD.n879 VDD.n875 0.145
R1510 VDD.n875 VDD.n870 0.145
R1511 VDD.n844 VDD.n840 0.145
R1512 VDD.n840 VDD.n835 0.145
R1513 VDD.n835 VDD.n831 0.145
R1514 VDD.n826 VDD.n822 0.145
R1515 VDD.n822 VDD.n818 0.145
R1516 VDD.n818 VDD.n813 0.145
R1517 VDD.n787 VDD.n783 0.145
R1518 VDD.n783 VDD.n778 0.145
R1519 VDD.n778 VDD.n774 0.145
R1520 VDD.n769 VDD.n765 0.145
R1521 VDD.n765 VDD.n761 0.145
R1522 VDD.n761 VDD.n756 0.145
R1523 VDD.n729 VDD.n725 0.145
R1524 VDD.n725 VDD.n721 0.145
R1525 VDD.n721 VDD.n717 0.145
R1526 VDD.n717 VDD.n713 0.145
R1527 VDD.n713 VDD.n707 0.145
R1528 VDD.n703 VDD.n699 0.145
R1529 VDD.n699 VDD.n693 0.145
R1530 VDD.n693 VDD.n689 0.145
R1531 VDD.n689 VDD.n684 0.145
R1532 VDD.n684 VDD.n680 0.145
R1533 VDD VDD.n657 0.086
R1534 VDD VDD.n1305 0.058
R1535 a_277_1050.n7 a_277_1050.t9 480.392
R1536 a_277_1050.n5 a_277_1050.t10 480.392
R1537 a_277_1050.n7 a_277_1050.t11 403.272
R1538 a_277_1050.n5 a_277_1050.t7 403.272
R1539 a_277_1050.n8 a_277_1050.t12 385.063
R1540 a_277_1050.n6 a_277_1050.t8 385.063
R1541 a_277_1050.n12 a_277_1050.n10 342.597
R1542 a_277_1050.n3 a_277_1050.n2 161.352
R1543 a_277_1050.n10 a_277_1050.n4 151.34
R1544 a_277_1050.n8 a_277_1050.n7 143.429
R1545 a_277_1050.n6 a_277_1050.n5 143.429
R1546 a_277_1050.n4 a_277_1050.n0 95.095
R1547 a_277_1050.n3 a_277_1050.n1 95.095
R1548 a_277_1050.n4 a_277_1050.n3 66.258
R1549 a_277_1050.n12 a_277_1050.n11 15.218
R1550 a_277_1050.n0 a_277_1050.t1 14.282
R1551 a_277_1050.n0 a_277_1050.t6 14.282
R1552 a_277_1050.n1 a_277_1050.t4 14.282
R1553 a_277_1050.n1 a_277_1050.t3 14.282
R1554 a_277_1050.n2 a_277_1050.t2 14.282
R1555 a_277_1050.n2 a_277_1050.t0 14.282
R1556 a_277_1050.n13 a_277_1050.n12 12.014
R1557 a_277_1050.n9 a_277_1050.n6 11.95
R1558 a_277_1050.n10 a_277_1050.n9 5.965
R1559 a_277_1050.n9 a_277_1050.n8 4.65
R1560 a_3177_1050.n1 a_3177_1050.t7 480.392
R1561 a_3177_1050.n1 a_3177_1050.t5 403.272
R1562 a_3177_1050.n2 a_3177_1050.t6 385.063
R1563 a_3177_1050.n4 a_3177_1050.n3 355.179
R1564 a_3177_1050.n6 a_3177_1050.n5 157.963
R1565 a_3177_1050.n2 a_3177_1050.n1 143.429
R1566 a_3177_1050.n5 a_3177_1050.n4 132.141
R1567 a_3177_1050.n5 a_3177_1050.n0 91.706
R1568 a_3177_1050.n0 a_3177_1050.t4 14.282
R1569 a_3177_1050.n0 a_3177_1050.t1 14.282
R1570 a_3177_1050.n6 a_3177_1050.t2 14.282
R1571 a_3177_1050.t3 a_3177_1050.n6 14.282
R1572 a_3177_1050.n4 a_3177_1050.n2 10.615
R1573 a_1845_1050.n3 a_1845_1050.t5 480.392
R1574 a_1845_1050.n3 a_1845_1050.t7 403.272
R1575 a_1845_1050.n4 a_1845_1050.t6 357.204
R1576 a_1845_1050.n7 a_1845_1050.n5 312.103
R1577 a_1845_1050.n4 a_1845_1050.n3 171.288
R1578 a_1845_1050.n5 a_1845_1050.n2 159.999
R1579 a_1845_1050.n2 a_1845_1050.n1 157.964
R1580 a_1845_1050.n2 a_1845_1050.n0 91.706
R1581 a_1845_1050.n7 a_1845_1050.n6 15.218
R1582 a_1845_1050.n0 a_1845_1050.t0 14.282
R1583 a_1845_1050.n0 a_1845_1050.t1 14.282
R1584 a_1845_1050.n1 a_1845_1050.t3 14.282
R1585 a_1845_1050.n1 a_1845_1050.t4 14.282
R1586 a_1845_1050.n8 a_1845_1050.n7 12.014
R1587 a_1845_1050.n5 a_1845_1050.n4 10.615
R1588 a_147_187.n5 a_147_187.t13 512.525
R1589 a_147_187.n3 a_147_187.t11 472.359
R1590 a_147_187.n1 a_147_187.t6 472.359
R1591 a_147_187.n6 a_147_187.t10 417.109
R1592 a_147_187.n3 a_147_187.t7 384.527
R1593 a_147_187.n1 a_147_187.t8 384.527
R1594 a_147_187.n10 a_147_187.n9 383.037
R1595 a_147_187.n5 a_147_187.t9 371.139
R1596 a_147_187.n4 a_147_187.t12 370.613
R1597 a_147_187.n2 a_147_187.t5 370.613
R1598 a_147_187.n6 a_147_187.n5 179.837
R1599 a_147_187.n12 a_147_187.n11 157.963
R1600 a_147_187.n4 a_147_187.n3 127.096
R1601 a_147_187.n2 a_147_187.n1 127.096
R1602 a_147_187.n11 a_147_187.n10 104.282
R1603 a_147_187.n11 a_147_187.n0 91.706
R1604 a_147_187.n0 a_147_187.t4 14.282
R1605 a_147_187.n0 a_147_187.t3 14.282
R1606 a_147_187.t1 a_147_187.n12 14.282
R1607 a_147_187.n12 a_147_187.t0 14.282
R1608 a_147_187.n7 a_147_187.n6 11.134
R1609 a_147_187.n8 a_147_187.n2 8.957
R1610 a_147_187.n7 a_147_187.n4 4.65
R1611 a_147_187.n10 a_147_187.n8 4.65
R1612 a_147_187.n8 a_147_187.n7 2.947
R1613 a_3303_411.n1 a_3303_411.t8 512.525
R1614 a_3303_411.n0 a_3303_411.t11 512.525
R1615 a_3303_411.n5 a_3303_411.t13 472.359
R1616 a_3303_411.n5 a_3303_411.t7 384.527
R1617 a_3303_411.n1 a_3303_411.t12 371.139
R1618 a_3303_411.n0 a_3303_411.t9 371.139
R1619 a_3303_411.n2 a_3303_411.n1 343.521
R1620 a_3303_411.n6 a_3303_411.t10 287.037
R1621 a_3303_411.n12 a_3303_411.n11 277.722
R1622 a_3303_411.n4 a_3303_411.n0 259.945
R1623 a_3303_411.n6 a_3303_411.n5 210.673
R1624 a_3303_411.n14 a_3303_411.n12 187.858
R1625 a_3303_411.n2 a_3303_411.t6 172.106
R1626 a_3303_411.n3 a_3303_411.t5 165.68
R1627 a_3303_411.n14 a_3303_411.n13 157.964
R1628 a_3303_411.n15 a_3303_411.n14 91.705
R1629 a_3303_411.n4 a_3303_411.n3 83.576
R1630 a_3303_411.n7 a_3303_411.n4 41.06
R1631 a_3303_411.n11 a_3303_411.n10 30
R1632 a_3303_411.n9 a_3303_411.n8 24.383
R1633 a_3303_411.n11 a_3303_411.n9 23.684
R1634 a_3303_411.n13 a_3303_411.t3 14.282
R1635 a_3303_411.n13 a_3303_411.t4 14.282
R1636 a_3303_411.t1 a_3303_411.n15 14.282
R1637 a_3303_411.n15 a_3303_411.t0 14.282
R1638 a_3303_411.n3 a_3303_411.n2 10.343
R1639 a_3303_411.n7 a_3303_411.n6 7.597
R1640 a_3303_411.n12 a_3303_411.n7 4.65
R1641 a_13654_101.t0 a_13654_101.n0 93.333
R1642 a_13654_101.n3 a_13654_101.n1 79.062
R1643 a_13654_101.n3 a_13654_101.n2 2.084
R1644 a_13654_101.t0 a_13654_101.n3 0.182
R1645 a_13268_209.n3 a_13268_209.t9 512.525
R1646 a_13268_209.n3 a_13268_209.t7 371.139
R1647 a_13268_209.n4 a_13268_209.t8 338.57
R1648 a_13268_209.n13 a_13268_209.n5 227.387
R1649 a_13268_209.n4 a_13268_209.n3 191.629
R1650 a_13268_209.n2 a_13268_209.n1 165.613
R1651 a_13268_209.n5 a_13268_209.n2 132.893
R1652 a_13268_209.n12 a_13268_209.n11 128.294
R1653 a_13268_209.n12 a_13268_209.n8 126.225
R1654 a_13268_209.n15 a_13268_209.n13 112.91
R1655 a_13268_209.n2 a_13268_209.n0 99.355
R1656 a_13268_209.n8 a_13268_209.n7 22.578
R1657 a_13268_209.n11 a_13268_209.n10 22.578
R1658 a_13268_209.n15 a_13268_209.n14 15.001
R1659 a_13268_209.n0 a_13268_209.t5 14.282
R1660 a_13268_209.n0 a_13268_209.t6 14.282
R1661 a_13268_209.n1 a_13268_209.t2 14.282
R1662 a_13268_209.n1 a_13268_209.t3 14.282
R1663 a_13268_209.n16 a_13268_209.n15 12.632
R1664 a_13268_209.n5 a_13268_209.n4 10.343
R1665 a_13268_209.n8 a_13268_209.n6 8.58
R1666 a_13268_209.n11 a_13268_209.n9 8.58
R1667 a_13268_209.n13 a_13268_209.n12 7.053
R1668 GND.n34 GND.n33 237.558
R1669 GND.n67 GND.n66 237.558
R1670 GND.n415 GND.n414 237.558
R1671 GND.n448 GND.n447 237.558
R1672 GND.n480 GND.n479 237.558
R1673 GND.n513 GND.n512 237.558
R1674 GND.n546 GND.n545 237.558
R1675 GND.n579 GND.n578 237.558
R1676 GND.n623 GND.n622 237.558
R1677 GND.n655 GND.n654 237.558
R1678 GND.n687 GND.n686 237.558
R1679 GND.n364 GND.n363 237.558
R1680 GND.n717 GND.n716 237.558
R1681 GND.n334 GND.n333 237.558
R1682 GND.n289 GND.n288 237.558
R1683 GND.n256 GND.n255 237.558
R1684 GND.n226 GND.n225 237.558
R1685 GND.n194 GND.n193 237.558
R1686 GND.n161 GND.n160 237.558
R1687 GND.n129 GND.n128 237.558
R1688 GND.n97 GND.n96 237.558
R1689 GND.n31 GND.n30 210.82
R1690 GND.n64 GND.n63 210.82
R1691 GND.n94 GND.n93 210.82
R1692 GND.n417 GND.n416 210.82
R1693 GND.n450 GND.n449 210.82
R1694 GND.n482 GND.n481 210.82
R1695 GND.n515 GND.n514 210.82
R1696 GND.n548 GND.n547 210.82
R1697 GND.n581 GND.n580 210.82
R1698 GND.n625 GND.n624 210.82
R1699 GND.n657 GND.n656 210.82
R1700 GND.n689 GND.n688 210.82
R1701 GND.n719 GND.n718 210.82
R1702 GND.n361 GND.n360 210.82
R1703 GND.n331 GND.n330 210.82
R1704 GND.n286 GND.n285 210.82
R1705 GND.n253 GND.n252 210.82
R1706 GND.n223 GND.n222 210.82
R1707 GND.n191 GND.n190 210.82
R1708 GND.n158 GND.n157 210.82
R1709 GND.n126 GND.n125 210.82
R1710 GND.n83 GND.n82 172.612
R1711 GND.n242 GND.n241 172.612
R1712 GND.n350 GND.n349 172.612
R1713 GND.n697 GND.n696 172.612
R1714 GND.n592 GND.n591 167.358
R1715 GND.n115 GND.n114 166.605
R1716 GND.n147 GND.n146 166.605
R1717 GND.n212 GND.n211 166.605
R1718 GND.n667 GND.n666 166.605
R1719 GND.n635 GND.n634 166.605
R1720 GND.n460 GND.n459 166.605
R1721 GND.n321 GND.n320 152.358
R1722 GND.n384 GND.n383 152.358
R1723 GND.n180 GND.n179 151.605
R1724 GND.n275 GND.n274 151.605
R1725 GND.n730 GND.n729 151.605
R1726 GND.n559 GND.n558 151.605
R1727 GND.n526 GND.n525 151.605
R1728 GND.n493 GND.n492 151.605
R1729 GND.n428 GND.n427 151.605
R1730 GND.n53 GND.n52 151.605
R1731 GND.n5 GND.n4 120.01
R1732 GND.n3 GND.n2 92.5
R1733 GND.n12 GND.n11 92.5
R1734 GND.n21 GND.t0 45.413
R1735 GND.n21 GND.n20 39.307
R1736 GND.n179 GND.n178 28.421
R1737 GND.n274 GND.n273 28.421
R1738 GND.n320 GND.n319 28.421
R1739 GND.n729 GND.n728 28.421
R1740 GND.n558 GND.n557 28.421
R1741 GND.n525 GND.n524 28.421
R1742 GND.n492 GND.n491 28.421
R1743 GND.n427 GND.n426 28.421
R1744 GND.n383 GND.n382 28.421
R1745 GND.n52 GND.n51 28.421
R1746 GND.n179 GND.n177 25.263
R1747 GND.n274 GND.n272 25.263
R1748 GND.n320 GND.n318 25.263
R1749 GND.n729 GND.n727 25.263
R1750 GND.n558 GND.n556 25.263
R1751 GND.n525 GND.n523 25.263
R1752 GND.n492 GND.n490 25.263
R1753 GND.n427 GND.n425 25.263
R1754 GND.n383 GND.n381 25.263
R1755 GND.n52 GND.n50 25.263
R1756 GND.n177 GND.n176 24.383
R1757 GND.n272 GND.n271 24.383
R1758 GND.n318 GND.n317 24.383
R1759 GND.n727 GND.n726 24.383
R1760 GND.n556 GND.n555 24.383
R1761 GND.n523 GND.n522 24.383
R1762 GND.n490 GND.n489 24.383
R1763 GND.n425 GND.n424 24.383
R1764 GND.n381 GND.n380 24.383
R1765 GND.n50 GND.n49 24.383
R1766 GND.n22 GND.n21 23.77
R1767 GND.n114 GND.n112 23.03
R1768 GND.n146 GND.n144 23.03
R1769 GND.n211 GND.n209 23.03
R1770 GND.n666 GND.n664 23.03
R1771 GND.n634 GND.n632 23.03
R1772 GND.n591 GND.n589 23.03
R1773 GND.n459 GND.n457 23.03
R1774 GND.n6 GND.n5 20.705
R1775 GND.n14 GND.n13 20.705
R1776 GND.n23 GND.n22 20.705
R1777 GND.n5 GND.n3 19.952
R1778 GND.n32 GND.n31 18.953
R1779 GND.n65 GND.n64 18.953
R1780 GND.n95 GND.n94 18.953
R1781 GND.n418 GND.n417 18.953
R1782 GND.n451 GND.n450 18.953
R1783 GND.n483 GND.n482 18.953
R1784 GND.n516 GND.n515 18.953
R1785 GND.n549 GND.n548 18.953
R1786 GND.n582 GND.n581 18.953
R1787 GND.n626 GND.n625 18.953
R1788 GND.n658 GND.n657 18.953
R1789 GND.n690 GND.n689 18.953
R1790 GND.n720 GND.n719 18.953
R1791 GND.n362 GND.n361 18.953
R1792 GND.n332 GND.n331 18.953
R1793 GND.n287 GND.n286 18.953
R1794 GND.n254 GND.n253 18.953
R1795 GND.n224 GND.n223 18.953
R1796 GND.n192 GND.n191 18.953
R1797 GND.n159 GND.n158 18.953
R1798 GND.n127 GND.n126 18.953
R1799 GND.n35 GND.n32 14.864
R1800 GND.n68 GND.n65 14.864
R1801 GND.n98 GND.n95 14.864
R1802 GND.n130 GND.n127 14.864
R1803 GND.n162 GND.n159 14.864
R1804 GND.n195 GND.n192 14.864
R1805 GND.n227 GND.n224 14.864
R1806 GND.n257 GND.n254 14.864
R1807 GND.n290 GND.n287 14.864
R1808 GND.n335 GND.n332 14.864
R1809 GND.n365 GND.n362 14.864
R1810 GND.n721 GND.n720 14.864
R1811 GND.n691 GND.n690 14.864
R1812 GND.n659 GND.n658 14.864
R1813 GND.n627 GND.n626 14.864
R1814 GND.n583 GND.n582 14.864
R1815 GND.n550 GND.n549 14.864
R1816 GND.n517 GND.n516 14.864
R1817 GND.n484 GND.n483 14.864
R1818 GND.n452 GND.n451 14.864
R1819 GND.n419 GND.n418 14.864
R1820 GND.n377 GND.n376 9.154
R1821 GND.n385 GND.n379 9.154
R1822 GND.n388 GND.n387 9.154
R1823 GND.n391 GND.n390 9.154
R1824 GND.n394 GND.n393 9.154
R1825 GND.n397 GND.n396 9.154
R1826 GND.n400 GND.n399 9.154
R1827 GND.n403 GND.n402 9.154
R1828 GND.n406 GND.n405 9.154
R1829 GND.n409 GND.n408 9.154
R1830 GND.n412 GND.n411 9.154
R1831 GND.n419 GND.n415 9.154
R1832 GND.n422 GND.n421 9.154
R1833 GND.n430 GND.n429 9.154
R1834 GND.n433 GND.n432 9.154
R1835 GND.n436 GND.n435 9.154
R1836 GND.n439 GND.n438 9.154
R1837 GND.n442 GND.n441 9.154
R1838 GND.n445 GND.n444 9.154
R1839 GND.n452 GND.n448 9.154
R1840 GND.n455 GND.n454 9.154
R1841 GND.n462 GND.n461 9.154
R1842 GND.n465 GND.n464 9.154
R1843 GND.n468 GND.n467 9.154
R1844 GND.n471 GND.n470 9.154
R1845 GND.n474 GND.n473 9.154
R1846 GND.n477 GND.n476 9.154
R1847 GND.n484 GND.n480 9.154
R1848 GND.n487 GND.n486 9.154
R1849 GND.n495 GND.n494 9.154
R1850 GND.n498 GND.n497 9.154
R1851 GND.n501 GND.n500 9.154
R1852 GND.n504 GND.n503 9.154
R1853 GND.n507 GND.n506 9.154
R1854 GND.n510 GND.n509 9.154
R1855 GND.n517 GND.n513 9.154
R1856 GND.n520 GND.n519 9.154
R1857 GND.n528 GND.n527 9.154
R1858 GND.n531 GND.n530 9.154
R1859 GND.n534 GND.n533 9.154
R1860 GND.n537 GND.n536 9.154
R1861 GND.n540 GND.n539 9.154
R1862 GND.n543 GND.n542 9.154
R1863 GND.n550 GND.n546 9.154
R1864 GND.n553 GND.n552 9.154
R1865 GND.n561 GND.n560 9.154
R1866 GND.n564 GND.n563 9.154
R1867 GND.n567 GND.n566 9.154
R1868 GND.n570 GND.n569 9.154
R1869 GND.n573 GND.n572 9.154
R1870 GND.n576 GND.n575 9.154
R1871 GND.n583 GND.n579 9.154
R1872 GND.n586 GND.n585 9.154
R1873 GND.n593 GND.n588 9.154
R1874 GND.n596 GND.n595 9.154
R1875 GND.n599 GND.n598 9.154
R1876 GND.n602 GND.n601 9.154
R1877 GND.n605 GND.n604 9.154
R1878 GND.n608 GND.n607 9.154
R1879 GND.n611 GND.n610 9.154
R1880 GND.n614 GND.n613 9.154
R1881 GND.n617 GND.n616 9.154
R1882 GND.n620 GND.n619 9.154
R1883 GND.n627 GND.n623 9.154
R1884 GND.n630 GND.n629 9.154
R1885 GND.n637 GND.n636 9.154
R1886 GND.n640 GND.n639 9.154
R1887 GND.n643 GND.n642 9.154
R1888 GND.n646 GND.n645 9.154
R1889 GND.n649 GND.n648 9.154
R1890 GND.n652 GND.n651 9.154
R1891 GND.n659 GND.n655 9.154
R1892 GND.n662 GND.n661 9.154
R1893 GND.n669 GND.n668 9.154
R1894 GND.n672 GND.n671 9.154
R1895 GND.n675 GND.n674 9.154
R1896 GND.n678 GND.n677 9.154
R1897 GND.n681 GND.n680 9.154
R1898 GND.n684 GND.n683 9.154
R1899 GND.n691 GND.n687 9.154
R1900 GND.n694 GND.n693 9.154
R1901 GND.n699 GND.n698 9.154
R1902 GND.n702 GND.n701 9.154
R1903 GND.n705 GND.n704 9.154
R1904 GND.n708 GND.n707 9.154
R1905 GND.n711 GND.n710 9.154
R1906 GND.n714 GND.n713 9.154
R1907 GND.n721 GND.n717 9.154
R1908 GND.n724 GND.n723 9.154
R1909 GND.n732 GND.n731 9.154
R1910 GND.n735 GND.n734 9.154
R1911 GND.n738 GND.n737 9.154
R1912 GND.n371 GND.n370 9.154
R1913 GND.n368 GND.n367 9.154
R1914 GND.n365 GND.n364 9.154
R1915 GND.n358 GND.n357 9.154
R1916 GND.n355 GND.n354 9.154
R1917 GND.n352 GND.n351 9.154
R1918 GND.n347 GND.n346 9.154
R1919 GND.n344 GND.n343 9.154
R1920 GND.n341 GND.n340 9.154
R1921 GND.n338 GND.n337 9.154
R1922 GND.n335 GND.n334 9.154
R1923 GND.n328 GND.n327 9.154
R1924 GND.n325 GND.n324 9.154
R1925 GND.n322 GND.n316 9.154
R1926 GND.n314 GND.n313 9.154
R1927 GND.n311 GND.n310 9.154
R1928 GND.n308 GND.n307 9.154
R1929 GND.n305 GND.n304 9.154
R1930 GND.n302 GND.n301 9.154
R1931 GND.n299 GND.n298 9.154
R1932 GND.n296 GND.n295 9.154
R1933 GND.n293 GND.n292 9.154
R1934 GND.n290 GND.n289 9.154
R1935 GND.n283 GND.n282 9.154
R1936 GND.n280 GND.n279 9.154
R1937 GND.n277 GND.n276 9.154
R1938 GND.n269 GND.n268 9.154
R1939 GND.n266 GND.n265 9.154
R1940 GND.n263 GND.n262 9.154
R1941 GND.n260 GND.n259 9.154
R1942 GND.n257 GND.n256 9.154
R1943 GND.n250 GND.n249 9.154
R1944 GND.n247 GND.n246 9.154
R1945 GND.n244 GND.n243 9.154
R1946 GND.n239 GND.n238 9.154
R1947 GND.n236 GND.n235 9.154
R1948 GND.n233 GND.n232 9.154
R1949 GND.n230 GND.n229 9.154
R1950 GND.n227 GND.n226 9.154
R1951 GND.n220 GND.n219 9.154
R1952 GND.n217 GND.n216 9.154
R1953 GND.n214 GND.n213 9.154
R1954 GND.n207 GND.n206 9.154
R1955 GND.n204 GND.n203 9.154
R1956 GND.n201 GND.n200 9.154
R1957 GND.n198 GND.n197 9.154
R1958 GND.n195 GND.n194 9.154
R1959 GND.n188 GND.n187 9.154
R1960 GND.n185 GND.n184 9.154
R1961 GND.n182 GND.n181 9.154
R1962 GND.n174 GND.n173 9.154
R1963 GND.n171 GND.n170 9.154
R1964 GND.n168 GND.n167 9.154
R1965 GND.n165 GND.n164 9.154
R1966 GND.n162 GND.n161 9.154
R1967 GND.n155 GND.n154 9.154
R1968 GND.n152 GND.n151 9.154
R1969 GND.n149 GND.n148 9.154
R1970 GND.n142 GND.n141 9.154
R1971 GND.n139 GND.n138 9.154
R1972 GND.n136 GND.n135 9.154
R1973 GND.n133 GND.n132 9.154
R1974 GND.n130 GND.n129 9.154
R1975 GND.n123 GND.n122 9.154
R1976 GND.n120 GND.n119 9.154
R1977 GND.n117 GND.n116 9.154
R1978 GND.n110 GND.n109 9.154
R1979 GND.n107 GND.n106 9.154
R1980 GND.n104 GND.n103 9.154
R1981 GND.n101 GND.n100 9.154
R1982 GND.n98 GND.n97 9.154
R1983 GND.n91 GND.n90 9.154
R1984 GND.n88 GND.n87 9.154
R1985 GND.n85 GND.n84 9.154
R1986 GND.n80 GND.n79 9.154
R1987 GND.n77 GND.n76 9.154
R1988 GND.n8 GND.n7 9.154
R1989 GND.n16 GND.n15 9.154
R1990 GND.n25 GND.n24 9.154
R1991 GND.n28 GND.n27 9.154
R1992 GND.n35 GND.n34 9.154
R1993 GND.n38 GND.n37 9.154
R1994 GND.n41 GND.n40 9.154
R1995 GND.n44 GND.n43 9.154
R1996 GND.n47 GND.n46 9.154
R1997 GND.n55 GND.n54 9.154
R1998 GND.n58 GND.n57 9.154
R1999 GND.n61 GND.n60 9.154
R2000 GND.n68 GND.n67 9.154
R2001 GND.n71 GND.n70 9.154
R2002 GND.n74 GND.n73 9.154
R2003 GND.n114 GND.n113 8.128
R2004 GND.n146 GND.n145 8.128
R2005 GND.n211 GND.n210 8.128
R2006 GND.n666 GND.n665 8.128
R2007 GND.n634 GND.n633 8.128
R2008 GND.n591 GND.n590 8.128
R2009 GND.n459 GND.n458 8.128
R2010 GND.n9 GND.n1 4.795
R2011 GND.n375 GND.n374 4.65
R2012 GND.n78 GND.n77 4.65
R2013 GND.n81 GND.n80 4.65
R2014 GND.n86 GND.n85 4.65
R2015 GND.n89 GND.n88 4.65
R2016 GND.n92 GND.n91 4.65
R2017 GND.n99 GND.n98 4.65
R2018 GND.n102 GND.n101 4.65
R2019 GND.n105 GND.n104 4.65
R2020 GND.n108 GND.n107 4.65
R2021 GND.n111 GND.n110 4.65
R2022 GND.n118 GND.n117 4.65
R2023 GND.n121 GND.n120 4.65
R2024 GND.n124 GND.n123 4.65
R2025 GND.n131 GND.n130 4.65
R2026 GND.n134 GND.n133 4.65
R2027 GND.n137 GND.n136 4.65
R2028 GND.n140 GND.n139 4.65
R2029 GND.n143 GND.n142 4.65
R2030 GND.n150 GND.n149 4.65
R2031 GND.n153 GND.n152 4.65
R2032 GND.n156 GND.n155 4.65
R2033 GND.n163 GND.n162 4.65
R2034 GND.n166 GND.n165 4.65
R2035 GND.n169 GND.n168 4.65
R2036 GND.n172 GND.n171 4.65
R2037 GND.n175 GND.n174 4.65
R2038 GND.n183 GND.n182 4.65
R2039 GND.n186 GND.n185 4.65
R2040 GND.n189 GND.n188 4.65
R2041 GND.n196 GND.n195 4.65
R2042 GND.n199 GND.n198 4.65
R2043 GND.n202 GND.n201 4.65
R2044 GND.n205 GND.n204 4.65
R2045 GND.n208 GND.n207 4.65
R2046 GND.n215 GND.n214 4.65
R2047 GND.n218 GND.n217 4.65
R2048 GND.n221 GND.n220 4.65
R2049 GND.n228 GND.n227 4.65
R2050 GND.n231 GND.n230 4.65
R2051 GND.n234 GND.n233 4.65
R2052 GND.n237 GND.n236 4.65
R2053 GND.n240 GND.n239 4.65
R2054 GND.n245 GND.n244 4.65
R2055 GND.n248 GND.n247 4.65
R2056 GND.n251 GND.n250 4.65
R2057 GND.n258 GND.n257 4.65
R2058 GND.n261 GND.n260 4.65
R2059 GND.n264 GND.n263 4.65
R2060 GND.n267 GND.n266 4.65
R2061 GND.n270 GND.n269 4.65
R2062 GND.n278 GND.n277 4.65
R2063 GND.n281 GND.n280 4.65
R2064 GND.n284 GND.n283 4.65
R2065 GND.n291 GND.n290 4.65
R2066 GND.n294 GND.n293 4.65
R2067 GND.n297 GND.n296 4.65
R2068 GND.n300 GND.n299 4.65
R2069 GND.n303 GND.n302 4.65
R2070 GND.n306 GND.n305 4.65
R2071 GND.n309 GND.n308 4.65
R2072 GND.n312 GND.n311 4.65
R2073 GND.n315 GND.n314 4.65
R2074 GND.n323 GND.n322 4.65
R2075 GND.n326 GND.n325 4.65
R2076 GND.n329 GND.n328 4.65
R2077 GND.n336 GND.n335 4.65
R2078 GND.n339 GND.n338 4.65
R2079 GND.n342 GND.n341 4.65
R2080 GND.n345 GND.n344 4.65
R2081 GND.n348 GND.n347 4.65
R2082 GND.n353 GND.n352 4.65
R2083 GND.n356 GND.n355 4.65
R2084 GND.n359 GND.n358 4.65
R2085 GND.n366 GND.n365 4.65
R2086 GND.n369 GND.n368 4.65
R2087 GND.n372 GND.n371 4.65
R2088 GND.n739 GND.n738 4.65
R2089 GND.n736 GND.n735 4.65
R2090 GND.n733 GND.n732 4.65
R2091 GND.n725 GND.n724 4.65
R2092 GND.n722 GND.n721 4.65
R2093 GND.n715 GND.n714 4.65
R2094 GND.n712 GND.n711 4.65
R2095 GND.n709 GND.n708 4.65
R2096 GND.n706 GND.n705 4.65
R2097 GND.n703 GND.n702 4.65
R2098 GND.n700 GND.n699 4.65
R2099 GND.n695 GND.n694 4.65
R2100 GND.n692 GND.n691 4.65
R2101 GND.n685 GND.n684 4.65
R2102 GND.n682 GND.n681 4.65
R2103 GND.n679 GND.n678 4.65
R2104 GND.n676 GND.n675 4.65
R2105 GND.n673 GND.n672 4.65
R2106 GND.n670 GND.n669 4.65
R2107 GND.n663 GND.n662 4.65
R2108 GND.n660 GND.n659 4.65
R2109 GND.n653 GND.n652 4.65
R2110 GND.n650 GND.n649 4.65
R2111 GND.n647 GND.n646 4.65
R2112 GND.n644 GND.n643 4.65
R2113 GND.n641 GND.n640 4.65
R2114 GND.n638 GND.n637 4.65
R2115 GND.n631 GND.n630 4.65
R2116 GND.n628 GND.n627 4.65
R2117 GND.n621 GND.n620 4.65
R2118 GND.n618 GND.n617 4.65
R2119 GND.n615 GND.n614 4.65
R2120 GND.n612 GND.n611 4.65
R2121 GND.n609 GND.n608 4.65
R2122 GND.n606 GND.n605 4.65
R2123 GND.n603 GND.n602 4.65
R2124 GND.n600 GND.n599 4.65
R2125 GND.n597 GND.n596 4.65
R2126 GND.n594 GND.n593 4.65
R2127 GND.n587 GND.n586 4.65
R2128 GND.n584 GND.n583 4.65
R2129 GND.n577 GND.n576 4.65
R2130 GND.n574 GND.n573 4.65
R2131 GND.n571 GND.n570 4.65
R2132 GND.n568 GND.n567 4.65
R2133 GND.n565 GND.n564 4.65
R2134 GND.n562 GND.n561 4.65
R2135 GND.n554 GND.n553 4.65
R2136 GND.n551 GND.n550 4.65
R2137 GND.n544 GND.n543 4.65
R2138 GND.n541 GND.n540 4.65
R2139 GND.n538 GND.n537 4.65
R2140 GND.n535 GND.n534 4.65
R2141 GND.n532 GND.n531 4.65
R2142 GND.n529 GND.n528 4.65
R2143 GND.n521 GND.n520 4.65
R2144 GND.n518 GND.n517 4.65
R2145 GND.n511 GND.n510 4.65
R2146 GND.n508 GND.n507 4.65
R2147 GND.n505 GND.n504 4.65
R2148 GND.n502 GND.n501 4.65
R2149 GND.n499 GND.n498 4.65
R2150 GND.n496 GND.n495 4.65
R2151 GND.n488 GND.n487 4.65
R2152 GND.n485 GND.n484 4.65
R2153 GND.n478 GND.n477 4.65
R2154 GND.n475 GND.n474 4.65
R2155 GND.n472 GND.n471 4.65
R2156 GND.n469 GND.n468 4.65
R2157 GND.n466 GND.n465 4.65
R2158 GND.n463 GND.n462 4.65
R2159 GND.n456 GND.n455 4.65
R2160 GND.n453 GND.n452 4.65
R2161 GND.n446 GND.n445 4.65
R2162 GND.n443 GND.n442 4.65
R2163 GND.n440 GND.n439 4.65
R2164 GND.n437 GND.n436 4.65
R2165 GND.n434 GND.n433 4.65
R2166 GND.n431 GND.n430 4.65
R2167 GND.n423 GND.n422 4.65
R2168 GND.n420 GND.n419 4.65
R2169 GND.n413 GND.n412 4.65
R2170 GND.n410 GND.n409 4.65
R2171 GND.n407 GND.n406 4.65
R2172 GND.n404 GND.n403 4.65
R2173 GND.n401 GND.n400 4.65
R2174 GND.n398 GND.n397 4.65
R2175 GND.n395 GND.n394 4.65
R2176 GND.n392 GND.n391 4.65
R2177 GND.n389 GND.n388 4.65
R2178 GND.n386 GND.n385 4.65
R2179 GND.n378 GND.n377 4.65
R2180 GND.n9 GND.n8 4.65
R2181 GND.n17 GND.n16 4.65
R2182 GND.n26 GND.n25 4.65
R2183 GND.n29 GND.n28 4.65
R2184 GND.n36 GND.n35 4.65
R2185 GND.n39 GND.n38 4.65
R2186 GND.n42 GND.n41 4.65
R2187 GND.n45 GND.n44 4.65
R2188 GND.n48 GND.n47 4.65
R2189 GND.n56 GND.n55 4.65
R2190 GND.n59 GND.n58 4.65
R2191 GND.n62 GND.n61 4.65
R2192 GND.n69 GND.n68 4.65
R2193 GND.n72 GND.n71 4.65
R2194 GND.n75 GND.n74 4.65
R2195 GND.n19 GND.n18 4.504
R2196 GND.n8 GND.n6 4.129
R2197 GND.n55 GND.n53 4.129
R2198 GND.n85 GND.n83 4.129
R2199 GND.n117 GND.n115 4.129
R2200 GND.n149 GND.n147 4.129
R2201 GND.n182 GND.n180 4.129
R2202 GND.n214 GND.n212 4.129
R2203 GND.n244 GND.n242 4.129
R2204 GND.n277 GND.n275 4.129
R2205 GND.n352 GND.n350 4.129
R2206 GND.n732 GND.n730 4.129
R2207 GND.n699 GND.n697 4.129
R2208 GND.n669 GND.n667 4.129
R2209 GND.n637 GND.n635 4.129
R2210 GND.n561 GND.n559 4.129
R2211 GND.n528 GND.n526 4.129
R2212 GND.n495 GND.n493 4.129
R2213 GND.n462 GND.n460 4.129
R2214 GND.n430 GND.n428 4.129
R2215 GND.n25 GND.n23 3.716
R2216 GND.t0 GND.n19 2.452
R2217 GND.n11 GND.n10 1.935
R2218 GND.n1 GND.n0 0.475
R2219 GND.n374 GND.n373 0.474
R2220 GND.n13 GND.n12 0.376
R2221 GND.n36 GND.n29 0.29
R2222 GND.n69 GND.n62 0.29
R2223 GND.n99 GND.n92 0.29
R2224 GND.n131 GND.n124 0.29
R2225 GND.n163 GND.n156 0.29
R2226 GND.n196 GND.n189 0.29
R2227 GND.n228 GND.n221 0.29
R2228 GND.n258 GND.n251 0.29
R2229 GND.n291 GND.n284 0.29
R2230 GND.n336 GND.n329 0.29
R2231 GND.n366 GND.n359 0.29
R2232 GND.n722 GND.n715 0.29
R2233 GND.n692 GND.n685 0.29
R2234 GND.n660 GND.n653 0.29
R2235 GND.n628 GND.n621 0.29
R2236 GND.n584 GND.n577 0.29
R2237 GND.n551 GND.n544 0.29
R2238 GND.n518 GND.n511 0.29
R2239 GND.n485 GND.n478 0.29
R2240 GND.n453 GND.n446 0.29
R2241 GND.n420 GND.n413 0.29
R2242 GND.n375 GND 0.207
R2243 GND.n16 GND.n14 0.206
R2244 GND.n322 GND.n321 0.206
R2245 GND.n593 GND.n592 0.206
R2246 GND.n385 GND.n384 0.206
R2247 GND.n309 GND.n306 0.197
R2248 GND.n606 GND.n603 0.197
R2249 GND.n398 GND.n395 0.197
R2250 GND.n48 GND.n45 0.181
R2251 GND.n81 GND.n78 0.181
R2252 GND.n111 GND.n108 0.181
R2253 GND.n143 GND.n140 0.181
R2254 GND.n175 GND.n172 0.181
R2255 GND.n208 GND.n205 0.181
R2256 GND.n240 GND.n237 0.181
R2257 GND.n270 GND.n267 0.181
R2258 GND.n348 GND.n345 0.181
R2259 GND.n739 GND.n736 0.181
R2260 GND.n706 GND.n703 0.181
R2261 GND.n676 GND.n673 0.181
R2262 GND.n644 GND.n641 0.181
R2263 GND.n568 GND.n565 0.181
R2264 GND.n535 GND.n532 0.181
R2265 GND.n502 GND.n499 0.181
R2266 GND.n469 GND.n466 0.181
R2267 GND.n437 GND.n434 0.181
R2268 GND.n17 GND.n9 0.157
R2269 GND.n26 GND.n17 0.157
R2270 GND.n29 GND.n26 0.145
R2271 GND.n39 GND.n36 0.145
R2272 GND.n42 GND.n39 0.145
R2273 GND.n45 GND.n42 0.145
R2274 GND.n56 GND.n48 0.145
R2275 GND.n59 GND.n56 0.145
R2276 GND.n62 GND.n59 0.145
R2277 GND.n72 GND.n69 0.145
R2278 GND.n75 GND.n72 0.145
R2279 GND.n78 GND.n75 0.145
R2280 GND.n86 GND.n81 0.145
R2281 GND.n89 GND.n86 0.145
R2282 GND.n92 GND.n89 0.145
R2283 GND.n102 GND.n99 0.145
R2284 GND.n105 GND.n102 0.145
R2285 GND.n108 GND.n105 0.145
R2286 GND.n118 GND.n111 0.145
R2287 GND.n121 GND.n118 0.145
R2288 GND.n124 GND.n121 0.145
R2289 GND.n134 GND.n131 0.145
R2290 GND.n137 GND.n134 0.145
R2291 GND.n140 GND.n137 0.145
R2292 GND.n150 GND.n143 0.145
R2293 GND.n153 GND.n150 0.145
R2294 GND.n156 GND.n153 0.145
R2295 GND.n166 GND.n163 0.145
R2296 GND.n169 GND.n166 0.145
R2297 GND.n172 GND.n169 0.145
R2298 GND.n183 GND.n175 0.145
R2299 GND.n186 GND.n183 0.145
R2300 GND.n189 GND.n186 0.145
R2301 GND.n199 GND.n196 0.145
R2302 GND.n202 GND.n199 0.145
R2303 GND.n205 GND.n202 0.145
R2304 GND.n215 GND.n208 0.145
R2305 GND.n218 GND.n215 0.145
R2306 GND.n221 GND.n218 0.145
R2307 GND.n231 GND.n228 0.145
R2308 GND.n234 GND.n231 0.145
R2309 GND.n237 GND.n234 0.145
R2310 GND.n245 GND.n240 0.145
R2311 GND.n248 GND.n245 0.145
R2312 GND.n251 GND.n248 0.145
R2313 GND.n261 GND.n258 0.145
R2314 GND.n264 GND.n261 0.145
R2315 GND.n267 GND.n264 0.145
R2316 GND.n278 GND.n270 0.145
R2317 GND.n281 GND.n278 0.145
R2318 GND.n284 GND.n281 0.145
R2319 GND.n294 GND.n291 0.145
R2320 GND.n297 GND.n294 0.145
R2321 GND.n300 GND.n297 0.145
R2322 GND.n303 GND.n300 0.145
R2323 GND.n306 GND.n303 0.145
R2324 GND.n312 GND.n309 0.145
R2325 GND.n315 GND.n312 0.145
R2326 GND.n323 GND.n315 0.145
R2327 GND.n326 GND.n323 0.145
R2328 GND.n329 GND.n326 0.145
R2329 GND.n339 GND.n336 0.145
R2330 GND.n342 GND.n339 0.145
R2331 GND.n345 GND.n342 0.145
R2332 GND.n353 GND.n348 0.145
R2333 GND.n356 GND.n353 0.145
R2334 GND.n359 GND.n356 0.145
R2335 GND.n369 GND.n366 0.145
R2336 GND.n372 GND.n369 0.145
R2337 GND.n736 GND.n733 0.145
R2338 GND.n733 GND.n725 0.145
R2339 GND.n725 GND.n722 0.145
R2340 GND.n715 GND.n712 0.145
R2341 GND.n712 GND.n709 0.145
R2342 GND.n709 GND.n706 0.145
R2343 GND.n703 GND.n700 0.145
R2344 GND.n700 GND.n695 0.145
R2345 GND.n695 GND.n692 0.145
R2346 GND.n685 GND.n682 0.145
R2347 GND.n682 GND.n679 0.145
R2348 GND.n679 GND.n676 0.145
R2349 GND.n673 GND.n670 0.145
R2350 GND.n670 GND.n663 0.145
R2351 GND.n663 GND.n660 0.145
R2352 GND.n653 GND.n650 0.145
R2353 GND.n650 GND.n647 0.145
R2354 GND.n647 GND.n644 0.145
R2355 GND.n641 GND.n638 0.145
R2356 GND.n638 GND.n631 0.145
R2357 GND.n631 GND.n628 0.145
R2358 GND.n621 GND.n618 0.145
R2359 GND.n618 GND.n615 0.145
R2360 GND.n615 GND.n612 0.145
R2361 GND.n612 GND.n609 0.145
R2362 GND.n609 GND.n606 0.145
R2363 GND.n603 GND.n600 0.145
R2364 GND.n600 GND.n597 0.145
R2365 GND.n597 GND.n594 0.145
R2366 GND.n594 GND.n587 0.145
R2367 GND.n587 GND.n584 0.145
R2368 GND.n577 GND.n574 0.145
R2369 GND.n574 GND.n571 0.145
R2370 GND.n571 GND.n568 0.145
R2371 GND.n565 GND.n562 0.145
R2372 GND.n562 GND.n554 0.145
R2373 GND.n554 GND.n551 0.145
R2374 GND.n544 GND.n541 0.145
R2375 GND.n541 GND.n538 0.145
R2376 GND.n538 GND.n535 0.145
R2377 GND.n532 GND.n529 0.145
R2378 GND.n529 GND.n521 0.145
R2379 GND.n521 GND.n518 0.145
R2380 GND.n511 GND.n508 0.145
R2381 GND.n508 GND.n505 0.145
R2382 GND.n505 GND.n502 0.145
R2383 GND.n499 GND.n496 0.145
R2384 GND.n496 GND.n488 0.145
R2385 GND.n488 GND.n485 0.145
R2386 GND.n478 GND.n475 0.145
R2387 GND.n475 GND.n472 0.145
R2388 GND.n472 GND.n469 0.145
R2389 GND.n466 GND.n463 0.145
R2390 GND.n463 GND.n456 0.145
R2391 GND.n456 GND.n453 0.145
R2392 GND.n446 GND.n443 0.145
R2393 GND.n443 GND.n440 0.145
R2394 GND.n440 GND.n437 0.145
R2395 GND.n434 GND.n431 0.145
R2396 GND.n431 GND.n423 0.145
R2397 GND.n423 GND.n420 0.145
R2398 GND.n413 GND.n410 0.145
R2399 GND.n410 GND.n407 0.145
R2400 GND.n407 GND.n404 0.145
R2401 GND.n404 GND.n401 0.145
R2402 GND.n401 GND.n398 0.145
R2403 GND.n395 GND.n392 0.145
R2404 GND.n392 GND.n389 0.145
R2405 GND.n389 GND.n386 0.145
R2406 GND.n386 GND.n378 0.145
R2407 GND.n378 GND.n375 0.145
R2408 GND GND.n372 0.086
R2409 GND GND.n739 0.058
R2410 a_11761_1050.n1 a_11761_1050.t6 480.392
R2411 a_11761_1050.n2 a_11761_1050.t7 440.954
R2412 a_11761_1050.n4 a_11761_1050.n3 410.896
R2413 a_11761_1050.n1 a_11761_1050.t5 403.272
R2414 a_11761_1050.n6 a_11761_1050.n5 157.963
R2415 a_11761_1050.n5 a_11761_1050.n0 91.706
R2416 a_11761_1050.n5 a_11761_1050.n4 76.423
R2417 a_11761_1050.n2 a_11761_1050.n1 20.835
R2418 a_11761_1050.n0 a_11761_1050.t0 14.282
R2419 a_11761_1050.n0 a_11761_1050.t1 14.282
R2420 a_11761_1050.n6 a_11761_1050.t2 14.282
R2421 a_11761_1050.t3 a_11761_1050.n6 14.282
R2422 a_11761_1050.n4 a_11761_1050.n2 8.044
R2423 a_11887_411.n3 a_11887_411.t8 512.525
R2424 a_11887_411.n1 a_11887_411.t13 477.179
R2425 a_11887_411.n6 a_11887_411.t5 472.359
R2426 a_11887_411.n2 a_11887_411.t9 440.954
R2427 a_11887_411.n1 a_11887_411.t7 406.485
R2428 a_11887_411.n6 a_11887_411.t6 384.527
R2429 a_11887_411.n5 a_11887_411.t10 378.636
R2430 a_11887_411.n3 a_11887_411.t12 371.139
R2431 a_11887_411.n7 a_11887_411.t11 342.755
R2432 a_11887_411.n13 a_11887_411.n12 333.44
R2433 a_11887_411.n15 a_11887_411.n14 157.963
R2434 a_11887_411.n7 a_11887_411.n6 154.955
R2435 a_11887_411.n14 a_11887_411.n13 132.141
R2436 a_11887_411.n14 a_11887_411.n0 91.706
R2437 a_11887_411.n4 a_11887_411.n3 77.972
R2438 a_11887_411.n5 a_11887_411.n4 55.891
R2439 a_11887_411.n12 a_11887_411.n11 30
R2440 a_11887_411.n10 a_11887_411.n9 24.383
R2441 a_11887_411.n12 a_11887_411.n10 23.684
R2442 a_11887_411.n2 a_11887_411.n1 21.4
R2443 a_11887_411.n0 a_11887_411.t3 14.282
R2444 a_11887_411.n0 a_11887_411.t4 14.282
R2445 a_11887_411.n15 a_11887_411.t0 14.282
R2446 a_11887_411.t1 a_11887_411.n15 14.282
R2447 a_11887_411.n8 a_11887_411.n7 7.597
R2448 a_11887_411.n4 a_11887_411.n2 6.833
R2449 a_11887_411.n8 a_11887_411.n5 5.693
R2450 a_11887_411.n13 a_11887_411.n8 4.65
R2451 D.n5 D.t4 472.359
R2452 D.n2 D.t1 472.359
R2453 D.n0 D.t0 472.359
R2454 D.n5 D.t7 384.527
R2455 D.n2 D.t5 384.527
R2456 D.n0 D.t2 384.527
R2457 D.n6 D.n5 294.249
R2458 D.n3 D.n2 294.249
R2459 D.n1 D.n0 294.249
R2460 D.n6 D.t3 136.225
R2461 D.n3 D.t8 136.225
R2462 D.n1 D.t6 136.225
R2463 D.n4 D.n1 20.384
R2464 D.n7 D.n4 15.734
R2465 D.n4 D.n3 4.65
R2466 D.n7 D.n6 4.65
R2467 D.n7 D 0.046
R2468 a_9183_989.n0 a_9183_989.t5 480.392
R2469 a_9183_989.n2 a_9183_989.t6 454.685
R2470 a_9183_989.n2 a_9183_989.t10 428.979
R2471 a_9183_989.n0 a_9183_989.t7 403.272
R2472 a_9183_989.n1 a_9183_989.t8 357.204
R2473 a_9183_989.n3 a_9183_989.t9 311.683
R2474 a_9183_989.n9 a_9183_989.n8 305.581
R2475 a_9183_989.n3 a_9183_989.n2 171.288
R2476 a_9183_989.n1 a_9183_989.n0 171.288
R2477 a_9183_989.n11 a_9183_989.n9 159.999
R2478 a_9183_989.n11 a_9183_989.n10 157.964
R2479 a_9183_989.n12 a_9183_989.n11 91.705
R2480 a_9183_989.n8 a_9183_989.n7 30
R2481 a_9183_989.n6 a_9183_989.n5 24.383
R2482 a_9183_989.n8 a_9183_989.n6 23.684
R2483 a_9183_989.n10 a_9183_989.t3 14.282
R2484 a_9183_989.n10 a_9183_989.t4 14.282
R2485 a_9183_989.t1 a_9183_989.n12 14.282
R2486 a_9183_989.n12 a_9183_989.t0 14.282
R2487 a_9183_989.n4 a_9183_989.n3 7.597
R2488 a_9183_989.n4 a_9183_989.n1 5.965
R2489 a_9183_989.n9 a_9183_989.n4 4.65
R2490 a_6137_1050.n4 a_6137_1050.t7 480.392
R2491 a_6137_1050.n4 a_6137_1050.t6 403.272
R2492 a_6137_1050.n5 a_6137_1050.t5 357.204
R2493 a_6137_1050.n8 a_6137_1050.n6 305.581
R2494 a_6137_1050.n5 a_6137_1050.n4 171.288
R2495 a_6137_1050.n6 a_6137_1050.n3 159.999
R2496 a_6137_1050.n3 a_6137_1050.n2 157.964
R2497 a_6137_1050.n3 a_6137_1050.n1 91.706
R2498 a_6137_1050.n8 a_6137_1050.n7 30
R2499 a_6137_1050.n9 a_6137_1050.n0 24.383
R2500 a_6137_1050.n9 a_6137_1050.n8 23.684
R2501 a_6137_1050.n1 a_6137_1050.t1 14.282
R2502 a_6137_1050.n1 a_6137_1050.t0 14.282
R2503 a_6137_1050.n2 a_6137_1050.t4 14.282
R2504 a_6137_1050.n2 a_6137_1050.t3 14.282
R2505 a_6137_1050.n6 a_6137_1050.n5 10.615
R2506 a_6698_101.n11 a_6698_101.n10 68.43
R2507 a_6698_101.n3 a_6698_101.n2 62.817
R2508 a_6698_101.n7 a_6698_101.n6 38.626
R2509 a_6698_101.n6 a_6698_101.n5 35.955
R2510 a_6698_101.n3 a_6698_101.n1 26.202
R2511 a_6698_101.t0 a_6698_101.n3 19.737
R2512 a_6698_101.t1 a_6698_101.n8 8.137
R2513 a_6698_101.t0 a_6698_101.n4 7.273
R2514 a_6698_101.t0 a_6698_101.n0 6.109
R2515 a_6698_101.t1 a_6698_101.n7 4.864
R2516 a_6698_101.t0 a_6698_101.n12 2.074
R2517 a_6698_101.n12 a_6698_101.t1 0.937
R2518 a_6698_101.t1 a_6698_101.n11 0.763
R2519 a_6698_101.n11 a_6698_101.n9 0.185
R2520 a_7595_411.n4 a_7595_411.t6 475.572
R2521 a_7595_411.n8 a_7595_411.t9 472.359
R2522 a_7595_411.n3 a_7595_411.t8 469.145
R2523 a_7595_411.n8 a_7595_411.t13 384.527
R2524 a_7595_411.n4 a_7595_411.t12 384.527
R2525 a_7595_411.n3 a_7595_411.t11 384.527
R2526 a_7595_411.n5 a_7595_411.t10 370.613
R2527 a_7595_411.n9 a_7595_411.n8 266.39
R2528 a_7595_411.n11 a_7595_411.n2 243.576
R2529 a_7595_411.n9 a_7595_411.t7 231.319
R2530 a_7595_411.n7 a_7595_411.t5 231.319
R2531 a_7595_411.n13 a_7595_411.n11 228.526
R2532 a_7595_411.n2 a_7595_411.n1 157.964
R2533 a_7595_411.n7 a_7595_411.n6 139.294
R2534 a_7595_411.n5 a_7595_411.n4 128.028
R2535 a_7595_411.n6 a_7595_411.n3 126.97
R2536 a_7595_411.n2 a_7595_411.n0 91.706
R2537 a_7595_411.n10 a_7595_411.n7 22.288
R2538 a_7595_411.n13 a_7595_411.n12 15.218
R2539 a_7595_411.n0 a_7595_411.t2 14.282
R2540 a_7595_411.n0 a_7595_411.t3 14.282
R2541 a_7595_411.n1 a_7595_411.t1 14.282
R2542 a_7595_411.n1 a_7595_411.t0 14.282
R2543 a_7595_411.n6 a_7595_411.n5 14.151
R2544 a_7595_411.n14 a_7595_411.n13 12.014
R2545 a_7595_411.n10 a_7595_411.n9 7.597
R2546 a_7595_411.n11 a_7595_411.n10 4.65
R2547 a_12988_101.n3 a_12988_101.n2 62.817
R2548 a_12988_101.n11 a_12988_101.n10 46.054
R2549 a_12988_101.n7 a_12988_101.n6 38.626
R2550 a_12988_101.n6 a_12988_101.n5 35.955
R2551 a_12988_101.n12 a_12988_101.n11 27.923
R2552 a_12988_101.n3 a_12988_101.n1 26.202
R2553 a_12988_101.t0 a_12988_101.n3 19.737
R2554 a_12988_101.t0 a_12988_101.n4 7.273
R2555 a_12988_101.n9 a_12988_101.n8 6.883
R2556 a_12988_101.t0 a_12988_101.n0 6.109
R2557 a_12988_101.t1 a_12988_101.n7 4.864
R2558 a_12988_101.t0 a_12988_101.n13 2.074
R2559 a_12988_101.t1 a_12988_101.n9 1.179
R2560 a_12988_101.t1 a_12988_101.n12 0.958
R2561 a_12988_101.n13 a_12988_101.t1 0.937
R2562 a_3072_101.n11 a_3072_101.n10 68.43
R2563 a_3072_101.n3 a_3072_101.n2 62.817
R2564 a_3072_101.n7 a_3072_101.n6 38.626
R2565 a_3072_101.n6 a_3072_101.n5 35.955
R2566 a_3072_101.n3 a_3072_101.n1 26.202
R2567 a_3072_101.t0 a_3072_101.n3 19.737
R2568 a_3072_101.t1 a_3072_101.n8 8.137
R2569 a_3072_101.t0 a_3072_101.n4 7.273
R2570 a_3072_101.t0 a_3072_101.n0 6.109
R2571 a_3072_101.t1 a_3072_101.n7 4.864
R2572 a_3072_101.t0 a_3072_101.n12 2.074
R2573 a_3072_101.n12 a_3072_101.t1 0.937
R2574 a_3072_101.t1 a_3072_101.n11 0.763
R2575 a_3072_101.n11 a_3072_101.n9 0.185
R2576 a_4891_989.n0 a_4891_989.t9 480.392
R2577 a_4891_989.n2 a_4891_989.t6 454.685
R2578 a_4891_989.n2 a_4891_989.t8 428.979
R2579 a_4891_989.n0 a_4891_989.t10 403.272
R2580 a_4891_989.n1 a_4891_989.t5 357.204
R2581 a_4891_989.n3 a_4891_989.t7 311.683
R2582 a_4891_989.n9 a_4891_989.n8 305.581
R2583 a_4891_989.n3 a_4891_989.n2 171.288
R2584 a_4891_989.n1 a_4891_989.n0 171.288
R2585 a_4891_989.n11 a_4891_989.n9 159.999
R2586 a_4891_989.n11 a_4891_989.n10 157.964
R2587 a_4891_989.n12 a_4891_989.n11 91.705
R2588 a_4891_989.n8 a_4891_989.n7 30
R2589 a_4891_989.n6 a_4891_989.n5 24.383
R2590 a_4891_989.n8 a_4891_989.n6 23.684
R2591 a_4891_989.n10 a_4891_989.t4 14.282
R2592 a_4891_989.n10 a_4891_989.t3 14.282
R2593 a_4891_989.t1 a_4891_989.n12 14.282
R2594 a_4891_989.n12 a_4891_989.t0 14.282
R2595 a_4891_989.n4 a_4891_989.n3 7.597
R2596 a_4891_989.n4 a_4891_989.n1 5.965
R2597 a_4891_989.n9 a_4891_989.n4 4.65
R2598 a_7469_1050.n0 a_7469_1050.t5 480.392
R2599 a_7469_1050.n0 a_7469_1050.t7 403.272
R2600 a_7469_1050.n1 a_7469_1050.t6 385.063
R2601 a_7469_1050.n6 a_7469_1050.n5 333.44
R2602 a_7469_1050.n8 a_7469_1050.n7 157.964
R2603 a_7469_1050.n1 a_7469_1050.n0 143.429
R2604 a_7469_1050.n8 a_7469_1050.n6 132.141
R2605 a_7469_1050.n9 a_7469_1050.n8 91.705
R2606 a_7469_1050.n5 a_7469_1050.n4 30
R2607 a_7469_1050.n3 a_7469_1050.n2 24.383
R2608 a_7469_1050.n5 a_7469_1050.n3 23.684
R2609 a_7469_1050.n7 a_7469_1050.t0 14.282
R2610 a_7469_1050.n7 a_7469_1050.t1 14.282
R2611 a_7469_1050.t3 a_7469_1050.n9 14.282
R2612 a_7469_1050.n9 a_7469_1050.t2 14.282
R2613 a_7469_1050.n6 a_7469_1050.n1 10.615
R2614 a_6032_101.n3 a_6032_101.n1 42.788
R2615 a_6032_101.t0 a_6032_101.n0 8.137
R2616 a_6032_101.n3 a_6032_101.n2 4.665
R2617 a_6032_101.t0 a_6032_101.n3 0.06
R2618 CLK.n15 CLK.t1 472.359
R2619 CLK.n6 CLK.t2 472.359
R2620 CLK.n0 CLK.t12 472.359
R2621 CLK.n20 CLK.t0 459.505
R2622 CLK.n11 CLK.t5 459.505
R2623 CLK.n2 CLK.t14 459.505
R2624 CLK.n21 CLK.t10 399.181
R2625 CLK.n12 CLK.t13 399.181
R2626 CLK.n3 CLK.t7 399.181
R2627 CLK.n1 CLK.t15 398.558
R2628 CLK.n17 CLK.t11 397.101
R2629 CLK.n8 CLK.t6 397.101
R2630 CLK.n20 CLK.t8 384.527
R2631 CLK.n15 CLK.t9 384.527
R2632 CLK.n11 CLK.t16 384.527
R2633 CLK.n6 CLK.t3 384.527
R2634 CLK.n2 CLK.t17 384.527
R2635 CLK.n0 CLK.t4 384.527
R2636 CLK.n21 CLK.n20 33.832
R2637 CLK.n3 CLK.n2 33.832
R2638 CLK.n12 CLK.n11 33.832
R2639 CLK.n1 CLK.n0 32.394
R2640 CLK.n16 CLK.n15 30.822
R2641 CLK.n7 CLK.n6 30.822
R2642 CLK.n4 CLK.n1 9.575
R2643 CLK.n13 CLK.n10 8.078
R2644 CLK.n22 CLK.n19 8.078
R2645 CLK.n14 CLK.n13 7.797
R2646 CLK.n5 CLK.n4 7.564
R2647 CLK.n17 CLK.n16 4.577
R2648 CLK.n8 CLK.n7 4.577
R2649 CLK.n9 CLK.n8 4.282
R2650 CLK.n18 CLK.n17 4.282
R2651 CLK.n4 CLK.n3 2.079
R2652 CLK.n13 CLK.n12 2.079
R2653 CLK.n22 CLK.n21 2.079
R2654 CLK.n22 CLK 0.046
R2655 CLK.n10 CLK.n9 0.038
R2656 CLK.n19 CLK.n18 0.038
R2657 CLK.n9 CLK.n5 0.008
R2658 CLK.n18 CLK.n14 0.008
R2659 a_14320_101.n3 a_14320_101.n1 42.788
R2660 a_14320_101.t0 a_14320_101.n0 8.137
R2661 a_14320_101.n3 a_14320_101.n2 4.665
R2662 a_14320_101.t0 a_14320_101.n3 0.06
R2663 a_13757_1051.t3 a_13757_1051.n5 179.898
R2664 a_13757_1051.n3 a_13757_1051.n2 165.613
R2665 a_13757_1051.n3 a_13757_1051.n1 142.653
R2666 a_13757_1051.n5 a_13757_1051.n4 106.183
R2667 a_13757_1051.n5 a_13757_1051.n0 99.355
R2668 a_13757_1051.n4 a_13757_1051.n3 82.665
R2669 a_13757_1051.n4 a_13757_1051.t4 73.712
R2670 a_13757_1051.n1 a_13757_1051.t7 14.282
R2671 a_13757_1051.n1 a_13757_1051.t6 14.282
R2672 a_13757_1051.n2 a_13757_1051.t1 14.282
R2673 a_13757_1051.n2 a_13757_1051.t0 14.282
R2674 a_13757_1051.n0 a_13757_1051.t2 14.282
R2675 a_13757_1051.n0 a_13757_1051.t5 14.282
R2676 a_7364_101.n11 a_7364_101.n10 68.43
R2677 a_7364_101.n3 a_7364_101.n2 62.817
R2678 a_7364_101.n7 a_7364_101.n6 38.626
R2679 a_7364_101.n6 a_7364_101.n5 35.955
R2680 a_7364_101.n3 a_7364_101.n1 26.202
R2681 a_7364_101.t0 a_7364_101.n3 19.737
R2682 a_7364_101.t1 a_7364_101.n8 8.137
R2683 a_7364_101.t0 a_7364_101.n4 7.273
R2684 a_7364_101.t0 a_7364_101.n0 6.109
R2685 a_7364_101.t1 a_7364_101.n7 4.864
R2686 a_7364_101.t0 a_7364_101.n12 2.074
R2687 a_7364_101.n12 a_7364_101.t1 0.937
R2688 a_7364_101.t1 a_7364_101.n11 0.763
R2689 a_7364_101.n11 a_7364_101.n9 0.185
R2690 a_3738_101.n3 a_3738_101.n1 42.788
R2691 a_3738_101.t0 a_3738_101.n0 8.137
R2692 a_3738_101.n3 a_3738_101.n2 4.665
R2693 a_3738_101.t0 a_3738_101.n3 0.06
R2694 a_10324_101.n5 a_10324_101.n4 62.817
R2695 a_10324_101.n2 a_10324_101.n0 41.528
R2696 a_10324_101.n5 a_10324_101.n3 26.202
R2697 a_10324_101.t0 a_10324_101.n5 19.737
R2698 a_10324_101.t0 a_10324_101.n6 8.137
R2699 a_10324_101.n2 a_10324_101.n1 3.644
R2700 a_10324_101.t0 a_10324_101.n2 1.093
R2701 a_10429_1050.n1 a_10429_1050.t7 480.392
R2702 a_10429_1050.n1 a_10429_1050.t5 403.272
R2703 a_10429_1050.n2 a_10429_1050.t6 357.204
R2704 a_10429_1050.n4 a_10429_1050.n3 327.32
R2705 a_10429_1050.n2 a_10429_1050.n1 171.288
R2706 a_10429_1050.n5 a_10429_1050.n4 159.999
R2707 a_10429_1050.n6 a_10429_1050.n5 157.963
R2708 a_10429_1050.n5 a_10429_1050.n0 91.706
R2709 a_10429_1050.n0 a_10429_1050.t3 14.282
R2710 a_10429_1050.n0 a_10429_1050.t2 14.282
R2711 a_10429_1050.t1 a_10429_1050.n6 14.282
R2712 a_10429_1050.n6 a_10429_1050.t0 14.282
R2713 a_10429_1050.n4 a_10429_1050.n2 10.615
R2714 a_4439_187.n5 a_4439_187.t5 512.525
R2715 a_4439_187.n3 a_4439_187.t12 472.359
R2716 a_4439_187.n1 a_4439_187.t13 472.359
R2717 a_4439_187.n6 a_4439_187.t8 417.109
R2718 a_4439_187.n3 a_4439_187.t6 384.527
R2719 a_4439_187.n1 a_4439_187.t10 384.527
R2720 a_4439_187.n10 a_4439_187.n9 383.037
R2721 a_4439_187.n5 a_4439_187.t11 371.139
R2722 a_4439_187.n4 a_4439_187.t7 370.613
R2723 a_4439_187.n2 a_4439_187.t9 370.613
R2724 a_4439_187.n6 a_4439_187.n5 179.837
R2725 a_4439_187.n12 a_4439_187.n11 157.963
R2726 a_4439_187.n4 a_4439_187.n3 127.096
R2727 a_4439_187.n2 a_4439_187.n1 127.096
R2728 a_4439_187.n11 a_4439_187.n10 104.282
R2729 a_4439_187.n11 a_4439_187.n0 91.706
R2730 a_4439_187.n0 a_4439_187.t3 14.282
R2731 a_4439_187.n0 a_4439_187.t2 14.282
R2732 a_4439_187.n12 a_4439_187.t0 14.282
R2733 a_4439_187.t1 a_4439_187.n12 14.282
R2734 a_4439_187.n7 a_4439_187.n6 11.134
R2735 a_4439_187.n8 a_4439_187.n2 8.957
R2736 a_4439_187.n7 a_4439_187.n4 4.65
R2737 a_4439_187.n10 a_4439_187.n8 4.65
R2738 a_4439_187.n8 a_4439_187.n7 2.947
R2739 a_8675_103.t0 a_8675_103.n7 59.616
R2740 a_8675_103.n4 a_8675_103.n2 54.496
R2741 a_8675_103.n4 a_8675_103.n3 54.496
R2742 a_8675_103.n1 a_8675_103.n0 24.679
R2743 a_8675_103.n6 a_8675_103.n4 7.859
R2744 a_8675_103.t0 a_8675_103.n1 7.505
R2745 a_8675_103.t0 a_8675_103.n6 3.034
R2746 a_8675_103.n6 a_8675_103.n5 0.443
R2747 a_599_989.n0 a_599_989.t7 480.392
R2748 a_599_989.n2 a_599_989.t9 454.685
R2749 a_599_989.n2 a_599_989.t5 428.979
R2750 a_599_989.n0 a_599_989.t10 403.272
R2751 a_599_989.n1 a_599_989.t8 357.204
R2752 a_599_989.n3 a_599_989.t6 311.683
R2753 a_599_989.n9 a_599_989.n8 305.581
R2754 a_599_989.n3 a_599_989.n2 171.288
R2755 a_599_989.n1 a_599_989.n0 171.288
R2756 a_599_989.n11 a_599_989.n9 159.999
R2757 a_599_989.n11 a_599_989.n10 157.964
R2758 a_599_989.n12 a_599_989.n11 91.705
R2759 a_599_989.n8 a_599_989.n7 30
R2760 a_599_989.n6 a_599_989.n5 24.383
R2761 a_599_989.n8 a_599_989.n6 23.684
R2762 a_599_989.n10 a_599_989.t4 14.282
R2763 a_599_989.n10 a_599_989.t3 14.282
R2764 a_599_989.t1 a_599_989.n12 14.282
R2765 a_599_989.n12 a_599_989.t0 14.282
R2766 a_599_989.n4 a_599_989.n3 7.597
R2767 a_599_989.n4 a_599_989.n1 5.965
R2768 a_599_989.n9 a_599_989.n4 4.65
R2769 a_8030_101.n11 a_8030_101.n10 68.43
R2770 a_8030_101.n3 a_8030_101.n2 62.817
R2771 a_8030_101.n7 a_8030_101.n6 38.626
R2772 a_8030_101.n6 a_8030_101.n5 35.955
R2773 a_8030_101.n3 a_8030_101.n1 26.202
R2774 a_8030_101.t0 a_8030_101.n3 19.737
R2775 a_8030_101.t1 a_8030_101.n8 8.137
R2776 a_8030_101.t0 a_8030_101.n4 7.273
R2777 a_8030_101.t0 a_8030_101.n0 6.109
R2778 a_8030_101.t1 a_8030_101.n7 4.864
R2779 a_8030_101.t0 a_8030_101.n12 2.074
R2780 a_8030_101.n12 a_8030_101.t1 0.937
R2781 a_8030_101.t1 a_8030_101.n11 0.763
R2782 a_8030_101.n11 a_8030_101.n9 0.185
R2783 a_1074_101.n3 a_1074_101.n1 42.788
R2784 a_1074_101.t0 a_1074_101.n0 8.137
R2785 a_1074_101.n3 a_1074_101.n2 4.665
R2786 a_1074_101.t0 a_1074_101.n3 0.06
R2787 a_4569_1050.n3 a_4569_1050.t12 480.392
R2788 a_4569_1050.n1 a_4569_1050.t7 480.392
R2789 a_4569_1050.n3 a_4569_1050.t9 403.272
R2790 a_4569_1050.n1 a_4569_1050.t10 403.272
R2791 a_4569_1050.n4 a_4569_1050.t8 385.063
R2792 a_4569_1050.n2 a_4569_1050.t11 385.063
R2793 a_4569_1050.n10 a_4569_1050.n9 336.075
R2794 a_4569_1050.n13 a_4569_1050.n12 161.352
R2795 a_4569_1050.n11 a_4569_1050.n10 151.34
R2796 a_4569_1050.n4 a_4569_1050.n3 143.429
R2797 a_4569_1050.n2 a_4569_1050.n1 143.429
R2798 a_4569_1050.n11 a_4569_1050.n0 95.095
R2799 a_4569_1050.n14 a_4569_1050.n13 95.094
R2800 a_4569_1050.n13 a_4569_1050.n11 66.258
R2801 a_4569_1050.n9 a_4569_1050.n8 30
R2802 a_4569_1050.n7 a_4569_1050.n6 24.383
R2803 a_4569_1050.n9 a_4569_1050.n7 23.684
R2804 a_4569_1050.n0 a_4569_1050.t2 14.282
R2805 a_4569_1050.n0 a_4569_1050.t3 14.282
R2806 a_4569_1050.n12 a_4569_1050.t6 14.282
R2807 a_4569_1050.n12 a_4569_1050.t5 14.282
R2808 a_4569_1050.t1 a_4569_1050.n14 14.282
R2809 a_4569_1050.n14 a_4569_1050.t0 14.282
R2810 a_4569_1050.n5 a_4569_1050.n2 11.95
R2811 a_4569_1050.n10 a_4569_1050.n5 5.965
R2812 a_4569_1050.n5 a_4569_1050.n4 4.65
R2813 Q.n2 Q.n1 349.908
R2814 Q.n2 Q.n0 215.564
R2815 Q.n0 Q.t0 14.282
R2816 Q.n0 Q.t1 14.282
R2817 Q.n3 Q.n2 4.65
R2818 Q.n3 Q 0.046
R2819 a_12322_101.n11 a_12322_101.n10 68.43
R2820 a_12322_101.n3 a_12322_101.n2 62.817
R2821 a_12322_101.n7 a_12322_101.n6 38.626
R2822 a_12322_101.n6 a_12322_101.n5 35.955
R2823 a_12322_101.n3 a_12322_101.n1 26.202
R2824 a_12322_101.t0 a_12322_101.n3 19.737
R2825 a_12322_101.t1 a_12322_101.n8 8.137
R2826 a_12322_101.t0 a_12322_101.n4 7.273
R2827 a_12322_101.t0 a_12322_101.n0 6.109
R2828 a_12322_101.t1 a_12322_101.n7 4.864
R2829 a_12322_101.t0 a_12322_101.n12 2.074
R2830 a_12322_101.n12 a_12322_101.t1 0.937
R2831 a_12322_101.t1 a_12322_101.n11 0.763
R2832 a_12322_101.n11 a_12322_101.n9 0.185
R2833 a_2406_101.n11 a_2406_101.n10 68.43
R2834 a_2406_101.n3 a_2406_101.n2 62.817
R2835 a_2406_101.n7 a_2406_101.n6 38.626
R2836 a_2406_101.n6 a_2406_101.n5 35.955
R2837 a_2406_101.n3 a_2406_101.n1 26.202
R2838 a_2406_101.t0 a_2406_101.n3 19.737
R2839 a_2406_101.t1 a_2406_101.n8 8.137
R2840 a_2406_101.t0 a_2406_101.n4 7.273
R2841 a_2406_101.t0 a_2406_101.n0 6.109
R2842 a_2406_101.t1 a_2406_101.n7 4.864
R2843 a_2406_101.t0 a_2406_101.n12 2.074
R2844 a_2406_101.n12 a_2406_101.t1 0.937
R2845 a_2406_101.t1 a_2406_101.n11 0.763
R2846 a_2406_101.n11 a_2406_101.n9 0.185
R2847 a_372_210.n10 a_372_210.n8 171.558
R2848 a_372_210.n8 a_372_210.t1 75.764
R2849 a_372_210.n3 a_372_210.n2 27.476
R2850 a_372_210.n10 a_372_210.n9 27.2
R2851 a_372_210.n11 a_372_210.n0 23.498
R2852 a_372_210.n11 a_372_210.n10 22.4
R2853 a_372_210.t1 a_372_210.n5 20.241
R2854 a_372_210.n7 a_372_210.n6 19.952
R2855 a_372_210.t1 a_372_210.n3 13.984
R2856 a_372_210.n5 a_372_210.n4 13.494
R2857 a_372_210.t1 a_372_210.n1 7.04
R2858 a_372_210.n8 a_372_210.n7 1.505
R2859 a_9658_101.n3 a_9658_101.n1 42.788
R2860 a_9658_101.t0 a_9658_101.n0 8.137
R2861 a_9658_101.n3 a_9658_101.n2 4.665
R2862 a_9658_101.t0 a_9658_101.n3 0.06
R2863 a_13093_1051.n2 a_13093_1051.t7 179.895
R2864 a_13093_1051.n5 a_13093_1051.n4 157.021
R2865 a_13093_1051.n4 a_13093_1051.n0 124.955
R2866 a_13093_1051.n3 a_13093_1051.n2 106.183
R2867 a_13093_1051.n2 a_13093_1051.n1 99.355
R2868 a_13093_1051.n4 a_13093_1051.n3 82.65
R2869 a_13093_1051.n3 a_13093_1051.t3 73.712
R2870 a_13093_1051.n0 a_13093_1051.t5 14.282
R2871 a_13093_1051.n0 a_13093_1051.t4 14.282
R2872 a_13093_1051.n1 a_13093_1051.t6 14.282
R2873 a_13093_1051.n1 a_13093_1051.t2 14.282
R2874 a_13093_1051.t1 a_13093_1051.n5 14.282
R2875 a_13093_1051.n5 a_13093_1051.t0 14.282
R2876 a_4664_210.n10 a_4664_210.n8 171.558
R2877 a_4664_210.n8 a_4664_210.t1 75.764
R2878 a_4664_210.n3 a_4664_210.n2 27.476
R2879 a_4664_210.n10 a_4664_210.n9 27.2
R2880 a_4664_210.n11 a_4664_210.n0 23.498
R2881 a_4664_210.n11 a_4664_210.n10 22.4
R2882 a_4664_210.t1 a_4664_210.n5 20.241
R2883 a_4664_210.n7 a_4664_210.n6 19.952
R2884 a_4664_210.t1 a_4664_210.n3 13.984
R2885 a_4664_210.n5 a_4664_210.n4 13.494
R2886 a_4664_210.t1 a_4664_210.n1 7.04
R2887 a_4664_210.n8 a_4664_210.n7 1.505
R2888 a_8956_210.n8 a_8956_210.n6 185.173
R2889 a_8956_210.t0 a_8956_210.n8 75.765
R2890 a_8956_210.n3 a_8956_210.n1 74.827
R2891 a_8956_210.n3 a_8956_210.n2 27.476
R2892 a_8956_210.n6 a_8956_210.n5 22.349
R2893 a_8956_210.t0 a_8956_210.n10 20.241
R2894 a_8956_210.t0 a_8956_210.n3 13.984
R2895 a_8956_210.n10 a_8956_210.n9 13.494
R2896 a_8956_210.n6 a_8956_210.n4 8.443
R2897 a_8956_210.t0 a_8956_210.n0 8.137
R2898 a_8956_210.n8 a_8956_210.n7 1.505
R2899 a_91_103.n5 a_91_103.n4 66.708
R2900 a_91_103.n2 a_91_103.n0 25.439
R2901 a_91_103.n5 a_91_103.n3 19.496
R2902 a_91_103.t0 a_91_103.n5 13.756
R2903 a_91_103.n2 a_91_103.n1 2.455
R2904 a_91_103.t0 a_91_103.n2 0.246
R2905 a_11656_101.n3 a_11656_101.n1 42.788
R2906 a_11656_101.t0 a_11656_101.n0 8.137
R2907 a_11656_101.n3 a_11656_101.n2 4.665
R2908 a_11656_101.t0 a_11656_101.n3 0.06
R2909 a_10990_101.n3 a_10990_101.n1 42.788
R2910 a_10990_101.t0 a_10990_101.n0 8.137
R2911 a_10990_101.n3 a_10990_101.n2 4.665
R2912 a_10990_101.t0 a_10990_101.n3 0.06
R2913 a_4383_103.t0 a_4383_103.n7 59.616
R2914 a_4383_103.n4 a_4383_103.n2 54.496
R2915 a_4383_103.n4 a_4383_103.n3 54.496
R2916 a_4383_103.n1 a_4383_103.n0 24.679
R2917 a_4383_103.t0 a_4383_103.n1 7.505
R2918 a_4383_103.n6 a_4383_103.n5 2.455
R2919 a_4383_103.n6 a_4383_103.n4 0.636
R2920 a_4383_103.t0 a_4383_103.n6 0.246
R2921 a_1740_101.n3 a_1740_101.n1 42.788
R2922 a_1740_101.t0 a_1740_101.n0 8.137
R2923 a_1740_101.n3 a_1740_101.n2 4.665
R2924 a_1740_101.t0 a_1740_101.n3 0.06
R2925 a_5366_101.n3 a_5366_101.n1 42.788
R2926 a_5366_101.t0 a_5366_101.n0 8.137
R2927 a_5366_101.n3 a_5366_101.n2 4.665
R2928 a_5366_101.t0 a_5366_101.n3 0.06
C4 VDD GND 24.52fF
C5 a_5366_101.n0 GND 0.05fF
C6 a_5366_101.n1 GND 0.12fF
C7 a_5366_101.n2 GND 0.04fF
C8 a_5366_101.n3 GND 0.17fF
C9 a_1740_101.n0 GND 0.05fF
C10 a_1740_101.n1 GND 0.12fF
C11 a_1740_101.n2 GND 0.04fF
C12 a_1740_101.n3 GND 0.17fF
C13 a_4383_103.n0 GND 0.08fF
C14 a_4383_103.n1 GND 0.07fF
C15 a_4383_103.n2 GND 0.04fF
C16 a_4383_103.n3 GND 0.06fF
C17 a_4383_103.n4 GND 0.03fF
C18 a_4383_103.n5 GND 0.04fF
C19 a_4383_103.n7 GND 0.08fF
C20 a_10990_101.n0 GND 0.05fF
C21 a_10990_101.n1 GND 0.12fF
C22 a_10990_101.n2 GND 0.04fF
C23 a_10990_101.n3 GND 0.17fF
C24 a_11656_101.n0 GND 0.05fF
C25 a_11656_101.n1 GND 0.12fF
C26 a_11656_101.n2 GND 0.04fF
C27 a_11656_101.n3 GND 0.17fF
C28 a_91_103.n0 GND 0.10fF
C29 a_91_103.n1 GND 0.03fF
C30 a_91_103.n2 GND 0.03fF
C31 a_91_103.n3 GND 0.07fF
C32 a_91_103.n4 GND 0.08fF
C33 a_91_103.n5 GND 0.03fF
C34 a_8956_210.n0 GND 0.07fF
C35 a_8956_210.n1 GND 0.09fF
C36 a_8956_210.n2 GND 0.12fF
C37 a_8956_210.n3 GND 0.08fF
C38 a_8956_210.n4 GND 0.02fF
C39 a_8956_210.n5 GND 0.03fF
C40 a_8956_210.n6 GND 0.05fF
C41 a_8956_210.n7 GND 0.02fF
C42 a_8956_210.n8 GND 0.14fF
C43 a_8956_210.n9 GND 0.08fF
C44 a_8956_210.n10 GND 0.02fF
C45 a_8956_210.t0 GND 0.31fF
C46 a_4664_210.n0 GND 0.02fF
C47 a_4664_210.n1 GND 0.09fF
C48 a_4664_210.n2 GND 0.12fF
C49 a_4664_210.n3 GND 0.08fF
C50 a_4664_210.n4 GND 0.08fF
C51 a_4664_210.n5 GND 0.02fF
C52 a_4664_210.t1 GND 0.29fF
C53 a_4664_210.n6 GND 0.09fF
C54 a_4664_210.n7 GND 0.02fF
C55 a_4664_210.n8 GND 0.13fF
C56 a_4664_210.n9 GND 0.02fF
C57 a_4664_210.n10 GND 0.03fF
C58 a_4664_210.n11 GND 0.03fF
C59 a_13093_1051.n0 GND 0.36fF
C60 a_13093_1051.n1 GND 0.32fF
C61 a_13093_1051.n2 GND 0.53fF
C62 a_13093_1051.n3 GND 0.30fF
C63 a_13093_1051.n4 GND 0.81fF
C64 a_13093_1051.n5 GND 0.43fF
C65 a_9658_101.n0 GND 0.05fF
C66 a_9658_101.n1 GND 0.12fF
C67 a_9658_101.n2 GND 0.04fF
C68 a_9658_101.n3 GND 0.17fF
C69 a_372_210.n0 GND 0.02fF
C70 a_372_210.n1 GND 0.09fF
C71 a_372_210.n2 GND 0.12fF
C72 a_372_210.n3 GND 0.08fF
C73 a_372_210.n4 GND 0.08fF
C74 a_372_210.n5 GND 0.02fF
C75 a_372_210.t1 GND 0.29fF
C76 a_372_210.n6 GND 0.09fF
C77 a_372_210.n7 GND 0.02fF
C78 a_372_210.n8 GND 0.13fF
C79 a_372_210.n9 GND 0.02fF
C80 a_372_210.n10 GND 0.03fF
C81 a_372_210.n11 GND 0.03fF
C82 a_2406_101.n0 GND 0.02fF
C83 a_2406_101.n1 GND 0.09fF
C84 a_2406_101.n2 GND 0.08fF
C85 a_2406_101.n3 GND 0.03fF
C86 a_2406_101.n4 GND 0.01fF
C87 a_2406_101.n5 GND 0.04fF
C88 a_2406_101.n6 GND 0.04fF
C89 a_2406_101.n7 GND 0.02fF
C90 a_2406_101.n8 GND 0.05fF
C91 a_2406_101.n9 GND 0.15fF
C92 a_2406_101.n10 GND 0.08fF
C93 a_2406_101.n11 GND 0.08fF
C94 a_2406_101.t1 GND 0.23fF
C95 a_2406_101.n12 GND 0.01fF
C96 a_12322_101.n0 GND 0.02fF
C97 a_12322_101.n1 GND 0.09fF
C98 a_12322_101.n2 GND 0.08fF
C99 a_12322_101.n3 GND 0.03fF
C100 a_12322_101.n4 GND 0.01fF
C101 a_12322_101.n5 GND 0.04fF
C102 a_12322_101.n6 GND 0.04fF
C103 a_12322_101.n7 GND 0.02fF
C104 a_12322_101.n8 GND 0.05fF
C105 a_12322_101.n9 GND 0.15fF
C106 a_12322_101.n10 GND 0.08fF
C107 a_12322_101.n11 GND 0.08fF
C108 a_12322_101.t1 GND 0.23fF
C109 a_12322_101.n12 GND 0.01fF
C110 Q.n0 GND 0.58fF
C111 Q.n1 GND 0.36fF
C112 Q.n2 GND 0.66fF
C113 Q.n3 GND 0.01fF
C114 a_4569_1050.n0 GND 0.57fF
C115 a_4569_1050.n1 GND 0.44fF
C116 a_4569_1050.n2 GND 1.38fF
C117 a_4569_1050.n3 GND 0.44fF
C118 a_4569_1050.n4 GND 0.63fF
C119 a_4569_1050.n5 GND 2.09fF
C120 a_4569_1050.n6 GND 0.06fF
C121 a_4569_1050.n7 GND 0.08fF
C122 a_4569_1050.n8 GND 0.05fF
C123 a_4569_1050.n9 GND 0.37fF
C124 a_4569_1050.n10 GND 0.82fF
C125 a_4569_1050.n11 GND 0.61fF
C126 a_4569_1050.n12 GND 0.72fF
C127 a_4569_1050.n13 GND 0.69fF
C128 a_4569_1050.n14 GND 0.57fF
C129 a_1074_101.n0 GND 0.05fF
C130 a_1074_101.n1 GND 0.12fF
C131 a_1074_101.n2 GND 0.04fF
C132 a_1074_101.n3 GND 0.17fF
C133 a_8030_101.n0 GND 0.02fF
C134 a_8030_101.n1 GND 0.09fF
C135 a_8030_101.n2 GND 0.08fF
C136 a_8030_101.n3 GND 0.03fF
C137 a_8030_101.n4 GND 0.01fF
C138 a_8030_101.n5 GND 0.04fF
C139 a_8030_101.n6 GND 0.04fF
C140 a_8030_101.n7 GND 0.02fF
C141 a_8030_101.n8 GND 0.05fF
C142 a_8030_101.n9 GND 0.15fF
C143 a_8030_101.n10 GND 0.08fF
C144 a_8030_101.n11 GND 0.08fF
C145 a_8030_101.t1 GND 0.23fF
C146 a_8030_101.n12 GND 0.01fF
C147 a_599_989.n0 GND 0.34fF
C148 a_599_989.n1 GND 0.49fF
C149 a_599_989.n2 GND 0.34fF
C150 a_599_989.t6 GND 0.55fF
C151 a_599_989.n3 GND 0.57fF
C152 a_599_989.n4 GND 0.89fF
C153 a_599_989.n5 GND 0.04fF
C154 a_599_989.n6 GND 0.06fF
C155 a_599_989.n7 GND 0.04fF
C156 a_599_989.n8 GND 0.23fF
C157 a_599_989.n9 GND 0.52fF
C158 a_599_989.n10 GND 0.52fF
C159 a_599_989.n11 GND 0.60fF
C160 a_599_989.n12 GND 0.40fF
C161 a_8675_103.n0 GND 0.08fF
C162 a_8675_103.n1 GND 0.07fF
C163 a_8675_103.n2 GND 0.04fF
C164 a_8675_103.n3 GND 0.06fF
C165 a_8675_103.n4 GND 0.11fF
C166 a_8675_103.n5 GND 0.04fF
C167 a_8675_103.n7 GND 0.08fF
C168 a_4439_187.n0 GND 0.65fF
C169 a_4439_187.n1 GND 0.47fF
C170 a_4439_187.t9 GND 0.98fF
C171 a_4439_187.n2 GND 1.08fF
C172 a_4439_187.n3 GND 0.47fF
C173 a_4439_187.t7 GND 0.98fF
C174 a_4439_187.n4 GND 0.66fF
C175 a_4439_187.n5 GND 0.48fF
C176 a_4439_187.n6 GND 1.55fF
C177 a_4439_187.n7 GND 2.34fF
C178 a_4439_187.n8 GND 1.85fF
C179 a_4439_187.n9 GND 0.67fF
C180 a_4439_187.n10 GND 0.88fF
C181 a_4439_187.n11 GND 0.88fF
C182 a_4439_187.n12 GND 0.84fF
C183 a_10429_1050.n0 GND 0.42fF
C184 a_10429_1050.n1 GND 0.36fF
C185 a_10429_1050.n2 GND 0.67fF
C186 a_10429_1050.n3 GND 0.37fF
C187 a_10429_1050.n4 GND 0.76fF
C188 a_10429_1050.n5 GND 0.64fF
C189 a_10429_1050.n6 GND 0.54fF
C190 a_10324_101.n0 GND 0.08fF
C191 a_10324_101.n1 GND 0.02fF
C192 a_10324_101.n2 GND 0.02fF
C193 a_10324_101.n3 GND 0.09fF
C194 a_10324_101.n4 GND 0.08fF
C195 a_10324_101.n5 GND 0.03fF
C196 a_10324_101.n6 GND 0.05fF
C197 a_3738_101.n0 GND 0.05fF
C198 a_3738_101.n1 GND 0.12fF
C199 a_3738_101.n2 GND 0.04fF
C200 a_3738_101.n3 GND 0.17fF
C201 a_7364_101.n0 GND 0.02fF
C202 a_7364_101.n1 GND 0.09fF
C203 a_7364_101.n2 GND 0.08fF
C204 a_7364_101.n3 GND 0.03fF
C205 a_7364_101.n4 GND 0.01fF
C206 a_7364_101.n5 GND 0.04fF
C207 a_7364_101.n6 GND 0.04fF
C208 a_7364_101.n7 GND 0.02fF
C209 a_7364_101.n8 GND 0.05fF
C210 a_7364_101.n9 GND 0.15fF
C211 a_7364_101.n10 GND 0.08fF
C212 a_7364_101.n11 GND 0.08fF
C213 a_7364_101.t1 GND 0.23fF
C214 a_7364_101.n12 GND 0.01fF
C215 a_13757_1051.n0 GND 0.29fF
C216 a_13757_1051.n1 GND 0.28fF
C217 a_13757_1051.n2 GND 0.37fF
C218 a_13757_1051.n3 GND 0.71fF
C219 a_13757_1051.n4 GND 0.27fF
C220 a_13757_1051.n5 GND 0.46fF
C221 a_14320_101.n0 GND 0.06fF
C222 a_14320_101.n1 GND 0.13fF
C223 a_14320_101.n2 GND 0.04fF
C224 a_14320_101.n3 GND 0.19fF
C225 a_6032_101.n0 GND 0.05fF
C226 a_6032_101.n1 GND 0.12fF
C227 a_6032_101.n2 GND 0.04fF
C228 a_6032_101.n3 GND 0.17fF
C229 a_7469_1050.n0 GND 0.31fF
C230 a_7469_1050.n1 GND 0.63fF
C231 a_7469_1050.n2 GND 0.04fF
C232 a_7469_1050.n3 GND 0.06fF
C233 a_7469_1050.n4 GND 0.04fF
C234 a_7469_1050.n5 GND 0.26fF
C235 a_7469_1050.n6 GND 0.69fF
C236 a_7469_1050.n7 GND 0.51fF
C237 a_7469_1050.n8 GND 0.56fF
C238 a_7469_1050.n9 GND 0.40fF
C239 a_4891_989.n0 GND 0.42fF
C240 a_4891_989.n1 GND 0.60fF
C241 a_4891_989.n2 GND 0.42fF
C242 a_4891_989.t7 GND 0.67fF
C243 a_4891_989.n3 GND 0.70fF
C244 a_4891_989.n4 GND 1.09fF
C245 a_4891_989.n5 GND 0.05fF
C246 a_4891_989.n6 GND 0.07fF
C247 a_4891_989.n7 GND 0.04fF
C248 a_4891_989.n8 GND 0.29fF
C249 a_4891_989.n9 GND 0.63fF
C250 a_4891_989.n10 GND 0.63fF
C251 a_4891_989.n11 GND 0.74fF
C252 a_4891_989.n12 GND 0.49fF
C253 a_3072_101.n0 GND 0.02fF
C254 a_3072_101.n1 GND 0.09fF
C255 a_3072_101.n2 GND 0.08fF
C256 a_3072_101.n3 GND 0.03fF
C257 a_3072_101.n4 GND 0.01fF
C258 a_3072_101.n5 GND 0.04fF
C259 a_3072_101.n6 GND 0.04fF
C260 a_3072_101.n7 GND 0.02fF
C261 a_3072_101.n8 GND 0.05fF
C262 a_3072_101.n9 GND 0.15fF
C263 a_3072_101.n10 GND 0.08fF
C264 a_3072_101.n11 GND 0.08fF
C265 a_3072_101.t1 GND 0.23fF
C266 a_3072_101.n12 GND 0.01fF
C267 a_12988_101.n0 GND 0.02fF
C268 a_12988_101.n1 GND 0.09fF
C269 a_12988_101.n2 GND 0.07fF
C270 a_12988_101.n3 GND 0.03fF
C271 a_12988_101.n4 GND 0.01fF
C272 a_12988_101.n5 GND 0.03fF
C273 a_12988_101.n6 GND 0.04fF
C274 a_12988_101.n7 GND 0.02fF
C275 a_12988_101.n8 GND 0.04fF
C276 a_12988_101.n9 GND 0.08fF
C277 a_12988_101.n10 GND 0.04fF
C278 a_12988_101.n11 GND 0.12fF
C279 a_12988_101.n12 GND 0.14fF
C280 a_12988_101.t1 GND 0.16fF
C281 a_12988_101.n13 GND 0.01fF
C282 a_7595_411.n0 GND 0.49fF
C283 a_7595_411.n1 GND 0.63fF
C284 a_7595_411.n2 GND 0.86fF
C285 a_7595_411.n3 GND 0.35fF
C286 a_7595_411.n4 GND 0.37fF
C287 a_7595_411.t10 GND 0.74fF
C288 a_7595_411.n5 GND 1.27fF
C289 a_7595_411.n6 GND 1.00fF
C290 a_7595_411.t5 GND 0.60fF
C291 a_7595_411.n7 GND 2.36fF
C292 a_7595_411.n8 GND 0.50fF
C293 a_7595_411.t7 GND 0.60fF
C294 a_7595_411.n9 GND 0.67fF
C295 a_7595_411.n10 GND 3.74fF
C296 a_7595_411.n11 GND 0.63fF
C297 a_7595_411.n12 GND 0.11fF
C298 a_7595_411.n13 GND 0.17fF
C299 a_7595_411.n14 GND 0.06fF
C300 a_6698_101.n0 GND 0.02fF
C301 a_6698_101.n1 GND 0.09fF
C302 a_6698_101.n2 GND 0.08fF
C303 a_6698_101.n3 GND 0.03fF
C304 a_6698_101.n4 GND 0.01fF
C305 a_6698_101.n5 GND 0.04fF
C306 a_6698_101.n6 GND 0.04fF
C307 a_6698_101.n7 GND 0.02fF
C308 a_6698_101.n8 GND 0.05fF
C309 a_6698_101.n9 GND 0.15fF
C310 a_6698_101.n10 GND 0.08fF
C311 a_6698_101.n11 GND 0.08fF
C312 a_6698_101.t1 GND 0.23fF
C313 a_6698_101.n12 GND 0.01fF
C314 a_6137_1050.n0 GND 0.04fF
C315 a_6137_1050.n1 GND 0.42fF
C316 a_6137_1050.n2 GND 0.54fF
C317 a_6137_1050.n3 GND 0.64fF
C318 a_6137_1050.n4 GND 0.36fF
C319 a_6137_1050.n5 GND 0.67fF
C320 a_6137_1050.n6 GND 0.74fF
C321 a_6137_1050.n7 GND 0.04fF
C322 a_6137_1050.n8 GND 0.25fF
C323 a_6137_1050.n9 GND 0.06fF
C324 a_9183_989.n0 GND 0.43fF
C325 a_9183_989.n1 GND 0.61fF
C326 a_9183_989.n2 GND 0.43fF
C327 a_9183_989.t9 GND 0.69fF
C328 a_9183_989.n3 GND 0.72fF
C329 a_9183_989.n4 GND 1.11fF
C330 a_9183_989.n5 GND 0.05fF
C331 a_9183_989.n6 GND 0.07fF
C332 a_9183_989.n7 GND 0.04fF
C333 a_9183_989.n8 GND 0.29fF
C334 a_9183_989.n9 GND 0.65fF
C335 a_9183_989.n10 GND 0.64fF
C336 a_9183_989.n11 GND 0.76fF
C337 a_9183_989.n12 GND 0.50fF
C338 a_11887_411.n0 GND 0.37fF
C339 a_11887_411.n1 GND 0.24fF
C340 a_11887_411.n2 GND 0.75fF
C341 a_11887_411.n3 GND 0.24fF
C342 a_11887_411.n4 GND 0.49fF
C343 a_11887_411.n5 GND 0.39fF
C344 a_11887_411.n6 GND 0.29fF
C345 a_11887_411.t11 GND 0.54fF
C346 a_11887_411.n7 GND 0.52fF
C347 a_11887_411.n8 GND 0.78fF
C348 a_11887_411.n9 GND 0.04fF
C349 a_11887_411.n10 GND 0.05fF
C350 a_11887_411.n11 GND 0.03fF
C351 a_11887_411.n12 GND 0.25fF
C352 a_11887_411.n13 GND 0.48fF
C353 a_11887_411.n14 GND 0.53fF
C354 a_11887_411.n15 GND 0.48fF
C355 a_11761_1050.n0 GND 0.37fF
C356 a_11761_1050.n1 GND 0.24fF
C357 a_11761_1050.n2 GND 0.65fF
C358 a_11761_1050.n3 GND 0.40fF
C359 a_11761_1050.n4 GND 0.61fF
C360 a_11761_1050.n5 GND 0.46fF
C361 a_11761_1050.n6 GND 0.47fF
C362 a_13268_209.n0 GND 0.26fF
C363 a_13268_209.n1 GND 0.34fF
C364 a_13268_209.n2 GND 0.41fF
C365 a_13268_209.n3 GND 0.24fF
C366 a_13268_209.n4 GND 0.47fF
C367 a_13268_209.n5 GND 0.43fF
C368 a_13268_209.n6 GND 0.03fF
C369 a_13268_209.n7 GND 0.04fF
C370 a_13268_209.n8 GND 0.05fF
C371 a_13268_209.n9 GND 0.03fF
C372 a_13268_209.n10 GND 0.04fF
C373 a_13268_209.n11 GND 0.06fF
C374 a_13268_209.n12 GND 0.96fF
C375 a_13268_209.n13 GND 0.33fF
C376 a_13268_209.n14 GND 0.06fF
C377 a_13268_209.n15 GND 0.03fF
C378 a_13268_209.n16 GND 0.04fF
C379 a_13654_101.n0 GND 0.02fF
C380 a_13654_101.n1 GND 0.13fF
C381 a_13654_101.n2 GND 0.15fF
C382 a_13654_101.n3 GND 0.16fF
C383 a_3303_411.n0 GND 0.55fF
C384 a_3303_411.n1 GND 0.67fF
C385 a_3303_411.n2 GND 0.93fF
C386 a_3303_411.t5 GND 0.66fF
C387 a_3303_411.n3 GND 0.56fF
C388 a_3303_411.n4 GND 5.97fF
C389 a_3303_411.n5 GND 0.51fF
C390 a_3303_411.t10 GND 0.77fF
C391 a_3303_411.n6 GND 0.82fF
C392 a_3303_411.n7 GND 7.69fF
C393 a_3303_411.n8 GND 0.06fF
C394 a_3303_411.n9 GND 0.08fF
C395 a_3303_411.n10 GND 0.05fF
C396 a_3303_411.n11 GND 0.30fF
C397 a_3303_411.n12 GND 0.75fF
C398 a_3303_411.n13 GND 0.75fF
C399 a_3303_411.n14 GND 0.93fF
C400 a_3303_411.n15 GND 0.59fF
C401 a_147_187.n0 GND 0.60fF
C402 a_147_187.n1 GND 0.44fF
C403 a_147_187.t5 GND 0.91fF
C404 a_147_187.n2 GND 0.99fF
C405 a_147_187.n3 GND 0.44fF
C406 a_147_187.t12 GND 0.91fF
C407 a_147_187.n4 GND 0.61fF
C408 a_147_187.n5 GND 0.45fF
C409 a_147_187.n6 GND 1.43fF
C410 a_147_187.n7 GND 2.16fF
C411 a_147_187.n8 GND 1.71fF
C412 a_147_187.n9 GND 0.62fF
C413 a_147_187.n10 GND 0.81fF
C414 a_147_187.n11 GND 0.81fF
C415 a_147_187.n12 GND 0.77fF
C416 a_1845_1050.n0 GND 0.38fF
C417 a_1845_1050.n1 GND 0.49fF
C418 a_1845_1050.n2 GND 0.57fF
C419 a_1845_1050.n3 GND 0.33fF
C420 a_1845_1050.n4 GND 0.60fF
C421 a_1845_1050.n5 GND 0.67fF
C422 a_1845_1050.n6 GND 0.08fF
C423 a_1845_1050.n7 GND 0.22fF
C424 a_1845_1050.n8 GND 0.04fF
C425 a_3177_1050.n0 GND 0.38fF
C426 a_3177_1050.n1 GND 0.30fF
C427 a_3177_1050.n2 GND 0.61fF
C428 a_3177_1050.n3 GND 0.36fF
C429 a_3177_1050.n4 GND 0.69fF
C430 a_3177_1050.n5 GND 0.55fF
C431 a_3177_1050.n6 GND 0.49fF
C432 a_277_1050.n0 GND 0.52fF
C433 a_277_1050.n1 GND 0.52fF
C434 a_277_1050.n2 GND 0.66fF
C435 a_277_1050.n3 GND 0.62fF
C436 a_277_1050.n4 GND 0.55fF
C437 a_277_1050.n5 GND 0.40fF
C438 a_277_1050.n6 GND 1.25fF
C439 a_277_1050.n7 GND 0.40fF
C440 a_277_1050.n8 GND 0.57fF
C441 a_277_1050.n9 GND 1.90fF
C442 a_277_1050.n10 GND 0.75fF
C443 a_277_1050.n11 GND 0.11fF
C444 a_277_1050.n12 GND 0.33fF
C445 a_277_1050.n13 GND 0.06fF
C446 VDD.n1 GND 0.03fF
C447 VDD.n2 GND 0.10fF
C448 VDD.n3 GND 0.03fF
C449 VDD.n4 GND 0.02fF
C450 VDD.n5 GND 0.06fF
C451 VDD.n6 GND 0.02fF
C452 VDD.n7 GND 0.02fF
C453 VDD.n8 GND 0.02fF
C454 VDD.n9 GND 0.02fF
C455 VDD.n10 GND 0.02fF
C456 VDD.n11 GND 0.02fF
C457 VDD.n12 GND 0.02fF
C458 VDD.n13 GND 0.02fF
C459 VDD.n14 GND 0.04fF
C460 VDD.n15 GND 0.01fF
C461 VDD.n20 GND 0.48fF
C462 VDD.n21 GND 0.29fF
C463 VDD.n22 GND 0.02fF
C464 VDD.n23 GND 0.03fF
C465 VDD.n24 GND 0.07fF
C466 VDD.n25 GND 0.21fF
C467 VDD.n26 GND 0.01fF
C468 VDD.n27 GND 0.01fF
C469 VDD.n28 GND 0.07fF
C470 VDD.n29 GND 0.18fF
C471 VDD.n30 GND 0.01fF
C472 VDD.n31 GND 0.03fF
C473 VDD.n32 GND 0.03fF
C474 VDD.n33 GND 0.21fF
C475 VDD.n34 GND 0.01fF
C476 VDD.n35 GND 0.07fF
C477 VDD.n36 GND 0.01fF
C478 VDD.n37 GND 0.02fF
C479 VDD.n38 GND 0.29fF
C480 VDD.n39 GND 0.01fF
C481 VDD.n40 GND 0.02fF
C482 VDD.n41 GND 0.04fF
C483 VDD.n42 GND 0.06fF
C484 VDD.n43 GND 0.02fF
C485 VDD.n44 GND 0.02fF
C486 VDD.n45 GND 0.02fF
C487 VDD.n46 GND 0.02fF
C488 VDD.n47 GND 0.02fF
C489 VDD.n48 GND 0.02fF
C490 VDD.n49 GND 0.02fF
C491 VDD.n50 GND 0.02fF
C492 VDD.n51 GND 0.02fF
C493 VDD.n52 GND 0.02fF
C494 VDD.n53 GND 0.02fF
C495 VDD.n54 GND 0.03fF
C496 VDD.n55 GND 0.02fF
C497 VDD.n56 GND 0.19fF
C498 VDD.n57 GND 0.02fF
C499 VDD.n58 GND 0.02fF
C500 VDD.n60 GND 0.02fF
C501 VDD.n64 GND 0.29fF
C502 VDD.n65 GND 0.29fF
C503 VDD.n66 GND 0.01fF
C504 VDD.n67 GND 0.02fF
C505 VDD.n68 GND 0.04fF
C506 VDD.n69 GND 0.25fF
C507 VDD.n70 GND 0.01fF
C508 VDD.n71 GND 0.02fF
C509 VDD.n72 GND 0.02fF
C510 VDD.n73 GND 0.18fF
C511 VDD.n74 GND 0.01fF
C512 VDD.n75 GND 0.02fF
C513 VDD.n76 GND 0.02fF
C514 VDD.n77 GND 0.01fF
C515 VDD.n78 GND 0.03fF
C516 VDD.n79 GND 0.03fF
C517 VDD.n80 GND 0.15fF
C518 VDD.n81 GND 0.01fF
C519 VDD.n82 GND 0.03fF
C520 VDD.n83 GND 0.03fF
C521 VDD.n84 GND 0.17fF
C522 VDD.n85 GND 0.01fF
C523 VDD.n86 GND 0.02fF
C524 VDD.n87 GND 0.02fF
C525 VDD.n88 GND 0.26fF
C526 VDD.n89 GND 0.01fF
C527 VDD.n90 GND 0.02fF
C528 VDD.n91 GND 0.02fF
C529 VDD.n92 GND 0.29fF
C530 VDD.n93 GND 0.01fF
C531 VDD.n94 GND 0.02fF
C532 VDD.n95 GND 0.04fF
C533 VDD.n96 GND 0.22fF
C534 VDD.n97 GND 0.02fF
C535 VDD.n98 GND 0.02fF
C536 VDD.n99 GND 0.02fF
C537 VDD.n100 GND 0.06fF
C538 VDD.n101 GND 0.02fF
C539 VDD.n102 GND 0.02fF
C540 VDD.n103 GND 0.02fF
C541 VDD.n104 GND 0.02fF
C542 VDD.n105 GND 0.02fF
C543 VDD.n106 GND 0.02fF
C544 VDD.n107 GND 0.02fF
C545 VDD.n108 GND 0.02fF
C546 VDD.n109 GND 0.02fF
C547 VDD.n110 GND 0.02fF
C548 VDD.n111 GND 0.03fF
C549 VDD.n112 GND 0.02fF
C550 VDD.n113 GND 0.02fF
C551 VDD.n117 GND 0.29fF
C552 VDD.n118 GND 0.29fF
C553 VDD.n119 GND 0.01fF
C554 VDD.n120 GND 0.02fF
C555 VDD.n121 GND 0.04fF
C556 VDD.n122 GND 0.26fF
C557 VDD.n123 GND 0.01fF
C558 VDD.n124 GND 0.02fF
C559 VDD.n125 GND 0.02fF
C560 VDD.n126 GND 0.17fF
C561 VDD.n127 GND 0.01fF
C562 VDD.n128 GND 0.02fF
C563 VDD.n129 GND 0.02fF
C564 VDD.n130 GND 0.15fF
C565 VDD.n131 GND 0.01fF
C566 VDD.n132 GND 0.03fF
C567 VDD.n133 GND 0.03fF
C568 VDD.n134 GND 0.01fF
C569 VDD.n135 GND 0.03fF
C570 VDD.n136 GND 0.03fF
C571 VDD.n137 GND 0.18fF
C572 VDD.n138 GND 0.01fF
C573 VDD.n139 GND 0.02fF
C574 VDD.n140 GND 0.02fF
C575 VDD.n141 GND 0.25fF
C576 VDD.n142 GND 0.01fF
C577 VDD.n143 GND 0.02fF
C578 VDD.n144 GND 0.02fF
C579 VDD.n145 GND 0.29fF
C580 VDD.n146 GND 0.01fF
C581 VDD.n147 GND 0.02fF
C582 VDD.n148 GND 0.04fF
C583 VDD.n149 GND 0.22fF
C584 VDD.n150 GND 0.02fF
C585 VDD.n151 GND 0.02fF
C586 VDD.n152 GND 0.02fF
C587 VDD.n153 GND 0.06fF
C588 VDD.n154 GND 0.02fF
C589 VDD.n155 GND 0.02fF
C590 VDD.n156 GND 0.02fF
C591 VDD.n157 GND 0.02fF
C592 VDD.n158 GND 0.02fF
C593 VDD.n159 GND 0.02fF
C594 VDD.n160 GND 0.02fF
C595 VDD.n161 GND 0.02fF
C596 VDD.n162 GND 0.02fF
C597 VDD.n163 GND 0.02fF
C598 VDD.n164 GND 0.03fF
C599 VDD.n165 GND 0.02fF
C600 VDD.n166 GND 0.02fF
C601 VDD.n170 GND 0.29fF
C602 VDD.n171 GND 0.29fF
C603 VDD.n172 GND 0.01fF
C604 VDD.n173 GND 0.02fF
C605 VDD.n174 GND 0.04fF
C606 VDD.n175 GND 0.07fF
C607 VDD.n176 GND 0.25fF
C608 VDD.n177 GND 0.01fF
C609 VDD.n178 GND 0.01fF
C610 VDD.n179 GND 0.02fF
C611 VDD.n180 GND 0.18fF
C612 VDD.n181 GND 0.01fF
C613 VDD.n182 GND 0.02fF
C614 VDD.n183 GND 0.02fF
C615 VDD.n184 GND 0.08fF
C616 VDD.n185 GND 0.05fF
C617 VDD.n186 GND 0.01fF
C618 VDD.n187 GND 0.02fF
C619 VDD.n188 GND 0.03fF
C620 VDD.n189 GND 0.15fF
C621 VDD.n190 GND 0.01fF
C622 VDD.n191 GND 0.02fF
C623 VDD.n192 GND 0.03fF
C624 VDD.n193 GND 0.17fF
C625 VDD.n194 GND 0.01fF
C626 VDD.n195 GND 0.02fF
C627 VDD.n196 GND 0.02fF
C628 VDD.n197 GND 0.07fF
C629 VDD.n198 GND 0.26fF
C630 VDD.n199 GND 0.01fF
C631 VDD.n200 GND 0.01fF
C632 VDD.n201 GND 0.02fF
C633 VDD.n202 GND 0.29fF
C634 VDD.n203 GND 0.01fF
C635 VDD.n204 GND 0.02fF
C636 VDD.n205 GND 0.04fF
C637 VDD.n206 GND 0.22fF
C638 VDD.n207 GND 0.02fF
C639 VDD.n208 GND 0.02fF
C640 VDD.n209 GND 0.02fF
C641 VDD.n210 GND 0.06fF
C642 VDD.n211 GND 0.02fF
C643 VDD.n212 GND 0.02fF
C644 VDD.n213 GND 0.02fF
C645 VDD.n214 GND 0.02fF
C646 VDD.n215 GND 0.02fF
C647 VDD.n216 GND 0.02fF
C648 VDD.n217 GND 0.02fF
C649 VDD.n218 GND 0.02fF
C650 VDD.n219 GND 0.02fF
C651 VDD.n220 GND 0.02fF
C652 VDD.n221 GND 0.03fF
C653 VDD.n222 GND 0.02fF
C654 VDD.n223 GND 0.02fF
C655 VDD.n227 GND 0.29fF
C656 VDD.n228 GND 0.29fF
C657 VDD.n229 GND 0.01fF
C658 VDD.n230 GND 0.02fF
C659 VDD.n231 GND 0.04fF
C660 VDD.n232 GND 0.06fF
C661 VDD.n233 GND 0.25fF
C662 VDD.n234 GND 0.01fF
C663 VDD.n235 GND 0.01fF
C664 VDD.n236 GND 0.02fF
C665 VDD.n237 GND 0.18fF
C666 VDD.n238 GND 0.01fF
C667 VDD.n239 GND 0.02fF
C668 VDD.n240 GND 0.02fF
C669 VDD.n241 GND 0.08fF
C670 VDD.n242 GND 0.05fF
C671 VDD.n243 GND 0.01fF
C672 VDD.n244 GND 0.02fF
C673 VDD.n245 GND 0.03fF
C674 VDD.n246 GND 0.15fF
C675 VDD.n247 GND 0.01fF
C676 VDD.n248 GND 0.02fF
C677 VDD.n249 GND 0.03fF
C678 VDD.n250 GND 0.17fF
C679 VDD.n251 GND 0.01fF
C680 VDD.n252 GND 0.02fF
C681 VDD.n253 GND 0.02fF
C682 VDD.n254 GND 0.07fF
C683 VDD.n255 GND 0.26fF
C684 VDD.n256 GND 0.01fF
C685 VDD.n257 GND 0.01fF
C686 VDD.n258 GND 0.02fF
C687 VDD.n259 GND 0.29fF
C688 VDD.n260 GND 0.01fF
C689 VDD.n261 GND 0.02fF
C690 VDD.n262 GND 0.04fF
C691 VDD.n263 GND 0.22fF
C692 VDD.n264 GND 0.02fF
C693 VDD.n265 GND 0.02fF
C694 VDD.n266 GND 0.02fF
C695 VDD.n267 GND 0.06fF
C696 VDD.n268 GND 0.02fF
C697 VDD.n269 GND 0.02fF
C698 VDD.n270 GND 0.02fF
C699 VDD.n271 GND 0.02fF
C700 VDD.n272 GND 0.02fF
C701 VDD.n273 GND 0.02fF
C702 VDD.n274 GND 0.02fF
C703 VDD.n275 GND 0.02fF
C704 VDD.n276 GND 0.02fF
C705 VDD.n277 GND 0.02fF
C706 VDD.n278 GND 0.03fF
C707 VDD.n279 GND 0.02fF
C708 VDD.n280 GND 0.02fF
C709 VDD.n284 GND 0.29fF
C710 VDD.n285 GND 0.29fF
C711 VDD.n286 GND 0.01fF
C712 VDD.n287 GND 0.02fF
C713 VDD.n288 GND 0.04fF
C714 VDD.n289 GND 0.06fF
C715 VDD.n290 GND 0.25fF
C716 VDD.n291 GND 0.01fF
C717 VDD.n292 GND 0.01fF
C718 VDD.n293 GND 0.02fF
C719 VDD.n294 GND 0.18fF
C720 VDD.n295 GND 0.01fF
C721 VDD.n296 GND 0.02fF
C722 VDD.n297 GND 0.02fF
C723 VDD.n298 GND 0.08fF
C724 VDD.n299 GND 0.05fF
C725 VDD.n300 GND 0.01fF
C726 VDD.n301 GND 0.02fF
C727 VDD.n302 GND 0.03fF
C728 VDD.n303 GND 0.15fF
C729 VDD.n304 GND 0.01fF
C730 VDD.n305 GND 0.02fF
C731 VDD.n306 GND 0.03fF
C732 VDD.n307 GND 0.17fF
C733 VDD.n308 GND 0.01fF
C734 VDD.n309 GND 0.02fF
C735 VDD.n310 GND 0.02fF
C736 VDD.n311 GND 0.07fF
C737 VDD.n312 GND 0.26fF
C738 VDD.n313 GND 0.01fF
C739 VDD.n314 GND 0.01fF
C740 VDD.n315 GND 0.02fF
C741 VDD.n316 GND 0.29fF
C742 VDD.n317 GND 0.01fF
C743 VDD.n318 GND 0.02fF
C744 VDD.n319 GND 0.04fF
C745 VDD.n320 GND 0.22fF
C746 VDD.n321 GND 0.02fF
C747 VDD.n322 GND 0.02fF
C748 VDD.n323 GND 0.02fF
C749 VDD.n324 GND 0.06fF
C750 VDD.n325 GND 0.02fF
C751 VDD.n326 GND 0.02fF
C752 VDD.n327 GND 0.02fF
C753 VDD.n328 GND 0.02fF
C754 VDD.n329 GND 0.02fF
C755 VDD.n330 GND 0.02fF
C756 VDD.n331 GND 0.02fF
C757 VDD.n332 GND 0.02fF
C758 VDD.n333 GND 0.02fF
C759 VDD.n334 GND 0.02fF
C760 VDD.n335 GND 0.03fF
C761 VDD.n336 GND 0.02fF
C762 VDD.n337 GND 0.02fF
C763 VDD.n341 GND 0.29fF
C764 VDD.n342 GND 0.29fF
C765 VDD.n343 GND 0.01fF
C766 VDD.n344 GND 0.02fF
C767 VDD.n345 GND 0.04fF
C768 VDD.n346 GND 0.06fF
C769 VDD.n347 GND 0.25fF
C770 VDD.n348 GND 0.01fF
C771 VDD.n349 GND 0.01fF
C772 VDD.n350 GND 0.02fF
C773 VDD.n351 GND 0.18fF
C774 VDD.n352 GND 0.01fF
C775 VDD.n353 GND 0.02fF
C776 VDD.n354 GND 0.02fF
C777 VDD.n355 GND 0.08fF
C778 VDD.n356 GND 0.05fF
C779 VDD.n357 GND 0.01fF
C780 VDD.n358 GND 0.02fF
C781 VDD.n359 GND 0.03fF
C782 VDD.n360 GND 0.15fF
C783 VDD.n361 GND 0.01fF
C784 VDD.n362 GND 0.02fF
C785 VDD.n363 GND 0.03fF
C786 VDD.n364 GND 0.17fF
C787 VDD.n365 GND 0.01fF
C788 VDD.n366 GND 0.02fF
C789 VDD.n367 GND 0.02fF
C790 VDD.n368 GND 0.07fF
C791 VDD.n369 GND 0.26fF
C792 VDD.n370 GND 0.01fF
C793 VDD.n371 GND 0.01fF
C794 VDD.n372 GND 0.02fF
C795 VDD.n373 GND 0.29fF
C796 VDD.n374 GND 0.01fF
C797 VDD.n375 GND 0.02fF
C798 VDD.n376 GND 0.04fF
C799 VDD.n377 GND 0.22fF
C800 VDD.n378 GND 0.02fF
C801 VDD.n379 GND 0.02fF
C802 VDD.n380 GND 0.02fF
C803 VDD.n381 GND 0.06fF
C804 VDD.n382 GND 0.02fF
C805 VDD.n383 GND 0.02fF
C806 VDD.n384 GND 0.02fF
C807 VDD.n385 GND 0.02fF
C808 VDD.n386 GND 0.02fF
C809 VDD.n387 GND 0.02fF
C810 VDD.n388 GND 0.02fF
C811 VDD.n389 GND 0.02fF
C812 VDD.n390 GND 0.02fF
C813 VDD.n391 GND 0.02fF
C814 VDD.n392 GND 0.03fF
C815 VDD.n393 GND 0.02fF
C816 VDD.n394 GND 0.02fF
C817 VDD.n398 GND 0.29fF
C818 VDD.n399 GND 0.29fF
C819 VDD.n400 GND 0.01fF
C820 VDD.n401 GND 0.02fF
C821 VDD.n402 GND 0.04fF
C822 VDD.n403 GND 0.06fF
C823 VDD.n404 GND 0.25fF
C824 VDD.n405 GND 0.01fF
C825 VDD.n406 GND 0.01fF
C826 VDD.n407 GND 0.02fF
C827 VDD.n408 GND 0.18fF
C828 VDD.n409 GND 0.01fF
C829 VDD.n410 GND 0.02fF
C830 VDD.n411 GND 0.02fF
C831 VDD.n412 GND 0.08fF
C832 VDD.n413 GND 0.05fF
C833 VDD.n414 GND 0.01fF
C834 VDD.n415 GND 0.02fF
C835 VDD.n416 GND 0.03fF
C836 VDD.n417 GND 0.15fF
C837 VDD.n418 GND 0.01fF
C838 VDD.n419 GND 0.02fF
C839 VDD.n420 GND 0.03fF
C840 VDD.n421 GND 0.17fF
C841 VDD.n422 GND 0.01fF
C842 VDD.n423 GND 0.02fF
C843 VDD.n424 GND 0.02fF
C844 VDD.n425 GND 0.07fF
C845 VDD.n426 GND 0.26fF
C846 VDD.n427 GND 0.01fF
C847 VDD.n428 GND 0.01fF
C848 VDD.n429 GND 0.02fF
C849 VDD.n430 GND 0.29fF
C850 VDD.n431 GND 0.01fF
C851 VDD.n432 GND 0.02fF
C852 VDD.n433 GND 0.04fF
C853 VDD.n434 GND 0.22fF
C854 VDD.n435 GND 0.02fF
C855 VDD.n436 GND 0.02fF
C856 VDD.n437 GND 0.02fF
C857 VDD.n438 GND 0.06fF
C858 VDD.n439 GND 0.02fF
C859 VDD.n440 GND 0.02fF
C860 VDD.n441 GND 0.02fF
C861 VDD.n442 GND 0.02fF
C862 VDD.n443 GND 0.02fF
C863 VDD.n444 GND 0.02fF
C864 VDD.n445 GND 0.02fF
C865 VDD.n446 GND 0.02fF
C866 VDD.n447 GND 0.02fF
C867 VDD.n448 GND 0.02fF
C868 VDD.n449 GND 0.03fF
C869 VDD.n450 GND 0.02fF
C870 VDD.n451 GND 0.02fF
C871 VDD.n455 GND 0.29fF
C872 VDD.n456 GND 0.29fF
C873 VDD.n457 GND 0.01fF
C874 VDD.n458 GND 0.02fF
C875 VDD.n459 GND 0.04fF
C876 VDD.n460 GND 0.06fF
C877 VDD.n461 GND 0.25fF
C878 VDD.n462 GND 0.01fF
C879 VDD.n463 GND 0.01fF
C880 VDD.n464 GND 0.02fF
C881 VDD.n465 GND 0.18fF
C882 VDD.n466 GND 0.01fF
C883 VDD.n467 GND 0.02fF
C884 VDD.n468 GND 0.02fF
C885 VDD.n469 GND 0.08fF
C886 VDD.n470 GND 0.05fF
C887 VDD.n471 GND 0.01fF
C888 VDD.n472 GND 0.02fF
C889 VDD.n473 GND 0.03fF
C890 VDD.n474 GND 0.15fF
C891 VDD.n475 GND 0.01fF
C892 VDD.n476 GND 0.02fF
C893 VDD.n477 GND 0.03fF
C894 VDD.n478 GND 0.17fF
C895 VDD.n479 GND 0.01fF
C896 VDD.n480 GND 0.02fF
C897 VDD.n481 GND 0.02fF
C898 VDD.n482 GND 0.07fF
C899 VDD.n483 GND 0.26fF
C900 VDD.n484 GND 0.01fF
C901 VDD.n485 GND 0.01fF
C902 VDD.n486 GND 0.02fF
C903 VDD.n487 GND 0.29fF
C904 VDD.n488 GND 0.01fF
C905 VDD.n489 GND 0.02fF
C906 VDD.n490 GND 0.04fF
C907 VDD.n491 GND 0.27fF
C908 VDD.n492 GND 0.02fF
C909 VDD.n493 GND 0.02fF
C910 VDD.n494 GND 0.02fF
C911 VDD.n495 GND 0.06fF
C912 VDD.n496 GND 0.02fF
C913 VDD.n497 GND 0.02fF
C914 VDD.n498 GND 0.02fF
C915 VDD.n499 GND 0.02fF
C916 VDD.n500 GND 0.02fF
C917 VDD.n501 GND 0.02fF
C918 VDD.n502 GND 0.02fF
C919 VDD.n503 GND 0.02fF
C920 VDD.n504 GND 0.02fF
C921 VDD.n505 GND 0.02fF
C922 VDD.n506 GND 0.03fF
C923 VDD.n507 GND 0.02fF
C924 VDD.n508 GND 0.02fF
C925 VDD.n512 GND 0.29fF
C926 VDD.n513 GND 0.29fF
C927 VDD.n514 GND 0.01fF
C928 VDD.n515 GND 0.02fF
C929 VDD.n516 GND 0.04fF
C930 VDD.n517 GND 0.29fF
C931 VDD.n518 GND 0.01fF
C932 VDD.n519 GND 0.02fF
C933 VDD.n520 GND 0.02fF
C934 VDD.n521 GND 0.23fF
C935 VDD.n522 GND 0.01fF
C936 VDD.n523 GND 0.07fF
C937 VDD.n524 GND 0.02fF
C938 VDD.n525 GND 0.18fF
C939 VDD.n526 GND 0.01fF
C940 VDD.n527 GND 0.02fF
C941 VDD.n528 GND 0.02fF
C942 VDD.n529 GND 0.17fF
C943 VDD.n530 GND 0.01fF
C944 VDD.n531 GND 0.08fF
C945 VDD.n532 GND 0.05fF
C946 VDD.n533 GND 0.02fF
C947 VDD.n534 GND 0.02fF
C948 VDD.n535 GND 0.15fF
C949 VDD.n536 GND 0.02fF
C950 VDD.n537 GND 0.02fF
C951 VDD.n538 GND 0.03fF
C952 VDD.n539 GND 0.16fF
C953 VDD.n540 GND 0.02fF
C954 VDD.n541 GND 0.02fF
C955 VDD.n542 GND 0.03fF
C956 VDD.n543 GND 0.08fF
C957 VDD.n544 GND 0.05fF
C958 VDD.n545 GND 0.16fF
C959 VDD.n546 GND 0.01fF
C960 VDD.n547 GND 0.02fF
C961 VDD.n548 GND 0.02fF
C962 VDD.n549 GND 0.18fF
C963 VDD.n550 GND 0.01fF
C964 VDD.n551 GND 0.02fF
C965 VDD.n552 GND 0.02fF
C966 VDD.n553 GND 0.07fF
C967 VDD.n554 GND 0.23fF
C968 VDD.n555 GND 0.01fF
C969 VDD.n556 GND 0.01fF
C970 VDD.n557 GND 0.02fF
C971 VDD.n558 GND 0.29fF
C972 VDD.n559 GND 0.01fF
C973 VDD.n560 GND 0.02fF
C974 VDD.n561 GND 0.02fF
C975 VDD.n562 GND 0.29fF
C976 VDD.n563 GND 0.01fF
C977 VDD.n564 GND 0.02fF
C978 VDD.n565 GND 0.04fF
C979 VDD.n566 GND 0.27fF
C980 VDD.n567 GND 0.02fF
C981 VDD.n568 GND 0.02fF
C982 VDD.n569 GND 0.02fF
C983 VDD.n570 GND 0.06fF
C984 VDD.n571 GND 0.02fF
C985 VDD.n572 GND 0.02fF
C986 VDD.n573 GND 0.02fF
C987 VDD.n574 GND 0.02fF
C988 VDD.n575 GND 0.02fF
C989 VDD.n576 GND 0.02fF
C990 VDD.n577 GND 0.02fF
C991 VDD.n578 GND 0.02fF
C992 VDD.n579 GND 0.02fF
C993 VDD.n580 GND 0.02fF
C994 VDD.n581 GND 0.03fF
C995 VDD.n582 GND 0.02fF
C996 VDD.n583 GND 0.02fF
C997 VDD.n587 GND 0.29fF
C998 VDD.n588 GND 0.29fF
C999 VDD.n589 GND 0.01fF
C1000 VDD.n590 GND 0.02fF
C1001 VDD.n591 GND 0.04fF
C1002 VDD.n592 GND 0.06fF
C1003 VDD.n593 GND 0.25fF
C1004 VDD.n594 GND 0.01fF
C1005 VDD.n595 GND 0.01fF
C1006 VDD.n596 GND 0.02fF
C1007 VDD.n597 GND 0.18fF
C1008 VDD.n598 GND 0.01fF
C1009 VDD.n599 GND 0.02fF
C1010 VDD.n600 GND 0.02fF
C1011 VDD.n601 GND 0.08fF
C1012 VDD.n602 GND 0.05fF
C1013 VDD.n603 GND 0.01fF
C1014 VDD.n604 GND 0.02fF
C1015 VDD.n605 GND 0.03fF
C1016 VDD.n606 GND 0.15fF
C1017 VDD.n607 GND 0.01fF
C1018 VDD.n608 GND 0.02fF
C1019 VDD.n609 GND 0.03fF
C1020 VDD.n610 GND 0.17fF
C1021 VDD.n611 GND 0.01fF
C1022 VDD.n612 GND 0.02fF
C1023 VDD.n613 GND 0.02fF
C1024 VDD.n614 GND 0.07fF
C1025 VDD.n615 GND 0.26fF
C1026 VDD.n616 GND 0.01fF
C1027 VDD.n617 GND 0.01fF
C1028 VDD.n618 GND 0.02fF
C1029 VDD.n619 GND 0.29fF
C1030 VDD.n620 GND 0.01fF
C1031 VDD.n621 GND 0.02fF
C1032 VDD.n622 GND 0.04fF
C1033 VDD.n623 GND 0.22fF
C1034 VDD.n624 GND 0.02fF
C1035 VDD.n625 GND 0.02fF
C1036 VDD.n626 GND 0.02fF
C1037 VDD.n627 GND 0.06fF
C1038 VDD.n628 GND 0.02fF
C1039 VDD.n629 GND 0.02fF
C1040 VDD.n630 GND 0.02fF
C1041 VDD.n631 GND 0.02fF
C1042 VDD.n632 GND 0.02fF
C1043 VDD.n633 GND 0.02fF
C1044 VDD.n634 GND 0.02fF
C1045 VDD.n635 GND 0.02fF
C1046 VDD.n636 GND 0.02fF
C1047 VDD.n637 GND 0.02fF
C1048 VDD.n638 GND 0.03fF
C1049 VDD.n639 GND 0.02fF
C1050 VDD.n640 GND 0.02fF
C1051 VDD.n644 GND 0.29fF
C1052 VDD.n645 GND 0.29fF
C1053 VDD.n646 GND 0.01fF
C1054 VDD.n647 GND 0.02fF
C1055 VDD.n648 GND 0.04fF
C1056 VDD.n649 GND 0.06fF
C1057 VDD.n650 GND 0.25fF
C1058 VDD.n651 GND 0.01fF
C1059 VDD.n652 GND 0.01fF
C1060 VDD.n653 GND 0.02fF
C1061 VDD.n654 GND 0.18fF
C1062 VDD.n655 GND 0.01fF
C1063 VDD.n656 GND 0.02fF
C1064 VDD.n657 GND 0.02fF
C1065 VDD.n658 GND 0.19fF
C1066 VDD.n659 GND 0.02fF
C1067 VDD.n660 GND 0.02fF
C1068 VDD.n661 GND 0.06fF
C1069 VDD.n662 GND 0.02fF
C1070 VDD.n663 GND 0.02fF
C1071 VDD.n664 GND 0.02fF
C1072 VDD.n665 GND 0.02fF
C1073 VDD.n666 GND 0.02fF
C1074 VDD.n667 GND 0.02fF
C1075 VDD.n668 GND 0.02fF
C1076 VDD.n669 GND 0.02fF
C1077 VDD.n670 GND 0.03fF
C1078 VDD.n671 GND 0.04fF
C1079 VDD.n672 GND 0.02fF
C1080 VDD.n676 GND 0.48fF
C1081 VDD.n677 GND 0.29fF
C1082 VDD.n678 GND 0.02fF
C1083 VDD.n679 GND 0.03fF
C1084 VDD.n680 GND 0.03fF
C1085 VDD.n681 GND 0.29fF
C1086 VDD.n682 GND 0.01fF
C1087 VDD.n683 GND 0.02fF
C1088 VDD.n684 GND 0.02fF
C1089 VDD.n685 GND 0.07fF
C1090 VDD.n686 GND 0.23fF
C1091 VDD.n687 GND 0.01fF
C1092 VDD.n688 GND 0.01fF
C1093 VDD.n689 GND 0.02fF
C1094 VDD.n690 GND 0.18fF
C1095 VDD.n691 GND 0.01fF
C1096 VDD.n692 GND 0.02fF
C1097 VDD.n693 GND 0.02fF
C1098 VDD.n694 GND 0.08fF
C1099 VDD.n695 GND 0.05fF
C1100 VDD.n696 GND 0.16fF
C1101 VDD.n697 GND 0.01fF
C1102 VDD.n698 GND 0.02fF
C1103 VDD.n699 GND 0.02fF
C1104 VDD.n700 GND 0.16fF
C1105 VDD.n701 GND 0.02fF
C1106 VDD.n702 GND 0.02fF
C1107 VDD.n703 GND 0.03fF
C1108 VDD.n704 GND 0.15fF
C1109 VDD.n705 GND 0.02fF
C1110 VDD.n706 GND 0.02fF
C1111 VDD.n707 GND 0.03fF
C1112 VDD.n708 GND 0.17fF
C1113 VDD.n709 GND 0.01fF
C1114 VDD.n710 GND 0.08fF
C1115 VDD.n711 GND 0.05fF
C1116 VDD.n712 GND 0.02fF
C1117 VDD.n713 GND 0.02fF
C1118 VDD.n714 GND 0.18fF
C1119 VDD.n715 GND 0.01fF
C1120 VDD.n716 GND 0.02fF
C1121 VDD.n717 GND 0.02fF
C1122 VDD.n718 GND 0.23fF
C1123 VDD.n719 GND 0.01fF
C1124 VDD.n720 GND 0.07fF
C1125 VDD.n721 GND 0.02fF
C1126 VDD.n722 GND 0.29fF
C1127 VDD.n723 GND 0.01fF
C1128 VDD.n724 GND 0.02fF
C1129 VDD.n725 GND 0.02fF
C1130 VDD.n726 GND 0.29fF
C1131 VDD.n727 GND 0.01fF
C1132 VDD.n728 GND 0.02fF
C1133 VDD.n729 GND 0.04fF
C1134 VDD.n730 GND 0.06fF
C1135 VDD.n731 GND 0.02fF
C1136 VDD.n732 GND 0.02fF
C1137 VDD.n733 GND 0.02fF
C1138 VDD.n734 GND 0.02fF
C1139 VDD.n735 GND 0.02fF
C1140 VDD.n736 GND 0.02fF
C1141 VDD.n737 GND 0.02fF
C1142 VDD.n738 GND 0.02fF
C1143 VDD.n739 GND 0.02fF
C1144 VDD.n740 GND 0.02fF
C1145 VDD.n741 GND 0.02fF
C1146 VDD.n742 GND 0.03fF
C1147 VDD.n743 GND 0.02fF
C1148 VDD.n746 GND 0.02fF
C1149 VDD.n748 GND 0.02fF
C1150 VDD.n749 GND 0.28fF
C1151 VDD.n750 GND 0.02fF
C1152 VDD.n752 GND 0.29fF
C1153 VDD.n753 GND 0.29fF
C1154 VDD.n754 GND 0.01fF
C1155 VDD.n755 GND 0.02fF
C1156 VDD.n756 GND 0.04fF
C1157 VDD.n757 GND 0.07fF
C1158 VDD.n758 GND 0.26fF
C1159 VDD.n759 GND 0.01fF
C1160 VDD.n760 GND 0.01fF
C1161 VDD.n761 GND 0.02fF
C1162 VDD.n762 GND 0.17fF
C1163 VDD.n763 GND 0.01fF
C1164 VDD.n764 GND 0.02fF
C1165 VDD.n765 GND 0.02fF
C1166 VDD.n766 GND 0.15fF
C1167 VDD.n767 GND 0.01fF
C1168 VDD.n768 GND 0.02fF
C1169 VDD.n769 GND 0.03fF
C1170 VDD.n770 GND 0.08fF
C1171 VDD.n771 GND 0.05fF
C1172 VDD.n772 GND 0.01fF
C1173 VDD.n773 GND 0.02fF
C1174 VDD.n774 GND 0.03fF
C1175 VDD.n775 GND 0.18fF
C1176 VDD.n776 GND 0.01fF
C1177 VDD.n777 GND 0.02fF
C1178 VDD.n778 GND 0.02fF
C1179 VDD.n779 GND 0.06fF
C1180 VDD.n780 GND 0.25fF
C1181 VDD.n781 GND 0.01fF
C1182 VDD.n782 GND 0.01fF
C1183 VDD.n783 GND 0.02fF
C1184 VDD.n784 GND 0.29fF
C1185 VDD.n785 GND 0.01fF
C1186 VDD.n786 GND 0.02fF
C1187 VDD.n787 GND 0.04fF
C1188 VDD.n788 GND 0.22fF
C1189 VDD.n789 GND 0.02fF
C1190 VDD.n790 GND 0.02fF
C1191 VDD.n791 GND 0.02fF
C1192 VDD.n792 GND 0.06fF
C1193 VDD.n793 GND 0.02fF
C1194 VDD.n794 GND 0.02fF
C1195 VDD.n795 GND 0.02fF
C1196 VDD.n796 GND 0.02fF
C1197 VDD.n797 GND 0.02fF
C1198 VDD.n798 GND 0.02fF
C1199 VDD.n799 GND 0.02fF
C1200 VDD.n800 GND 0.02fF
C1201 VDD.n801 GND 0.02fF
C1202 VDD.n802 GND 0.02fF
C1203 VDD.n803 GND 0.03fF
C1204 VDD.n804 GND 0.02fF
C1205 VDD.n805 GND 0.02fF
C1206 VDD.n809 GND 0.29fF
C1207 VDD.n810 GND 0.29fF
C1208 VDD.n811 GND 0.01fF
C1209 VDD.n812 GND 0.02fF
C1210 VDD.n813 GND 0.04fF
C1211 VDD.n814 GND 0.07fF
C1212 VDD.n815 GND 0.26fF
C1213 VDD.n816 GND 0.01fF
C1214 VDD.n817 GND 0.01fF
C1215 VDD.n818 GND 0.02fF
C1216 VDD.n819 GND 0.17fF
C1217 VDD.n820 GND 0.01fF
C1218 VDD.n821 GND 0.02fF
C1219 VDD.n822 GND 0.02fF
C1220 VDD.n823 GND 0.15fF
C1221 VDD.n824 GND 0.01fF
C1222 VDD.n825 GND 0.02fF
C1223 VDD.n826 GND 0.03fF
C1224 VDD.n827 GND 0.08fF
C1225 VDD.n828 GND 0.05fF
C1226 VDD.n829 GND 0.01fF
C1227 VDD.n830 GND 0.02fF
C1228 VDD.n831 GND 0.03fF
C1229 VDD.n832 GND 0.18fF
C1230 VDD.n833 GND 0.01fF
C1231 VDD.n834 GND 0.02fF
C1232 VDD.n835 GND 0.02fF
C1233 VDD.n836 GND 0.06fF
C1234 VDD.n837 GND 0.25fF
C1235 VDD.n838 GND 0.01fF
C1236 VDD.n839 GND 0.01fF
C1237 VDD.n840 GND 0.02fF
C1238 VDD.n841 GND 0.29fF
C1239 VDD.n842 GND 0.01fF
C1240 VDD.n843 GND 0.02fF
C1241 VDD.n844 GND 0.04fF
C1242 VDD.n845 GND 0.22fF
C1243 VDD.n846 GND 0.02fF
C1244 VDD.n847 GND 0.02fF
C1245 VDD.n848 GND 0.02fF
C1246 VDD.n849 GND 0.06fF
C1247 VDD.n850 GND 0.02fF
C1248 VDD.n851 GND 0.02fF
C1249 VDD.n852 GND 0.02fF
C1250 VDD.n853 GND 0.02fF
C1251 VDD.n854 GND 0.02fF
C1252 VDD.n855 GND 0.02fF
C1253 VDD.n856 GND 0.02fF
C1254 VDD.n857 GND 0.02fF
C1255 VDD.n858 GND 0.02fF
C1256 VDD.n859 GND 0.02fF
C1257 VDD.n860 GND 0.03fF
C1258 VDD.n861 GND 0.02fF
C1259 VDD.n862 GND 0.02fF
C1260 VDD.n866 GND 0.29fF
C1261 VDD.n867 GND 0.29fF
C1262 VDD.n868 GND 0.01fF
C1263 VDD.n869 GND 0.02fF
C1264 VDD.n870 GND 0.04fF
C1265 VDD.n871 GND 0.07fF
C1266 VDD.n872 GND 0.26fF
C1267 VDD.n873 GND 0.01fF
C1268 VDD.n874 GND 0.01fF
C1269 VDD.n875 GND 0.02fF
C1270 VDD.n876 GND 0.17fF
C1271 VDD.n877 GND 0.01fF
C1272 VDD.n878 GND 0.02fF
C1273 VDD.n879 GND 0.02fF
C1274 VDD.n880 GND 0.15fF
C1275 VDD.n881 GND 0.01fF
C1276 VDD.n882 GND 0.02fF
C1277 VDD.n883 GND 0.03fF
C1278 VDD.n884 GND 0.08fF
C1279 VDD.n885 GND 0.05fF
C1280 VDD.n886 GND 0.01fF
C1281 VDD.n887 GND 0.02fF
C1282 VDD.n888 GND 0.03fF
C1283 VDD.n889 GND 0.18fF
C1284 VDD.n890 GND 0.01fF
C1285 VDD.n891 GND 0.02fF
C1286 VDD.n892 GND 0.02fF
C1287 VDD.n893 GND 0.06fF
C1288 VDD.n894 GND 0.25fF
C1289 VDD.n895 GND 0.01fF
C1290 VDD.n896 GND 0.01fF
C1291 VDD.n897 GND 0.02fF
C1292 VDD.n898 GND 0.29fF
C1293 VDD.n899 GND 0.01fF
C1294 VDD.n900 GND 0.02fF
C1295 VDD.n901 GND 0.04fF
C1296 VDD.n902 GND 0.22fF
C1297 VDD.n903 GND 0.02fF
C1298 VDD.n904 GND 0.02fF
C1299 VDD.n905 GND 0.02fF
C1300 VDD.n906 GND 0.06fF
C1301 VDD.n907 GND 0.02fF
C1302 VDD.n908 GND 0.02fF
C1303 VDD.n909 GND 0.02fF
C1304 VDD.n910 GND 0.02fF
C1305 VDD.n911 GND 0.02fF
C1306 VDD.n912 GND 0.02fF
C1307 VDD.n913 GND 0.02fF
C1308 VDD.n914 GND 0.02fF
C1309 VDD.n915 GND 0.02fF
C1310 VDD.n916 GND 0.02fF
C1311 VDD.n917 GND 0.03fF
C1312 VDD.n918 GND 0.02fF
C1313 VDD.n919 GND 0.02fF
C1314 VDD.n923 GND 0.29fF
C1315 VDD.n924 GND 0.29fF
C1316 VDD.n925 GND 0.01fF
C1317 VDD.n926 GND 0.02fF
C1318 VDD.n927 GND 0.04fF
C1319 VDD.n928 GND 0.07fF
C1320 VDD.n929 GND 0.26fF
C1321 VDD.n930 GND 0.01fF
C1322 VDD.n931 GND 0.01fF
C1323 VDD.n932 GND 0.02fF
C1324 VDD.n933 GND 0.17fF
C1325 VDD.n934 GND 0.01fF
C1326 VDD.n935 GND 0.02fF
C1327 VDD.n936 GND 0.02fF
C1328 VDD.n937 GND 0.15fF
C1329 VDD.n938 GND 0.01fF
C1330 VDD.n939 GND 0.02fF
C1331 VDD.n940 GND 0.03fF
C1332 VDD.n941 GND 0.08fF
C1333 VDD.n942 GND 0.05fF
C1334 VDD.n943 GND 0.01fF
C1335 VDD.n944 GND 0.02fF
C1336 VDD.n945 GND 0.03fF
C1337 VDD.n946 GND 0.18fF
C1338 VDD.n947 GND 0.01fF
C1339 VDD.n948 GND 0.02fF
C1340 VDD.n949 GND 0.02fF
C1341 VDD.n950 GND 0.06fF
C1342 VDD.n951 GND 0.25fF
C1343 VDD.n952 GND 0.01fF
C1344 VDD.n953 GND 0.01fF
C1345 VDD.n954 GND 0.02fF
C1346 VDD.n955 GND 0.29fF
C1347 VDD.n956 GND 0.01fF
C1348 VDD.n957 GND 0.02fF
C1349 VDD.n958 GND 0.04fF
C1350 VDD.n959 GND 0.22fF
C1351 VDD.n960 GND 0.02fF
C1352 VDD.n961 GND 0.02fF
C1353 VDD.n962 GND 0.02fF
C1354 VDD.n963 GND 0.06fF
C1355 VDD.n964 GND 0.02fF
C1356 VDD.n965 GND 0.02fF
C1357 VDD.n966 GND 0.02fF
C1358 VDD.n967 GND 0.02fF
C1359 VDD.n968 GND 0.02fF
C1360 VDD.n969 GND 0.02fF
C1361 VDD.n970 GND 0.02fF
C1362 VDD.n971 GND 0.02fF
C1363 VDD.n972 GND 0.02fF
C1364 VDD.n973 GND 0.02fF
C1365 VDD.n974 GND 0.03fF
C1366 VDD.n975 GND 0.02fF
C1367 VDD.n976 GND 0.02fF
C1368 VDD.n980 GND 0.29fF
C1369 VDD.n981 GND 0.29fF
C1370 VDD.n982 GND 0.01fF
C1371 VDD.n983 GND 0.02fF
C1372 VDD.n984 GND 0.04fF
C1373 VDD.n985 GND 0.07fF
C1374 VDD.n986 GND 0.26fF
C1375 VDD.n987 GND 0.01fF
C1376 VDD.n988 GND 0.01fF
C1377 VDD.n989 GND 0.02fF
C1378 VDD.n990 GND 0.17fF
C1379 VDD.n991 GND 0.01fF
C1380 VDD.n992 GND 0.02fF
C1381 VDD.n993 GND 0.02fF
C1382 VDD.n994 GND 0.15fF
C1383 VDD.n995 GND 0.01fF
C1384 VDD.n996 GND 0.02fF
C1385 VDD.n997 GND 0.03fF
C1386 VDD.n998 GND 0.08fF
C1387 VDD.n999 GND 0.05fF
C1388 VDD.n1000 GND 0.01fF
C1389 VDD.n1001 GND 0.02fF
C1390 VDD.n1002 GND 0.03fF
C1391 VDD.n1003 GND 0.18fF
C1392 VDD.n1004 GND 0.01fF
C1393 VDD.n1005 GND 0.02fF
C1394 VDD.n1006 GND 0.02fF
C1395 VDD.n1007 GND 0.06fF
C1396 VDD.n1008 GND 0.25fF
C1397 VDD.n1009 GND 0.01fF
C1398 VDD.n1010 GND 0.01fF
C1399 VDD.n1011 GND 0.02fF
C1400 VDD.n1012 GND 0.29fF
C1401 VDD.n1013 GND 0.01fF
C1402 VDD.n1014 GND 0.02fF
C1403 VDD.n1015 GND 0.04fF
C1404 VDD.n1016 GND 0.27fF
C1405 VDD.n1017 GND 0.02fF
C1406 VDD.n1018 GND 0.02fF
C1407 VDD.n1019 GND 0.02fF
C1408 VDD.n1020 GND 0.06fF
C1409 VDD.n1021 GND 0.02fF
C1410 VDD.n1022 GND 0.02fF
C1411 VDD.n1023 GND 0.02fF
C1412 VDD.n1024 GND 0.02fF
C1413 VDD.n1025 GND 0.02fF
C1414 VDD.n1026 GND 0.02fF
C1415 VDD.n1027 GND 0.02fF
C1416 VDD.n1028 GND 0.02fF
C1417 VDD.n1029 GND 0.02fF
C1418 VDD.n1030 GND 0.02fF
C1419 VDD.n1031 GND 0.03fF
C1420 VDD.n1032 GND 0.02fF
C1421 VDD.n1033 GND 0.02fF
C1422 VDD.n1037 GND 0.29fF
C1423 VDD.n1038 GND 0.29fF
C1424 VDD.n1039 GND 0.01fF
C1425 VDD.n1040 GND 0.02fF
C1426 VDD.n1041 GND 0.04fF
C1427 VDD.n1042 GND 0.29fF
C1428 VDD.n1043 GND 0.01fF
C1429 VDD.n1044 GND 0.02fF
C1430 VDD.n1045 GND 0.02fF
C1431 VDD.n1046 GND 0.07fF
C1432 VDD.n1047 GND 0.23fF
C1433 VDD.n1048 GND 0.01fF
C1434 VDD.n1049 GND 0.01fF
C1435 VDD.n1050 GND 0.02fF
C1436 VDD.n1051 GND 0.18fF
C1437 VDD.n1052 GND 0.01fF
C1438 VDD.n1053 GND 0.02fF
C1439 VDD.n1054 GND 0.02fF
C1440 VDD.n1055 GND 0.08fF
C1441 VDD.n1056 GND 0.05fF
C1442 VDD.n1057 GND 0.16fF
C1443 VDD.n1058 GND 0.01fF
C1444 VDD.n1059 GND 0.02fF
C1445 VDD.n1060 GND 0.02fF
C1446 VDD.n1061 GND 0.16fF
C1447 VDD.n1062 GND 0.02fF
C1448 VDD.n1063 GND 0.02fF
C1449 VDD.n1064 GND 0.03fF
C1450 VDD.n1065 GND 0.15fF
C1451 VDD.n1066 GND 0.02fF
C1452 VDD.n1067 GND 0.02fF
C1453 VDD.n1068 GND 0.03fF
C1454 VDD.n1069 GND 0.17fF
C1455 VDD.n1070 GND 0.01fF
C1456 VDD.n1071 GND 0.08fF
C1457 VDD.n1072 GND 0.05fF
C1458 VDD.n1073 GND 0.02fF
C1459 VDD.n1074 GND 0.02fF
C1460 VDD.n1075 GND 0.18fF
C1461 VDD.n1076 GND 0.01fF
C1462 VDD.n1077 GND 0.02fF
C1463 VDD.n1078 GND 0.02fF
C1464 VDD.n1079 GND 0.23fF
C1465 VDD.n1080 GND 0.01fF
C1466 VDD.n1081 GND 0.07fF
C1467 VDD.n1082 GND 0.02fF
C1468 VDD.n1083 GND 0.29fF
C1469 VDD.n1084 GND 0.01fF
C1470 VDD.n1085 GND 0.02fF
C1471 VDD.n1086 GND 0.02fF
C1472 VDD.n1087 GND 0.29fF
C1473 VDD.n1088 GND 0.01fF
C1474 VDD.n1089 GND 0.02fF
C1475 VDD.n1090 GND 0.04fF
C1476 VDD.n1091 GND 0.27fF
C1477 VDD.n1092 GND 0.02fF
C1478 VDD.n1093 GND 0.02fF
C1479 VDD.n1094 GND 0.02fF
C1480 VDD.n1095 GND 0.06fF
C1481 VDD.n1096 GND 0.02fF
C1482 VDD.n1097 GND 0.02fF
C1483 VDD.n1098 GND 0.02fF
C1484 VDD.n1099 GND 0.02fF
C1485 VDD.n1100 GND 0.02fF
C1486 VDD.n1101 GND 0.02fF
C1487 VDD.n1102 GND 0.02fF
C1488 VDD.n1103 GND 0.02fF
C1489 VDD.n1104 GND 0.02fF
C1490 VDD.n1105 GND 0.02fF
C1491 VDD.n1106 GND 0.03fF
C1492 VDD.n1107 GND 0.02fF
C1493 VDD.n1108 GND 0.02fF
C1494 VDD.n1112 GND 0.29fF
C1495 VDD.n1113 GND 0.29fF
C1496 VDD.n1114 GND 0.01fF
C1497 VDD.n1115 GND 0.02fF
C1498 VDD.n1116 GND 0.04fF
C1499 VDD.n1117 GND 0.07fF
C1500 VDD.n1118 GND 0.26fF
C1501 VDD.n1119 GND 0.01fF
C1502 VDD.n1120 GND 0.01fF
C1503 VDD.n1121 GND 0.02fF
C1504 VDD.n1122 GND 0.17fF
C1505 VDD.n1123 GND 0.01fF
C1506 VDD.n1124 GND 0.02fF
C1507 VDD.n1125 GND 0.02fF
C1508 VDD.n1126 GND 0.15fF
C1509 VDD.n1127 GND 0.01fF
C1510 VDD.n1128 GND 0.02fF
C1511 VDD.n1129 GND 0.03fF
C1512 VDD.n1130 GND 0.08fF
C1513 VDD.n1131 GND 0.05fF
C1514 VDD.n1132 GND 0.01fF
C1515 VDD.n1133 GND 0.02fF
C1516 VDD.n1134 GND 0.03fF
C1517 VDD.n1135 GND 0.18fF
C1518 VDD.n1136 GND 0.01fF
C1519 VDD.n1137 GND 0.02fF
C1520 VDD.n1138 GND 0.02fF
C1521 VDD.n1139 GND 0.06fF
C1522 VDD.n1140 GND 0.25fF
C1523 VDD.n1141 GND 0.01fF
C1524 VDD.n1142 GND 0.01fF
C1525 VDD.n1143 GND 0.02fF
C1526 VDD.n1144 GND 0.29fF
C1527 VDD.n1145 GND 0.01fF
C1528 VDD.n1146 GND 0.02fF
C1529 VDD.n1147 GND 0.04fF
C1530 VDD.n1148 GND 0.22fF
C1531 VDD.n1149 GND 0.02fF
C1532 VDD.n1150 GND 0.02fF
C1533 VDD.n1151 GND 0.02fF
C1534 VDD.n1152 GND 0.06fF
C1535 VDD.n1153 GND 0.02fF
C1536 VDD.n1154 GND 0.02fF
C1537 VDD.n1155 GND 0.02fF
C1538 VDD.n1156 GND 0.02fF
C1539 VDD.n1157 GND 0.02fF
C1540 VDD.n1158 GND 0.02fF
C1541 VDD.n1159 GND 0.02fF
C1542 VDD.n1160 GND 0.02fF
C1543 VDD.n1161 GND 0.02fF
C1544 VDD.n1162 GND 0.02fF
C1545 VDD.n1163 GND 0.03fF
C1546 VDD.n1164 GND 0.02fF
C1547 VDD.n1165 GND 0.02fF
C1548 VDD.n1169 GND 0.29fF
C1549 VDD.n1170 GND 0.29fF
C1550 VDD.n1171 GND 0.01fF
C1551 VDD.n1172 GND 0.02fF
C1552 VDD.n1173 GND 0.04fF
C1553 VDD.n1174 GND 0.07fF
C1554 VDD.n1175 GND 0.26fF
C1555 VDD.n1176 GND 0.01fF
C1556 VDD.n1177 GND 0.01fF
C1557 VDD.n1178 GND 0.02fF
C1558 VDD.n1179 GND 0.17fF
C1559 VDD.n1180 GND 0.01fF
C1560 VDD.n1181 GND 0.02fF
C1561 VDD.n1182 GND 0.02fF
C1562 VDD.n1183 GND 0.15fF
C1563 VDD.n1184 GND 0.01fF
C1564 VDD.n1185 GND 0.02fF
C1565 VDD.n1186 GND 0.03fF
C1566 VDD.n1187 GND 0.08fF
C1567 VDD.n1188 GND 0.05fF
C1568 VDD.n1189 GND 0.01fF
C1569 VDD.n1190 GND 0.02fF
C1570 VDD.n1191 GND 0.03fF
C1571 VDD.n1192 GND 0.18fF
C1572 VDD.n1193 GND 0.01fF
C1573 VDD.n1194 GND 0.02fF
C1574 VDD.n1195 GND 0.02fF
C1575 VDD.n1196 GND 0.06fF
C1576 VDD.n1197 GND 0.25fF
C1577 VDD.n1198 GND 0.01fF
C1578 VDD.n1199 GND 0.01fF
C1579 VDD.n1200 GND 0.02fF
C1580 VDD.n1201 GND 0.29fF
C1581 VDD.n1202 GND 0.01fF
C1582 VDD.n1203 GND 0.02fF
C1583 VDD.n1204 GND 0.04fF
C1584 VDD.n1205 GND 0.22fF
C1585 VDD.n1206 GND 0.02fF
C1586 VDD.n1207 GND 0.02fF
C1587 VDD.n1208 GND 0.02fF
C1588 VDD.n1209 GND 0.06fF
C1589 VDD.n1210 GND 0.02fF
C1590 VDD.n1211 GND 0.02fF
C1591 VDD.n1212 GND 0.02fF
C1592 VDD.n1213 GND 0.02fF
C1593 VDD.n1214 GND 0.02fF
C1594 VDD.n1215 GND 0.02fF
C1595 VDD.n1216 GND 0.02fF
C1596 VDD.n1217 GND 0.02fF
C1597 VDD.n1218 GND 0.02fF
C1598 VDD.n1219 GND 0.02fF
C1599 VDD.n1220 GND 0.03fF
C1600 VDD.n1221 GND 0.02fF
C1601 VDD.n1222 GND 0.02fF
C1602 VDD.n1226 GND 0.29fF
C1603 VDD.n1227 GND 0.29fF
C1604 VDD.n1228 GND 0.01fF
C1605 VDD.n1229 GND 0.02fF
C1606 VDD.n1230 GND 0.04fF
C1607 VDD.n1231 GND 0.07fF
C1608 VDD.n1232 GND 0.26fF
C1609 VDD.n1233 GND 0.01fF
C1610 VDD.n1234 GND 0.01fF
C1611 VDD.n1235 GND 0.02fF
C1612 VDD.n1236 GND 0.17fF
C1613 VDD.n1237 GND 0.01fF
C1614 VDD.n1238 GND 0.02fF
C1615 VDD.n1239 GND 0.02fF
C1616 VDD.n1240 GND 0.15fF
C1617 VDD.n1241 GND 0.01fF
C1618 VDD.n1242 GND 0.02fF
C1619 VDD.n1243 GND 0.03fF
C1620 VDD.n1244 GND 0.08fF
C1621 VDD.n1245 GND 0.05fF
C1622 VDD.n1246 GND 0.01fF
C1623 VDD.n1247 GND 0.02fF
C1624 VDD.n1248 GND 0.03fF
C1625 VDD.n1249 GND 0.18fF
C1626 VDD.n1250 GND 0.01fF
C1627 VDD.n1251 GND 0.02fF
C1628 VDD.n1252 GND 0.02fF
C1629 VDD.n1253 GND 0.06fF
C1630 VDD.n1254 GND 0.25fF
C1631 VDD.n1255 GND 0.01fF
C1632 VDD.n1256 GND 0.01fF
C1633 VDD.n1257 GND 0.02fF
C1634 VDD.n1258 GND 0.29fF
C1635 VDD.n1259 GND 0.01fF
C1636 VDD.n1260 GND 0.02fF
C1637 VDD.n1261 GND 0.04fF
C1638 VDD.n1262 GND 0.22fF
C1639 VDD.n1263 GND 0.02fF
C1640 VDD.n1264 GND 0.02fF
C1641 VDD.n1265 GND 0.02fF
C1642 VDD.n1266 GND 0.06fF
C1643 VDD.n1267 GND 0.02fF
C1644 VDD.n1268 GND 0.02fF
C1645 VDD.n1269 GND 0.02fF
C1646 VDD.n1270 GND 0.02fF
C1647 VDD.n1271 GND 0.02fF
C1648 VDD.n1272 GND 0.02fF
C1649 VDD.n1273 GND 0.02fF
C1650 VDD.n1274 GND 0.02fF
C1651 VDD.n1275 GND 0.02fF
C1652 VDD.n1276 GND 0.02fF
C1653 VDD.n1277 GND 0.03fF
C1654 VDD.n1278 GND 0.02fF
C1655 VDD.n1279 GND 0.02fF
C1656 VDD.n1283 GND 0.29fF
C1657 VDD.n1284 GND 0.29fF
C1658 VDD.n1285 GND 0.01fF
C1