magic
tech sky130A
magscale 1 2
timestamp 1642371692
<< error_p >>
rect 85 322 86 323
rect 86 321 87 322
rect 101 291 102 292
rect 136 291 137 292
rect 101 188 102 189
rect 136 188 137 189
<< nwell >>
rect -36 591 354 1353
<< nmos >>
rect 56 322 86 375
rect 56 292 152 322
tri 152 292 182 322 sw
rect 56 188 86 292
tri 86 276 102 292 nw
tri 136 276 152 292 ne
tri 86 188 102 204 sw
tri 136 188 152 204 se
rect 152 188 182 292
tri 56 158 86 188 ne
rect 86 158 152 188
tri 152 158 182 188 nw
<< pmos >>
rect 56 629 86 1229
rect 144 629 174 1229
rect 232 629 262 1229
<< ndiff >>
rect 0 298 56 375
rect 86 322 236 375
rect 0 264 10 298
rect 44 264 56 298
tri 152 292 182 322 ne
rect 182 298 236 322
rect 0 215 56 264
rect 0 181 10 215
rect 44 181 56 215
tri 86 276 102 292 se
rect 102 276 136 292
tri 136 276 152 292 sw
rect 86 244 152 276
rect 86 210 98 244
rect 132 210 152 244
rect 86 204 152 210
tri 86 188 102 204 ne
rect 102 188 136 204
tri 136 188 152 204 nw
rect 182 264 194 298
rect 228 264 236 298
rect 182 215 236 264
rect 0 158 56 181
tri 56 158 86 188 sw
tri 152 158 182 188 se
rect 182 181 194 215
rect 228 181 236 215
rect 182 158 236 181
rect 0 147 236 158
rect 0 113 10 147
rect 44 113 98 147
rect 132 113 194 147
rect 228 113 236 147
rect 0 101 236 113
<< pdiff >>
rect 0 1213 56 1229
rect 0 1179 10 1213
rect 44 1179 56 1213
rect 0 1145 56 1179
rect 0 1111 10 1145
rect 44 1111 56 1145
rect 0 1077 56 1111
rect 0 1043 10 1077
rect 44 1043 56 1077
rect 0 1009 56 1043
rect 0 975 10 1009
rect 44 975 56 1009
rect 0 941 56 975
rect 0 907 10 941
rect 44 907 56 941
rect 0 873 56 907
rect 0 839 10 873
rect 44 839 56 873
rect 0 805 56 839
rect 0 771 10 805
rect 44 771 56 805
rect 0 737 56 771
rect 0 703 10 737
rect 44 703 56 737
rect 0 629 56 703
rect 86 1213 144 1229
rect 86 1179 98 1213
rect 132 1179 144 1213
rect 86 1145 144 1179
rect 86 1111 98 1145
rect 132 1111 144 1145
rect 86 1077 144 1111
rect 86 1043 98 1077
rect 132 1043 144 1077
rect 86 1009 144 1043
rect 86 975 98 1009
rect 132 975 144 1009
rect 86 941 144 975
rect 86 907 98 941
rect 132 907 144 941
rect 86 873 144 907
rect 86 839 98 873
rect 132 839 144 873
rect 86 805 144 839
rect 86 771 98 805
rect 132 771 144 805
rect 86 737 144 771
rect 86 703 98 737
rect 132 703 144 737
rect 86 629 144 703
rect 174 1213 232 1229
rect 174 1179 186 1213
rect 220 1179 232 1213
rect 174 1145 232 1179
rect 174 1111 186 1145
rect 220 1111 232 1145
rect 174 1077 232 1111
rect 174 1043 186 1077
rect 220 1043 232 1077
rect 174 1009 232 1043
rect 174 975 186 1009
rect 220 975 232 1009
rect 174 941 232 975
rect 174 907 186 941
rect 220 907 232 941
rect 174 873 232 907
rect 174 839 186 873
rect 220 839 232 873
rect 174 805 232 839
rect 174 771 186 805
rect 220 771 232 805
rect 174 737 232 771
rect 174 703 186 737
rect 220 703 232 737
rect 174 629 232 703
rect 262 1213 318 1229
rect 262 1179 274 1213
rect 308 1179 318 1213
rect 262 1145 318 1179
rect 262 1111 274 1145
rect 308 1111 318 1145
rect 262 1077 318 1111
rect 262 1043 274 1077
rect 308 1043 318 1077
rect 262 1009 318 1043
rect 262 975 274 1009
rect 308 975 318 1009
rect 262 941 318 975
rect 262 907 274 941
rect 308 907 318 941
rect 262 873 318 907
rect 262 839 274 873
rect 308 839 318 873
rect 262 805 318 839
rect 262 771 274 805
rect 308 771 318 805
rect 262 737 318 771
rect 262 703 274 737
rect 308 703 318 737
rect 262 629 318 703
<< ndiffc >>
rect 10 264 44 298
rect 10 181 44 215
rect 98 210 132 244
rect 194 264 228 298
rect 194 181 228 215
rect 10 113 44 147
rect 98 113 132 147
rect 194 113 228 147
<< pdiffc >>
rect 10 1179 44 1213
rect 10 1111 44 1145
rect 10 1043 44 1077
rect 10 975 44 1009
rect 10 907 44 941
rect 10 839 44 873
rect 10 771 44 805
rect 10 703 44 737
rect 98 1179 132 1213
rect 98 1111 132 1145
rect 98 1043 132 1077
rect 98 975 132 1009
rect 98 907 132 941
rect 98 839 132 873
rect 98 771 132 805
rect 98 703 132 737
rect 186 1179 220 1213
rect 186 1111 220 1145
rect 186 1043 220 1077
rect 186 975 220 1009
rect 186 907 220 941
rect 186 839 220 873
rect 186 771 220 805
rect 186 703 220 737
rect 274 1179 308 1213
rect 274 1111 308 1145
rect 274 1043 308 1077
rect 274 975 308 1009
rect 274 907 308 941
rect 274 839 308 873
rect 274 771 308 805
rect 274 703 308 737
<< psubdiff >>
rect 0 13 24 47
rect 58 13 93 47
rect 127 13 169 47
rect 203 13 237 47
rect 271 13 319 47
<< nsubdiff >>
rect 0 1283 24 1317
rect 58 1283 92 1317
rect 126 1283 160 1317
rect 195 1283 229 1317
rect 263 1283 318 1317
<< psubdiffcont >>
rect 24 13 58 47
rect 93 13 127 47
rect 169 13 203 47
rect 237 13 271 47
<< nsubdiffcont >>
rect 24 1283 58 1317
rect 92 1283 126 1317
rect 160 1283 195 1317
rect 229 1283 263 1317
<< poly >>
rect 56 1229 86 1255
rect 144 1229 174 1255
rect 232 1229 262 1255
rect 56 612 86 629
rect 144 612 174 629
rect 232 612 262 629
rect 56 582 262 612
rect 56 494 86 582
rect 20 478 86 494
rect 20 444 30 478
rect 64 444 86 478
rect 20 428 86 444
rect 56 375 86 428
<< polycont >>
rect 30 444 64 478
<< locali >>
rect 0 1317 318 1332
rect 0 1283 24 1317
rect 58 1283 92 1317
rect 126 1283 160 1317
rect 195 1283 229 1317
rect 263 1283 318 1317
rect 0 1270 318 1283
rect 10 1213 44 1270
rect 10 1145 44 1179
rect 10 1077 44 1111
rect 10 1009 44 1043
rect 10 941 44 975
rect 10 873 44 907
rect 10 805 44 839
rect 10 737 44 771
rect 10 627 44 703
rect 98 1213 132 1229
rect 98 1145 132 1179
rect 98 1077 132 1111
rect 98 1009 132 1043
rect 98 941 132 975
rect 98 873 132 907
rect 98 805 132 839
rect 98 737 132 771
rect 98 672 132 703
rect 30 478 64 494
rect 30 428 64 444
rect 10 298 44 343
rect 10 215 44 264
rect 98 244 132 638
rect 186 1213 220 1270
rect 186 1145 220 1179
rect 186 1077 220 1111
rect 186 1009 220 1043
rect 186 941 220 975
rect 186 873 220 907
rect 186 805 220 839
rect 186 737 220 771
rect 186 627 220 703
rect 274 1213 308 1229
rect 274 1145 308 1179
rect 274 1077 308 1111
rect 274 1009 308 1043
rect 274 941 308 975
rect 274 873 308 907
rect 274 805 308 839
rect 274 737 308 771
rect 274 673 308 703
rect 98 194 132 210
rect 194 298 228 343
rect 194 215 228 264
rect 10 147 44 181
rect 194 147 228 181
rect 44 113 98 147
rect 132 113 194 147
rect 10 62 44 113
rect 194 62 228 113
rect 0 47 319 62
rect 0 13 24 47
rect 58 13 93 47
rect 127 13 169 47
rect 203 13 237 47
rect 271 13 319 47
rect 0 0 319 13
<< viali >>
rect 24 1283 58 1317
rect 92 1283 126 1317
rect 160 1283 195 1317
rect 229 1283 263 1317
rect 98 638 132 672
rect 30 444 64 478
rect 274 639 308 673
rect 24 13 58 47
rect 93 13 127 47
rect 169 13 203 47
rect 237 13 271 47
<< metal1 >>
rect 0 1317 318 1332
rect 0 1283 24 1317
rect 58 1283 92 1317
rect 126 1283 160 1317
rect 195 1283 229 1317
rect 263 1283 318 1317
rect 0 1270 318 1283
rect 86 672 143 678
rect 262 673 320 679
rect 262 672 274 673
rect 86 638 98 672
rect 132 639 274 672
rect 308 639 320 673
rect 132 638 320 639
rect 86 632 143 638
rect 262 632 320 638
rect 98 628 132 632
rect 30 485 64 502
rect 24 478 70 485
rect 24 444 30 478
rect 64 444 70 478
rect 24 437 70 444
rect 30 421 64 437
rect 0 47 319 62
rect 0 13 24 47
rect 58 13 93 47
rect 127 13 169 47
rect 203 13 237 47
rect 271 13 319 47
rect 0 0 319 13
<< labels >>
rlabel metal1 161 1325 161 1325 1 VDD
rlabel metal1 30 444 64 478 1 A
rlabel metal1 148 31 148 31 1 VSS
rlabel metal1 98 638 132 672 1 Y
<< end >>
