magic
tech sky130A
magscale 1 2
timestamp 1648064525
<< nwell >>
rect 528 1554 1026 1575
rect 1194 1554 1692 1575
rect 475 1492 1079 1554
rect 1141 1492 1745 1554
rect 528 1486 1026 1492
rect 528 1015 539 1486
rect 585 1377 619 1411
rect 1015 1015 1026 1486
rect 528 832 1026 1015
rect 1194 1487 1692 1492
rect 1194 1015 1205 1487
rect 1681 1015 1692 1487
rect 1194 832 1692 1015
<< pdiffc >>
rect 585 1377 619 1411
rect 761 1377 795 1411
rect 937 1377 971 1411
rect 1251 1377 1285 1411
rect 1427 1377 1461 1411
rect 1603 1377 1637 1411
rect 585 1105 619 1139
rect 761 1105 795 1139
rect 849 1105 883 1139
rect 1251 1105 1285 1139
rect 1427 1105 1461 1139
rect 1515 1105 1549 1139
<< psubdiff >>
rect 475 510 1079 572
rect 1141 510 1745 572
rect 475 13 499 47
rect 533 13 571 47
rect 605 13 643 47
rect 677 13 715 47
rect 749 13 805 47
rect 839 13 877 47
rect 911 13 949 47
rect 983 13 1021 47
rect 1055 13 1079 47
rect 1141 13 1165 47
rect 1199 13 1237 47
rect 1271 13 1309 47
rect 1343 13 1381 47
rect 1415 13 1471 47
rect 1505 13 1543 47
rect 1577 13 1615 47
rect 1649 13 1687 47
rect 1721 13 1745 47
<< nsubdiff >>
rect 475 1505 499 1539
rect 533 1505 571 1539
rect 605 1505 643 1539
rect 677 1505 715 1539
rect 749 1505 805 1539
rect 839 1505 877 1539
rect 911 1505 949 1539
rect 983 1505 1021 1539
rect 1055 1505 1079 1539
rect 1141 1505 1165 1539
rect 1199 1505 1237 1539
rect 1271 1505 1309 1539
rect 1343 1505 1381 1539
rect 1415 1505 1471 1539
rect 1505 1505 1543 1539
rect 1577 1505 1615 1539
rect 1649 1505 1687 1539
rect 1721 1505 1745 1539
rect 475 868 1079 930
rect 1141 868 1745 930
<< psubdiffcont >>
rect 499 13 533 47
rect 571 13 605 47
rect 643 13 677 47
rect 715 13 749 47
rect 805 13 839 47
rect 877 13 911 47
rect 949 13 983 47
rect 1021 13 1055 47
rect 1165 13 1199 47
rect 1237 13 1271 47
rect 1309 13 1343 47
rect 1381 13 1415 47
rect 1471 13 1505 47
rect 1543 13 1577 47
rect 1615 13 1649 47
rect 1687 13 1721 47
<< nsubdiffcont >>
rect 499 1505 533 1539
rect 571 1505 605 1539
rect 643 1505 677 1539
rect 715 1505 749 1539
rect 805 1505 839 1539
rect 877 1505 911 1539
rect 949 1505 983 1539
rect 1021 1505 1055 1539
rect 1165 1505 1199 1539
rect 1237 1505 1271 1539
rect 1309 1505 1343 1539
rect 1381 1505 1415 1539
rect 1471 1505 1505 1539
rect 1543 1505 1577 1539
rect 1615 1505 1649 1539
rect 1687 1505 1721 1539
<< poly >>
rect 612 411 639 441
rect 806 411 861 441
rect 1278 411 1305 441
rect 1472 411 1527 441
rect 612 403 642 411
rect 806 410 836 411
rect 1278 403 1308 411
rect 1472 410 1502 411
<< locali >>
rect 475 1539 1079 1554
rect 475 1505 499 1539
rect 533 1505 571 1539
rect 605 1505 643 1539
rect 677 1505 715 1539
rect 749 1505 805 1539
rect 839 1505 877 1539
rect 911 1505 949 1539
rect 983 1505 1021 1539
rect 1055 1505 1079 1539
rect 475 1492 1079 1505
rect 1141 1539 1745 1554
rect 1141 1505 1165 1539
rect 1199 1505 1237 1539
rect 1271 1505 1309 1539
rect 1343 1505 1381 1539
rect 1415 1505 1471 1539
rect 1505 1505 1543 1539
rect 1577 1505 1615 1539
rect 1649 1505 1687 1539
rect 1721 1505 1745 1539
rect 1141 1492 1745 1505
rect 585 1411 619 1427
rect 585 1359 619 1377
rect 673 1359 707 1492
rect 761 1411 971 1445
rect 761 1359 795 1377
rect 937 1359 971 1377
rect 1251 1411 1285 1427
rect 1251 1359 1285 1377
rect 1339 1359 1373 1492
rect 1427 1411 1637 1445
rect 1427 1359 1461 1377
rect 1603 1359 1637 1377
rect 585 1139 619 1157
rect 761 1139 795 1157
rect 585 1071 795 1105
rect 849 1139 883 1157
rect 1251 1139 1285 1157
rect 1427 1139 1461 1157
rect 849 1071 979 1105
rect 1251 1071 1461 1105
rect 1515 1139 1549 1157
rect 1515 1071 1645 1105
rect 649 475 683 954
rect 871 847 905 954
rect 871 477 905 617
rect 945 375 979 1071
rect 1315 475 1349 954
rect 1537 913 1571 954
rect 1389 551 1423 856
rect 1536 782 1571 913
rect 1537 476 1571 545
rect 1611 375 1645 1071
rect 857 341 979 375
rect 1523 341 1645 375
rect 857 244 891 341
rect 1523 244 1557 341
rect 663 62 697 202
rect 1329 62 1363 202
rect 475 47 1079 62
rect 475 13 499 47
rect 533 13 571 47
rect 605 13 643 47
rect 677 13 715 47
rect 749 13 805 47
rect 839 13 877 47
rect 911 13 949 47
rect 983 13 1021 47
rect 1055 13 1079 47
rect 475 0 1079 13
rect 1141 47 1745 62
rect 1141 13 1165 47
rect 1199 13 1237 47
rect 1271 13 1309 47
rect 1343 13 1381 47
rect 1415 13 1471 47
rect 1505 13 1543 47
rect 1577 13 1615 47
rect 1649 13 1687 47
rect 1721 13 1745 47
rect 1141 0 1745 13
<< viali >>
rect 499 1505 533 1539
rect 571 1505 605 1539
rect 643 1505 677 1539
rect 715 1505 749 1539
rect 805 1505 839 1539
rect 877 1505 911 1539
rect 949 1505 983 1539
rect 1021 1505 1055 1539
rect 1165 1505 1199 1539
rect 1237 1505 1271 1539
rect 1309 1505 1343 1539
rect 1381 1505 1415 1539
rect 1471 1505 1505 1539
rect 1543 1505 1577 1539
rect 1615 1505 1649 1539
rect 1687 1505 1721 1539
rect 499 13 533 47
rect 571 13 605 47
rect 643 13 677 47
rect 715 13 749 47
rect 805 13 839 47
rect 877 13 911 47
rect 949 13 983 47
rect 1021 13 1055 47
rect 1165 13 1199 47
rect 1237 13 1271 47
rect 1309 13 1343 47
rect 1381 13 1415 47
rect 1471 13 1505 47
rect 1543 13 1577 47
rect 1615 13 1649 47
rect 1687 13 1721 47
<< metal1 >>
rect 475 1539 1079 1554
rect 475 1505 499 1539
rect 533 1505 571 1539
rect 605 1505 643 1539
rect 677 1505 715 1539
rect 749 1505 805 1539
rect 839 1505 877 1539
rect 911 1505 949 1539
rect 983 1505 1021 1539
rect 1055 1505 1079 1539
rect 475 1492 1079 1505
rect 1141 1539 1745 1554
rect 1141 1505 1165 1539
rect 1199 1505 1237 1539
rect 1271 1505 1309 1539
rect 1343 1505 1381 1539
rect 1415 1505 1471 1539
rect 1505 1505 1543 1539
rect 1577 1505 1615 1539
rect 1649 1505 1687 1539
rect 1721 1505 1745 1539
rect 1141 1492 1745 1505
rect 315 871 1359 905
rect 683 797 1871 831
rect 981 723 1586 757
rect 1425 501 1501 535
rect 475 47 1079 62
rect 475 13 499 47
rect 533 13 571 47
rect 605 13 643 47
rect 677 13 715 47
rect 749 13 805 47
rect 839 13 877 47
rect 911 13 949 47
rect 983 13 1021 47
rect 1055 13 1079 47
rect 475 0 1079 13
rect 1141 47 1745 62
rect 1141 13 1165 47
rect 1199 13 1237 47
rect 1271 13 1309 47
rect 1343 13 1381 47
rect 1415 13 1471 47
rect 1505 13 1543 47
rect 1577 13 1615 47
rect 1649 13 1687 47
rect 1721 13 1745 47
rect 1141 0 1745 13
use invx1_pcell  invx1_pcell_0
timestamp 1648064504
transform 1 0 0 0 1 0
box -84 0 528 1575
use diff_ring_side  diff_ring_side_1
timestamp 1648063806
transform 1 0 444 0 1 0
box -84 0 84 1575
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform -1 0 296 0 -1 888
box -53 -33 29 33
use poly_li1_contact  poly_li1_contact_0
timestamp 1648060378
transform 0 1 667 -1 0 988
box -32 -28 34 26
use poly_li1_contact  poly_li1_contact_1
timestamp 1648060378
transform 0 1 667 -1 0 445
box -32 -28 34 26
use nmos_top_trim1  nmos_top_trim1_0
timestamp 1648061897
transform -1 0 998 0 1 101
box 0 0 248 309
use nmos_bottom  nmos_bottom_0
timestamp 1648062456
transform -1 0 804 0 1 101
box 0 0 248 302
use li1_M1_contact  li1_M1_contact_3
timestamp 1648061256
transform -1 0 666 0 -1 814
box -53 -33 29 33
use pmos2_1  pmos2_1_0
timestamp 1647326732
transform 1 0 487 0 1 1450
box 52 -460 352 37
use pmos2_1  pmos2_1_1
timestamp 1647326732
transform 1 0 663 0 1 1450
box 52 -460 352 37
use diff_ring_side  diff_ring_side_0
timestamp 1648063806
transform 1 0 1110 0 1 0
box -84 0 84 1575
use poly_li1_contact  poly_li1_contact_3
timestamp 1648060378
transform 0 1 889 -1 0 988
box -32 -28 34 26
use poly_li1_contact  poly_li1_contact_2
timestamp 1648060378
transform 0 1 889 -1 0 445
box -32 -28 34 26
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform 1 0 888 0 1 888
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_7
timestamp 1648061256
transform -1 0 962 0 -1 740
box -53 -33 29 33
use poly_li1_contact  poly_li1_contact_5
timestamp 1648060378
transform 0 1 1333 -1 0 988
box -32 -28 34 26
use poly_li1_contact  poly_li1_contact_4
timestamp 1648060378
transform 0 1 1333 -1 0 445
box -32 -28 34 26
use nmos_top_trim1  nmos_top_trim1_1
timestamp 1648061897
transform -1 0 1664 0 1 101
box 0 0 248 309
use nmos_bottom  nmos_bottom_1
timestamp 1648062456
transform -1 0 1470 0 1 101
box 0 0 248 302
use li1_M1_contact  li1_M1_contact_5
timestamp 1648061256
transform -1 0 1406 0 -1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_4
timestamp 1648061256
transform 1 0 1406 0 1 888
box -53 -33 29 33
use pmos2_1  pmos2_1_3
timestamp 1647326732
transform 1 0 1329 0 1 1450
box 52 -460 352 37
use pmos2_1  pmos2_1_2
timestamp 1647326732
transform 1 0 1153 0 1 1450
box 52 -460 352 37
use diff_ring_side  diff_ring_side_3
timestamp 1648063806
transform 1 0 1776 0 1 0
box -84 0 84 1575
use poly_li1_contact  poly_li1_contact_7
timestamp 1648060378
transform 0 1 1555 -1 0 988
box -32 -28 34 26
use poly_li1_contact  poly_li1_contact_6
timestamp 1648060378
transform 0 1 1555 -1 0 445
box -32 -28 34 26
use li1_M1_contact  li1_M1_contact_6
timestamp 1648061256
transform 1 0 1554 0 1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_8
timestamp 1648061256
transform 1 0 1628 0 1 740
box -53 -33 29 33
use invx1_pcell  invx1_pcell_1
timestamp 1648064504
transform 1 0 1776 0 1 0
box -84 0 528 1575
use li1_M1_contact  li1_M1_contact_2
timestamp 1648061256
transform 1 0 1924 0 1 814
box -53 -33 29 33
<< end >>
