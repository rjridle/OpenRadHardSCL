* HSPICE file created from tmp.ext - technology: sky130A

.option scale=5000u

.subckt tmp A B Y VDD VSS
X0 VDD A Y VDD sky130_fd_pr__pfet_01v8 ad=33600 pd=1368 as=23200 ps=916 w=400 l=30 M=2
X1 VDD B Y VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=400 l=30 M=2
X2 VSS A a_112_101 VSS sky130_fd_pr__nfet_01v8 ad=7088 pd=312 as=0 ps=0 w=598 l=30
X3 Y B a_112_101 VSS sky130_fd_pr__nfet_01v8 ad=7088 pd=312 as=0 ps=0 w=598 l=30
.ends

** hspice subcircuit dictionary
