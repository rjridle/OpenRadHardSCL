magic
tech sky130A
magscale 1 2
timestamp 1643181757
<< nwell >>
rect -36 1344 464 1353
rect -38 1332 464 1344
rect 536 1332 569 1334
rect -116 1278 569 1332
rect -54 1270 569 1278
rect -38 1245 464 1270
rect 536 1265 569 1270
rect 234 1055 464 1245
rect -150 759 558 1055
rect 234 758 464 759
<< psubdiff >>
rect -116 490 476 552
rect -54 13 24 47
rect 58 13 92 47
rect 126 13 160 47
rect 194 13 228 47
rect 262 13 296 47
rect 330 13 364 47
rect 398 13 476 47
<< nsubdiff >>
rect -69 1283 24 1317
rect 58 1283 92 1317
rect 126 1283 160 1317
rect 195 1283 229 1317
rect 263 1283 297 1317
rect 331 1283 365 1317
rect 399 1283 503 1317
rect -116 795 534 857
<< psubdiffcont >>
rect 24 13 58 47
rect 92 13 126 47
rect 160 13 194 47
rect 228 13 262 47
rect 296 13 330 47
rect 364 13 398 47
<< nsubdiffcont >>
rect 24 1283 58 1317
rect 92 1283 126 1317
rect 160 1283 195 1317
rect 229 1283 263 1317
rect 297 1283 331 1317
rect 365 1283 399 1317
<< poly >>
rect 184 916 242 946
rect 86 401 270 431
<< locali >>
rect -116 1317 536 1332
rect -116 1283 24 1317
rect 58 1283 92 1317
rect 126 1283 160 1317
rect 195 1283 229 1317
rect 263 1283 297 1317
rect 331 1283 365 1317
rect 399 1283 536 1317
rect -116 1278 536 1283
rect -54 1270 536 1278
rect 370 1269 404 1270
rect 10 62 44 101
rect 194 62 228 101
rect 378 62 412 101
rect -54 47 476 62
rect -54 13 24 47
rect 58 13 92 47
rect 126 13 160 47
rect 194 13 228 47
rect 262 13 296 47
rect 330 13 364 47
rect 398 13 476 47
rect -54 0 476 13
<< viali >>
rect 24 1283 58 1317
rect 92 1283 126 1317
rect 160 1283 195 1317
rect 229 1283 263 1317
rect 297 1283 331 1317
rect 365 1283 399 1317
rect 24 13 58 47
rect 92 13 126 47
rect 160 13 194 47
rect 228 13 262 47
rect 296 13 330 47
rect 364 13 398 47
<< metal1 >>
rect -116 1317 536 1332
rect -116 1283 24 1317
rect 58 1283 92 1317
rect 126 1283 160 1317
rect 195 1283 229 1317
rect 263 1283 297 1317
rect 331 1283 365 1317
rect 399 1283 536 1317
rect -116 1278 536 1283
rect -54 1270 536 1278
rect 42 462 76 876
rect -54 47 476 62
rect -54 13 24 47
rect 58 13 92 47
rect 126 13 160 47
rect 194 13 228 47
rect 262 13 296 47
rect 330 13 364 47
rect 398 13 476 47
rect -54 0 476 13
use diff_ring_side  diff_ring_side_1 ./pcells
timestamp 1643181737
transform 1 0 582 0 1 0
box -159 0 9 1353
use diff_ring_side  diff_ring_side_0
timestamp 1643181737
transform 1 0 -10 0 1 0
box -159 0 9 1353
use M1_M2_contact  M1_M2_contact_0 pcells
timestamp 1643168619
transform 1 0 -38 0 1 481
box 64 391 130 473
use pmos  pmos_0 pcells
timestamp 1643179034
transform 1 0 10 0 1 1228
box -36 -312 264 42
use pmos  pmos_1
timestamp 1643179034
transform 1 0 186 0 1 1228
box -36 -312 264 42
use nmos_top_left  nmos_top_left_1 pcells
timestamp 1643177486
transform 1 0 229 0 1 165
box -45 -64 193 238
use nmos_top_left  nmos_top_left_0
timestamp 1643177486
transform 1 0 45 0 1 165
box -45 -64 193 238
use M1_M2_contact  M1_M2_contact_1
timestamp 1643168619
transform -1 0 156 0 -1 866
box 64 391 130 473
<< labels >>
rlabel metal1 278 26 278 26 1 VSS
port 4 n
rlabel metal1 281 1301 281 1301 1 VDD
port 1 n
<< end >>
