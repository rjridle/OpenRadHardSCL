* HSPICE file created from tmp.ext - technology: sky130A

.option scale=5000u

.subckt tmp A B Y VDD VSS
X0 a_131_1051 A VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=11600 ps=458 w=400 l=30 M=2
X1 Y A VSS VSS sky130_fd_pr__nfet_01v8 ad=14176 pd=624 as=77676 ps=2588 w=598 l=30
X2 a_131_1051 B Y VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=11600 ps=458 w=400 l=30 M=2
X3 Y B VSS VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=598 l=30
.ends

** hspice subcircuit dictionary
