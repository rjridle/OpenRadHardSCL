** sch_path: /home/rjridle/OpenRadHardSCL/lib/xschem/NOR2X2.sch
.subckt NOR2X2 Y B A
*.PININFO Y:O B:I A:I
M1 Y A GND GND nmos w=3u l=0.15u m=1
M3 Y B GND GND nmos w=3u l=0.15u m=1
M4 net1 A VDD VDD pmos w=2u l=0.15u m=1
M5 Y B net1 VDD pmos w=2u l=0.15u m=1
M2 Y B net2 VDD pmos w=2u l=0.15u m=1
M6 net2 A VDD VDD pmos w=2u l=0.15u m=1
.ends
.GLOBAL GND
.GLOBAL VDD
.end
