* SPICE3 file created from INVX1_square_elt.ext - technology: sky130A

.subckt INVX1_square_elt VSS VDD A Y
M1000 Y A VSS VSS nshort w=2.285u l=0.15u
+  ad=0.19p pd=1.76u as=1.12745p ps=8.86u
M1001 VDD A Y VDD pshort w=1.26u l=0.15u
+  ad=1.0584p pd=9.24u as=0.7308p ps=6.2u
M1002 Y A VDD VDD pshort w=1.26u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 VDD A Y VDD pshort w=1.26u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A VDD VDD pshort w=1.26u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
.ends
