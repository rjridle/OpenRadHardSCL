magic
tech sky130A
magscale 1 2
timestamp 1642387122
<< error_p >>
rect 91 318 92 319
rect 275 318 276 319
rect 92 317 93 318
rect 276 317 277 318
rect 107 287 108 288
rect 142 287 143 288
rect 291 287 292 288
rect 326 287 327 288
rect 107 184 108 185
rect 142 184 143 185
rect 291 184 292 185
rect 326 184 327 185
<< nwell >>
rect -36 591 470 1353
<< nmos >>
rect 62 318 92 368
rect 62 288 158 318
tri 158 288 188 318 sw
rect 246 318 276 368
rect 62 184 92 288
tri 92 272 108 288 nw
tri 142 272 158 288 ne
tri 92 184 108 200 sw
tri 142 184 158 200 se
rect 158 184 188 288
rect 246 288 342 318
tri 342 288 372 318 sw
tri 62 154 92 184 ne
rect 92 154 158 184
tri 158 154 188 184 nw
rect 246 184 276 288
tri 276 272 292 288 nw
tri 326 272 342 288 ne
tri 276 184 292 200 sw
tri 326 184 342 200 se
rect 342 184 372 288
tri 246 154 276 184 ne
rect 276 154 342 184
tri 342 154 372 184 nw
<< pmos >>
rect 62 629 92 1229
rect 150 629 180 1229
rect 246 629 276 1229
rect 334 629 364 1229
<< ndiff >>
rect 0 347 62 368
rect 0 313 16 347
rect 50 313 62 347
rect 92 347 246 368
rect 92 318 200 347
rect 0 279 62 313
tri 158 288 188 318 ne
rect 188 313 200 318
rect 234 313 246 347
rect 276 347 434 368
rect 276 318 384 347
rect 0 245 16 279
rect 50 245 62 279
rect 0 211 62 245
rect 0 177 16 211
rect 50 177 62 211
tri 92 272 108 288 se
rect 108 272 142 288
tri 142 272 158 288 sw
rect 92 240 158 272
rect 92 206 104 240
rect 138 206 158 240
rect 92 200 158 206
tri 92 184 108 200 ne
rect 108 184 142 200
tri 142 184 158 200 nw
rect 188 279 246 313
tri 342 288 372 318 ne
rect 372 313 384 318
rect 418 313 434 347
rect 188 245 200 279
rect 234 245 246 279
rect 188 211 246 245
rect 0 154 62 177
tri 62 154 92 184 sw
tri 158 154 188 184 se
rect 188 177 200 211
rect 234 177 246 211
tri 276 272 292 288 se
rect 292 272 326 288
tri 326 272 342 288 sw
rect 276 240 342 272
rect 276 206 288 240
rect 322 206 342 240
rect 276 200 342 206
tri 276 184 292 200 ne
rect 292 184 326 200
tri 326 184 342 200 nw
rect 372 279 434 313
rect 372 245 384 279
rect 418 245 434 279
rect 372 211 434 245
rect 188 154 246 177
tri 246 154 276 184 sw
tri 342 154 372 184 se
rect 372 177 384 211
rect 418 177 434 211
rect 372 154 434 177
rect 0 143 434 154
rect 0 109 16 143
rect 50 109 108 143
rect 142 109 200 143
rect 234 109 384 143
rect 418 109 434 143
rect 0 101 434 109
<< pdiff >>
rect 6 1213 62 1229
rect 6 1179 16 1213
rect 50 1179 62 1213
rect 6 1145 62 1179
rect 6 1111 16 1145
rect 50 1111 62 1145
rect 6 1077 62 1111
rect 6 1043 16 1077
rect 50 1043 62 1077
rect 6 1009 62 1043
rect 6 975 16 1009
rect 50 975 62 1009
rect 6 941 62 975
rect 6 907 16 941
rect 50 907 62 941
rect 6 873 62 907
rect 6 839 16 873
rect 50 839 62 873
rect 6 805 62 839
rect 6 771 16 805
rect 50 771 62 805
rect 6 737 62 771
rect 6 703 16 737
rect 50 703 62 737
rect 6 629 62 703
rect 92 1213 150 1229
rect 92 1179 104 1213
rect 138 1179 150 1213
rect 92 1145 150 1179
rect 92 1111 104 1145
rect 138 1111 150 1145
rect 92 1077 150 1111
rect 92 1043 104 1077
rect 138 1043 150 1077
rect 92 1009 150 1043
rect 92 975 104 1009
rect 138 975 150 1009
rect 92 941 150 975
rect 92 907 104 941
rect 138 907 150 941
rect 92 873 150 907
rect 92 839 104 873
rect 138 839 150 873
rect 92 805 150 839
rect 92 771 104 805
rect 138 771 150 805
rect 92 737 150 771
rect 92 703 104 737
rect 138 703 150 737
rect 92 629 150 703
rect 180 1213 246 1229
rect 180 1179 200 1213
rect 234 1179 246 1213
rect 180 1145 246 1179
rect 180 1111 200 1145
rect 234 1111 246 1145
rect 180 1077 246 1111
rect 180 1043 200 1077
rect 234 1043 246 1077
rect 180 1009 246 1043
rect 180 975 200 1009
rect 234 975 246 1009
rect 180 941 246 975
rect 180 907 200 941
rect 234 907 246 941
rect 180 873 246 907
rect 180 839 200 873
rect 234 839 246 873
rect 180 805 246 839
rect 180 771 200 805
rect 234 771 246 805
rect 180 737 246 771
rect 180 703 200 737
rect 234 703 246 737
rect 180 629 246 703
rect 276 1213 334 1229
rect 276 1179 288 1213
rect 322 1179 334 1213
rect 276 1145 334 1179
rect 276 1111 288 1145
rect 322 1111 334 1145
rect 276 1077 334 1111
rect 276 1043 288 1077
rect 322 1043 334 1077
rect 276 1009 334 1043
rect 276 975 288 1009
rect 322 975 334 1009
rect 276 941 334 975
rect 276 907 288 941
rect 322 907 334 941
rect 276 873 334 907
rect 276 839 288 873
rect 322 839 334 873
rect 276 805 334 839
rect 276 771 288 805
rect 322 771 334 805
rect 276 737 334 771
rect 276 703 288 737
rect 322 703 334 737
rect 276 629 334 703
rect 364 1213 418 1229
rect 364 1179 376 1213
rect 410 1179 418 1213
rect 364 1145 418 1179
rect 364 1111 376 1145
rect 410 1111 418 1145
rect 364 1077 418 1111
rect 364 1043 376 1077
rect 410 1043 418 1077
rect 364 1009 418 1043
rect 364 975 376 1009
rect 410 975 418 1009
rect 364 941 418 975
rect 364 907 376 941
rect 410 907 418 941
rect 364 873 418 907
rect 364 839 376 873
rect 410 839 418 873
rect 364 805 418 839
rect 364 771 376 805
rect 410 771 418 805
rect 364 737 418 771
rect 364 703 376 737
rect 410 703 418 737
rect 364 629 418 703
<< ndiffc >>
rect 16 313 50 347
rect 200 313 234 347
rect 16 245 50 279
rect 16 177 50 211
rect 104 206 138 240
rect 384 313 418 347
rect 200 245 234 279
rect 200 177 234 211
rect 288 206 322 240
rect 384 245 418 279
rect 384 177 418 211
rect 16 109 50 143
rect 108 109 142 143
rect 200 109 234 143
rect 384 109 418 143
<< pdiffc >>
rect 16 1179 50 1213
rect 16 1111 50 1145
rect 16 1043 50 1077
rect 16 975 50 1009
rect 16 907 50 941
rect 16 839 50 873
rect 16 771 50 805
rect 16 703 50 737
rect 104 1179 138 1213
rect 104 1111 138 1145
rect 104 1043 138 1077
rect 104 975 138 1009
rect 104 907 138 941
rect 104 839 138 873
rect 104 771 138 805
rect 104 703 138 737
rect 200 1179 234 1213
rect 200 1111 234 1145
rect 200 1043 234 1077
rect 200 975 234 1009
rect 200 907 234 941
rect 200 839 234 873
rect 200 771 234 805
rect 200 703 234 737
rect 288 1179 322 1213
rect 288 1111 322 1145
rect 288 1043 322 1077
rect 288 975 322 1009
rect 288 907 322 941
rect 288 839 322 873
rect 288 771 322 805
rect 288 703 322 737
rect 376 1179 410 1213
rect 376 1111 410 1145
rect 376 1043 410 1077
rect 376 975 410 1009
rect 376 907 410 941
rect 376 839 410 873
rect 376 771 410 805
rect 376 703 410 737
<< psubdiff >>
rect 0 13 24 47
rect 58 13 93 47
rect 127 13 169 47
rect 203 13 237 47
rect 271 13 306 47
rect 340 13 374 47
rect 408 13 434 47
<< nsubdiff >>
rect 0 1283 24 1317
rect 58 1283 92 1317
rect 126 1283 160 1317
rect 195 1283 229 1317
rect 263 1283 297 1317
rect 331 1283 434 1317
<< psubdiffcont >>
rect 24 13 58 47
rect 93 13 127 47
rect 169 13 203 47
rect 237 13 271 47
rect 306 13 340 47
rect 374 13 408 47
<< nsubdiffcont >>
rect 24 1283 58 1317
rect 92 1283 126 1317
rect 160 1283 195 1317
rect 229 1283 263 1317
rect 297 1283 331 1317
<< poly >>
rect 62 1229 92 1255
rect 150 1229 180 1255
rect 246 1229 276 1255
rect 334 1229 364 1255
rect 62 612 92 629
rect 150 612 180 629
rect 62 582 180 612
rect 246 612 276 629
rect 334 612 364 629
rect 246 582 364 612
rect 62 568 92 582
rect 26 552 92 568
rect 26 518 36 552
rect 70 518 92 552
rect 26 502 92 518
rect 62 368 92 502
rect 246 494 276 582
rect 213 478 276 494
rect 213 444 223 478
rect 257 444 276 478
rect 213 428 276 444
rect 246 368 276 428
<< polycont >>
rect 36 518 70 552
rect 223 444 257 478
<< locali >>
rect 0 1317 434 1332
rect 0 1283 24 1317
rect 58 1283 92 1317
rect 126 1283 160 1317
rect 195 1283 229 1317
rect 263 1283 297 1317
rect 331 1283 434 1317
rect 0 1270 434 1283
rect 16 1213 50 1270
rect 16 1145 50 1179
rect 16 1077 50 1111
rect 16 1009 50 1043
rect 16 941 50 975
rect 16 873 50 907
rect 16 805 50 839
rect 16 737 50 771
rect 16 687 50 703
rect 104 1213 138 1229
rect 104 1145 138 1179
rect 104 1077 138 1111
rect 104 1009 138 1043
rect 104 941 138 975
rect 104 873 138 907
rect 104 805 138 839
rect 104 737 138 771
rect 104 684 138 703
rect 200 1213 234 1270
rect 200 1145 234 1179
rect 200 1077 234 1111
rect 200 1009 234 1043
rect 200 941 234 975
rect 200 873 234 907
rect 200 805 234 839
rect 200 737 234 771
rect 200 687 234 703
rect 288 1213 322 1229
rect 288 1145 322 1179
rect 288 1077 322 1111
rect 288 1009 322 1043
rect 288 941 322 975
rect 288 873 322 907
rect 288 805 322 839
rect 288 737 322 771
rect 288 684 322 703
rect 376 1213 410 1270
rect 376 1145 410 1179
rect 376 1077 410 1111
rect 376 1009 410 1043
rect 376 941 410 975
rect 376 873 410 907
rect 376 805 410 839
rect 376 737 410 771
rect 36 552 70 568
rect 36 502 70 518
rect 16 347 50 363
rect 16 279 50 313
rect 16 211 50 245
rect 104 240 138 650
rect 376 627 410 703
rect 223 478 257 494
rect 223 428 257 444
rect 104 190 138 206
rect 200 347 418 363
rect 234 329 384 347
rect 200 279 234 313
rect 200 211 234 245
rect 16 143 50 177
rect 200 143 234 177
rect 288 240 322 280
rect 0 109 16 143
rect 50 109 108 143
rect 142 109 200 143
rect 234 109 250 143
rect 288 62 322 206
rect 384 279 418 313
rect 384 211 418 245
rect 384 143 418 177
rect 368 109 384 143
rect 418 109 434 143
rect 0 47 434 62
rect 0 13 24 47
rect 58 13 93 47
rect 127 13 169 47
rect 203 13 237 47
rect 271 13 306 47
rect 340 13 374 47
rect 408 13 434 47
rect 0 0 434 13
<< viali >>
rect 24 1283 58 1317
rect 92 1283 126 1317
rect 160 1283 195 1317
rect 229 1283 263 1317
rect 297 1283 331 1317
rect 104 650 138 684
rect 288 650 322 684
rect 36 518 70 552
rect 223 444 257 478
rect 24 13 58 47
rect 93 13 127 47
rect 169 13 203 47
rect 237 13 271 47
rect 306 13 340 47
rect 374 13 408 47
<< metal1 >>
rect 0 1317 434 1332
rect 0 1283 24 1317
rect 58 1283 92 1317
rect 126 1283 160 1317
rect 195 1283 229 1317
rect 263 1283 297 1317
rect 331 1283 434 1317
rect 0 1270 434 1283
rect 98 684 144 690
rect 282 684 328 690
rect 92 650 104 684
rect 138 650 288 684
rect 322 650 334 684
rect 98 649 328 650
rect 98 644 144 649
rect 282 644 328 649
rect 36 559 70 573
rect 26 552 76 559
rect 26 518 36 552
rect 70 518 76 552
rect 26 511 76 518
rect 36 497 70 511
rect 223 485 257 499
rect 213 478 263 485
rect 213 444 223 478
rect 257 444 263 478
rect 213 437 263 444
rect 223 423 257 437
rect 0 47 434 62
rect 0 13 24 47
rect 58 13 93 47
rect 127 13 169 47
rect 203 13 237 47
rect 271 13 306 47
rect 340 13 374 47
rect 408 13 434 47
rect 0 0 434 13
<< labels >>
rlabel metal1 161 1325 161 1325 1 VDD
rlabel metal1 148 31 148 31 1 VSS
rlabel metal1 36 518 70 552 1 A
rlabel metal1 223 444 257 478 1 B
rlabel metal1 104 650 138 684 1 YN
<< end >>
