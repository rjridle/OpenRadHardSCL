magic
tech sky130A
magscale 1 2
timestamp 1649530803
<< metal1 >>
rect 55 1505 89 1539
rect 2091 945 5719 979
rect 131 871 165 905
rect 1315 871 1349 905
rect 4098 871 4679 905
rect 1474 723 2349 757
rect 3691 723 3865 757
rect 6232 649 6367 683
rect 6530 649 7016 683
rect 7605 649 7639 683
rect 5421 575 6861 609
rect 2387 427 4822 461
rect 649 387 683 400
rect 5903 387 5937 401
rect 649 353 5937 387
rect 55 13 89 47
use li1_M1_contact  li1_M1_contact_3 pcells
timestamp 1648061256
transform 0 -1 666 1 0 444
box -53 -33 29 33
use xor2X1_pcell  xor2X1_pcell_0 pcells
timestamp 1648314317
transform 1 0 0 0 1 0
box -84 0 2304 1575
use xor2X1_pcell  xor2X1_pcell_1
timestamp 1648314317
transform 1 0 2220 0 1 0
box -84 0 2304 1575
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform -1 0 2072 0 -1 962
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_11
timestamp 1648061256
transform 1 0 2368 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_10
timestamp 1648061256
transform -1 0 2368 0 -1 444
box -53 -33 29 33
use and2x1_pcell  and2x1_pcell_0 pcells
timestamp 1648064711
transform 1 0 4440 0 1 0
box -84 0 1194 1575
use li1_M1_contact  li1_M1_contact_6
timestamp 1648061256
transform 1 0 4662 0 1 888
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_2
timestamp 1648061256
transform 1 0 5772 0 1 962
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_4
timestamp 1648061256
transform 0 -1 5920 1 0 444
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_12
timestamp 1648061256
transform -1 0 6512 0 -1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform 1 0 4810 0 1 444
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_8
timestamp 1648061256
transform 1 0 6882 0 1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_7
timestamp 1648061256
transform 1 0 7030 0 1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_5
timestamp 1648061256
transform -1 0 5402 0 -1 592
box -53 -33 29 33
use and2x1_pcell  and2x1_pcell_1
timestamp 1648064711
transform 1 0 5550 0 1 0
box -84 0 1194 1575
use or2x1_pcell  or2x1_pcell_0 pcells
timestamp 1648066488
transform 1 0 6660 0 1 0
box -84 0 1194 1575
use li1_M1_contact  li1_M1_contact_9
timestamp 1648061256
transform -1 0 7622 0 -1 666
box -53 -33 29 33
<< labels >>
rlabel metal1 3831 723 3865 757 1 SUM
port 1 n
rlabel metal1 7605 649 7639 683 1 COUT
port 2 n
rlabel metal1 131 871 165 905 1 A
port 3 n
rlabel metal1 1315 871 1349 905 1 B
port 4 n
rlabel metal1 4645 871 4679 905 1 CIN
port 5 n
rlabel metal1 55 1505 89 1539 1 VDD
port 6 n
rlabel metal1 55 13 89 47 1 VSS
port 7 n
<< end >>
