* SPICE3 file created from DLATCHN.ext - technology: sky130A

.subckt DLATCHN Q D GATE_N VDD GND
X0 GND a_185_209.t3 a_556_101.t0 GND sky130_fd_pr__nfet_01v8 ad=8.7946p pd=6.142u as=0p ps=0u w=0u l=0u
X1 VDD.t41 a_1771_1050.t5 a_2405_209.t2 C�Y�U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X2 VDD.t15 D.t0 a_1771_1050.t0 �eZ�U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X3 a_185_209.t2 D.t1 VDD.t7  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X4 a_1295_209.t2 a_661_1050.t5 VDD.t31  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X5 a_661_1050.t2 a_n259_209.t3 VDD.t17 VDD.t16 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X6 a_1771_1050.t4 D.t3 VDD.t35  L1�0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X7 Q.t1 a_3007_411.t5 a_2795_1051.t3 VDD.t42 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X8 a_3461_1051.t3 a_2405_209.t3 a_3007_411.t2  L1�0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X9 a_661_1050.t1 a_185_209.t4 VDD.t5 �K1�0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X10 a_1771_1050.t1 a_n259_209.t4 VDD.t19  L1�0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X11 a_2795_1051.t1 a_1295_209.t3 VDD.t1 �K1�0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X12 VDD.t21 Q.t4 a_3461_1051.t1  L1�0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X13 VDD.t13 GATE_N.t0 a_n259_209.t1 �K1�0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X14 a_2405_209.t1 a_1771_1050.t6 VDD.t39  L1�0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X15 GND a_n259_209.t7 a_1666_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X16 VDD.t11 a_185_209.t5 a_661_1050.t0 �K1�0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X17 VDD.t25 a_n259_209.t6 a_1771_1050.t2  L1�0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X18 VDD.t33 D.t5 a_185_209.t1 �K1�0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X19 VDD.t29 a_661_1050.t6 a_1295_209.t1  L1�0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X20 a_3007_411.t3 a_2405_209.t4 a_3461_1051.t2 �K1�0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X21 Q a_1295_209.t4 GND.t1 GND sky130_fd_pr__nfet_01v8 ad=3.582p pd=3.15u as=0p ps=0u w=0u l=0u
X22 a_2795_1051.t2 a_3007_411.t6 Q.t2  L1�0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X23 a_3461_1051.t0 Q.t6 VDD.t9 �K1�0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X24 Q a_3007_411.t4 GND.t3 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X25 a_n259_209.t2 GATE_N.t2 VDD.t27  L1�0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X26 VDD.t23 a_n259_209.t8 a_661_1050.t4 �K1�0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X27 VDD.t3 a_1295_209.t5 a_2795_1051.t0  L1�0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
C0 VDD GATE_N 0.38fF
C1 Q VDD 0.85fF
C2 VDD D 0.73fF
C3 D GATE_N 0.01fF
R0 a_1771_1050.n3 a_1771_1050.t5 512.525
R1 a_1771_1050.n3 a_1771_1050.t6 371.139
R2 a_1771_1050.n7 a_1771_1050.n5 284.244
R3 a_1771_1050.n4 a_1771_1050.t7 282.852
R4 a_1771_1050.n4 a_1771_1050.n3 247.347
R5 a_1771_1050.n5 a_1771_1050.n2 187.858
R6 a_1771_1050.n2 a_1771_1050.n1 157.964
R7 a_1771_1050.n2 a_1771_1050.n0 91.706
R8 a_1771_1050.n7 a_1771_1050.n6 15.218
R9 a_1771_1050.n0 a_1771_1050.t0 14.282
R10 a_1771_1050.n0 a_1771_1050.t4 14.282
R11 a_1771_1050.n1 a_1771_1050.t2 14.282
R12 a_1771_1050.n1 a_1771_1050.t1 14.282
R13 a_1771_1050.n8 a_1771_1050.n7 12.014
R14 a_1771_1050.n5 a_1771_1050.n4 10.343
R15 a_2405_209.n2 a_2405_209.t3 470.752
R16 a_2405_209.n2 a_2405_209.t4 384.527
R17 a_2405_209.n3 a_2405_209.t5 342.755
R18 a_2405_209.n6 a_2405_209.n4 328.169
R19 a_2405_209.n4 a_2405_209.n1 215.564
R20 a_2405_209.n3 a_2405_209.n2 155.073
R21 a_2405_209.n6 a_2405_209.n5 30
R22 a_2405_209.n7 a_2405_209.n0 24.383
R23 a_2405_209.n7 a_2405_209.n6 23.684
R24 a_2405_209.n1 a_2405_209.t2 14.282
R25 a_2405_209.n1 a_2405_209.t1 14.282
R26 a_2405_209.n4 a_2405_209.n3 13.607
R27 VDD.n249 VDD.n238 144.705
R28 VDD.n306 VDD.n299 144.705
R29 VDD.n363 VDD.n356 144.705
R30 VDD.n176 VDD.n169 144.705
R31 VDD.n391 VDD.n384 144.705
R32 VDD.n132 VDD.n125 144.705
R33 VDD.n77 VDD.n66 144.705
R34 VDD.n331 VDD.t23 143.754
R35 VDD.n181 VDD.t15 143.754
R36 VDD.n222 VDD.t27 135.17
R37 VDD.n229 VDD.t13 135.17
R38 VDD.n265 VDD.t7 135.17
R39 VDD.n274 VDD.t33 135.17
R40 VDD.n309 VDD.t5 135.17
R41 VDD.n368 VDD.t31 135.17
R42 VDD.n375 VDD.t29 135.17
R43 VDD.n410 VDD.t19 135.17
R44 VDD.n144 VDD.t39 135.17
R45 VDD.n135 VDD.t41 135.17
R46 VDD.n96 VDD.n95 129.849
R47 VDD.n40 VDD.n39 129.849
R48 VDD.n323 VDD.n322 129.472
R49 VDD.n190 VDD.n189 129.472
R50 VDD.n62 VDD.n61 92.5
R51 VDD.n60 VDD.n59 92.5
R52 VDD.n58 VDD.n57 92.5
R53 VDD.n56 VDD.n55 92.5
R54 VDD.n64 VDD.n63 92.5
R55 VDD.n121 VDD.n120 92.5
R56 VDD.n119 VDD.n118 92.5
R57 VDD.n117 VDD.n116 92.5
R58 VDD.n115 VDD.n114 92.5
R59 VDD.n123 VDD.n122 92.5
R60 VDD.n165 VDD.n164 92.5
R61 VDD.n163 VDD.n162 92.5
R62 VDD.n161 VDD.n160 92.5
R63 VDD.n159 VDD.n158 92.5
R64 VDD.n167 VDD.n166 92.5
R65 VDD.n404 VDD.n403 92.5
R66 VDD.n402 VDD.n401 92.5
R67 VDD.n400 VDD.n399 92.5
R68 VDD.n398 VDD.n397 92.5
R69 VDD.n406 VDD.n405 92.5
R70 VDD.n352 VDD.n351 92.5
R71 VDD.n350 VDD.n349 92.5
R72 VDD.n348 VDD.n347 92.5
R73 VDD.n346 VDD.n345 92.5
R74 VDD.n354 VDD.n353 92.5
R75 VDD.n295 VDD.n294 92.5
R76 VDD.n293 VDD.n292 92.5
R77 VDD.n291 VDD.n290 92.5
R78 VDD.n289 VDD.n288 92.5
R79 VDD.n297 VDD.n296 92.5
R80 VDD.n259 VDD.n258 92.5
R81 VDD.n257 VDD.n256 92.5
R82 VDD.n255 VDD.n254 92.5
R83 VDD.n253 VDD.n252 92.5
R84 VDD.n261 VDD.n260 92.5
R85 VDD.n208 VDD.n207 92.5
R86 VDD.n206 VDD.n205 92.5
R87 VDD.n204 VDD.n203 92.5
R88 VDD.n202 VDD.n201 92.5
R89 VDD.n210 VDD.n209 92.5
R90 VDD.n14 VDD.n1 92.5
R91 VDD.n5 VDD.n4 92.5
R92 VDD.n7 VDD.n6 92.5
R93 VDD.n9 VDD.n8 92.5
R94 VDD.n11 VDD.n10 92.5
R95 VDD.n13 VDD.n12 92.5
R96 VDD.n21 VDD.n20 92.059
R97 VDD.n76 VDD.n75 92.059
R98 VDD.n131 VDD.n130 92.059
R99 VDD.n175 VDD.n174 92.059
R100 VDD.n390 VDD.n389 92.059
R101 VDD.n362 VDD.n361 92.059
R102 VDD.n305 VDD.n304 92.059
R103 VDD.n248 VDD.n247 92.059
R104 VDD.n216 VDD.n215 92.059
R105 VDD.n20 VDD.n16 67.194
R106 VDD.n20 VDD.n17 67.194
R107 VDD.n20 VDD.n18 67.194
R108 VDD.n20 VDD.n19 67.194
R109 VDD.n200 VDD.n199 44.141
R110 VDD.n287 VDD.n286 44.141
R111 VDD.n344 VDD.n343 44.141
R112 VDD.n396 VDD.n395 44.141
R113 VDD.n157 VDD.n156 44.141
R114 VDD.n113 VDD.n112 44.141
R115 VDD.n5 VDD.n3 44.141
R116 VDD.n286 VDD.n284 44.107
R117 VDD.n343 VDD.n341 44.107
R118 VDD.n395 VDD.n393 44.107
R119 VDD.n156 VDD.n154 44.107
R120 VDD.n112 VDD.n110 44.107
R121 VDD.n199 VDD.n197 44.107
R122 VDD.n3 VDD.n2 44.107
R123 VDD.n136 C�Y�U 43.472
R124 VDD.n145  L1�0 43.472
R125 VDD.n376  L1�0 43.472
R126 VDD.n366 �c�Z�U 43.472
R127 VDD.n275 �K1�0 43.472
R128 VDD.n266  43.472
R129 VDD.n230 �K1�0 43.472
R130 VDD.n220  L1�0 43.472
R131 VDD.n20 VDD.n15 41.052
R132 VDD.n70 VDD.n68 39.742
R133 VDD.n70 VDD.n69 39.742
R134 VDD.n72 VDD.n71 39.742
R135 VDD.n127 VDD.n126 39.742
R136 VDD.n171 VDD.n170 39.742
R137 VDD.n386 VDD.n385 39.742
R138 VDD.n358 VDD.n357 39.742
R139 VDD.n301 VDD.n300 39.742
R140 VDD.n212 VDD.n211 39.742
R141 VDD.n246 VDD.n243 39.742
R142 VDD.n246 VDD.n245 39.742
R143 VDD.n242 VDD.n241 39.742
R144 VDD.n112 VDD.n111 38
R145 VDD.n156 VDD.n155 38
R146 VDD.n395 VDD.n394 38
R147 VDD.n343 VDD.n342 38
R148 VDD.n286 VDD.n285 38
R149 VDD.n199 VDD.n198 38
R150 VDD.n284 VDD.n283 36.774
R151 VDD.n341 VDD.n340 36.774
R152 VDD.n393 VDD.n392 36.774
R153 VDD.n154 VDD.n153 36.774
R154 VDD.n110 VDD.n109 36.774
R155 VDD.n68 VDD.n67 36.774
R156 VDD.n245 VDD.n244 36.774
R157 VDD.n1 VDD.n0 30.923
R158 VDD.n75 VDD.n73 26.38
R159 VDD.n75 VDD.n72 26.38
R160 VDD.n75 VDD.n70 26.38
R161 VDD.n75 VDD.n74 26.38
R162 VDD.n130 VDD.n128 26.38
R163 VDD.n130 VDD.n127 26.38
R164 VDD.n130 VDD.n129 26.38
R165 VDD.n174 VDD.n172 26.38
R166 VDD.n174 VDD.n171 26.38
R167 VDD.n174 VDD.n173 26.38
R168 VDD.n389 VDD.n387 26.38
R169 VDD.n389 VDD.n386 26.38
R170 VDD.n389 VDD.n388 26.38
R171 VDD.n361 VDD.n359 26.38
R172 VDD.n361 VDD.n358 26.38
R173 VDD.n361 VDD.n360 26.38
R174 VDD.n304 VDD.n302 26.38
R175 VDD.n304 VDD.n301 26.38
R176 VDD.n304 VDD.n303 26.38
R177 VDD.n215 VDD.n213 26.38
R178 VDD.n215 VDD.n212 26.38
R179 VDD.n215 VDD.n214 26.38
R180 VDD.n247 VDD.n246 26.38
R181 VDD.n247 VDD.n242 26.38
R182 VDD.n247 VDD.n240 26.38
R183 VDD.n247 VDD.n239 26.38
R184 VDD.n218 VDD.n210 22.915
R185 VDD.n23 VDD.n14 22.915
R186 VDD.n28  L1�0 20.457
R187 VDD.n84  L1�0 20.457
R188 VDD.n184 �eZ�U 20.457
R189 VDD.n327 �K1�0 20.457
R190 VDD.n41  L1�0 17.9
R191 VDD.n97  L1�0 17.9
R192 VDD.n415  L1�0 17.9
R193 VDD.n314 �K1�0 17.9
R194 VDD.n210 VDD.n208 14.864
R195 VDD.n208 VDD.n206 14.864
R196 VDD.n206 VDD.n204 14.864
R197 VDD.n204 VDD.n202 14.864
R198 VDD.n202 VDD.n200 14.864
R199 VDD.n297 VDD.n295 14.864
R200 VDD.n295 VDD.n293 14.864
R201 VDD.n293 VDD.n291 14.864
R202 VDD.n291 VDD.n289 14.864
R203 VDD.n289 VDD.n287 14.864
R204 VDD.n354 VDD.n352 14.864
R205 VDD.n352 VDD.n350 14.864
R206 VDD.n350 VDD.n348 14.864
R207 VDD.n348 VDD.n346 14.864
R208 VDD.n346 VDD.n344 14.864
R209 VDD.n406 VDD.n404 14.864
R210 VDD.n404 VDD.n402 14.864
R211 VDD.n402 VDD.n400 14.864
R212 VDD.n400 VDD.n398 14.864
R213 VDD.n398 VDD.n396 14.864
R214 VDD.n167 VDD.n165 14.864
R215 VDD.n165 VDD.n163 14.864
R216 VDD.n163 VDD.n161 14.864
R217 VDD.n161 VDD.n159 14.864
R218 VDD.n159 VDD.n157 14.864
R219 VDD.n123 VDD.n121 14.864
R220 VDD.n121 VDD.n119 14.864
R221 VDD.n119 VDD.n117 14.864
R222 VDD.n117 VDD.n115 14.864
R223 VDD.n115 VDD.n113 14.864
R224 VDD.n64 VDD.n62 14.864
R225 VDD.n62 VDD.n60 14.864
R226 VDD.n60 VDD.n58 14.864
R227 VDD.n58 VDD.n56 14.864
R228 VDD.n56 VDD.n54 14.864
R229 VDD.n54 VDD.n53 14.864
R230 VDD.n261 VDD.n259 14.864
R231 VDD.n259 VDD.n257 14.864
R232 VDD.n257 VDD.n255 14.864
R233 VDD.n255 VDD.n253 14.864
R234 VDD.n253 VDD.n251 14.864
R235 VDD.n251 VDD.n250 14.864
R236 VDD.n14 VDD.n13 14.864
R237 VDD.n13 VDD.n11 14.864
R238 VDD.n11 VDD.n9 14.864
R239 VDD.n9 VDD.n7 14.864
R240 VDD.n7 VDD.n5 14.864
R241 VDD.n78 VDD.n65 14.864
R242 VDD.n133 VDD.n124 14.864
R243 VDD.n177 VDD.n168 14.864
R244 VDD.n408 VDD.n407 14.864
R245 VDD.n364 VDD.n355 14.864
R246 VDD.n307 VDD.n298 14.864
R247 VDD.n263 VDD.n262 14.864
R248 VDD.n322 VDD.t17 14.282
R249 VDD.n322 VDD.t11 14.282
R250 VDD.n189 VDD.t35 14.282
R251 VDD.n189 VDD.t25 14.282
R252 VDD.n95 VDD.t1 14.282
R253 VDD.n95 VDD.t3 14.282
R254 VDD.n39 VDD.t9 14.282
R255 VDD.n39 VDD.t21 14.282
R256 VDD.n191 VDD.n190 9.083
R257 VDD.n325 VDD.n323 9.083
R258 VDD.n23 VDD.n22 8.855
R259 VDD.n22 VDD.n21 8.855
R260 VDD.n26 VDD.n25 8.855
R261 VDD.n25 VDD.n24 8.855
R262 VDD.n30 VDD.n29 8.855
R263 VDD.n29 VDD.n28 8.855
R264 VDD.n33 VDD.n32 8.855
R265 VDD.n32 �K1�0 8.855
R266 VDD.n37 VDD.n36 8.855
R267 VDD.n36 VDD.n35 8.855
R268 VDD.n43 VDD.n42 8.855
R269 VDD.n42 VDD.n41 8.855
R270 VDD.n47 VDD.n46 8.855
R271 VDD.n46 VDD.n45 8.855
R272 VDD.n51 VDD.n50 8.855
R273 VDD.n50 VDD.n49 8.855
R274 VDD.n78 VDD.n77 8.855
R275 VDD.n77 VDD.n76 8.855
R276 VDD.n82 VDD.n81 8.855
R277 VDD.n81 VDD.n80 8.855
R278 VDD.n86 VDD.n85 8.855
R279 VDD.n85 VDD.n84 8.855
R280 VDD.n89 VDD.n88 8.855
R281 VDD.n88 VDD.t42 8.855
R282 VDD.n93 VDD.n92 8.855
R283 VDD.n92 VDD.n91 8.855
R284 VDD.n99 VDD.n98 8.855
R285 VDD.n98 VDD.n97 8.855
R286 VDD.n103 VDD.n102 8.855
R287 VDD.n102 VDD.n101 8.855
R288 VDD.n107 VDD.n106 8.855
R289 VDD.n106 VDD.n105 8.855
R290 VDD.n133 VDD.n132 8.855
R291 VDD.n132 VDD.n131 8.855
R292 VDD.n138 VDD.n137 8.855
R293 VDD.n137 VDD.n136 8.855
R294 VDD.n142 VDD.n141 8.855
R295 VDD.n141 VDD.n140 8.855
R296 VDD.n147 VDD.n146 8.855
R297 VDD.n146 VDD.n145 8.855
R298 VDD.n151 VDD.n150 8.855
R299 VDD.n150 VDD.n149 8.855
R300 VDD.n177 VDD.n176 8.855
R301 VDD.n176 VDD.n175 8.855
R302 VDD.n182 VDD.n180 8.855
R303 VDD.n180 VDD.n179 8.855
R304 VDD.n186 VDD.n185 8.855
R305 VDD.n185 VDD.n184 8.855
R306 VDD.n191 VDD.n188 8.855
R307 VDD.n188  L1�0 8.855
R308 VDD.n195 VDD.n194 8.855
R309 VDD.n194 VDD.n193 8.855
R310 VDD.n417 VDD.n416 8.855
R311 VDD.n416 VDD.n415 8.855
R312 VDD.n413 VDD.n412 8.855
R313 VDD.n412 VDD.n411 8.855
R314 VDD.n408 VDD.n391 8.855
R315 VDD.n391 VDD.n390 8.855
R316 VDD.n382 VDD.n381 8.855
R317 VDD.n381 VDD.n380 8.855
R318 VDD.n378 VDD.n377 8.855
R319 VDD.n377 VDD.n376 8.855
R320 VDD.n373 VDD.n372 8.855
R321 VDD.n372 VDD.n371 8.855
R322 VDD.n369 VDD.n367 8.855
R323 VDD.n367 VDD.n366 8.855
R324 VDD.n364 VDD.n363 8.855
R325 VDD.n363 VDD.n362 8.855
R326 VDD.n338 VDD.n337 8.855
R327 VDD.n337 VDD.n336 8.855
R328 VDD.n334 VDD.n333 8.855
R329 VDD.n333 VDD.n332 8.855
R330 VDD.n329 VDD.n328 8.855
R331 VDD.n328 VDD.n327 8.855
R332 VDD.n325 VDD.n324 8.855
R333 VDD.n324 VDD.t16 8.855
R334 VDD.n320 VDD.n319 8.855
R335 VDD.n319 VDD.n318 8.855
R336 VDD.n316 VDD.n315 8.855
R337 VDD.n315 VDD.n314 8.855
R338 VDD.n312 VDD.n311 8.855
R339 VDD.n311 VDD.n310 8.855
R340 VDD.n307 VDD.n306 8.855
R341 VDD.n306 VDD.n305 8.855
R342 VDD.n281 VDD.n280 8.855
R343 VDD.n280 VDD.n279 8.855
R344 VDD.n277 VDD.n276 8.855
R345 VDD.n276 VDD.n275 8.855
R346 VDD.n272 VDD.n271 8.855
R347 VDD.n271 VDD.n270 8.855
R348 VDD.n268 VDD.n267 8.855
R349 VDD.n267 VDD.n266 8.855
R350 VDD.n263 VDD.n249 8.855
R351 VDD.n249 VDD.n248 8.855
R352 VDD.n236 VDD.n235 8.855
R353 VDD.n235 VDD.n234 8.855
R354 VDD.n232 VDD.n231 8.855
R355 VDD.n231 VDD.n230 8.855
R356 VDD.n227 VDD.n226 8.855
R357 VDD.n226 VDD.n225 8.855
R358 VDD.n223 VDD.n221 8.855
R359 VDD.n221 VDD.n220 8.855
R360 VDD.n218 VDD.n217 8.855
R361 VDD.n217 VDD.n216 8.855
R362 VDD.n298 VDD.n297 8.051
R363 VDD.n355 VDD.n354 8.051
R364 VDD.n407 VDD.n406 8.051
R365 VDD.n168 VDD.n167 8.051
R366 VDD.n124 VDD.n123 8.051
R367 VDD.n65 VDD.n64 8.051
R368 VDD.n262 VDD.n261 8.051
R369 VDD.n43 VDD.n40 6.193
R370 VDD.n99 VDD.n96 6.193
R371 VDD.n31 VDD.n30 4.65
R372 VDD.n34 VDD.n33 4.65
R373 VDD.n38 VDD.n37 4.65
R374 VDD.n44 VDD.n43 4.65
R375 VDD.n48 VDD.n47 4.65
R376 VDD.n52 VDD.n51 4.65
R377 VDD.n79 VDD.n78 4.65
R378 VDD.n83 VDD.n82 4.65
R379 VDD.n87 VDD.n86 4.65
R380 VDD.n90 VDD.n89 4.65
R381 VDD.n94 VDD.n93 4.65
R382 VDD.n100 VDD.n99 4.65
R383 VDD.n104 VDD.n103 4.65
R384 VDD.n108 VDD.n107 4.65
R385 VDD.n134 VDD.n133 4.65
R386 VDD.n139 VDD.n138 4.65
R387 VDD.n143 VDD.n142 4.65
R388 VDD.n148 VDD.n147 4.65
R389 VDD.n152 VDD.n151 4.65
R390 VDD.n178 VDD.n177 4.65
R391 VDD.n183 VDD.n182 4.65
R392 VDD.n187 VDD.n186 4.65
R393 VDD.n192 VDD.n191 4.65
R394 VDD.n196 VDD.n195 4.65
R395 VDD.n418 VDD.n417 4.65
R396 VDD.n414 VDD.n413 4.65
R397 VDD.n409 VDD.n408 4.65
R398 VDD.n383 VDD.n382 4.65
R399 VDD.n379 VDD.n378 4.65
R400 VDD.n374 VDD.n373 4.65
R401 VDD.n370 VDD.n369 4.65
R402 VDD.n365 VDD.n364 4.65
R403 VDD.n339 VDD.n338 4.65
R404 VDD.n335 VDD.n334 4.65
R405 VDD.n330 VDD.n329 4.65
R406 VDD.n326 VDD.n325 4.65
R407 VDD.n321 VDD.n320 4.65
R408 VDD.n317 VDD.n316 4.65
R409 VDD.n313 VDD.n312 4.65
R410 VDD.n308 VDD.n307 4.65
R411 VDD.n282 VDD.n281 4.65
R412 VDD.n278 VDD.n277 4.65
R413 VDD.n273 VDD.n272 4.65
R414 VDD.n269 VDD.n268 4.65
R415 VDD.n264 VDD.n263 4.65
R416 VDD.n237 VDD.n236 4.65
R417 VDD.n233 VDD.n232 4.65
R418 VDD.n228 VDD.n227 4.65
R419 VDD.n224 VDD.n223 4.65
R420 VDD.n219 VDD.n218 4.65
R421 VDD.n27 VDD.n23 2.933
R422 VDD.n413 VDD.n410 2.89
R423 VDD.n312 VDD.n309 2.89
R424 VDD.n27 VDD.n26 2.844
R425 VDD.n35 �K1�0 2.557
R426 VDD.n91 �K1�0 2.557
R427 VDD.n193  L1�0 2.557
R428 VDD.n318 �K1�0 2.557
R429 VDD.n182 VDD.n181 2.477
R430 VDD.n334 VDD.n331 2.477
R431 VDD.n138 VDD.n135 2.064
R432 VDD.n147 VDD.n144 2.064
R433 VDD.n378 VDD.n375 2.064
R434 VDD.n369 VDD.n368 2.064
R435 VDD.n277 VDD.n274 2.064
R436 VDD.n268 VDD.n265 2.064
R437 VDD.n232 VDD.n229 2.064
R438 VDD.n223 VDD.n222 2.064
R439 VDD.n31 VDD.n27 1.063
R440 VDD.n79 VDD.n52 0.29
R441 VDD.n134 VDD.n108 0.29
R442 VDD.n178 VDD.n152 0.29
R443 VDD.n409 VDD.n383 0.29
R444 VDD.n365 VDD.n339 0.29
R445 VDD.n308 VDD.n282 0.29
R446 VDD.n264 VDD.n237 0.29
R447 VDD.n219 VDD 0.207
R448 VDD.n38 VDD.n34 0.181
R449 VDD.n94 VDD.n90 0.181
R450 VDD.n196 VDD.n192 0.181
R451 VDD.n326 VDD.n321 0.181
R452 VDD.n143 VDD.n139 0.157
R453 VDD.n148 VDD.n143 0.157
R454 VDD.n379 VDD.n374 0.157
R455 VDD.n374 VDD.n370 0.157
R456 VDD.n278 VDD.n273 0.157
R457 VDD.n273 VDD.n269 0.157
R458 VDD.n233 VDD.n228 0.157
R459 VDD.n228 VDD.n224 0.157
R460 VDD.n34 VDD.n31 0.145
R461 VDD.n44 VDD.n38 0.145
R462 VDD.n48 VDD.n44 0.145
R463 VDD.n52 VDD.n48 0.145
R464 VDD.n83 VDD.n79 0.145
R465 VDD.n87 VDD.n83 0.145
R466 VDD.n90 VDD.n87 0.145
R467 VDD.n100 VDD.n94 0.145
R468 VDD.n104 VDD.n100 0.145
R469 VDD.n108 VDD.n104 0.145
R470 VDD.n139 VDD.n134 0.145
R471 VDD.n152 VDD.n148 0.145
R472 VDD.n183 VDD.n178 0.145
R473 VDD.n187 VDD.n183 0.145
R474 VDD.n192 VDD.n187 0.145
R475 VDD.n418 VDD.n414 0.145
R476 VDD.n414 VDD.n409 0.145
R477 VDD.n383 VDD.n379 0.145
R478 VDD.n370 VDD.n365 0.145
R479 VDD.n339 VDD.n335 0.145
R480 VDD.n335 VDD.n330 0.145
R481 VDD.n330 VDD.n326 0.145
R482 VDD.n321 VDD.n317 0.145
R483 VDD.n317 VDD.n313 0.145
R484 VDD.n313 VDD.n308 0.145
R485 VDD.n282 VDD.n278 0.145
R486 VDD.n269 VDD.n264 0.145
R487 VDD.n237 VDD.n233 0.145
R488 VDD.n224 VDD.n219 0.145
R489 VDD VDD.n196 0.133
R490 VDD VDD.n418 0.012
R491 a_3007_411.n2 a_3007_411.t6 470.752
R492 a_3007_411.n2 a_3007_411.t5 384.527
R493 a_3007_411.n3 a_3007_411.t4 314.896
R494 a_3007_411.n4 a_3007_411.n1 260.107
R495 a_3007_411.n9 a_3007_411.n8 208.452
R496 a_3007_411.n3 a_3007_411.n2 182.932
R497 a_3007_411.n9 a_3007_411.n4 170.164
R498 a_3007_411.n11 a_3007_411.n9 135.417
R499 a_3007_411.n12 a_3007_411.n0 55.263
R500 a_3007_411.n8 a_3007_411.n7 30
R501 a_3007_411.n11 a_3007_411.n10 30
R502 a_3007_411.n12 a_3007_411.n11 25.263
R503 a_3007_411.n6 a_3007_411.n5 24.383
R504 a_3007_411.n8 a_3007_411.n6 23.684
R505 a_3007_411.n1 a_3007_411.t2 14.282
R506 a_3007_411.n1 a_3007_411.t3 14.282
R507 a_3007_411.n4 a_3007_411.n3 12.247
R508 GND.n170 GND.n169 237.558
R509 GND.n203 GND.n202 237.558
R510 GND.n233 GND.n232 237.558
R511 GND.n123 GND.n122 237.558
R512 GND.n266 GND.n265 237.558
R513 GND.n90 GND.n89 237.558
R514 GND.n43 GND.n42 237.558
R515 GND.n40 GND.n39 210.82
R516 GND.n172 GND.n171 210.82
R517 GND.n205 GND.n204 210.82
R518 GND.n235 GND.n234 210.82
R519 GND.n268 GND.n267 210.82
R520 GND.n120 GND.n119 210.82
R521 GND.n87 GND.n86 210.82
R522 GND.n213 GND.n212 172.612
R523 GND.n279 GND.n278 151.605
R524 GND.n161 GND.n160 120.01
R525 GND.n55 GND.n54 92.5
R526 GND.n71 GND.n70 92.5
R527 GND.n159 GND.n158 92.5
R528 GND.n152 GND.n151 92.5
R529 GND.n78 GND.t1 45.413
R530 GND.n145 GND.t2 45.413
R531 GND.n19 GND.n18 40.431
R532 GND.n65 GND.n64 40.431
R533 GND.n4 GND.n3 40.003
R534 GND.n78 GND.n77 39.307
R535 GND.n145 GND.n144 39.307
R536 GND.n32 GND.n31 37.582
R537 GND.n112 GND.n111 37.582
R538 GND.n246 GND.n245 37.582
R539 GND.n183 GND.n182 37.582
R540 GND.n47 GND.n46 35.865
R541 GND.t11 GND.n109 32.601
R542 GND.t8 GND.n243 32.601
R543 GND.t9 GND.n180 32.601
R544 GND.n48 GND.n47 28.503
R545 GND.n278 GND.n277 28.421
R546 GND.n278 GND.n276 25.263
R547 GND.n276 GND.n275 24.383
R548 GND.n79 GND.n78 23.77
R549 GND.n146 GND.n145 23.77
R550 GND.n109 GND.n108 21.734
R551 GND.n243 GND.n242 21.734
R552 GND.n180 GND.n179 21.734
R553 GND.n25 GND.n24 20.705
R554 GND.n20 GND.n19 20.705
R555 GND.n11 GND.n10 20.705
R556 GND.n5 GND.n4 20.705
R557 GND.n33 GND.n32 20.705
R558 GND.n72 GND.n71 20.705
R559 GND.n66 GND.n65 20.705
R560 GND.n56 GND.n55 20.705
R561 GND.n49 GND.n48 20.705
R562 GND.n80 GND.n79 20.705
R563 GND.n95 GND.n94 20.705
R564 GND.n101 GND.n100 20.705
R565 GND.n113 GND.n112 20.705
R566 GND.n258 GND.n257 20.705
R567 GND.n252 GND.n251 20.705
R568 GND.n247 GND.n246 20.705
R569 GND.n195 GND.n194 20.705
R570 GND.n189 GND.n188 20.705
R571 GND.n184 GND.n183 20.705
R572 GND.n162 GND.n161 20.705
R573 GND.n154 GND.n153 20.705
R574 GND.n147 GND.n146 20.705
R575 GND.n94 GND.n93 19.952
R576 GND.n257 GND.n256 19.952
R577 GND.n194 GND.n193 19.952
R578 GND.n161 GND.n159 19.952
R579 GND.n41 GND.n40 18.953
R580 GND.n173 GND.n172 18.953
R581 GND.n206 GND.n205 18.953
R582 GND.n236 GND.n235 18.953
R583 GND.n269 GND.n268 18.953
R584 GND.n121 GND.n120 18.953
R585 GND.n88 GND.n87 18.953
R586 GND.n3 GND.n2 17.258
R587 GND.n31 GND.t0 15.644
R588 GND.n111 GND.t11 15.644
R589 GND.n245 GND.t8 15.644
R590 GND.n182 GND.t9 15.644
R591 GND.n44 GND.n41 14.864
R592 GND.n91 GND.n88 14.864
R593 GND.n124 GND.n121 14.864
R594 GND.n270 GND.n269 14.864
R595 GND.n237 GND.n236 14.864
R596 GND.n207 GND.n206 14.864
R597 GND.n174 GND.n173 14.864
R598 GND.n18 GND.t10 13.654
R599 GND.n64 GND.t3 13.654
R600 GND.n64 GND.n63 13.654
R601 GND.n31 GND.n30 13.541
R602 GND.n111 GND.n110 13.541
R603 GND.n245 GND.n244 13.541
R604 GND.n182 GND.n181 13.541
R605 GND.n22 GND.n20 9.29
R606 GND.n68 GND.n66 9.29
R607 GND.n148 GND.n141 9.154
R608 GND.n156 GND.n155 9.154
R609 GND.n164 GND.n163 9.154
R610 GND.n167 GND.n166 9.154
R611 GND.n174 GND.n170 9.154
R612 GND.n185 GND.n176 9.154
R613 GND.n191 GND.n190 9.154
R614 GND.n197 GND.n196 9.154
R615 GND.n200 GND.n199 9.154
R616 GND.n207 GND.n203 9.154
R617 GND.n210 GND.n209 9.154
R618 GND.n215 GND.n214 9.154
R619 GND.n218 GND.n217 9.154
R620 GND.n221 GND.n220 9.154
R621 GND.n224 GND.n223 9.154
R622 GND.n227 GND.n226 9.154
R623 GND.n230 GND.n229 9.154
R624 GND.n237 GND.n233 9.154
R625 GND.n248 GND.n239 9.154
R626 GND.n254 GND.n253 9.154
R627 GND.n260 GND.n259 9.154
R628 GND.n263 GND.n262 9.154
R629 GND.n270 GND.n266 9.154
R630 GND.n273 GND.n272 9.154
R631 GND.n281 GND.n280 9.154
R632 GND.n136 GND.n135 9.154
R633 GND.n133 GND.n132 9.154
R634 GND.n130 GND.n129 9.154
R635 GND.n127 GND.n126 9.154
R636 GND.n124 GND.n123 9.154
R637 GND.n117 GND.n116 9.154
R638 GND.n114 GND.n105 9.154
R639 GND.n103 GND.n102 9.154
R640 GND.n97 GND.n96 9.154
R641 GND.n91 GND.n90 9.154
R642 GND.n84 GND.n83 9.154
R643 GND.n81 GND.n76 9.154
R644 GND.n74 GND.n73 9.154
R645 GND.n68 GND.n67 9.154
R646 GND.n60 GND.n59 9.154
R647 GND.n57 GND.n53 9.154
R648 GND.n51 GND.n50 9.154
R649 GND.n44 GND.n43 9.154
R650 GND.n37 GND.n36 9.154
R651 GND.n34 GND.n29 9.154
R652 GND.n27 GND.n26 9.154
R653 GND.n22 GND.n21 9.154
R654 GND.n15 GND.n14 9.154
R655 GND.n12 GND.n9 9.154
R656 GND.n7 GND.n6 9.154
R657 GND.t10 GND.n17 7.04
R658 GND.t3 GND.n62 7.04
R659 GND.n8 GND.n1 4.795
R660 GND.n140 GND.n139 4.65
R661 GND.n8 GND.n7 4.65
R662 GND.n13 GND.n12 4.65
R663 GND.n16 GND.n15 4.65
R664 GND.n23 GND.n22 4.65
R665 GND.n28 GND.n27 4.65
R666 GND.n35 GND.n34 4.65
R667 GND.n38 GND.n37 4.65
R668 GND.n45 GND.n44 4.65
R669 GND.n52 GND.n51 4.65
R670 GND.n58 GND.n57 4.65
R671 GND.n61 GND.n60 4.65
R672 GND.n69 GND.n68 4.65
R673 GND.n75 GND.n74 4.65
R674 GND.n82 GND.n81 4.65
R675 GND.n85 GND.n84 4.65
R676 GND.n92 GND.n91 4.65
R677 GND.n98 GND.n97 4.65
R678 GND.n104 GND.n103 4.65
R679 GND.n115 GND.n114 4.65
R680 GND.n118 GND.n117 4.65
R681 GND.n125 GND.n124 4.65
R682 GND.n128 GND.n127 4.65
R683 GND.n131 GND.n130 4.65
R684 GND.n134 GND.n133 4.65
R685 GND.n137 GND.n136 4.65
R686 GND.n282 GND.n281 4.65
R687 GND.n274 GND.n273 4.65
R688 GND.n271 GND.n270 4.65
R689 GND.n264 GND.n263 4.65
R690 GND.n261 GND.n260 4.65
R691 GND.n255 GND.n254 4.65
R692 GND.n249 GND.n248 4.65
R693 GND.n238 GND.n237 4.65
R694 GND.n231 GND.n230 4.65
R695 GND.n228 GND.n227 4.65
R696 GND.n225 GND.n224 4.65
R697 GND.n222 GND.n221 4.65
R698 GND.n219 GND.n218 4.65
R699 GND.n216 GND.n215 4.65
R700 GND.n211 GND.n210 4.65
R701 GND.n208 GND.n207 4.65
R702 GND.n201 GND.n200 4.65
R703 GND.n198 GND.n197 4.65
R704 GND.n192 GND.n191 4.65
R705 GND.n186 GND.n185 4.65
R706 GND.n175 GND.n174 4.65
R707 GND.n168 GND.n167 4.65
R708 GND.n165 GND.n164 4.65
R709 GND.n157 GND.n156 4.65
R710 GND.n149 GND.n148 4.65
R711 GND.n107 GND.n106 4.504
R712 GND.n241 GND.n240 4.504
R713 GND.n178 GND.n177 4.504
R714 GND.n143 GND.n142 4.504
R715 GND.n12 GND.n11 4.129
R716 GND.n27 GND.n25 4.129
R717 GND.n57 GND.n56 4.129
R718 GND.n74 GND.n72 4.129
R719 GND.n97 GND.n95 4.129
R720 GND.n281 GND.n279 4.129
R721 GND.n260 GND.n258 4.129
R722 GND.n215 GND.n213 4.129
R723 GND.n197 GND.n195 4.129
R724 GND.n164 GND.n162 4.129
R725 GND.n114 GND.n113 3.716
R726 GND.n248 GND.n247 3.716
R727 GND.n185 GND.n184 3.716
R728 GND.n148 GND.n147 3.716
R729 GND.t11 GND.n107 2.452
R730 GND.t8 GND.n241 2.452
R731 GND.t9 GND.n178 2.452
R732 GND.t2 GND.n143 2.452
R733 GND.n151 GND.n150 1.935
R734 GND.n7 GND.n5 1.032
R735 GND.n34 GND.n33 1.032
R736 GND.n51 GND.n49 1.032
R737 GND.n81 GND.n80 1.032
R738 GND.n1 GND.n0 0.474
R739 GND.n139 GND.n138 0.474
R740 GND.n100 GND.n99 0.376
R741 GND.n251 GND.n250 0.376
R742 GND.n188 GND.n187 0.376
R743 GND.n153 GND.n152 0.376
R744 GND.n45 GND.n38 0.29
R745 GND.n92 GND.n85 0.29
R746 GND.n125 GND.n118 0.29
R747 GND.n271 GND.n264 0.29
R748 GND.n238 GND.n231 0.29
R749 GND.n208 GND.n201 0.29
R750 GND.n175 GND.n168 0.29
R751 GND.n140 GND 0.207
R752 GND.n103 GND.n101 0.206
R753 GND.n254 GND.n252 0.206
R754 GND.n191 GND.n189 0.206
R755 GND.n156 GND.n154 0.206
R756 GND.n23 GND.n16 0.181
R757 GND.n69 GND.n61 0.181
R758 GND.n137 GND.n134 0.181
R759 GND.n222 GND.n219 0.181
R760 GND.n104 GND.n98 0.157
R761 GND.n115 GND.n104 0.157
R762 GND.n261 GND.n255 0.157
R763 GND.n255 GND.n249 0.157
R764 GND.n198 GND.n192 0.157
R765 GND.n192 GND.n186 0.157
R766 GND.n165 GND.n157 0.157
R767 GND.n157 GND.n149 0.157
R768 GND.n13 GND.n8 0.145
R769 GND.n16 GND.n13 0.145
R770 GND.n28 GND.n23 0.145
R771 GND.n35 GND.n28 0.145
R772 GND.n38 GND.n35 0.145
R773 GND.n52 GND.n45 0.145
R774 GND.n58 GND.n52 0.145
R775 GND.n61 GND.n58 0.145
R776 GND.n75 GND.n69 0.145
R777 GND.n82 GND.n75 0.145
R778 GND.n85 GND.n82 0.145
R779 GND.n98 GND.n92 0.145
R780 GND.n118 GND.n115 0.145
R781 GND.n128 GND.n125 0.145
R782 GND.n131 GND.n128 0.145
R783 GND.n134 GND.n131 0.145
R784 GND.n282 GND.n274 0.145
R785 GND.n274 GND.n271 0.145
R786 GND.n264 GND.n261 0.145
R787 GND.n249 GND.n238 0.145
R788 GND.n231 GND.n228 0.145
R789 GND.n228 GND.n225 0.145
R790 GND.n225 GND.n222 0.145
R791 GND.n219 GND.n216 0.145
R792 GND.n216 GND.n211 0.145
R793 GND.n211 GND.n208 0.145
R794 GND.n201 GND.n198 0.145
R795 GND.n186 GND.n175 0.145
R796 GND.n168 GND.n165 0.145
R797 GND.n149 GND.n140 0.145
R798 GND GND.n137 0.133
R799 GND GND.n282 0.012
R800 Q.n0 Q.t6 486.819
R801 Q.n0 Q.t4 384.527
R802 Q.n1 Q.t5 322.919
R803 Q.n8 Q.n2 287.966
R804 Q.n7 Q.n6 223.975
R805 Q.n1 Q.n0 206.987
R806 Q.n7 Q.n3 157.274
R807 Q.n8 Q.n7 142.305
R808 Q.n6 Q.n5 22.578
R809 Q.n2 Q.t2 14.282
R810 Q.n2 Q.t1 14.282
R811 Q.n6 Q.n4 8.58
R812 Q.n9 Q.n1 5.965
R813 Q.n9 Q.n8 4.65
R814 Q.n9 Q 0.046
R815 D.n2 D.t5 512.525
R816 D.n0 D.t0 472.359
R817 D.n0 D.t3 384.527
R818 D.n2 D.t1 371.139
R819 D.n1 D.t2 342.755
R820 D.n3 D.t4 338.57
R821 D.n3 D.n2 191.629
R822 D.n1 D.n0 154.955
R823 D.n4 D.n1 11.134
R824 D.n4 D.n3 4.65
R825 D.n4 D 0.046
R826 a_185_209.n0 a_185_209.t5 480.392
R827 a_185_209.n0 a_185_209.t4 403.272
R828 a_185_209.n1 a_185_209.t3 357.204
R829 a_185_209.n3 a_185_209.n2 322.049
R830 a_185_209.n4 a_185_209.n3 243.422
R831 a_185_209.n1 a_185_209.n0 171.288
R832 a_185_209.n4 a_185_209.t1 14.282
R833 a_185_209.t2 a_185_209.n4 14.282
R834 a_185_209.n3 a_185_209.n1 10.615
R835 a_661_1050.n1 a_661_1050.t6 512.525
R836 a_661_1050.n1 a_661_1050.t5 371.139
R837 a_661_1050.n4 a_661_1050.n3 299.461
R838 a_661_1050.n2 a_661_1050.t7 282.852
R839 a_661_1050.n2 a_661_1050.n1 247.347
R840 a_661_1050.n5 a_661_1050.n4 187.858
R841 a_661_1050.n6 a_661_1050.n5 157.963
R842 a_661_1050.n5 a_661_1050.n0 91.706
R843 a_661_1050.n0 a_661_1050.t4 14.282
R844 a_661_1050.n0 a_661_1050.t2 14.282
R845 a_661_1050.n6 a_661_1050.t0 14.282
R846 a_661_1050.t1 a_661_1050.n6 14.282
R847 a_661_1050.n4 a_661_1050.n2 10.343
R848 a_1295_209.n0 a_1295_209.t3 486.819
R849 a_1295_209.n0 a_1295_209.t5 384.527
R850 a_1295_209.n1 a_1295_209.t4 350.778
R851 a_1295_209.n3 a_1295_209.n2 322.049
R852 a_1295_209.n4 a_1295_209.n3 243.422
R853 a_1295_209.n1 a_1295_209.n0 179.128
R854 a_1295_209.n3 a_1295_209.n1 14.696
R855 a_1295_209.n4 a_1295_209.t1 14.282
R856 a_1295_209.t2 a_1295_209.n4 14.282
R857 a_1666_101.n11 a_1666_101.n10 68.43
R858 a_1666_101.n3 a_1666_101.n2 62.817
R859 a_1666_101.n7 a_1666_101.n6 38.626
R860 a_1666_101.n6 a_1666_101.n5 35.955
R861 a_1666_101.n3 a_1666_101.n1 26.202
R862 a_1666_101.t0 a_1666_101.n3 19.737
R863 a_1666_101.t1 a_1666_101.n8 8.137
R864 a_1666_101.t0 a_1666_101.n4 7.273
R865 a_1666_101.t0 a_1666_101.n0 6.109
R866 a_1666_101.t1 a_1666_101.n7 4.864
R867 a_1666_101.t0 a_1666_101.n12 2.074
R868 a_1666_101.n12 a_1666_101.t1 0.937
R869 a_1666_101.t1 a_1666_101.n11 0.763
R870 a_1666_101.n11 a_1666_101.n9 0.185
R871 a_n259_209.n1 a_n259_209.t6 480.392
R872 a_n259_209.n3 a_n259_209.t8 472.359
R873 a_n259_209.n1 a_n259_209.t4 403.272
R874 a_n259_209.n3 a_n259_209.t3 384.527
R875 a_n259_209.n2 a_n259_209.t7 301.486
R876 a_n259_209.n6 a_n259_209.n0 299.141
R877 a_n259_209.n4 a_n259_209.t5 259.178
R878 a_n259_209.n8 a_n259_209.n6 251.114
R879 a_n259_209.n4 a_n259_209.n3 238.531
R880 a_n259_209.n2 a_n259_209.n1 227.006
R881 a_n259_209.n8 a_n259_209.n7 15.218
R882 a_n259_209.n0 a_n259_209.t1 14.282
R883 a_n259_209.n0 a_n259_209.t2 14.282
R884 a_n259_209.n9 a_n259_209.n8 12.014
R885 a_n259_209.n5 a_n259_209.n2 8.141
R886 a_n259_209.n6 a_n259_209.n5 8.141
R887 a_n259_209.n5 a_n259_209.n4 4.65
R888 a_556_101.n3 a_556_101.n1 42.788
R889 a_556_101.t0 a_556_101.n0 8.137
R890 a_556_101.n3 a_556_101.n2 4.665
R891 a_556_101.t0 a_556_101.n3 0.06
R892 a_2795_1051.n0 a_2795_1051.t2 228.369
R893 a_2795_1051.n0 a_2795_1051.t0 219.778
R894 a_2795_1051.n1 a_2795_1051.n0 42.29
R895 a_2795_1051.n1 a_2795_1051.t3 14.282
R896 a_2795_1051.t1 a_2795_1051.n1 14.282
R897 a_3461_1051.n1 a_3461_1051.t3 228.368
R898 a_3461_1051.t1 a_3461_1051.n1 219.777
R899 a_3461_1051.n1 a_3461_1051.n0 42.29
R900 a_3461_1051.n0 a_3461_1051.t2 14.282
R901 a_3461_1051.n0 a_3461_1051.t0 14.282
R902 GATE_N.n0 GATE_N.t0 512.525
R903 GATE_N.n0 GATE_N.t2 371.139
R904 GATE_N.n1 GATE_N.n0 275.206
R905 GATE_N.n1 GATE_N.t1 254.993
R906 GATE_N.n2 GATE_N.n1 4.65
R907 GATE_N.n2 GATE_N 0.046
C4 VDD GND 7.47fF
C5 a_3461_1051.n0 GND 0.21fF
C6 a_3461_1051.n1 GND 0.50fF
C7 a_2795_1051.n0 GND 0.52fF
C8 a_2795_1051.n1 GND 0.22fF
C9 a_556_101.n0 GND 0.05fF
C10 a_556_101.n1 GND 0.12fF
C11 a_556_101.n2 GND 0.04fF
C12 a_556_101.n3 GND 0.17fF
C13 a_n259_209.n0 GND 0.62fF
C14 a_n259_209.n1 GND 0.35fF
C15 a_n259_209.n2 GND 0.55fF
C16 a_n259_209.n3 GND 0.33fF
C17 a_n259_209.t5 GND 0.45fF
C18 a_n259_209.n4 GND 0.36fF
C19 a_n259_209.n5 GND 1.17fF
C20 a_n259_209.n6 GND 0.74fF
C21 a_n259_209.n7 GND 0.08fF
C22 a_n259_209.n8 GND 0.14fF
C23 a_n259_209.n9 GND 0.04fF
C24 a_1666_101.n0 GND 0.02fF
C25 a_1666_101.n1 GND 0.09fF
C26 a_1666_101.n2 GND 0.08fF
C27 a_1666_101.n3 GND 0.03fF
C28 a_1666_101.n4 GND 0.01fF
C29 a_1666_101.n5 GND 0.04fF
C30 a_1666_101.n6 GND 0.04fF
C31 a_1666_101.n7 GND 0.02fF
C32 a_1666_101.n8 GND 0.05fF
C33 a_1666_101.n9 GND 0.15fF
C34 a_1666_101.n10 GND 0.08fF
C35 a_1666_101.n11 GND 0.08fF
C36 a_1666_101.t1 GND 0.23fF
C37 a_1666_101.n12 GND 0.01fF
C38 a_1295_209.n0 GND 0.39fF
C39 a_1295_209.n1 GND 1.25fF
C40 a_1295_209.n2 GND 0.39fF
C41 a_1295_209.n3 GND 1.51fF
C42 a_1295_209.n4 GND 0.72fF
C43 a_661_1050.n0 GND 0.34fF
C44 a_661_1050.n1 GND 0.31fF
C45 a_661_1050.t7 GND 0.45fF
C46 a_661_1050.n2 GND 0.52fF
C47 a_661_1050.n3 GND 0.27fF
C48 a_661_1050.n4 GND 0.58fF
C49 a_661_1050.n5 GND 0.54fF
C50 a_661_1050.n6 GND 0.44fF
C51 a_185_209.n0 GND 0.33fF
C52 a_185_209.n1 GND 0.60fF
C53 a_185_209.n2 GND 0.32fF
C54 a_185_209.n3 GND 0.81fF
C55 a_185_209.n4 GND 0.60fF
C56 Q.n0 GND 0.34fF
C57 Q.t5 GND 0.50fF
C58 Q.n1 GND 0.45fF
C59 Q.n2 GND 0.57fF
C60 Q.n3 GND 0.17fF
C61 Q.n4 GND 0.04fF
C62 Q.n5 GND 0.05fF
C63 Q.n6 GND 0.14fF
C64 Q.n7 GND 0.47fF
C65 Q.n8 GND 0.48fF
C66 Q.n9 GND 0.30fF
C67 a_3007_411.n0 GND 0.05fF
C68 a_3007_411.n1 GND 0.60fF
C69 a_3007_411.n2 GND 0.34fF
C70 a_3007_411.n3 GND 0.83fF
C71 a_3007_411.n4 GND 0.93fF
C72 a_3007_411.n5 GND 0.04fF
C73 a_3007_411.n6 GND 0.06fF
C74 a_3007_411.n7 GND 0.04fF
C75 a_3007_411.n8 GND 0.13fF
C76 a_3007_411.n9 GND 0.54fF
C77 a_3007_411.n10 GND 0.04fF
C78 a_3007_411.n11 GND 0.06fF
C79 a_3007_411.n12 GND 0.05fF
C80 VDD.n1 GND 0.03fF
C81 VDD.n2 GND 0.11fF
C82 VDD.n3 GND 0.02fF
C83 VDD.n4 GND 0.02fF
C84 VDD.n5 GND 0.05fF
C85 VDD.n6 GND 0.02fF
C86 VDD.n7 GND 0.02fF
C87 VDD.n8 GND 0.02fF
C88 VDD.n9 GND 0.02fF
C89 VDD.n10 GND 0.02fF
C90 VDD.n11 GND 0.02fF
C91 VDD.n12 GND 0.02fF
C92 VDD.n13 GND 0.02fF
C93 VDD.n14 GND 0.03fF
C94 VDD.n15 GND 0.01fF
C95 VDD.n20 GND 0.38fF
C96 VDD.n21 GND 0.23fF
C97 VDD.n22 GND 0.02fF
C98 VDD.n23 GND 0.03fF
C99 VDD.n24 GND 0.20fF
C100 VDD.n25 GND 0.01fF
C101 VDD.n26 GND 0.02fF
C102 VDD.n27 GND 0.01fF
C103 VDD.n28 GND 0.14fF
C104 VDD.n29 GND 0.01fF
C105 VDD.n30 GND 0.02fF
C106 VDD.n31 GND 0.07fF
C107 VDD.n32 GND 0.01fF
C108 VDD.n33 GND 0.02fF
C109 VDD.n34 GND 0.02fF
C110 VDD.n35 GND 0.12fF
C111 VDD.n36 GND 0.01fF
C112 VDD.n37 GND 0.02fF
C113 VDD.n38 GND 0.02fF
C114 VDD.n39 GND 0.07fF
C115 VDD.n40 GND 0.04fF
C116 VDD.n41 GND 0.13fF
C117 VDD.n42 GND 0.01fF
C118 VDD.n43 GND 0.01fF
C119 VDD.n44 GND 0.02fF
C120 VDD.n45 GND 0.20fF
C121 VDD.n46 GND 0.01fF
C122 VDD.n47 GND 0.02fF
C123 VDD.n48 GND 0.02fF
C124 VDD.n49 GND 0.23fF
C125 VDD.n50 GND 0.01fF
C126 VDD.n51 GND 0.02fF
C127 VDD.n52 GND 0.03fF
C128 VDD.n53 GND 0.05fF
C129 VDD.n54 GND 0.02fF
C130 VDD.n55 GND 0.02fF
C131 VDD.n56 GND 0.02fF
C132 VDD.n57 GND 0.02fF
C133 VDD.n58 GND 0.02fF
C134 VDD.n59 GND 0.02fF
C135 VDD.n60 GND 0.02fF
C136 VDD.n61 GND 0.02fF
C137 VDD.n62 GND 0.02fF
C138 VDD.n63 GND 0.02fF
C139 VDD.n64 GND 0.01fF
C140 VDD.n65 GND 0.02fF
C141 VDD.n66 GND 0.02fF
C142 VDD.n67 GND 0.18fF
C143 VDD.n68 GND 0.02fF
C144 VDD.n69 GND 0.02fF
C145 VDD.n71 GND 0.02fF
C146 VDD.n75 GND 0.23fF
C147 VDD.n76 GND 0.23fF
C148 VDD.n77 GND 0.01fF
C149 VDD.n78 GND 0.02fF
C150 VDD.n79 GND 0.03fF
C151 VDD.n80 GND 0.20fF
C152 VDD.n81 GND 0.01fF
C153 VDD.n82 GND 0.02fF
C154 VDD.n83 GND 0.02fF
C155 VDD.n84 GND 0.14fF
C156 VDD.n85 GND 0.01fF
C157 VDD.n86 GND 0.02fF
C158 VDD.n87 GND 0.02fF
C159 VDD.n88 GND 0.01fF
C160 VDD.n89 GND 0.02fF
C161 VDD.n90 GND 0.02fF
C162 VDD.n91 GND 0.12fF
C163 VDD.n92 GND 0.01fF
C164 VDD.n93 GND 0.02fF
C165 VDD.n94 GND 0.02fF
C166 VDD.n95 GND 0.07fF
C167 VDD.n96 GND 0.04fF
C168 VDD.n97 GND 0.13fF
C169 VDD.n98 GND 0.01fF
C170 VDD.n99 GND 0.01fF
C171 VDD.n100 GND 0.02fF
C172 VDD.n101 GND 0.20fF
C173 VDD.n102 GND 0.01fF
C174 VDD.n103 GND 0.02fF
C175 VDD.n104 GND 0.02fF
C176 VDD.n105 GND 0.23fF
C177 VDD.n106 GND 0.01fF
C178 VDD.n107 GND 0.02fF
C179 VDD.n108 GND 0.03fF
C180 VDD.n109 GND 0.15fF
C181 VDD.n110 GND 0.02fF
C182 VDD.n111 GND 0.02fF
C183 VDD.n112 GND 0.02fF
C184 VDD.n113 GND 0.05fF
C185 VDD.n114 GND 0.02fF
C186 VDD.n115 GND 0.02fF
C187 VDD.n116 GND 0.02fF
C188 VDD.n117 GND 0.02fF
C189 VDD.n118 GND 0.02fF
C190 VDD.n119 GND 0.02fF
C191 VDD.n120 GND 0.02fF
C192 VDD.n121 GND 0.02fF
C193 VDD.n122 GND 0.02fF
C194 VDD.n123 GND 0.01fF
C195 VDD.n124 GND 0.02fF
C196 VDD.n125 GND 0.02fF
C197 VDD.n126 GND 0.02fF
C198 VDD.n130 GND 0.23fF
C199 VDD.n131 GND 0.23fF
C200 VDD.n132 GND 0.01fF
C201 VDD.n133 GND 0.02fF
C202 VDD.n134 GND 0.03fF
C203 VDD.n135 GND 0.05fF
C204 VDD.n136 GND 0.17fF
C205 VDD.n137 GND 0.01fF
C206 VDD.n138 GND 0.01fF
C207 VDD.n139 GND 0.02fF
C208 VDD.n140 GND 0.14fF
C209 VDD.n141 GND 0.01fF
C210 VDD.n142 GND 0.02fF
C211 VDD.n143 GND 0.02fF
C212 VDD.n144 GND 0.05fF
C213 VDD.n145 GND 0.17fF
C214 VDD.n146 GND 0.01fF
C215 VDD.n147 GND 0.01fF
C216 VDD.n148 GND 0.02fF
C217 VDD.n149 GND 0.23fF
C218 VDD.n150 GND 0.01fF
C219 VDD.n151 GND 0.02fF
C220 VDD.n152 GND 0.03fF
C221 VDD.n153 GND 0.15fF
C222 VDD.n154 GND 0.02fF
C223 VDD.n155 GND 0.02fF
C224 VDD.n156 GND 0.02fF
C225 VDD.n157 GND 0.05fF
C226 VDD.n158 GND 0.02fF
C227 VDD.n159 GND 0.02fF
C228 VDD.n160 GND 0.02fF
C229 VDD.n161 GND 0.02fF
C230 VDD.n162 GND 0.02fF
C231 VDD.n163 GND 0.02fF
C232 VDD.n164 GND 0.02fF
C233 VDD.n165 GND 0.02fF
C234 VDD.n166 GND 0.02fF
C235 VDD.n167 GND 0.01fF
C236 VDD.n168 GND 0.02fF
C237 VDD.n169 GND 0.02fF
C238 VDD.n170 GND 0.02fF
C239 VDD.n174 GND 0.23fF
C240 VDD.n175 GND 0.23fF
C241 VDD.n176 GND 0.01fF
C242 VDD.n177 GND 0.02fF
C243 VDD.n178 GND 0.03fF
C244 VDD.n179 GND 0.20fF
C245 VDD.n180 GND 0.01fF
C246 VDD.n181 GND 0.05fF
C247 VDD.n182 GND 0.01fF
C248 VDD.n183 GND 0.02fF
C249 VDD.n184 GND 0.14fF
C250 VDD.n185 GND 0.01fF
C251 VDD.n186 GND 0.02fF
C252 VDD.n187 GND 0.02fF
C253 VDD.n188 GND 0.01fF
C254 VDD.n189 GND 0.07fF
C255 VDD.n190 GND 0.04fF
C256 VDD.n191 GND 0.02fF
C257 VDD.n192 GND 0.02fF
C258 VDD.n193 GND 0.12fF
C259 VDD.n194 GND 0.01fF
C260 VDD.n195 GND 0.02fF
C261 VDD.n196 GND 0.02fF
C262 VDD.n197 GND 0.08fF
C263 VDD.n198 GND 0.02fF
C264 VDD.n199 GND 0.02fF
C265 VDD.n200 GND 0.05fF
C266 VDD.n201 GND 0.02fF
C267 VDD.n202 GND 0.02fF
C268 VDD.n203 GND 0.02fF
C269 VDD.n204 GND 0.02fF
C270 VDD.n205 GND 0.02fF
C271 VDD.n206 GND 0.02fF
C272 VDD.n207 GND 0.02fF
C273 VDD.n208 GND 0.02fF
C274 VDD.n209 GND 0.03fF
C275 VDD.n210 GND 0.03fF
C276 VDD.n211 GND 0.02fF
C277 VDD.n215 GND 0.38fF
C278 VDD.n216 GND 0.23fF
C279 VDD.n217 GND 0.02fF
C280 VDD.n218 GND 0.03fF
C281 VDD.n219 GND 0.02fF
C282 VDD.n220 GND 0.17fF
C283 VDD.n221 GND 0.01fF
C284 VDD.n222 GND 0.05fF
C285 VDD.n223 GND 0.01fF
C286 VDD.n224 GND 0.02fF
C287 VDD.n225 GND 0.14fF
C288 VDD.n226 GND 0.01fF
C289 VDD.n227 GND 0.02fF
C290 VDD.n228 GND 0.02fF
C291 VDD.n229 GND 0.05fF
C292 VDD.n230 GND 0.17fF
C293 VDD.n231 GND 0.01fF
C294 VDD.n232 GND 0.01fF
C295 VDD.n233 GND 0.02fF
C296 VDD.n234 GND 0.23fF
C297 VDD.n235 GND 0.01fF
C298 VDD.n236 GND 0.02fF
C299 VDD.n237 GND 0.03fF
C300 VDD.n238 GND 0.02fF
C301 VDD.n241 GND 0.02fF
C302 VDD.n243 GND 0.02fF
C303 VDD.n244 GND 0.12fF
C304 VDD.n245 GND 0.02fF
C305 VDD.n247 GND 0.23fF
C306 VDD.n248 GND 0.23fF
C307 VDD.n249 GND 0.01fF
C308 VDD.n250 GND 0.05fF
C309 VDD.n251 GND 0.02fF
C310 VDD.n252 GND 0.02fF
C311 VDD.n253 GND 0.02fF
C312 VDD.n254 GND 0.02fF
C313 VDD.n255 GND 0.02fF
C314 VDD.n256 GND 0.02fF
C315 VDD.n257 GND 0.02fF
C316 VDD.n258 GND 0.02fF
C317 VDD.n259 GND 0.02fF
C318 VDD.n260 GND 0.02fF
C319 VDD.n261 GND 0.01fF
C320 VDD.n262 GND 0.02fF
C321 VDD.n263 GND 0.02fF
C322 VDD.n264 GND 0.03fF
C323 VDD.n265 GND 0.05fF
C324 VDD.n266 GND 0.17fF
C325 VDD.n267 GND 0.01fF
C326 VDD.n268 GND 0.01fF
C327 VDD.n269 GND 0.02fF
C328 VDD.n270 GND 0.14fF
C329 VDD.n271 GND 0.01fF
C330 VDD.n272 GND 0.02fF
C331 VDD.n273 GND 0.02fF
C332 VDD.n274 GND 0.05fF
C333 VDD.n275 GND 0.17fF
C334 VDD.n276 GND 0.01fF
C335 VDD.n277 GND 0.01fF
C336 VDD.n278 GND 0.02fF
C337 VDD.n279 GND 0.23fF
C338 VDD.n280 GND 0.01fF
C339 VDD.n281 GND 0.02fF
C340 VDD.n282 GND 0.03fF
C341 VDD.n283 GND 0.15fF
C342 VDD.n284 GND 0.02fF
C343 VDD.n285 GND 0.02fF
C344 VDD.n286 GND 0.02fF
C345 VDD.n287 GND 0.05fF
C346 VDD.n288 GND 0.02fF
C347 VDD.n289 GND 0.02fF
C348 VDD.n290 GND 0.02fF
C349 VDD.n291 GND 0.02fF
C350 VDD.n292 GND 0.02fF
C351 VDD.n293 GND 0.02fF
C352 VDD.n294 GND 0.02fF
C353 VDD.n295 GND 0.02fF
C354 VDD.n296 GND 0.02fF
C355 VDD.n297 GND 0.01fF
C356 VDD.n298 GND 0.02fF
C357 VDD.n299 GND 0.02fF
C358 VDD.n300 GND 0.02fF
C359 VDD.n304 GND 0.23fF
C360 VDD.n305 GND 0.23fF
C361 VDD.n306 GND 0.01fF
C362 VDD.n307 GND 0.02fF
C363 VDD.n308 GND 0.03fF
C364 VDD.n309 GND 0.05fF
C365 VDD.n310 GND 0.20fF
C366 VDD.n311 GND 0.01fF
C367 VDD.n312 GND 0.01fF
C368 VDD.n313 GND 0.02fF
C369 VDD.n314 GND 0.13fF
C370 VDD.n315 GND 0.01fF
C371 VDD.n316 GND 0.02fF
C372 VDD.n317 GND 0.02fF
C373 VDD.n318 GND 0.12fF
C374 VDD.n319 GND 0.01fF
C375 VDD.n320 GND 0.02fF
C376 VDD.n321 GND 0.02fF
C377 VDD.n322 GND 0.07fF
C378 VDD.n323 GND 0.04fF
C379 VDD.n324 GND 0.01fF
C380 VDD.n325 GND 0.02fF
C381 VDD.n326 GND 0.02fF
C382 VDD.n327 GND 0.14fF
C383 VDD.n328 GND 0.01fF
C384 VDD.n329 GND 0.02fF
C385 VDD.n330 GND 0.02fF
C386 VDD.n331 GND 0.05fF
C387 VDD.n332 GND 0.20fF
C388 VDD.n333 GND 0.01fF
C389 VDD.n334 GND 0.01fF
C390 VDD.n335 GND 0.02fF
C391 VDD.n336 GND 0.23fF
C392 VDD.n337 GND 0.01fF
C393 VDD.n338 GND 0.02fF
C394 VDD.n339 GND 0.03fF
C395 VDD.n340 GND 0.15fF
C396 VDD.n341 GND 0.02fF
C397 VDD.n342 GND 0.02fF
C398 VDD.n343 GND 0.02fF
C399 VDD.n344 GND 0.05fF
C400 VDD.n345 GND 0.02fF
C401 VDD.n346 GND 0.02fF
C402 VDD.n347 GND 0.02fF
C403 VDD.n348 GND 0.02fF
C404 VDD.n349 GND 0.02fF
C405 VDD.n350 GND 0.02fF
C406 VDD.n351 GND 0.02fF
C407 VDD.n352 GND 0.02fF
C408 VDD.n353 GND 0.02fF
C409 VDD.n354 GND 0.01fF
C410 VDD.n355 GND 0.02fF
C411 VDD.n356 GND 0.02fF
C412 VDD.n357 GND 0.02fF
C413 VDD.n361 GND 0.23fF
C414 VDD.n362 GND 0.23fF
C415 VDD.n363 GND 0.01fF
C416 VDD.n364 GND 0.02fF
C417 VDD.n365 GND 0.03fF
C418 VDD.n366 GND 0.17fF
C419 VDD.n367 GND 0.01fF
C420 VDD.n368 GND 0.05fF
C421 VDD.n369 GND 0.01fF
C422 VDD.n370 GND 0.02fF
C423 VDD.n371 GND 0.14fF
C424 VDD.n372 GND 0.01fF
C425 VDD.n373 GND 0.02fF
C426 VDD.n374 GND 0.02fF
C427 VDD.n375 GND 0.05fF
C428 VDD.n376 GND 0.17fF
C429 VDD.n377 GND 0.01fF
C430 VDD.n378 GND 0.01fF
C431 VDD.n379 GND 0.02fF
C432 VDD.n380 GND 0.23fF
C433 VD