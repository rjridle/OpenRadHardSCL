magic
tech sky130
magscale 1 2
timestamp 1645050557
<< locali >>
rect -17 17 17 33
rect -17 -33 17 -17
<< viali >>
rect -17 -17 17 17
<< metal1 >>
rect -17 23 17 53
rect -23 17 23 23
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -23 23 -17
rect -17 -29 17 -23
<< end >>
