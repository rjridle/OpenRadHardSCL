* SPICE3 file created from NAND2X1.ext - technology: sky130A

.subckt NAND2X1 Y A B VDD VSS
X0 VDD A Y VDD sky130_fd_pr__pfet_01v8 ad=1.68p pd=1.368u as=1.16p ps=9.16u w=2u l=0.15u M=2
X1 VDD B Y VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X2 VSS A a_112_101# VSS sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=0p ps=0u w=3u l=0.15u
X3 Y B a_112_101# VSS sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=0p ps=0u w=3u l=0.15u
.ends
