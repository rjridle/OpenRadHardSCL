magic
tech sky130A
magscale 1 2
timestamp 1642971013
<< error_p >>
rect 85 322 86 323
rect 269 322 270 323
rect 86 321 87 322
rect 270 321 271 322
rect 101 291 102 292
rect 136 291 137 292
rect 285 291 286 292
rect 320 291 321 292
rect 101 188 102 189
rect 136 188 137 189
rect 285 188 286 189
rect 320 188 321 189
<< nmos >>
rect 56 322 86 375
rect 240 322 270 375
rect 56 292 152 322
tri 152 292 182 322 sw
rect 56 188 86 292
tri 86 276 102 292 nw
tri 136 276 152 292 ne
tri 86 188 102 204 sw
tri 136 188 152 204 se
rect 152 188 182 292
rect 240 292 336 322
tri 336 292 366 322 sw
tri 56 158 86 188 ne
rect 86 158 152 188
tri 152 158 182 188 nw
rect 240 188 270 292
tri 270 276 286 292 nw
tri 320 276 336 292 ne
tri 270 188 286 204 sw
tri 320 188 336 204 se
rect 336 188 366 292
tri 240 158 270 188 ne
rect 270 158 336 188
tri 336 158 366 188 nw
<< ndiff >>
rect 0 298 56 375
rect 86 322 240 375
rect 270 322 420 375
rect 0 264 10 298
rect 44 264 56 298
tri 152 292 182 322 ne
rect 182 298 240 322
rect 0 215 56 264
rect 0 181 10 215
rect 44 181 56 215
tri 86 276 102 292 se
rect 102 276 136 292
tri 136 276 152 292 sw
rect 86 242 152 276
rect 86 208 98 242
rect 132 208 152 242
rect 86 204 152 208
tri 86 188 102 204 ne
rect 102 188 136 204
tri 136 188 152 204 nw
rect 182 264 194 298
rect 228 264 240 298
tri 336 292 366 322 ne
rect 366 298 420 322
rect 182 215 240 264
rect 0 158 56 181
tri 56 158 86 188 sw
tri 152 158 182 188 se
rect 182 181 194 215
rect 228 181 240 215
tri 270 276 286 292 se
rect 286 276 320 292
tri 320 276 336 292 sw
rect 270 242 336 276
rect 270 208 282 242
rect 316 208 336 242
rect 270 204 336 208
tri 270 188 286 204 ne
rect 286 188 320 204
tri 320 188 336 204 nw
rect 366 264 378 298
rect 412 264 420 298
rect 366 215 420 264
rect 182 158 240 181
tri 240 158 270 188 sw
tri 336 158 366 188 se
rect 366 181 378 215
rect 412 181 420 215
rect 366 158 420 181
rect 0 147 420 158
rect 0 113 10 147
rect 44 113 98 147
rect 132 113 194 147
rect 228 113 282 147
rect 316 113 378 147
rect 412 113 420 147
rect 0 101 420 113
<< ndiffc >>
rect 10 264 44 298
rect 10 181 44 215
rect 98 208 132 242
rect 194 264 228 298
rect 194 181 228 215
rect 282 208 316 242
rect 378 264 412 298
rect 378 181 412 215
rect 10 113 44 147
rect 98 113 132 147
rect 194 113 228 147
rect 282 113 316 147
rect 378 113 412 147
<< psubdiff >>
rect -116 429 536 491
rect -116 47 -54 429
rect 474 47 536 429
rect -116 13 24 47
rect 58 13 92 47
rect 126 13 160 47
rect 194 13 228 47
rect 262 13 296 47
rect 330 13 364 47
rect 398 13 536 47
rect -116 0 536 13
<< psubdiffcont >>
rect 24 13 58 47
rect 92 13 126 47
rect 160 13 194 47
rect 228 13 262 47
rect 296 13 330 47
rect 364 13 398 47
<< poly >>
rect 56 375 86 404
rect 240 375 270 404
<< locali >>
rect -116 62 -54 491
rect 10 298 44 343
rect 194 298 228 343
rect 10 215 44 264
rect 98 278 132 287
rect 98 242 132 244
rect 98 192 132 208
rect 378 298 412 343
rect 194 215 228 264
rect 10 147 44 181
rect 282 278 316 288
rect 282 242 316 244
rect 282 192 316 208
rect 378 215 412 264
rect 194 147 228 181
rect 378 147 412 181
rect 44 113 98 147
rect 132 113 194 147
rect 228 113 282 147
rect 316 113 378 147
rect 10 62 44 113
rect 194 62 228 113
rect 378 62 412 113
rect 474 62 536 491
rect -116 47 536 62
rect -116 13 24 47
rect 58 13 92 47
rect 126 13 160 47
rect 194 13 228 47
rect 262 13 296 47
rect 330 13 364 47
rect 398 13 536 47
rect -116 0 536 13
<< viali >>
rect 98 244 132 278
rect 282 244 316 278
rect 24 13 58 47
rect 92 13 126 47
rect 160 13 194 47
rect 228 13 262 47
rect 296 13 330 47
rect 364 13 398 47
<< metal1 >>
rect -116 62 -54 491
rect 98 285 132 290
rect 282 285 316 290
rect 92 278 138 285
rect 276 278 322 285
rect 92 244 98 278
rect 132 244 282 278
rect 316 244 322 278
rect 92 237 138 244
rect 276 237 322 244
rect 98 232 132 237
rect 282 232 316 237
rect 474 62 536 491
rect -116 47 536 62
rect -116 13 24 47
rect 58 13 92 47
rect 126 13 160 47
rect 194 13 228 47
rect 262 13 296 47
rect 330 13 364 47
rect 398 13 536 47
rect -116 0 536 13
<< labels >>
rlabel metal1 98 244 132 278 1 A
rlabel metal1 278 26 278 26 1 VSS
<< end >>
