magic
tech sky130A
magscale 1 2
timestamp 1651071336
<< metal1 >>
rect -31 1492 2029 1554
rect 1685 797 1719 831
rect 1019 723 1053 757
rect 353 649 387 683
rect 205 575 239 609
rect 1833 575 1867 609
rect -31 0 2029 62
use aoai4x1_pcell  aoai4x1_pcell_0 pcells
timestamp 1648661172
transform 1 0 0 0 1 0
box -84 0 2082 1575
use li1_M1_contact  li1_M1_contact_1 pcells
timestamp 1648061256
transform 1 0 222 0 1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform 1 0 370 0 1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_2
timestamp 1648061256
transform 1 0 1036 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_3
timestamp 1648061256
transform 1 0 1702 0 1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_4
timestamp 1648061256
transform -1 0 1850 0 -1 592
box -53 -33 29 33
<< labels >>
rlabel metal1 1833 575 1867 609 1 YN
port 1 n
rlabel metal1 205 575 239 609 1 A
port 2 n
rlabel metal1 353 649 387 683 1 B
port 3 n
rlabel metal1 1019 723 1053 757 1 C
port 4 n
rlabel metal1 1685 797 1719 831 1 D
port 5 n
rlabel metal1 -31 1492 2029 1554 1 VDD
port 6 n
rlabel metal1 -31 0 2029 62 1 GND
port 7 n
<< end >>
