* SPICE3 file created from INVX1.ext - technology: sky130A

.subckt INVX1 Y A VDD VSS
X0 Y A VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=1.1e+12p ps=9.1e+06u w=2e+06u l=150000u M=2
X1 Y A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.791e+11p pd=1.57e+06u as=1.1408e+12p ps=8.1e+06u w=3e+06u l=150000u
.ends
