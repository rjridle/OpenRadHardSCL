* SPICE3 file created from NAND2X1.ext - technology: sky130A

.subckt NAND2X1 Y A B VDD VSS
X0 VDD A Y VDD sky130_fd_pr__pfet_01v8 ad=1.68e+12p pd=1.368e+07u as=1.16e+12p ps=9.16e+06u w=2e+06u l=150000u M=2
X1 VDD B Y VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X2 VSS A a_112_101 VSS sky130_fd_pr__nfet_01v8 ad=1.791e+11p pd=1.57e+06u as=0p ps=0u w=3e+06u l=150000u
X3 Y B a_112_101 VSS sky130_fd_pr__nfet_01v8 ad=1.791e+11p pd=1.57e+06u as=0p ps=0u w=3e+06u l=150000u
.ends
