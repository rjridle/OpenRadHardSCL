* SPICE3 file created from NAND3X1.ext - technology: sky130A

.subckt NAND3X1 Y A B VDD VSS
X0 VDD B Y VDD sky130_fd_pr__pfet_01v8 ad=2.26e+12p pd=1.826e+07u as=1.74e+12p ps=1.374e+07u w=2e+06u l=150000u M=2
X1 VDD a_599_989 Y VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X2 Y a_599_989 a_372_210 VSS sky130_fd_pr__nfet_01v8 ad=1.791e+11p pd=1.57e+06u as=0p ps=0u w=3e+06u l=150000u
X3 Y A VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X4 VSS A a_91_103 VSS sky130_fd_pr__nfet_01v8 ad=1.791e+11p pd=1.57e+06u as=0p ps=0u w=3e+06u l=150000u
X5 a_372_210 B a_91_103 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
C0 VDD Y 2.50fF
.ends
