magic
tech sky130A
magscale 1 2
timestamp 1645132717
<< nwell >>
rect 49 1352 949 1353
rect 49 1344 1106 1352
rect 47 1332 1106 1344
rect -31 1278 1106 1332
rect 31 1270 1106 1278
rect 47 1265 1106 1270
rect 47 1261 637 1265
rect 47 1245 549 1261
rect 319 1055 549 1245
rect 643 1055 1106 1265
rect -65 759 1106 1055
<< psubdiff >>
rect 12 499 915 561
rect 31 13 109 47
rect 143 13 177 47
rect 211 13 245 47
rect 279 13 313 47
rect 347 13 381 47
rect 415 13 449 47
rect 483 13 915 47
<< nsubdiff >>
rect 16 1283 109 1317
rect 143 1283 177 1317
rect 211 1283 245 1317
rect 280 1283 314 1317
rect 348 1283 382 1317
rect 416 1283 450 1317
rect 484 1283 991 1317
rect 12 795 915 857
<< psubdiffcont >>
rect 109 13 143 47
rect 177 13 211 47
rect 245 13 279 47
rect 313 13 347 47
rect 381 13 415 47
rect 449 13 483 47
<< nsubdiffcont >>
rect 109 1283 143 1317
rect 177 1283 211 1317
rect 245 1283 280 1317
rect 314 1283 348 1317
rect 382 1283 416 1317
rect 450 1283 484 1317
<< poly >>
rect 445 916 503 946
rect 181 429 532 459
rect 318 415 348 429
rect 502 415 532 429
<< locali >>
rect -31 1319 991 1332
rect -31 1317 995 1319
rect -31 1283 109 1317
rect 143 1283 177 1317
rect 211 1283 245 1317
rect 280 1283 314 1317
rect 348 1283 382 1317
rect 416 1283 450 1317
rect 484 1283 995 1317
rect -31 1281 995 1283
rect -31 1278 991 1281
rect 31 1270 991 1278
rect 455 1269 489 1270
rect 364 427 582 461
rect 364 272 398 427
rect 548 255 582 427
rect 279 101 306 102
rect 463 101 490 102
rect 272 62 306 101
rect 456 62 490 101
rect 640 62 674 101
rect 31 47 915 62
rect 31 13 109 47
rect 143 13 177 47
rect 211 13 245 47
rect 279 13 313 47
rect 347 13 381 47
rect 415 13 449 47
rect 483 13 915 47
rect 31 0 915 13
<< viali >>
rect 109 1283 143 1317
rect 177 1283 211 1317
rect 245 1283 280 1317
rect 314 1283 348 1317
rect 382 1283 416 1317
rect 450 1283 484 1317
rect 109 13 143 47
rect 177 13 211 47
rect 245 13 279 47
rect 313 13 347 47
rect 381 13 415 47
rect 449 13 483 47
<< metal1 >>
rect -31 1319 991 1332
rect -31 1317 995 1319
rect -31 1283 109 1317
rect 143 1283 177 1317
rect 211 1283 245 1317
rect 280 1283 314 1317
rect 348 1283 382 1317
rect 416 1283 450 1317
rect 484 1283 995 1317
rect -31 1281 995 1283
rect -31 1278 991 1281
rect 31 1270 991 1278
rect 131 497 165 876
rect 31 47 915 62
rect 31 13 109 47
rect 143 13 177 47
rect 211 13 245 47
rect 279 13 313 47
rect 347 13 381 47
rect 415 13 449 47
rect 483 13 915 47
rect 31 0 915 13
use poly_li1_contact_perp  poly_li1_contact_perp_1 pcells
timestamp 1645049645
transform 1 0 71 0 1 460
box 44 399 110 481
use nmos_top  nmos_top_1 pcells
timestamp 1643656459
transform -1 0 684 0 1 101
box 0 0 238 314
use nmos_top  nmos_top_0
timestamp 1643656459
transform -1 0 500 0 1 101
box 0 0 238 314
use diff_ring_side  diff_ring_side_1 pcells
timestamp 1643181737
transform 1 0 1021 0 1 0
box -159 0 9 1353
use pmos4  pmos4_1 pcells
timestamp 1645051079
transform 1 0 447 0 1 1228
box -36 -312 440 42
use poly_li1_contact_perp  poly_li1_contact_perp_0
timestamp 1645049645
transform -1 0 225 0 -1 896
box 44 399 110 481
use pmos4  pmos4_0
timestamp 1645051079
transform 1 0 95 0 1 1228
box -36 -312 440 42
use diff_ring_side  diff_ring_side_0
timestamp 1643181737
transform 1 0 75 0 1 0
box -159 0 9 1353
<< labels >>
rlabel metal1 363 26 363 26 1 VSS
port 1 n
rlabel metal1 366 1301 366 1301 1 VDD
port 2 n
<< end >>
