magic
tech sky130
magscale 1 2
timestamp 1651259535
<< metal1 >>
rect 1201 501 1443 535
use aoi3x1_pcell  aoi3x1_pcell_0
timestamp 1651259532
transform 1 0 0 0 1 0
box -84 0 1416 1575
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform -1 0 1184 0 -1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform 1 0 1480 0 1 518
box -53 -33 29 33
use invx1_pcell  invx1_pcell_0
timestamp 1651259471
transform 1 0 1332 0 1 0
box -84 0 528 1575
<< end >>
