* SPICE3 file created from AOI3X1.ext - technology: sky130A

.subckt AOI3X1 YN A B C VDD VSS
X0 VDD A a_217_1050# VDD sky130_fd_pr__pfet_01v8 ad=2.26p pd=1.826u as=0p ps=0u w=2u l=0.15u M=2
X1 VDD a_217_1050# a_797_1051# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X2 VDD B a_217_1050# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X3 a_797_1051# C YN VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8p ps=4.58u w=2u l=0.15u M=2
X4 VSS A a_112_101# VSS sky130_fd_pr__nfet_01v8 ad=2.1157p pd=1.451u as=0p ps=0u w=3u l=0.15u
X5 YN a_217_1050# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.582p pd=3.15u as=0p ps=0u w=3u l=0.15u
X6 a_217_1050# B a_112_101# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X7 YN C VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
C0 a_217_1050# VDD 2.17fF
.ends
