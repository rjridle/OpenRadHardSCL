magic
tech sky130A
magscale 1 2
timestamp 1648157493
<< metal1 >>
rect 55 1505 89 1539
rect 427 797 461 831
rect 205 723 239 757
rect 797 649 831 683
rect 55 13 89 47
use li1_M1_contact  li1_M1_contact_1 pcells
timestamp 1648061256
transform 1 0 222 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_4
timestamp 1648061256
transform -1 0 814 0 -1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform 1 0 444 0 1 814
box -53 -33 29 33
use nand3x1_pcell  nand3x1_pcell_0 pcells
timestamp 1648064657
transform 1 0 0 0 1 0
box -84 0 1046 1575
<< labels >>
rlabel metal1 797 649 831 683 1 Y
port 1 n
rlabel metal1 205 723 239 757 1 A
port 2 n
rlabel metal1 427 797 461 831 1 B
port 3 n
rlabel metal1 55 1505 89 1539 1 VDD
port 4 n
rlabel metal1 55 13 89 47 1 VSS
port 5 n
<< end >>
