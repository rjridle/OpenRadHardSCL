* SPICE3 file created from TMRDFFSNQX1.ext - technology: sky130A

.subckt TMRDFFSNQX1 Q D CLK SN VDD GND
X0 VDD.t101 a_8357_1050.t5 a_8483_411.t4 ��3	�U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X1 VDD.t113 D.t0 a_5101_1050.t4  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X2 a_5227_411.t4 CLK.t0 VDD.t85 VDD.t84 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X3 a_14869_1051.t5 a_3599_411.t7 a_15533_1051.t7 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X4 VDD.t197 D.t1 a_217_1050.t3  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X5 VDD.t138 a_1265_989.t5 a_1905_1050.t1 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X6 a_9985_1050.t3 a_10111_411.t7 VDD.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X7 GND a_9985_1050.t6 a_11487_103.t0 GND sky130_fd_pr__nfet_01v8 ad=4.9019p pd=4.107u as=0p ps=0u w=0u l=0u
X8 VDD.t50 a_5101_1050.t5 a_6789_1050.t0 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X9 a_15533_1051.t0 a_13367_411.t7 a_15044_209.t4  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X10 a_6789_1050.t1 a_6149_989.t5 VDD.t53 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X11 VDD.t36 a_11033_989.t5 a_11673_1050.t4  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X12 a_3599_411.t0 a_1265_989.t6 VDD.t55 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X13 a_13241_1050.t4 a_10111_411.t8 VDD.t127  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X14 a_1905_1050.t4 a_217_1050.t5 VDD.t97 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X15 VDD.t20 a_11673_1050.t7 a_11033_989.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X16 a_14869_1051.t1 a_8483_411.t8 a_15533_1051.t1 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X17 VDD.t150 a_343_411.t7 a_217_1050.t4  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X18 VDD.t93 a_5227_411.t7 a_5101_1050.t2 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X19 GND a_11673_1050.t8 a_12470_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X20 a_11673_1050.t3 a_11033_989.t6 VDD.t61  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X21 VDD.t87 a_217_1050.t6 a_343_411.t4 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X22 a_3473_1050.t4 a_3599_411.t9 VDD.t184  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X23 VDD.t174 a_13241_1050.t5 a_13367_411.t3 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X24 a_10111_411.t2 CLK.t2 VDD.t18  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X25 GND a_8483_411.t11 a_15430_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X26 a_5227_411.t1 a_6149_989.t7 VDD.t59 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X27 VDD.t186 a_11033_989.t7 a_10111_411.t6  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X28 VDD.t24 a_5227_411.t8 a_8357_1050.t1 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X29 a_13241_1050.t2 a_13367_411.t9 VDD.t148  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X30 a_6149_989.t2 CLK.t3 VDD.t14 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X31 a_14869_1051.t3 a_8483_411.t9 VDD.t110  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X32 VDD.t6 a_6149_989.t8 a_8483_411.t0 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X33 a_13367_411.t4 a_13241_1050.t6 VDD.t176  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X34 GND a_217_1050.t7 a_757_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X35 VDD.t136 a_13367_411.t10 a_14869_1051.t6 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X36 GND D.t3 a_112_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X37 VDD.t12 CLK.t5 a_343_411.t6  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X38 a_3473_1050.t1 a_343_411.t8 VDD.t28 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X39 VDD.t44 a_1905_1050.t7 a_1265_989.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X40 a_8483_411.t6 SN.t2 VDD.t172 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X41 VDD.t180 SN.t3 a_13367_411.t5  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X42 a_10111_411.t0 a_9985_1050.t7 VDD.t74 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X43 GND a_343_411.t9 a_3368_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X44 a_15533_1051.t2 a_8483_411.t10 a_14869_1051.t0  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X45 VDD.t79 a_10111_411.t9 a_9985_1050.t2 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X46 GND a_8357_1050.t7 a_8897_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X47 VDD.t170 SN.t4 a_11673_1050.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X48 a_6149_989.t4 a_6789_1050.t8 VDD.t178 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X49 VDD.t66 a_3473_1050.t5 a_3599_411.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X50 VDD.t131 a_1265_989.t9 a_3599_411.t3 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X51 VDD.t129 a_1265_989.t10 a_343_411.t2  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X52 VDD.t144 a_15044_209.t7 Q.t2 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X53 a_8483_411.t3 a_8357_1050.t6 VDD.t99  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X54 VDD.t42 a_11033_989.t9 a_13367_411.t0 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X55 VDD.t34 a_5101_1050.t6 a_5227_411.t6  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X56 a_8483_411.t1 a_6149_989.t10 VDD.t72 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X57 a_15533_1051.t4 a_3599_411.t10 a_14869_1051.t4  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X58 a_217_1050.t2 D.t4 VDD.t191 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X59 VDD.t77 D.t5 a_9985_1050.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X60 a_1905_1050.t0 a_1265_989.t11 VDD.t125 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X61 GND D.t6 a_9880_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X62 a_6789_1050.t4 a_5101_1050.t7 VDD.t134  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X63 VDD.t46 a_9985_1050.t8 a_11673_1050.t6 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X64 GND a_217_1050.t8 a_1719_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X65 a_15044_209.t3 a_13367_411.t12 a_15533_1051.t3  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X66 VDD.t168 SN.t7 a_3599_411.t5 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X67 VDD.t166 SN.t8 a_6789_1050.t6  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X68 a_11033_989.t1 a_11673_1050.t9 VDD.t26 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X69 a_1905_1050.t6 SN.t9 VDD.t164  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X70 a_5101_1050.t1 a_5227_411.t10 VDD.t91 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X71 a_217_1050.t1 a_343_411.t10 VDD.t32  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X72 GND a_10111_411.t12 a_13136_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X73 GND a_1905_1050.t8 a_2702_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X74 a_6789_1050.t5 SN.t10 VDD.t162 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X75 a_15044_209.t1 a_3599_411.t11 a_15533_1051.t6  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X76 VDD.t140 a_9985_1050.t9 a_10111_411.t3 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X77 GND a_13241_1050.t7 a_13781_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X78 a_343_411.t3 a_217_1050.t9 VDD.t8  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X79 VDD.t107 a_8483_411.t12 a_8357_1050.t2 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X80 GND a_5227_411.t12 a_8252_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X81 Q a_15044_209.t8 GND.t28 GND sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=0p ps=0u w=0u l=0u
X82 VDD.t70 a_6149_989.t12 a_6789_1050.t2  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X83 GND a_5101_1050.t8 a_5641_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X84 VDD.t119 a_10111_411.t11 a_13241_1050.t3 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X85 a_10111_411.t4 a_11033_989.t11 VDD.t142  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X86 VDD.t16 a_217_1050.t10 a_1905_1050.t3 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X87 a_8357_1050.t0 a_5227_411.t11 VDD.t22  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X88 VDD.t146 a_6789_1050.t9 a_6149_989.t3 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X89 a_11033_989.t4 CLK.t8 VDD.t3  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X90 GND a_8483_411.t15 a_14764_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X91 a_5101_1050.t3 D.t7 VDD.t123 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X92 a_343_411.t5 CLK.t10 VDD.t10  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X93 a_14869_1051.t7 a_13367_411.t13 VDD.t199 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X94 a_9985_1050.t0 D.t8 VDD.t63  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X95 a_13367_411.t2 SN.t12 VDD.t160 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X96 a_1265_989.t4 a_1905_1050.t9 VDD.t193  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X97 VDD.t117 a_3599_411.t13 a_3473_1050.t3 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X98 VDD.t40 CLK.t11 a_10111_411.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X99 a_11673_1050.t0 SN.t13 VDD.t158 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X100 VDD.t57 CLK.t12 a_1265_989.t2  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X101 GND a_5101_1050.t10 a_6603_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X102 VDD.t68 a_6149_989.t13 a_5227_411.t2 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X103 VDD.t48 a_13367_411.t14 a_13241_1050.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X104 a_8357_1050.t3 a_8483_411.t13 VDD.t105 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X105 a_3599_411.t6 a_3473_1050.t6 VDD.t182  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X106 VDD.t30 CLK.t13 a_6149_989.t1 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X107 GND a_3473_1050.t7 a_4013_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X108 VDD.t103 a_8483_411.t14 a_14869_1051.t2  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X109 Q.t1 a_15044_209.t9 VDD.t195 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X110 a_343_411.t1 a_1265_989.t13 VDD.t95  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X111 VDD.t38 a_343_411.t12 a_3473_1050.t0 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X112 a_5227_411.t5 a_5101_1050.t9 VDD.t81  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X113 VDD.t156 SN.t15 a_8483_411.t5 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X114 a_13367_411.t1 a_11033_989.t13 VDD.t115  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X115 GND a_6789_1050.t7 a_7586_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X116 a_1265_989.t1 CLK.t14 VDD.t189 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X117 VDD.t154 SN.t16 a_1905_1050.t5  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X118 GND a_9985_1050.t5 a_10525_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X119 GND a_3599_411.t8 a_16096_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X120 GND D.t2 a_4996_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X121 a_11673_1050.t5 a_9985_1050.t10 VDD.t89 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X122 VDD.t83 CLK.t15 a_5227_411.t3  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X123 a_15533_1051.t5 a_3599_411.t15 a_15044_209.t0 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X124 a_3599_411.t4 SN.t17 VDD.t152  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X125 VDD.t121 CLK.t17 a_11033_989.t3 0���0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
C0 SN VDD 1.76fF
C1 Q VDD 1.05fF
C2 SN D 9.38fF
C3 SN CLK 0.46fF
C4 VDD D 0.95fF
C5 VDD CLK 7.98fF
C6 D CLK 0.39fF
R0 a_8357_1050.n3 a_8357_1050.t5 512.525
R1 a_8357_1050.n4 a_8357_1050.t7 417.109
R2 a_8357_1050.n3 a_8357_1050.t6 371.139
R3 a_8357_1050.n7 a_8357_1050.n5 367.82
R4 a_8357_1050.n4 a_8357_1050.n3 179.837
R5 a_8357_1050.n2 a_8357_1050.n1 157.964
R6 a_8357_1050.n5 a_8357_1050.n2 104.282
R7 a_8357_1050.n2 a_8357_1050.n0 91.706
R8 a_8357_1050.n7 a_8357_1050.n6 15.218
R9 a_8357_1050.n0 a_8357_1050.t2 14.282
R10 a_8357_1050.n0 a_8357_1050.t3 14.282
R11 a_8357_1050.n1 a_8357_1050.t1 14.282
R12 a_8357_1050.n1 a_8357_1050.t0 14.282
R13 a_8357_1050.n8 a_8357_1050.n7 12.014
R14 a_8357_1050.n5 a_8357_1050.n4 10.615
R15 a_8483_411.n8 a_8483_411.t14 512.525
R16 a_8483_411.n6 a_8483_411.t8 477.179
R17 a_8483_411.n11 a_8483_411.t12 472.359
R18 a_8483_411.n7 a_8483_411.t11 440.954
R19 a_8483_411.n6 a_8483_411.t10 406.485
R20 a_8483_411.n11 a_8483_411.t13 384.527
R21 a_8483_411.n8 a_8483_411.t9 371.139
R22 a_8483_411.n10 a_8483_411.t15 350.777
R23 a_8483_411.n12 a_8483_411.t7 314.896
R24 a_8483_411.n16 a_8483_411.n14 308.216
R25 a_8483_411.n12 a_8483_411.n11 182.814
R26 a_8483_411.n14 a_8483_411.n5 179.199
R27 a_8483_411.n4 a_8483_411.n3 161.352
R28 a_8483_411.n5 a_8483_411.n1 95.095
R29 a_8483_411.n4 a_8483_411.n2 95.095
R30 a_8483_411.n10 a_8483_411.n9 83.75
R31 a_8483_411.n9 a_8483_411.n8 77.972
R32 a_8483_411.n5 a_8483_411.n4 66.258
R33 a_8483_411.n17 a_8483_411.n0 55.263
R34 a_8483_411.n16 a_8483_411.n15 30
R35 a_8483_411.n17 a_8483_411.n16 23.684
R36 a_8483_411.n13 a_8483_411.n10 23.649
R37 a_8483_411.n7 a_8483_411.n6 21.4
R38 a_8483_411.n1 a_8483_411.t0 14.282
R39 a_8483_411.n1 a_8483_411.t1 14.282
R40 a_8483_411.n2 a_8483_411.t5 14.282
R41 a_8483_411.n2 a_8483_411.t6 14.282
R42 a_8483_411.n3 a_8483_411.t4 14.282
R43 a_8483_411.n3 a_8483_411.t3 14.282
R44 a_8483_411.n13 a_8483_411.n12 8.685
R45 a_8483_411.n9 a_8483_411.n7 6.833
R46 a_8483_411.n14 a_8483_411.n13 4.65
R47 VDD.n790 VDD.n779 144.705
R48 VDD.n865 VDD.n858 144.705
R49 VDD.n940 VDD.n933 144.705
R50 VDD.n997 VDD.n990 144.705
R51 VDD.n1054 VDD.n1047 144.705
R52 VDD.n1129 VDD.n1122 144.705
R53 VDD.n1186 VDD.n1179 144.705
R54 VDD.n1261 VDD.n1254 144.705
R55 VDD.n1336 VDD.n1329 144.705
R56 VDD.n700 VDD.n693 144.705
R57 VDD.n1393 VDD.n1386 144.705
R58 VDD.n625 VDD.n618 144.705
R59 VDD.n568 VDD.n561 144.705
R60 VDD.n493 VDD.n486 144.705
R61 VDD.n418 VDD.n411 144.705
R62 VDD.n361 VDD.n354 144.705
R63 VDD.n304 VDD.n297 144.705
R64 VDD.n229 VDD.n222 144.705
R65 VDD.n172 VDD.n165 144.705
R66 VDD.n119 VDD.n112 144.705
R67 VDD.n66 VDD.n55 144.705
R68 VDD.n832 VDD.t129 143.754
R69 VDD.n907 VDD.t138 143.754
R70 VDD.n1096 VDD.t131 143.754
R71 VDD.n1228 VDD.t68 143.754
R72 VDD.n1303 VDD.t70 143.754
R73 VDD.n634 VDD.t6 143.754
R74 VDD.n502 VDD.t186 143.754
R75 VDD.n427 VDD.t36 143.754
R76 VDD.n238 VDD.t42 143.754
R77 VDD.n757 VDD.t150 143.754
R78 VDD.n965 VDD.t57 143.754
R79 VDD.n1022 VDD.t117 143.754
R80 VDD.n1154 VDD.t93 143.754
R81 VDD.n1361 VDD.t30 143.754
R82 VDD.n703 VDD.t107 143.754
R83 VDD.n571 VDD.t79 143.754
R84 VDD.n364 VDD.t121 143.754
R85 VDD.n307 VDD.t48 143.754
R86 VDD.n197 VDD.t110 135.539
R87 VDD.n175 VDD.t136 135.539
R88 VDD.n735 VDD.t191 135.17
R89 VDD.n797 VDD.t8 135.17
R90 VDD.n872 VDD.t97 135.17
R91 VDD.n943 VDD.t193 135.17
R92 VDD.n1000 VDD.t28 135.17
R93 VDD.n1061 VDD.t182 135.17
R94 VDD.n1132 VDD.t123 135.17
R95 VDD.n1193 VDD.t81 135.17
R96 VDD.n1268 VDD.t134 135.17
R97 VDD.n1339 VDD.t178 135.17
R98 VDD.n1396 VDD.t22 135.17
R99 VDD.n664 VDD.t99 135.17
R100 VDD.n593 VDD.t63 135.17
R101 VDD.n532 VDD.t74 135.17
R102 VDD.n457 VDD.t89 135.17
R103 VDD.n386 VDD.t26 135.17
R104 VDD.n329 VDD.t127 135.17
R105 VDD.n268 VDD.t176 135.17
R106 VDD.n35 VDD.t195 135.17
R107 VDD.n24 VDD.t144 135.17
R108 VDD.n185 VDD.n184 129.849
R109 VDD.n749 VDD.n748 129.472
R110 VDD.n807 VDD.n806 129.472
R111 VDD.n823 VDD.n822 129.472
R112 VDD.n882 VDD.n881 129.472
R113 VDD.n898 VDD.n897 129.472
R114 VDD.n957 VDD.n956 129.472
R115 VDD.n1014 VDD.n1013 129.472
R116 VDD.n1071 VDD.n1070 129.472
R117 VDD.n1087 VDD.n1086 129.472
R118 VDD.n1146 VDD.n1145 129.472
R119 VDD.n1203 VDD.n1202 129.472
R120 VDD.n1219 VDD.n1218 129.472
R121 VDD.n1278 VDD.n1277 129.472
R122 VDD.n1294 VDD.n1293 129.472
R123 VDD.n1353 VDD.n1352 129.472
R124 VDD.n1410 VDD.n1409 129.472
R125 VDD.n655 VDD.n654 129.472
R126 VDD.n643 VDD.n642 129.472
R127 VDD.n581 VDD.n580 129.472
R128 VDD.n523 VDD.n522 129.472
R129 VDD.n511 VDD.n510 129.472
R130 VDD.n448 VDD.n447 129.472
R131 VDD.n436 VDD.n435 129.472
R132 VDD.n374 VDD.n373 129.472
R133 VDD.n317 VDD.n316 129.472
R134 VDD.n259 VDD.n258 129.472
R135 VDD.n247 VDD.n246 129.472
R136 VDD.n51 VDD.n50 92.5
R137 VDD.n49 VDD.n48 92.5
R138 VDD.n47 VDD.n46 92.5
R139 VDD.n45 VDD.n44 92.5
R140 VDD.n53 VDD.n52 92.5
R141 VDD.n108 VDD.n107 92.5
R142 VDD.n106 VDD.n105 92.5
R143 VDD.n104 VDD.n103 92.5
R144 VDD.n102 VDD.n101 92.5
R145 VDD.n110 VDD.n109 92.5
R146 VDD.n161 VDD.n160 92.5
R147 VDD.n159 VDD.n158 92.5
R148 VDD.n157 VDD.n156 92.5
R149 VDD.n155 VDD.n154 92.5
R150 VDD.n163 VDD.n162 92.5
R151 VDD.n218 VDD.n217 92.5
R152 VDD.n216 VDD.n215 92.5
R153 VDD.n214 VDD.n213 92.5
R154 VDD.n212 VDD.n211 92.5
R155 VDD.n220 VDD.n219 92.5
R156 VDD.n293 VDD.n292 92.5
R157 VDD.n291 VDD.n290 92.5
R158 VDD.n289 VDD.n288 92.5
R159 VDD.n287 VDD.n286 92.5
R160 VDD.n295 VDD.n294 92.5
R161 VDD.n350 VDD.n349 92.5
R162 VDD.n348 VDD.n347 92.5
R163 VDD.n346 VDD.n345 92.5
R164 VDD.n344 VDD.n343 92.5
R165 VDD.n352 VDD.n351 92.5
R166 VDD.n407 VDD.n406 92.5
R167 VDD.n405 VDD.n404 92.5
R168 VDD.n403 VDD.n402 92.5
R169 VDD.n401 VDD.n400 92.5
R170 VDD.n409 VDD.n408 92.5
R171 VDD.n482 VDD.n481 92.5
R172 VDD.n480 VDD.n479 92.5
R173 VDD.n478 VDD.n477 92.5
R174 VDD.n476 VDD.n475 92.5
R175 VDD.n484 VDD.n483 92.5
R176 VDD.n557 VDD.n556 92.5
R177 VDD.n555 VDD.n554 92.5
R178 VDD.n553 VDD.n552 92.5
R179 VDD.n551 VDD.n550 92.5
R180 VDD.n559 VDD.n558 92.5
R181 VDD.n614 VDD.n613 92.5
R182 VDD.n612 VDD.n611 92.5
R183 VDD.n610 VDD.n609 92.5
R184 VDD.n608 VDD.n607 92.5
R185 VDD.n616 VDD.n615 92.5
R186 VDD.n689 VDD.n688 92.5
R187 VDD.n687 VDD.n686 92.5
R188 VDD.n685 VDD.n684 92.5
R189 VDD.n683 VDD.n682 92.5
R190 VDD.n691 VDD.n690 92.5
R191 VDD.n1382 VDD.n1381 92.5
R192 VDD.n1380 VDD.n1379 92.5
R193 VDD.n1378 VDD.n1377 92.5
R194 VDD.n1376 VDD.n1375 92.5
R195 VDD.n1384 VDD.n1383 92.5
R196 VDD.n1325 VDD.n1324 92.5
R197 VDD.n1323 VDD.n1322 92.5
R198 VDD.n1321 VDD.n1320 92.5
R199 VDD.n1319 VDD.n1318 92.5
R200 VDD.n1327 VDD.n1326 92.5
R201 VDD.n1250 VDD.n1249 92.5
R202 VDD.n1248 VDD.n1247 92.5
R203 VDD.n1246 VDD.n1245 92.5
R204 VDD.n1244 VDD.n1243 92.5
R205 VDD.n1252 VDD.n1251 92.5
R206 VDD.n1175 VDD.n1174 92.5
R207 VDD.n1173 VDD.n1172 92.5
R208 VDD.n1171 VDD.n1170 92.5
R209 VDD.n1169 VDD.n1168 92.5
R210 VDD.n1177 VDD.n1176 92.5
R211 VDD.n1118 VDD.n1117 92.5
R212 VDD.n1116 VDD.n1115 92.5
R213 VDD.n1114 VDD.n1113 92.5
R214 VDD.n1112 VDD.n1111 92.5
R215 VDD.n1120 VDD.n1119 92.5
R216 VDD.n1043 VDD.n1042 92.5
R217 VDD.n1041 VDD.n1040 92.5
R218 VDD.n1039 VDD.n1038 92.5
R219 VDD.n1037 VDD.n1036 92.5
R220 VDD.n1045 VDD.n1044 92.5
R221 VDD.n986 VDD.n985 92.5
R222 VDD.n984 VDD.n983 92.5
R223 VDD.n982 VDD.n981 92.5
R224 VDD.n980 VDD.n979 92.5
R225 VDD.n988 VDD.n987 92.5
R226 VDD.n929 VDD.n928 92.5
R227 VDD.n927 VDD.n926 92.5
R228 VDD.n925 VDD.n924 92.5
R229 VDD.n923 VDD.n922 92.5
R230 VDD.n931 VDD.n930 92.5
R231 VDD.n854 VDD.n853 92.5
R232 VDD.n852 VDD.n851 92.5
R233 VDD.n850 VDD.n849 92.5
R234 VDD.n848 VDD.n847 92.5
R235 VDD.n856 VDD.n855 92.5
R236 VDD.n775 VDD.n774 92.5
R237 VDD.n773 VDD.n772 92.5
R238 VDD.n771 VDD.n770 92.5
R239 VDD.n769 VDD.n768 92.5
R240 VDD.n777 VDD.n776 92.5
R241 VDD.n723 VDD.n722 92.5
R242 VDD.n721 VDD.n720 92.5
R243 VDD.n719 VDD.n718 92.5
R244 VDD.n717 VDD.n716 92.5
R245 VDD.n725 VDD.n724 92.5
R246 VDD.n14 VDD.n1 92.5
R247 VDD.n5 VDD.n4 92.5
R248 VDD.n7 VDD.n6 92.5
R249 VDD.n9 VDD.n8 92.5
R250 VDD.n11 VDD.n10 92.5
R251 VDD.n13 VDD.n12 92.5
R252 VDD.n21 VDD.n20 92.059
R253 VDD.n65 VDD.n64 92.059
R254 VDD.n118 VDD.n117 92.059
R255 VDD.n171 VDD.n170 92.059
R256 VDD.n228 VDD.n227 92.059
R257 VDD.n303 VDD.n302 92.059
R258 VDD.n360 VDD.n359 92.059
R259 VDD.n417 VDD.n416 92.059
R260 VDD.n492 VDD.n491 92.059
R261 VDD.n567 VDD.n566 92.059
R262 VDD.n624 VDD.n623 92.059
R263 VDD.n699 VDD.n698 92.059
R264 VDD.n1392 VDD.n1391 92.059
R265 VDD.n1335 VDD.n1334 92.059
R266 VDD.n1260 VDD.n1259 92.059
R267 VDD.n1185 VDD.n1184 92.059
R268 VDD.n1128 VDD.n1127 92.059
R269 VDD.n1053 VDD.n1052 92.059
R270 VDD.n996 VDD.n995 92.059
R271 VDD.n939 VDD.n938 92.059
R272 VDD.n864 VDD.n863 92.059
R273 VDD.n789 VDD.n788 92.059
R274 VDD.n731 VDD.n730 92.059
R275 VDD.n20 VDD.n16 67.194
R276 VDD.n20 VDD.n17 67.194
R277 VDD.n20 VDD.n18 67.194
R278 VDD.n20 VDD.n19 67.194
R279 VDD.n715 VDD.n714 44.141
R280 VDD.n846 VDD.n845 44.141
R281 VDD.n921 VDD.n920 44.141
R282 VDD.n978 VDD.n977 44.141
R283 VDD.n1035 VDD.n1034 44.141
R284 VDD.n1110 VDD.n1109 44.141
R285 VDD.n1167 VDD.n1166 44.141
R286 VDD.n1242 VDD.n1241 44.141
R287 VDD.n1317 VDD.n1316 44.141
R288 VDD.n1374 VDD.n1373 44.141
R289 VDD.n681 VDD.n680 44.141
R290 VDD.n606 VDD.n605 44.141
R291 VDD.n549 VDD.n548 44.141
R292 VDD.n474 VDD.n473 44.141
R293 VDD.n399 VDD.n398 44.141
R294 VDD.n342 VDD.n341 44.141
R295 VDD.n285 VDD.n284 44.141
R296 VDD.n210 VDD.n209 44.141
R297 VDD.n153 VDD.n152 44.141
R298 VDD.n100 VDD.n99 44.141
R299 VDD.n5 VDD.n3 44.141
R300 VDD.n845 VDD.n843 44.107
R301 VDD.n920 VDD.n918 44.107
R302 VDD.n977 VDD.n975 44.107
R303 VDD.n1034 VDD.n1032 44.107
R304 VDD.n1109 VDD.n1107 44.107
R305 VDD.n1166 VDD.n1164 44.107
R306 VDD.n1241 VDD.n1239 44.107
R307 VDD.n1316 VDD.n1314 44.107
R308 VDD.n1373 VDD.n1371 44.107
R309 VDD.n680 VDD.n678 44.107
R310 VDD.n605 VDD.n603 44.107
R311 VDD.n548 VDD.n546 44.107
R312 VDD.n473 VDD.n471 44.107
R313 VDD.n398 VDD.n396 44.107
R314 VDD.n341 VDD.n339 44.107
R315 VDD.n284 VDD.n282 44.107
R316 VDD.n209 VDD.n207 44.107
R317 VDD.n152 VDD.n150 44.107
R318 VDD.n99 VDD.n97 44.107
R319 VDD.n714 VDD.n712 44.107
R320 VDD.n3 VDD.n2 44.107
R321 VDD.n25 0���0 43.472
R322 VDD.n33 0���0 43.472
R323 VDD.n20 VDD.n15 41.052
R324 VDD.n59 VDD.n57 39.742
R325 VDD.n59 VDD.n58 39.742
R326 VDD.n61 VDD.n60 39.742
R327 VDD.n114 VDD.n113 39.742
R328 VDD.n167 VDD.n166 39.742
R329 VDD.n224 VDD.n223 39.742
R330 VDD.n299 VDD.n298 39.742
R331 VDD.n356 VDD.n355 39.742
R332 VDD.n413 VDD.n412 39.742
R333 VDD.n488 VDD.n487 39.742
R334 VDD.n563 VDD.n562 39.742
R335 VDD.n620 VDD.n619 39.742
R336 VDD.n695 VDD.n694 39.742
R337 VDD.n1388 VDD.n1387 39.742
R338 VDD.n1331 VDD.n1330 39.742
R339 VDD.n1256 VDD.n1255 39.742
R340 VDD.n1181 VDD.n1180 39.742
R341 VDD.n1124 VDD.n1123 39.742
R342 VDD.n1049 VDD.n1048 39.742
R343 VDD.n992 VDD.n991 39.742
R344 VDD.n935 VDD.n934 39.742
R345 VDD.n860 VDD.n859 39.742
R346 VDD.n727 VDD.n726 39.742
R347 VDD.n787 VDD.n784 39.742
R348 VDD.n787 VDD.n786 39.742
R349 VDD.n783 VDD.n782 39.742
R350 VDD.n99 VDD.n98 38
R351 VDD.n152 VDD.n151 38
R352 VDD.n209 VDD.n208 38
R353 VDD.n284 VDD.n283 38
R354 VDD.n341 VDD.n340 38
R355 VDD.n398 VDD.n397 38
R356 VDD.n473 VDD.n472 38
R357 VDD.n548 VDD.n547 38
R358 VDD.n605 VDD.n604 38
R359 VDD.n680 VDD.n679 38
R360 VDD.n1373 VDD.n1372 38
R361 VDD.n1316 VDD.n1315 38
R362 VDD.n1241 VDD.n1240 38
R363 VDD.n1166 VDD.n1165 38
R364 VDD.n1109 VDD.n1108 38
R365 VDD.n1034 VDD.n1033 38
R366 VDD.n977 VDD.n976 38
R367 VDD.n920 VDD.n919 38
R368 VDD.n845 VDD.n844 38
R369 VDD.n714 VDD.n713 38
R370 VDD.n843 VDD.n842 36.774
R371 VDD.n918 VDD.n917 36.774
R372 VDD.n975 VDD.n974 36.774
R373 VDD.n1032 VDD.n1031 36.774
R374 VDD.n1107 VDD.n1106 36.774
R375 VDD.n1164 VDD.n1163 36.774
R376 VDD.n1239 VDD.n1238 36.774
R377 VDD.n1314 VDD.n1313 36.774
R378 VDD.n1371 VDD.n1370 36.774
R379 VDD.n678 VDD.n677 36.774
R380 VDD.n603 VDD.n602 36.774
R381 VDD.n546 VDD.n545 36.774
R382 VDD.n471 VDD.n470 36.774
R383 VDD.n396 VDD.n395 36.774
R384 VDD.n339 VDD.n338 36.774
R385 VDD.n282 VDD.n281 36.774
R386 VDD.n207 VDD.n206 36.774
R387 VDD.n150 VDD.n149 36.774
R388 VDD.n97 VDD.n96 36.774
R389 VDD.n57 VDD.n56 36.774
R390 VDD.n786 VDD.n785 36.774
R391 VDD.n240 0���0 35.8
R392 VDD.n429  35.8
R393 VDD.n504  35.8
R394 VDD.n636 0���0 35.8
R395 VDD.n1297  35.8
R396 VDD.n1222 0���0 35.8
R397 VDD.n1090 0���0 35.8
R398 VDD.n901 0���0 35.8
R399 VDD.n826  35.8
R400 VDD.n264  33.243
R401 VDD.n453 0���0 33.243
R402 VDD.n528 0���0 33.243
R403 VDD.n660  33.243
R404 VDD.n1273  33.243
R405 VDD.n1198  33.243
R406 VDD.n1066  33.243
R407 VDD.n877 0���0 33.243
R408 VDD.n802  33.243
R409 VDD.n1 VDD.n0 30.923
R410 VDD.n64 VDD.n62 26.38
R411 VDD.n64 VDD.n61 26.38
R412 VDD.n64 VDD.n59 26.38
R413 VDD.n64 VDD.n63 26.38
R414 VDD.n117 VDD.n115 26.38
R415 VDD.n117 VDD.n114 26.38
R416 VDD.n117 VDD.n116 26.38
R417 VDD.n170 VDD.n168 26.38
R418 VDD.n170 VDD.n167 26.38
R419 VDD.n170 VDD.n169 26.38
R420 VDD.n227 VDD.n225 26.38
R421 VDD.n227 VDD.n224 26.38
R422 VDD.n227 VDD.n226 26.38
R423 VDD.n302 VDD.n300 26.38
R424 VDD.n302 VDD.n299 26.38
R425 VDD.n302 VDD.n301 26.38
R426 VDD.n359 VDD.n357 26.38
R427 VDD.n359 VDD.n356 26.38
R428 VDD.n359 VDD.n358 26.38
R429 VDD.n416 VDD.n414 26.38
R430 VDD.n416 VDD.n413 26.38
R431 VDD.n416 VDD.n415 26.38
R432 VDD.n491 VDD.n489 26.38
R433 VDD.n491 VDD.n488 26.38
R434 VDD.n491 VDD.n490 26.38
R435 VDD.n566 VDD.n564 26.38
R436 VDD.n566 VDD.n563 26.38
R437 VDD.n566 VDD.n565 26.38
R438 VDD.n623 VDD.n621 26.38
R439 VDD.n623 VDD.n620 26.38
R440 VDD.n623 VDD.n622 26.38
R441 VDD.n698 VDD.n696 26.38
R442 VDD.n698 VDD.n695 26.38
R443 VDD.n698 VDD.n697 26.38
R444 VDD.n1391 VDD.n1389 26.38
R445 VDD.n1391 VDD.n1388 26.38
R446 VDD.n1391 VDD.n1390 26.38
R447 VDD.n1334 VDD.n1332 26.38
R448 VDD.n1334 VDD.n1331 26.38
R449 VDD.n1334 VDD.n1333 26.38
R450 VDD.n1259 VDD.n1257 26.38
R451 VDD.n1259 VDD.n1256 26.38
R452 VDD.n1259 VDD.n1258 26.38
R453 VDD.n1184 VDD.n1182 26.38
R454 VDD.n1184 VDD.n1181 26.38
R455 VDD.n1184 VDD.n1183 26.38
R456 VDD.n1127 VDD.n1125 26.38
R457 VDD.n1127 VDD.n1124 26.38
R458 VDD.n1127 VDD.n1126 26.38
R459 VDD.n1052 VDD.n1050 26.38
R460 VDD.n1052 VDD.n1049 26.38
R461 VDD.n1052 VDD.n1051 26.38
R462 VDD.n995 VDD.n993 26.38
R463 VDD.n995 VDD.n992 26.38
R464 VDD.n995 VDD.n994 26.38
R465 VDD.n938 VDD.n936 26.38
R466 VDD.n938 VDD.n935 26.38
R467 VDD.n938 VDD.n937 26.38
R468 VDD.n863 VDD.n861 26.38
R469 VDD.n863 VDD.n860 26.38
R470 VDD.n863 VDD.n862 26.38
R471 VDD.n730 VDD.n728 26.38
R472 VDD.n730 VDD.n727 26.38
R473 VDD.n730 VDD.n729 26.38
R474 VDD.n788 VDD.n787 26.38
R475 VDD.n788 VDD.n783 26.38
R476 VDD.n788 VDD.n781 26.38
R477 VDD.n788 VDD.n780 26.38
R478 VDD.n733 VDD.n725 22.915
R479 VDD.n23 VDD.n14 22.915
R480 VDD.n73  20.457
R481 VDD.n137  20.457
R482 VDD.n180 0���0 20.457
R483 VDD.n312  20.457
R484 VDD.n369 0���0 20.457
R485 VDD.n576 0���0 20.457
R486 VDD.n708 0���0 20.457
R487 VDD.n1357 0���0 20.457
R488 VDD.n1150 0���0 20.457
R489 VDD.n1018 0���0 20.457
R490 VDD.n961  20.457
R491 VDD.n753  20.457
R492 VDD.n84  17.9
R493 VDD.n126 0���0 17.9
R494 VDD.n193  17.9
R495 VDD.n325  17.9
R496 VDD.n382 0���0 17.9
R497 VDD.n589  17.9
R498 VDD.n1401  17.9
R499 VDD.n1344 0���0 17.9
R500 VDD.n1137 0���0 17.9
R501 VDD.n1005 0���0 17.9
R502 VDD.n948  17.9
R503 VDD.n740 0���0 17.9
R504 VDD.n244  15.343
R505 VDD.n433  15.343
R506 VDD.n508  15.343
R507 VDD.n640 0���0 15.343
R508 VDD.n1291 0���0 15.343
R509 VDD.n1216 0���0 15.343
R510 VDD.n1084 0���0 15.343
R511 VDD.n895 0���0 15.343
R512 VDD.n820  15.343
R513 VDD.n725 VDD.n723 14.864
R514 VDD.n723 VDD.n721 14.864
R515 VDD.n721 VDD.n719 14.864
R516 VDD.n719 VDD.n717 14.864
R517 VDD.n717 VDD.n715 14.864
R518 VDD.n856 VDD.n854 14.864
R519 VDD.n854 VDD.n852 14.864
R520 VDD.n852 VDD.n850 14.864
R521 VDD.n850 VDD.n848 14.864
R522 VDD.n848 VDD.n846 14.864
R523 VDD.n931 VDD.n929 14.864
R524 VDD.n929 VDD.n927 14.864
R525 VDD.n927 VDD.n925 14.864
R526 VDD.n925 VDD.n923 14.864
R527 VDD.n923 VDD.n921 14.864
R528 VDD.n988 VDD.n986 14.864
R529 VDD.n986 VDD.n984 14.864
R530 VDD.n984 VDD.n982 14.864
R531 VDD.n982 VDD.n980 14.864
R532 VDD.n980 VDD.n978 14.864
R533 VDD.n1045 VDD.n1043 14.864
R534 VDD.n1043 VDD.n1041 14.864
R535 VDD.n1041 VDD.n1039 14.864
R536 VDD.n1039 VDD.n1037 14.864
R537 VDD.n1037 VDD.n1035 14.864
R538 VDD.n1120 VDD.n1118 14.864
R539 VDD.n1118 VDD.n1116 14.864
R540 VDD.n1116 VDD.n1114 14.864
R541 VDD.n1114 VDD.n1112 14.864
R542 VDD.n1112 VDD.n1110 14.864
R543 VDD.n1177 VDD.n1175 14.864
R544 VDD.n1175 VDD.n1173 14.864
R545 VDD.n1173 VDD.n1171 14.864
R546 VDD.n1171 VDD.n1169 14.864
R547 VDD.n1169 VDD.n1167 14.864
R548 VDD.n1252 VDD.n1250 14.864
R549 VDD.n1250 VDD.n1248 14.864
R550 VDD.n1248 VDD.n1246 14.864
R551 VDD.n1246 VDD.n1244 14.864
R552 VDD.n1244 VDD.n1242 14.864
R553 VDD.n1327 VDD.n1325 14.864
R554 VDD.n1325 VDD.n1323 14.864
R555 VDD.n1323 VDD.n1321 14.864
R556 VDD.n1321 VDD.n1319 14.864
R557 VDD.n1319 VDD.n1317 14.864
R558 VDD.n1384 VDD.n1382 14.864
R559 VDD.n1382 VDD.n1380 14.864
R560 VDD.n1380 VDD.n1378 14.864
R561 VDD.n1378 VDD.n1376 14.864
R562 VDD.n1376 VDD.n1374 14.864
R563 VDD.n691 VDD.n689 14.864
R564 VDD.n689 VDD.n687 14.864
R565 VDD.n687 VDD.n685 14.864
R566 VDD.n685 VDD.n683 14.864
R567 VDD.n683 VDD.n681 14.864
R568 VDD.n616 VDD.n614 14.864
R569 VDD.n614 VDD.n612 14.864
R570 VDD.n612 VDD.n610 14.864
R571 VDD.n610 VDD.n608 14.864
R572 VDD.n608 VDD.n606 14.864
R573 VDD.n559 VDD.n557 14.864
R574 VDD.n557 VDD.n555 14.864
R575 VDD.n555 VDD.n553 14.864
R576 VDD.n553 VDD.n551 14.864
R577 VDD.n551 VDD.n549 14.864
R578 VDD.n484 VDD.n482 14.864
R579 VDD.n482 VDD.n480 14.864
R580 VDD.n480 VDD.n478 14.864
R581 VDD.n478 VDD.n476 14.864
R582 VDD.n476 VDD.n474 14.864
R583 VDD.n409 VDD.n407 14.864
R584 VDD.n407 VDD.n405 14.864
R585 VDD.n405 VDD.n403 14.864
R586 VDD.n403 VDD.n401 14.864
R587 VDD.n401 VDD.n399 14.864
R588 VDD.n352 VDD.n350 14.864
R589 VDD.n350 VDD.n348 14.864
R590 VDD.n348 VDD.n346 14.864
R591 VDD.n346 VDD.n344 14.864
R592 VDD.n344 VDD.n342 14.864
R593 VDD.n295 VDD.n293 14.864
R594 VDD.n293 VDD.n291 14.864
R595 VDD.n291 VDD.n289 14.864
R596 VDD.n289 VDD.n287 14.864
R597 VDD.n287 VDD.n285 14.864
R598 VDD.n220 VDD.n218 14.864
R599 VDD.n218 VDD.n216 14.864
R600 VDD.n216 VDD.n214 14.864
R601 VDD.n214 VDD.n212 14.864
R602 VDD.n212 VDD.n210 14.864
R603 VDD.n163 VDD.n161 14.864
R604 VDD.n161 VDD.n159 14.864
R605 VDD.n159 VDD.n157 14.864
R606 VDD.n157 VDD.n155 14.864
R607 VDD.n155 VDD.n153 14.864
R608 VDD.n110 VDD.n108 14.864
R609 VDD.n108 VDD.n106 14.864
R610 VDD.n106 VDD.n104 14.864
R611 VDD.n104 VDD.n102 14.864
R612 VDD.n102 VDD.n100 14.864
R613 VDD.n53 VDD.n51 14.864
R614 VDD.n51 VDD.n49 14.864
R615 VDD.n49 VDD.n47 14.864
R616 VDD.n47 VDD.n45 14.864
R617 VDD.n45 VDD.n43 14.864
R618 VDD.n43 VDD.n42 14.864
R619 VDD.n777 VDD.n775 14.864
R620 VDD.n775 VDD.n773 14.864
R621 VDD.n773 VDD.n771 14.864
R622 VDD.n771 VDD.n769 14.864
R623 VDD.n769 VDD.n767 14.864
R624 VDD.n767 VDD.n766 14.864
R625 VDD.n14 VDD.n13 14.864
R626 VDD.n13 VDD.n11 14.864
R627 VDD.n11 VDD.n9 14.864
R628 VDD.n9 VDD.n7 14.864
R629 VDD.n7 VDD.n5 14.864
R630 VDD.n67 VDD.n54 14.864
R631 VDD.n120 VDD.n111 14.864
R632 VDD.n173 VDD.n164 14.864
R633 VDD.n230 VDD.n221 14.864
R634 VDD.n305 VDD.n296 14.864
R635 VDD.n362 VDD.n353 14.864
R636 VDD.n419 VDD.n410 14.864
R637 VDD.n494 VDD.n485 14.864
R638 VDD.n569 VDD.n560 14.864
R639 VDD.n626 VDD.n617 14.864
R640 VDD.n701 VDD.n692 14.864
R641 VDD.n1394 VDD.n1385 14.864
R642 VDD.n1337 VDD.n1328 14.864
R643 VDD.n1262 VDD.n1253 14.864
R644 VDD.n1187 VDD.n1178 14.864
R645 VDD.n1130 VDD.n1121 14.864
R646 VDD.n1055 VDD.n1046 14.864
R647 VDD.n998 VDD.n989 14.864
R648 VDD.n941 VDD.n932 14.864
R649 VDD.n866 VDD.n857 14.864
R650 VDD.n791 VDD.n778 14.864
R651 VDD.n748 VDD.t32 14.282
R652 VDD.n748 VDD.t197 14.282
R653 VDD.n806 VDD.t10 14.282
R654 VDD.n806 VDD.t87 14.282
R655 VDD.n822 VDD.t95 14.282
R656 VDD.n822 VDD.t12 14.282
R657 VDD.n881 VDD.t164 14.282
R658 VDD.n881 VDD.t16 14.282
R659 VDD.n897 VDD.t125 14.282
R660 VDD.n897 VDD.t154 14.282
R661 VDD.n956 VDD.t189 14.282
R662 VDD.n956 VDD.t44 14.282
R663 VDD.n1013 VDD.t184 14.282
R664 VDD.n1013 VDD.t38 14.282
R665 VDD.n1070 VDD.t152 14.282
R666 VDD.n1070 VDD.t66 14.282
R667 VDD.n1086 VDD.t55 14.282
R668 VDD.n1086 VDD.t168 14.282
R669 VDD.n1145 VDD.t91 14.282
R670 VDD.n1145 VDD.t113 14.282
R671 VDD.n1202 VDD.t85 14.282
R672 VDD.n1202 VDD.t34 14.282
R673 VDD.n1218 VDD.t59 14.282
R674 VDD.n1218 VDD.t83 14.282
R675 VDD.n1277 VDD.t162 14.282
R676 VDD.n1277 VDD.t50 14.282
R677 VDD.n1293 VDD.t53 14.282
R678 VDD.n1293 VDD.t166 14.282
R679 VDD.n1352 VDD.t14 14.282
R680 VDD.n1352 VDD.t146 14.282
R681 VDD.n1409 VDD.t105 14.282
R682 VDD.n1409 VDD.t24 14.282
R683 VDD.n654 VDD.t172 14.282
R684 VDD.n654 VDD.t101 14.282
R685 VDD.n642 VDD.t72 14.282
R686 VDD.n642 VDD.t156 14.282
R687 VDD.n580 VDD.t1 14.282
R688 VDD.n580 VDD.t77 14.282
R689 VDD.n522 VDD.t18 14.282
R690 VDD.n522 VDD.t140 14.282
R691 VDD.n510 VDD.t142 14.282
R692 VDD.n510 VDD.t40 14.282
R693 VDD.n447 VDD.t158 14.282
R694 VDD.n447 VDD.t46 14.282
R695 VDD.n435 VDD.t61 14.282
R696 VDD.n435 VDD.t170 14.282
R697 VDD.n373 VDD.t3 14.282
R698 VDD.n373 VDD.t20 14.282
R699 VDD.n316 VDD.t148 14.282
R700 VDD.n316 VDD.t119 14.282
R701 VDD.n258 VDD.t160 14.282
R702 VDD.n258 VDD.t174 14.282
R703 VDD.n246 VDD.t115 14.282
R704 VDD.n246 VDD.t180 14.282
R705 VDD.n184 VDD.t199 14.282
R706 VDD.n184 VDD.t103 14.282
R707 VDD.n260 0���0 12.786
R708 VDD.n449 0���0 12.786
R709 VDD.n524 0���0 12.786
R710 VDD.n656 ��3	�U 12.786
R711 VDD.n1279 0���0 12.786
R712 VDD.n1204  12.786
R713 VDD.n1072  12.786
R714 VDD.n883 0���0 12.786
R715 VDD.n808 0���0 12.786
R716 VDD.n187 VDD.n185 9.083
R717 VDD.n319 VDD.n317 9.083
R718 VDD.n376 VDD.n374 9.083
R719 VDD.n583 VDD.n581 9.083
R720 VDD.n1412 VDD.n1410 9.083
R721 VDD.n1355 VDD.n1353 9.083
R722 VDD.n1148 VDD.n1146 9.083
R723 VDD.n1016 VDD.n1014 9.083
R724 VDD.n959 VDD.n957 9.083
R725 VDD.n751 VDD.n749 9.083
R726 VDD.n23 VDD.n22 8.855
R727 VDD.n22 VDD.n21 8.855
R728 VDD.n27 VDD.n26 8.855
R729 VDD.n26 VDD.n25 8.855
R730 VDD.n31 VDD.n30 8.855
R731 VDD.n30 VDD.n29 8.855
R732 VDD.n36 VDD.n34 8.855
R733 VDD.n34 VDD.n33 8.855
R734 VDD.n40 VDD.n39 8.855
R735 VDD.n39 VDD.n38 8.855
R736 VDD.n67 VDD.n66 8.855
R737 VDD.n66 VDD.n65 8.855
R738 VDD.n71 VDD.n70 8.855
R739 VDD.n70 VDD.n69 8.855
R740 VDD.n75 VDD.n74 8.855
R741 VDD.n74 VDD.n73 8.855
R742 VDD.n78 VDD.n77 8.855
R743 VDD.n77  8.855
R744 VDD.n82 VDD.n81 8.855
R745 VDD.n81 VDD.n80 8.855
R746 VDD.n86 VDD.n85 8.855
R747 VDD.n85 VDD.n84 8.855
R748 VDD.n90 VDD.n89 8.855
R749 VDD.n89 VDD.n88 8.855
R750 VDD.n94 VDD.n93 8.855
R751 VDD.n93 VDD.n92 8.855
R752 VDD.n120 VDD.n119 8.855
R753 VDD.n119 VDD.n118 8.855
R754 VDD.n124 VDD.n123 8.855
R755 VDD.n123 VDD.n122 8.855
R756 VDD.n128 VDD.n127 8.855
R757 VDD.n127 VDD.n126 8.855
R758 VDD.n132 VDD.n131 8.855
R759 VDD.n131 VDD.n130 8.855
R760 VDD.n135 VDD.n134 8.855
R761 VDD.n134 0���0 8.855
R762 VDD.n139 VDD.n138 8.855
R763 VDD.n138 VDD.n137 8.855
R764 VDD.n143 VDD.n142 8.855
R765 VDD.n142 VDD.n141 8.855
R766 VDD.n147 VDD.n146 8.855
R767 VDD.n146 VDD.n145 8.855
R768 VDD.n173 VDD.n172 8.855
R769 VDD.n172 VDD.n171 8.855
R770 VDD.n178 VDD.n177 8.855
R771 VDD.n177 VDD.n176 8.855
R772 VDD.n182 VDD.n181 8.855
R773 VDD.n181 VDD.n180 8.855
R774 VDD.n187 VDD.n186 8.855
R775 VDD.n186 0���0 8.855
R776 VDD.n191 VDD.n190 8.855
R777 VDD.n190 VDD.n189 8.855
R778 VDD.n195 VDD.n194 8.855
R779 VDD.n194 VDD.n193 8.855
R780 VDD.n200 VDD.n199 8.855
R781 VDD.n199 VDD.n198 8.855
R782 VDD.n204 VDD.n203 8.855
R783 VDD.n203 VDD.n202 8.855
R784 VDD.n230 VDD.n229 8.855
R785 VDD.n229 VDD.n228 8.855
R786 VDD.n234 VDD.n233 8.855
R787 VDD.n233 VDD.n232 8.855
R788 VDD.n238 VDD.n237 8.855
R789 VDD.n237 VDD.n236 8.855
R790 VDD.n242 VDD.n241 8.855
R791 VDD.n241 VDD.n240 8.855
R792 VDD.n248 VDD.n245 8.855
R793 VDD.n245 VDD.n244 8.855
R794 VDD.n252 VDD.n251 8.855
R795 VDD.n251 VDD.n250 8.855
R796 VDD.n256 VDD.n255 8.855
R797 VDD.n255 VDD.n254 8.855
R798 VDD.n262 VDD.n261 8.855
R799 VDD.n261 VDD.n260 8.855
R800 VDD.n266 VDD.n265 8.855
R801 VDD.n265 VDD.n264 8.855
R802 VDD.n271 VDD.n270 8.855
R803 VDD.n270 VDD.n269 8.855
R804 VDD.n275 VDD.n274 8.855
R805 VDD.n274 VDD.n273 8.855
R806 VDD.n279 VDD.n278 8.855
R807 VDD.n278 VDD.n277 8.855
R808 VDD.n305 VDD.n304 8.855
R809 VDD.n304 VDD.n303 8.855
R810 VDD.n310 VDD.n309 8.855
R811 VDD.n309 VDD.n308 8.855
R812 VDD.n314 VDD.n313 8.855
R813 VDD.n313 VDD.n312 8.855
R814 VDD.n319 VDD.n318 8.855
R815 VDD.n318  8.855
R816 VDD.n323 VDD.n322 8.855
R817 VDD.n322 VDD.n321 8.855
R818 VDD.n327 VDD.n326 8.855
R819 VDD.n326 VDD.n325 8.855
R820 VDD.n332 VDD.n331 8.855
R821 VDD.n331 VDD.n330 8.855
R822 VDD.n336 VDD.n335 8.855
R823 VDD.n335 VDD.n334 8.855
R824 VDD.n362 VDD.n361 8.855
R825 VDD.n361 VDD.n360 8.855
R826 VDD.n367 VDD.n366 8.855
R827 VDD.n366 VDD.n365 8.855
R828 VDD.n371 VDD.n370 8.855
R829 VDD.n370 VDD.n369 8.855
R830 VDD.n376 VDD.n375 8.855
R831 VDD.n375  8.855
R832 VDD.n380 VDD.n379 8.855
R833 VDD.n379 VDD.n378 8.855
R834 VDD.n384 VDD.n383 8.855
R835 VDD.n383 VDD.n382 8.855
R836 VDD.n389 VDD.n388 8.855
R837 VDD.n388 VDD.n387 8.855
R838 VDD.n393 VDD.n392 8.855
R839 VDD.n392 VDD.n391 8.855
R840 VDD.n419 VDD.n418 8.855
R841 VDD.n418 VDD.n417 8.855
R842 VDD.n423 VDD.n422 8.855
R843 VDD.n422 VDD.n421 8.855
R844 VDD.n427 VDD.n426 8.855
R845 VDD.n426 VDD.n425 8.855
R846 VDD.n431 VDD.n430 8.855
R847 VDD.n430 VDD.n429 8.855
R848 VDD.n437 VDD.n434 8.855
R849 VDD.n434 VDD.n433 8.855
R850 VDD.n441 VDD.n440 8.855
R851 VDD.n440 VDD.n439 8.855
R852 VDD.n445 VDD.n444 8.855
R853 VDD.n444 VDD.n443 8.855
R854 VDD.n451 VDD.n450 8.855
R855 VDD.n450 VDD.n449 8.855
R856 VDD.n455 VDD.n454 8.855
R857 VDD.n454 VDD.n453 8.855
R858 VDD.n460 VDD.n459 8.855
R859 VDD.n459 VDD.n458 8.855
R860 VDD.n464 VDD.n463 8.855
R861 VDD.n463 VDD.n462 8.855
R862 VDD.n468 VDD.n467 8.855
R863 VDD.n467 VDD.n466 8.855
R864 VDD.n494 VDD.n493 8.855
R865 VDD.n493 VDD.n492 8.855
R866 VDD.n498 VDD.n497 8.855
R867 VDD.n497 VDD.n496 8.855
R868 VDD.n502 VDD.n501 8.855
R869 VDD.n501 VDD.n500 8.855
R870 VDD.n506 VDD.n505 8.855
R871 VDD.n505 VDD.n504 8.855
R872 VDD.n512 VDD.n509 8.855
R873 VDD.n509 VDD.n508 8.855
R874 VDD.n516 VDD.n515 8.855
R875 VDD.n515 VDD.n514 8.855
R876 VDD.n520 VDD.n519 8.855
R877 VDD.n519 VDD.n518 8.855
R878 VDD.n526 VDD.n525 8.855
R879 VDD.n525 VDD.n524 8.855
R880 VDD.n530 VDD.n529 8.855
R881 VDD.n529 VDD.n528 8.855
R882 VDD.n535 VDD.n534 8.855
R883 VDD.n534 VDD.n533 8.855
R884 VDD.n539 VDD.n538 8.855
R885 VDD.n538 VDD.n537 8.855
R886 VDD.n543 VDD.n542 8.855
R887 VDD.n542 VDD.n541 8.855
R888 VDD.n569 VDD.n568 8.855
R889 VDD.n568 VDD.n567 8.855
R890 VDD.n574 VDD.n573 8.855
R891 VDD.n573 VDD.n572 8.855
R892 VDD.n578 VDD.n577 8.855
R893 VDD.n577 VDD.n576 8.855
R894 VDD.n583 VDD.n582 8.855
R895 VDD.n582  8.855
R896 VDD.n587 VDD.n586 8.855
R897 VDD.n586 VDD.n585 8.855
R898 VDD.n591 VDD.n590 8.855
R899 VDD.n590 VDD.n589 8.855
R900 VDD.n596 VDD.n595 8.855
R901 VDD.n595 VDD.n594 8.855
R902 VDD.n600 VDD.n599 8.855
R903 VDD.n599 VDD.n598 8.855
R904 VDD.n626 VDD.n625 8.855
R905 VDD.n625 VDD.n624 8.855
R906 VDD.n630 VDD.n629 8.855
R907 VDD.n629 VDD.n628 8.855
R908 VDD.n634 VDD.n633 8.855
R909 VDD.n633 VDD.n632 8.855
R910 VDD.n638 VDD.n637 8.855
R911 VDD.n637 VDD.n636 8.855
R912 VDD.n644 VDD.n641 8.855
R913 VDD.n641 VDD.n640 8.855
R914 VDD.n648 VDD.n647 8.855
R915 VDD.n647 VDD.n646 8.855
R916 VDD.n652 VDD.n651 8.855
R917 VDD.n651 VDD.n650 8.855
R918 VDD.n658 VDD.n657 8.855
R919 VDD.n657 VDD.n656 8.855
R920 VDD.n662 VDD.n661 8.855
R921 VDD.n661 VDD.n660 8.855
R922 VDD.n667 VDD.n666 8.855
R923 VDD.n666 VDD.n665 8.855
R924 VDD.n671 VDD.n670 8.855
R925 VDD.n670 VDD.n669 8.855
R926 VDD.n675 VDD.n674 8.855
R927 VDD.n674 VDD.n673 8.855
R928 VDD.n701 VDD.n700 8.855
R929 VDD.n700 VDD.n699 8.855
R930 VDD.n706 VDD.n705 8.855
R931 VDD.n705 VDD.n704 8.855
R932 VDD.n710 VDD.n709 8.855
R933 VDD.n709 VDD.n708 8.855
R934 VDD.n1412 VDD.n1411 8.855
R935 VDD.n1411 0���0 8.855
R936 VDD.n1407 VDD.n1406 8.855
R937 VDD.n1406 VDD.n1405 8.855
R938 VDD.n1403 VDD.n1402 8.855
R939 VDD.n1402 VDD.n1401 8.855
R940 VDD.n1399 VDD.n1398 8.855
R941 VDD.n1398 VDD.n1397 8.855
R942 VDD.n1394 VDD.n1393 8.855
R943 VDD.n1393 VDD.n1392 8.855
R944 VDD.n1368 VDD.n1367 8.855
R945 VDD.n1367 VDD.n1366 8.855
R946 VDD.n1364 VDD.n1363 8.855
R947 VDD.n1363 VDD.n1362 8.855
R948 VDD.n1359 VDD.n1358 8.855
R949 VDD.n1358 VDD.n1357 8.855
R950 VDD.n1355 VDD.n1354 8.855
R951 VDD.n1354 0���0 8.855
R952 VDD.n1350 VDD.n1349 8.855
R953 VDD.n1349 VDD.n1348 8.855
R954 VDD.n1346 VDD.n1345 8.855
R955 VDD.n1345 VDD.n1344 8.855
R956 VDD.n1342 VDD.n1341 8.855
R957 VDD.n1341 VDD.n1340 8.855
R958 VDD.n1337 VDD.n1336 8.855
R959 VDD.n1336 VDD.n1335 8.855
R960 VDD.n1311 VDD.n1310 8.855
R961 VDD.n1310 VDD.n1309 8.855
R962 VDD.n1307 VDD.n1306 8.855
R963 VDD.n1306 VDD.n1305 8.855
R964 VDD.n1303 VDD.n1302 8.855
R965 VDD.n1302 VDD.n1301 8.855
R966 VDD.n1299 VDD.n1298 8.855
R967 VDD.n1298 VDD.n1297 8.855
R968 VDD.n1295 VDD.n1292 8.855
R969 VDD.n1292 VDD.n1291 8.855
R970 VDD.n1289 VDD.n1288 8.855
R971 VDD.n1288 VDD.n1287 8.855
R972 VDD.n1285 VDD.n1284 8.855
R973 VDD.n1284 VDD.n1283 8.855
R974 VDD.n1281 VDD.n1280 8.855
R975 VDD.n1280 VDD.n1279 8.855
R976 VDD.n1275 VDD.n1274 8.855
R977 VDD.n1274 VDD.n1273 8.855
R978 VDD.n1271 VDD.n1270 8.855
R979 VDD.n1270 VDD.n1269 8.855
R980 VDD.n1266 VDD.n1265 8.855
R981 VDD.n1265 VDD.n1264 8.855
R982 VDD.n1262 VDD.n1261 8.855
R983 VDD.n1261 VDD.n1260 8.855
R984 VDD.n1236 VDD.n1235 8.855
R985 VDD.n1235 VDD.n1234 8.855
R986 VDD.n1232 VDD.n1231 8.855
R987 VDD.n1231 VDD.n1230 8.855
R988 VDD.n1228 VDD.n1227 8.855
R989 VDD.n1227 VDD.n1226 8.855
R990 VDD.n1224 VDD.n1223 8.855
R991 VDD.n1223 VDD.n1222 8.855
R992 VDD.n1220 VDD.n1217 8.855
R993 VDD.n1217 VDD.n1216 8.855
R994 VDD.n1214 VDD.n1213 8.855
R995 VDD.n1213 VDD.n1212 8.855
R996 VDD.n1210 VDD.n1209 8.855
R997 VDD.n1209 VDD.n1208 8.855
R998 VDD.n1206 VDD.n1205 8.855
R999 VDD.n1205 VDD.n1204 8.855
R1000 VDD.n1200 VDD.n1199 8.855
R1001 VDD.n1199 VDD.n1198 8.855
R1002 VDD.n1196 VDD.n1195 8.855
R1003 VDD.n1195 VDD.n1194 8.855
R1004 VDD.n1191 VDD.n1190 8.855
R1005 VDD.n1190 VDD.n1189 8.855
R1006 VDD.n1187 VDD.n1186 8.855
R1007 VDD.n1186 VDD.n1185 8.855
R1008 VDD.n1161 VDD.n1160 8.855
R1009 VDD.n1160 VDD.n1159 8.855
R1010 VDD.n1157 VDD.n1156 8.855
R1011 VDD.n1156 VDD.n1155 8.855
R1012 VDD.n1152 VDD.n1151 8.855
R1013 VDD.n1151 VDD.n1150 8.855
R1014 VDD.n1148 VDD.n1147 8.855
R1015 VDD.n1147 0���0 8.855
R1016 VDD.n1143 VDD.n1142 8.855
R1017 VDD.n1142 VDD.n1141 8.855
R1018 VDD.n1139 VDD.n1138 8.855
R1019 VDD.n1138 VDD.n1137 8.855
R1020 VDD.n1135 VDD.n1134 8.855
R1021 VDD.n1134 VDD.n1133 8.855
R1022 VDD.n1130 VDD.n1129 8.855
R1023 VDD.n1129 VDD.n1128 8.855
R1024 VDD.n1104 VDD.n1103 8.855
R1025 VDD.n1103 VDD.n1102 8.855
R1026 VDD.n1100 VDD.n1099 8.855
R1027 VDD.n1099 VDD.n1098 8.855
R1028 VDD.n1096 VDD.n1095 8.855
R1029 VDD.n1095 VDD.n1094 8.855
R1030 VDD.n1092 VDD.n1091 8.855
R1031 VDD.n1091 VDD.n1090 8.855
R1032 VDD.n1088 VDD.n1085 8.855
R1033 VDD.n1085 VDD.n1084 8.855
R1034 VDD.n1082 VDD.n1081 8.855
R1035 VDD.n1081 VDD.n1080 8.855
R1036 VDD.n1078 VDD.n1077 8.855
R1037 VDD.n1077 VDD.n1076 8.855
R1038 VDD.n1074 VDD.n1073 8.855
R1039 VDD.n1073 VDD.n1072 8.855
R1040 VDD.n1068 VDD.n1067 8.855
R1041 VDD.n1067 VDD.n1066 8.855
R1042 VDD.n1064 VDD.n1063 8.855
R1043 VDD.n1063 VDD.n1062 8.855
R1044 VDD.n1059 VDD.n1058 8.855
R1045 VDD.n1058 VDD.n1057 8.855
R1046 VDD.n1055 VDD.n1054 8.855
R1047 VDD.n1054 VDD.n1053 8.855
R1048 VDD.n1029 VDD.n1028 8.855
R1049 VDD.n1028 VDD.n1027 8.855
R1050 VDD.n1025 VDD.n1024 8.855
R1051 VDD.n1024 VDD.n1023 8.855
R1052 VDD.n1020 VDD.n1019 8.855
R1053 VDD.n1019 VDD.n1018 8.855
R1054 VDD.n1016 VDD.n1015 8.855
R1055 VDD.n1015  8.855
R1056 VDD.n1011 VDD.n1010 8.855
R1057 VDD.n1010 VDD.n1009 8.855
R1058 VDD.n1007 VDD.n1006 8.855
R1059 VDD.n1006 VDD.n1005 8.855
R1060 VDD.n1003 VDD.n1002 8.855
R1061 VDD.n1002 VDD.n1001 8.855
R1062 VDD.n998 VDD.n997 8.855
R1063 VDD.n997 VDD.n996 8.855
R1064 VDD.n972 VDD.n971 8.855
R1065 VDD.n971 VDD.n970 8.855
R1066 VDD.n968 VDD.n967 8.855
R1067 VDD.n967 VDD.n966 8.855
R1068 VDD.n963 VDD.n962 8.855
R1069 VDD.n962 VDD.n961 8.855
R1070 VDD.n959 VDD.n958 8.855
R1071 VDD.n958 0���0 8.855
R1072 VDD.n954 VDD.n953 8.855
R1073 VDD.n953 VDD.n952 8.855
R1074 VDD.n950 VDD.n949 8.855
R1075 VDD.n949 VDD.n948 8.855
R1076 VDD.n946 VDD.n945 8.855
R1077 VDD.n945 VDD.n944 8.855
R1078 VDD.n941 VDD.n940 8.855
R1079 VDD.n940 VDD.n939 8.855
R1080 VDD.n915 VDD.n914 8.855
R1081 VDD.n914 VDD.n913 8.855
R1082 VDD.n911 VDD.n910 8.855
R1083 VDD.n910 VDD.n909 8.855
R1084 VDD.n907 VDD.n906 8.855
R1085 VDD.n906 VDD.n905 8.855
R1086 VDD.n903 VDD.n902 8.855
R1087 VDD.n902 VDD.n901 8.855
R1088 VDD.n899 VDD.n896 8.855
R1089 VDD.n896 VDD.n895 8.855
R1090 VDD.n893 VDD.n892 8.855
R1091 VDD.n892 VDD.n891 8.855
R1092 VDD.n889 VDD.n888 8.855
R1093 VDD.n888 VDD.n887 8.855
R1094 VDD.n885 VDD.n884 8.855
R1095 VDD.n884 VDD.n883 8.855
R1096 VDD.n879 VDD.n878 8.855
R1097 VDD.n878 VDD.n877 8.855
R1098 VDD.n875 VDD.n874 8.855
R1099 VDD.n874 VDD.n873 8.855
R1100 VDD.n870 VDD.n869 8.855
R1101 VDD.n869 VDD.n868 8.855
R1102 VDD.n866 VDD.n865 8.855
R1103 VDD.n865 VDD.n864 8.855
R1104 VDD.n840 VDD.n839 8.855
R1105 VDD.n839 VDD.n838 8.855
R1106 VDD.n836 VDD.n835 8.855
R1107 VDD.n835 VDD.n834 8.855
R1108 VDD.n832 VDD.n831 8.855
R1109 VDD.n831 VDD.n830 8.855
R1110 VDD.n828 VDD.n827 8.855
R1111 VDD.n827 VDD.n826 8.855
R1112 VDD.n824 VDD.n821 8.855
R1113 VDD.n821 VDD.n820 8.855
R1114 VDD.n818 VDD.n817 8.855
R1115 VDD.n817 VDD.n816 8.855
R1116 VDD.n814 VDD.n813 8.855
R1117 VDD.n813 VDD.n812 8.855
R1118 VDD.n810 VDD.n809 8.855
R1119 VDD.n809 VDD.n808 8.855
R1120 VDD.n804 VDD.n803 8.855
R1121 VDD.n803 VDD.n802 8.855
R1122 VDD.n800 VDD.n799 8.855
R1123 VDD.n799 VDD.n798 8.855
R1124 VDD.n795 VDD.n794 8.855
R1125 VDD.n794 VDD.n793 8.855
R1126 VDD.n791 VDD.n790 8.855
R1127 VDD.n790 VDD.n789 8.855
R1128 VDD.n764 VDD.n763 8.855
R1129 VDD.n763 VDD.n762 8.855
R1130 VDD.n760 VDD.n759 8.855
R1131 VDD.n759 VDD.n758 8.855
R1132 VDD.n755 VDD.n754 8.855
R1133 VDD.n754 VDD.n753 8.855
R1134 VDD.n751 VDD.n750 8.855
R1135 VDD.n750  8.855
R1136 VDD.n746 VDD.n745 8.855
R1137 VDD.n745 VDD.n744 8.855
R1138 VDD.n742 VDD.n741 8.855
R1139 VDD.n741 VDD.n740 8.855
R1140 VDD.n738 VDD.n737 8.855
R1141 VDD.n737 VDD.n736 8.855
R1142 VDD.n733 VDD.n732 8.855
R1143 VDD.n732 VDD.n731 8.855
R1144 VDD.n857 VDD.n856 8.051
R1145 VDD.n932 VDD.n931 8.051
R1146 VDD.n989 VDD.n988 8.051
R1147 VDD.n1046 VDD.n1045 8.051
R1148 VDD.n1121 VDD.n1120 8.051
R1149 VDD.n1178 VDD.n1177 8.051
R1150 VDD.n1253 VDD.n1252 8.051
R1151 VDD.n1328 VDD.n1327 8.051
R1152 VDD.n1385 VDD.n1384 8.051
R1153 VDD.n692 VDD.n691 8.051
R1154 VDD.n617 VDD.n616 8.051
R1155 VDD.n560 VDD.n559 8.051
R1156 VDD.n485 VDD.n484 8.051
R1157 VDD.n410 VDD.n409 8.051
R1158 VDD.n353 VDD.n352 8.051
R1159 VDD.n296 VDD.n295 8.051
R1160 VDD.n221 VDD.n220 8.051
R1161 VDD.n164 VDD.n163 8.051
R1162 VDD.n111 VDD.n110 8.051
R1163 VDD.n54 VDD.n53 8.051
R1164 VDD.n778 VDD.n777 8.051
R1165 VDD.n254 0���0 7.671
R1166 VDD.n443 0���0 7.671
R1167 VDD.n518  7.671
R1168 VDD.n650 0���0 7.671
R1169 VDD.n1283 0���0 7.671
R1170 VDD.n1208 VDD.t84 7.671
R1171 VDD.n1076  7.671
R1172 VDD.n887  7.671
R1173 VDD.n812  7.671
R1174 VDD.n262 VDD.n259 7.019
R1175 VDD.n451 VDD.n448 7.019
R1176 VDD.n526 VDD.n523 7.019
R1177 VDD.n658 VDD.n655 7.019
R1178 VDD.n1281 VDD.n1278 7.019
R1179 VDD.n1206 VDD.n1203 7.019
R1180 VDD.n1074 VDD.n1071 7.019
R1181 VDD.n885 VDD.n882 7.019
R1182 VDD.n810 VDD.n807 7.019
R1183 VDD.n248 VDD.n247 6.606
R1184 VDD.n437 VDD.n436 6.606
R1185 VDD.n512 VDD.n511 6.606
R1186 VDD.n644 VDD.n643 6.606
R1187 VDD.n1295 VDD.n1294 6.606
R1188 VDD.n1220 VDD.n1219 6.606
R1189 VDD.n1088 VDD.n1087 6.606
R1190 VDD.n899 VDD.n898 6.606
R1191 VDD.n824 VDD.n823 6.606
R1192 VDD.n250  5.114
R1193 VDD.n439  5.114
R1194 VDD.n514  5.114
R1195 VDD.n646 0���0 5.114
R1196 VDD.n1287  5.114
R1197 VDD.n1212  5.114
R1198 VDD.n1080 0���0 5.114
R1199 VDD.n891  5.114
R1200 VDD.n816  5.114
R1201 VDD.n28 VDD.n23 4.795
R1202 VDD.n28 VDD.n27 4.65
R1203 VDD.n32 VDD.n31 4.65
R1204 VDD.n37 VDD.n36 4.65
R1205 VDD.n41 VDD.n40 4.65
R1206 VDD.n68 VDD.n67 4.65
R1207 VDD.n72 VDD.n71 4.65
R1208 VDD.n76 VDD.n75 4.65
R1209 VDD.n79 VDD.n78 4.65
R1210 VDD.n83 VDD.n82 4.65
R1211 VDD.n87 VDD.n86 4.65
R1212 VDD.n91 VDD.n90 4.65
R1213 VDD.n95 VDD.n94 4.65
R1214 VDD.n121 VDD.n120 4.65
R1215 VDD.n125 VDD.n124 4.65
R1216 VDD.n129 VDD.n128 4.65
R1217 VDD.n133 VDD.n132 4.65
R1218 VDD.n136 VDD.n135 4.65
R1219 VDD.n140 VDD.n139 4.65
R1220 VDD.n144 VDD.n143 4.65
R1221 VDD.n148 VDD.n147 4.65
R1222 VDD.n174 VDD.n173 4.65
R1223 VDD.n179 VDD.n178 4.65
R1224 VDD.n183 VDD.n182 4.65
R1225 VDD.n188 VDD.n187 4.65
R1226 VDD.n192 VDD.n191 4.65
R1227 VDD.n196 VDD.n195 4.65
R1228 VDD.n201 VDD.n200 4.65
R1229 VDD.n205 VDD.n204 4.65
R1230 VDD.n231 VDD.n230 4.65
R1231 VDD.n235 VDD.n234 4.65
R1232 VDD.n239 VDD.n238 4.65
R1233 VDD.n243 VDD.n242 4.65
R1234 VDD.n249 VDD.n248 4.65
R1235 VDD.n253 VDD.n252 4.65
R1236 VDD.n257 VDD.n256 4.65
R1237 VDD.n263 VDD.n262 4.65
R1238 VDD.n267 VDD.n266 4.65
R1239 VDD.n272 VDD.n271 4.65
R1240 VDD.n276 VDD.n275 4.65
R1241 VDD.n280 VDD.n279 4.65
R1242 VDD.n306 VDD.n305 4.65
R1243 VDD.n311 VDD.n310 4.65
R1244 VDD.n315 VDD.n314 4.65
R1245 VDD.n320 VDD.n319 4.65
R1246 VDD.n324 VDD.n323 4.65
R1247 VDD.n328 VDD.n327 4.65
R1248 VDD.n333 VDD.n332 4.65
R1249 VDD.n337 VDD.n336 4.65
R1250 VDD.n363 VDD.n362 4.65
R1251 VDD.n368 VDD.n367 4.65
R1252 VDD.n372 VDD.n371 4.65
R1253 VDD.n377 VDD.n376 4.65
R1254 VDD.n381 VDD.n380 4.65
R1255 VDD.n385 VDD.n384 4.65
R1256 VDD.n390 VDD.n389 4.65
R1257 VDD.n394 VDD.n393 4.65
R1258 VDD.n420 VDD.n419 4.65
R1259 VDD.n424 VDD.n423 4.65
R1260 VDD.n428 VDD.n427 4.65
R1261 VDD.n432 VDD.n431 4.65
R1262 VDD.n438 VDD.n437 4.65
R1263 VDD.n442 VDD.n441 4.65
R1264 VDD.n446 VDD.n445 4.65
R1265 VDD.n452 VDD.n451 4.65
R1266 VDD.n456 VDD.n455 4.65
R1267 VDD.n461 VDD.n460 4.65
R1268 VDD.n465 VDD.n464 4.65
R1269 VDD.n469 VDD.n468 4.65
R1270 VDD.n495 VDD.n494 4.65
R1271 VDD.n499 VDD.n498 4.65
R1272 VDD.n503 VDD.n502 4.65
R1273 VDD.n507 VDD.n506 4.65
R1274 VDD.n513 VDD.n512 4.65
R1275 VDD.n517 VDD.n516 4.65
R1276 VDD.n521 VDD.n520 4.65
R1277 VDD.n527 VDD.n526 4.65
R1278 VDD.n531 VDD.n530 4.65
R1279 VDD.n536 VDD.n535 4.65
R1280 VDD.n540 VDD.n539 4.65
R1281 VDD.n544 VDD.n543 4.65
R1282 VDD.n570 VDD.n569 4.65
R1283 VDD.n575 VDD.n574 4.65
R1284 VDD.n579 VDD.n578 4.65
R1285 VDD.n584 VDD.n583 4.65
R1286 VDD.n588 VDD.n587 4.65
R1287 VDD.n592 VDD.n591 4.65
R1288 VDD.n597 VDD.n596 4.65
R1289 VDD.n601 VDD.n600 4.65
R1290 VDD.n627 VDD.n626 4.65
R1291 VDD.n631 VDD.n630 4.65
R1292 VDD.n635 VDD.n634 4.65
R1293 VDD.n639 VDD.n638 4.65
R1294 VDD.n645 VDD.n644 4.65
R1295 VDD.n649 VDD.n648 4.65
R1296 VDD.n653 VDD.n652 4.65
R1297 VDD.n659 VDD.n658 4.65
R1298 VDD.n663 VDD.n662 4.65
R1299 VDD.n668 VDD.n667 4.65
R1300 VDD.n672 VDD.n671 4.65
R1301 VDD.n676 VDD.n675 4.65
R1302 VDD.n702 VDD.n701 4.65
R1303 VDD.n707 VDD.n706 4.65
R1304 VDD.n711 VDD.n710 4.65
R1305 VDD.n1413 VDD.n1412 4.65
R1306 VDD.n1408 VDD.n1407 4.65
R1307 VDD.n1404 VDD.n1403 4.65
R1308 VDD.n1400 VDD.n1399 4.65
R1309 VDD.n1395 VDD.n1394 4.65
R1310 VDD.n1369 VDD.n1368 4.65
R1311 VDD.n1365 VDD.n1364 4.65
R1312 VDD.n1360 VDD.n1359 4.65
R1313 VDD.n1356 VDD.n1355 4.65
R1314 VDD.n1351 VDD.n1350 4.65
R1315 VDD.n1347 VDD.n1346 4.65
R1316 VDD.n1343 VDD.n1342 4.65
R1317 VDD.n1338 VDD.n1337 4.65
R1318 VDD.n1312 VDD.n1311 4.65
R1319 VDD.n1308 VDD.n1307 4.65
R1320 VDD.n1304 VDD.n1303 4.65
R1321 VDD.n1300 VDD.n1299 4.65
R1322 VDD.n1296 VDD.n1295 4.65
R1323 VDD.n1290 VDD.n1289 4.65
R1324 VDD.n1286 VDD.n1285 4.65
R1325 VDD.n1282 VDD.n1281 4.65
R1326 VDD.n1276 VDD.n1275 4.65
R1327 VDD.n1272 VDD.n1271 4.65
R1328 VDD.n1267 VDD.n1266 4.65
R1329 VDD.n1263 VDD.n1262 4.65
R1330 VDD.n1237 VDD.n1236 4.65
R1331 VDD.n1233 VDD.n1232 4.65
R1332 VDD.n1229 VDD.n1228 4.65
R1333 VDD.n1225 VDD.n1224 4.65
R1334 VDD.n1221 VDD.n1220 4.65
R1335 VDD.n1215 VDD.n1214 4.65
R1336 VDD.n1211 VDD.n1210 4.65
R1337 VDD.n1207 VDD.n1206 4.65
R1338 VDD.n1201 VDD.n1200 4.65
R1339 VDD.n1197 VDD.n1196 4.65
R1340 VDD.n1192 VDD.n1191 4.65
R1341 VDD.n1188 VDD.n1187 4.65
R1342 VDD.n1162 VDD.n1161 4.65
R1343 VDD.n1158 VDD.n1157 4.65
R1344 VDD.n1153 VDD.n1152 4.65
R1345 VDD.n1149 VDD.n1148 4.65
R1346 VDD.n1144 VDD.n1143 4.65
R1347 VDD.n1140 VDD.n1139 4.65
R1348 VDD.n1136 VDD.n1135 4.65
R1349 VDD.n1131 VDD.n1130 4.65
R1350 VDD.n1105 VDD.n1104 4.65
R1351 VDD.n1101 VDD.n1100 4.65
R1352 VDD.n1097 VDD.n1096 4.65
R1353 VDD.n1093 VDD.n1092 4.65
R1354 VDD.n1089 VDD.n1088 4.65
R1355 VDD.n1083 VDD.n1082 4.65
R1356 VDD.n1079 VDD.n1078 4.65
R1357 VDD.n1075 VDD.n1074 4.65
R1358 VDD.n1069 VDD.n1068 4.65
R1359 VDD.n1065 VDD.n1064 4.65
R1360 VDD.n1060 VDD.n1059 4.65
R1361 VDD.n1056 VDD.n1055 4.65
R1362 VDD.n1030 VDD.n1029 4.65
R1363 VDD.n1026 VDD.n1025 4.65
R1364 VDD.n1021 VDD.n1020 4.65
R1365 VDD.n1017 VDD.n1016 4.65
R1366 VDD.n1012 VDD.n1011 4.65
R1367 VDD.n1008 VDD.n1007 4.65
R1368 VDD.n1004 VDD.n1003 4.65
R1369 VDD.n999 VDD.n998 4.65
R1370 VDD.n973 VDD.n972 4.65
R1371 VDD.n969 VDD.n968 4.65
R1372 VDD.n964 VDD.n963 4.65
R1373 VDD.n960 VDD.n959 4.65
R1374 VDD.n955 VDD.n954 4.65
R1375 VDD.n951 VDD.n950 4.65
R1376 VDD.n947 VDD.n946 4.65
R1377 VDD.n942 VDD.n941 4.65
R1378 VDD.n916 VDD.n915 4.65
R1379 VDD.n912 VDD.n911 4.65
R1380 VDD.n908 VDD.n907 4.65
R1381 VDD.n904 VDD.n903 4.65
R1382 VDD.n900 VDD.n899 4.65
R1383 VDD.n894 VDD.n893 4.65
R1384 VDD.n890 VDD.n889 4.65
R1385 VDD.n886 VDD.n885 4.65
R1386 VDD.n880 VDD.n879 4.65
R1387 VDD.n876 VDD.n875 4.65
R1388 VDD.n871 VDD.n870 4.65
R1389 VDD.n867 VDD.n866 4.65
R1390 VDD.n841 VDD.n840 4.65
R1391 VDD.n837 VDD.n836 4.65
R1392 VDD.n833 VDD.n832 4.65
R1393 VDD.n829 VDD.n828 4.65
R1394 VDD.n825 VDD.n824 4.65
R1395 VDD.n819 VDD.n818 4.65
R1396 VDD.n815 VDD.n814 4.65
R1397 VDD.n811 VDD.n810 4.65
R1398 VDD.n805 VDD.n804 4.65
R1399 VDD.n801 VDD.n800 4.65
R1400 VDD.n796 VDD.n795 4.65
R1401 VDD.n792 VDD.n791 4.65
R1402 VDD.n765 VDD.n764 4.65
R1403 VDD.n761 VDD.n760 4.65
R1404 VDD.n756 VDD.n755 4.65
R1405 VDD.n752 VDD.n751 4.65
R1406 VDD.n747 VDD.n746 4.65
R1407 VDD.n743 VDD.n742 4.65
R1408 VDD.n739 VDD.n738 4.65
R1409 VDD.n734 VDD.n733 4.65
R1410 VDD.n200 VDD.n197 2.89
R1411 VDD.n332 VDD.n329 2.89
R1412 VDD.n389 VDD.n386 2.89
R1413 VDD.n596 VDD.n593 2.89
R1414 VDD.n1399 VDD.n1396 2.89
R1415 VDD.n1342 VDD.n1339 2.89
R1416 VDD.n1135 VDD.n1132 2.89
R1417 VDD.n1003 VDD.n1000 2.89
R1418 VDD.n946 VDD.n943 2.89
R1419 VDD.n738 VDD.n735 2.89
R1420 VDD.n80 0���0 2.557
R1421 VDD.n130  2.557
R1422 VDD.n189  2.557
R1423 VDD.n321 0���0 2.557
R1424 VDD.n378  2.557
R1425 VDD.n585  2.557
R1426 VDD.n1405 0���0 2.557
R1427 VDD.n1348 0���0 2.557
R1428 VDD.n1141 @b4	�U 2.557
R1429 VDD.n1009 0���0 2.557
R1430 VDD.n952  2.557
R1431 VDD.n744  2.557
R1432 VDD.n178 VDD.n175 2.477
R1433 VDD.n310 VDD.n307 2.477
R1434 VDD.n367 VDD.n364 2.477
R1435 VDD.n574 VDD.n571 2.477
R1436 VDD.n706 VDD.n703 2.477
R1437 VDD.n1364 VDD.n1361 2.477
R1438 VDD.n1157 VDD.n1154 2.477
R1439 VDD.n1025 VDD.n1022 2.477
R1440 VDD.n968 VDD.n965 2.477
R1441 VDD.n760 VDD.n757 2.477
R1442 VDD.n27 VDD.n24 2.064
R1443 VDD.n36 VDD.n35 2.064
R1444 VDD.n271 VDD.n268 0.412
R1445 VDD.n460 VDD.n457 0.412
R1446 VDD.n535 VDD.n532 0.412
R1447 VDD.n667 VDD.n664 0.412
R1448 VDD.n1271 VDD.n1268 0.412
R1449 VDD.n1196 VDD.n1193 0.412
R1450 VDD.n1064 VDD.n1061 0.412
R1451 VDD.n875 VDD.n872 0.412
R1452 VDD.n800 VDD.n797 0.412
R1453 VDD.n68 VDD.n41 0.29
R1454 VDD.n121 VDD.n95 0.29
R1455 VDD.n174 VDD.n148 0.29
R1456 VDD.n231 VDD.n205 0.29
R1457 VDD.n306 VDD.n280 0.29
R1458 VDD.n363 VDD.n337 0.29
R1459 VDD.n420 VDD.n394 0.29
R1460 VDD.n495 VDD.n469 0.29
R1461 VDD.n570 VDD.n544 0.29
R1462 VDD.n627 VDD.n601 0.29
R1463 VDD.n702 VDD.n676 0.29
R1464 VDD.n1395 VDD.n1369 0.29
R1465 VDD.n1338 VDD.n1312 0.29
R1466 VDD.n1263 VDD.n1237 0.29
R1467 VDD.n1188 VDD.n1162 0.29
R1468 VDD.n1131 VDD.n1105 0.29
R1469 VDD.n1056 VDD.n1030 0.29
R1470 VDD.n999 VDD.n973 0.29
R1471 VDD.n942 VDD.n916 0.29
R1472 VDD.n867 VDD.n841 0.29
R1473 VDD.n792 VDD.n765 0.29
R1474 VDD.n734 VDD 0.207
R1475 VDD.n257 VDD.n253 0.197
R1476 VDD.n446 VDD.n442 0.197
R1477 VDD.n521 VDD.n517 0.197
R1478 VDD.n653 VDD.n649 0.197
R1479 VDD.n1290 VDD.n1286 0.197
R1480 VDD.n1215 VDD.n1211 0.197
R1481 VDD.n1083 VDD.n1079 0.197
R1482 VDD.n894 VDD.n890 0.197
R1483 VDD.n819 VDD.n815 0.197
R1484 VDD.n83 VDD.n79 0.181
R1485 VDD.n136 VDD.n133 0.181
R1486 VDD.n192 VDD.n188 0.181
R1487 VDD.n324 VDD.n320 0.181
R1488 VDD.n381 VDD.n377 0.181
R1489 VDD.n588 VDD.n584 0.181
R1490 VDD.n1413 VDD.n1408 0.181
R1491 VDD.n1356 VDD.n1351 0.181
R1492 VDD.n1149 VDD.n1144 0.181
R1493 VDD.n1017 VDD.n1012 0.181
R1494 VDD.n960 VDD.n955 0.181
R1495 VDD.n752 VDD.n747 0.181
R1496 VDD.n32 VDD.n28 0.157
R1497 VDD.n37 VDD.n32 0.157
R1498 VDD.n41 VDD.n37 0.145
R1499 VDD.n72 VDD.n68 0.145
R1500 VDD.n76 VDD.n72 0.145
R1501 VDD.n79 VDD.n76 0.145
R1502 VDD.n87 VDD.n83 0.145
R1503 VDD.n91 VDD.n87 0.145
R1504 VDD.n95 VDD.n91 0.145
R1505 VDD.n125 VDD.n121 0.145
R1506 VDD.n129 VDD.n125 0.145
R1507 VDD.n133 VDD.n129 0.145
R1508 VDD.n140 VDD.n136 0.145
R1509 VDD.n144 VDD.n140 0.145
R1510 VDD.n148 VDD.n144 0.145
R1511 VDD.n179 VDD.n174 0.145
R1512 VDD.n183 VDD.n179 0.145
R1513 VDD.n188 VDD.n183 0.145
R1514 VDD.n196 VDD.n192 0.145
R1515 VDD.n201 VDD.n196 0.145
R1516 VDD.n205 VDD.n201 0.145
R1517 VDD.n235 VDD.n231 0.145
R1518 VDD.n239 VDD.n235 0.145
R1519 VDD.n243 VDD.n239 0.145
R1520 VDD.n249 VDD.n243 0.145
R1521 VDD.n253 VDD.n249 0.145
R1522 VDD.n263 VDD.n257 0.145
R1523 VDD.n267 VDD.n263 0.145
R1524 VDD.n272 VDD.n267 0.145
R1525 VDD.n276 VDD.n272 0.145
R1526 VDD.n280 VDD.n276 0.145
R1527 VDD.n311 VDD.n306 0.145
R1528 VDD.n315 VDD.n311 0.145
R1529 VDD.n320 VDD.n315 0.145
R1530 VDD.n328 VDD.n324 0.145
R1531 VDD.n333 VDD.n328 0.145
R1532 VDD.n337 VDD.n333 0.145
R1533 VDD.n368 VDD.n363 0.145
R1534 VDD.n372 VDD.n368 0.145
R1535 VDD.n377 VDD.n372 0.145
R1536 VDD.n385 VDD.n381 0.145
R1537 VDD.n390 VDD.n385 0.145
R1538 VDD.n394 VDD.n390 0.145
R1539 VDD.n424 VDD.n420 0.145
R1540 VDD.n428 VDD.n424 0.145
R1541 VDD.n432 VDD.n428 0.145
R1542 VDD.n438 VDD.n432 0.145
R1543 VDD.n442 VDD.n438 0.145
R1544 VDD.n452 VDD.n446 0.145
R1545 VDD.n456 VDD.n452 0.145
R1546 VDD.n461 VDD.n456 0.145
R1547 VDD.n465 VDD.n461 0.145
R1548 VDD.n469 VDD.n465 0.145
R1549 VDD.n499 VDD.n495 0.145
R1550 VDD.n503 VDD.n499 0.145
R1551 VDD.n507 VDD.n503 0.145
R1552 VDD.n513 VDD.n507 0.145
R1553 VDD.n517 VDD.n513 0.145
R1554 VDD.n527 VDD.n521 0.145
R1555 VDD.n531 VDD.n527 0.145
R1556 VDD.n536 VDD.n531 0.145
R1557 VDD.n540 VDD.n536 0.145
R1558 VDD.n544 VDD.n540 0.145
R1559 VDD.n575 VDD.n570 0.145
R1560 VDD.n579 VDD.n575 0.145
R1561 VDD.n584 VDD.n579 0.145
R1562 VDD.n592 VDD.n588 0.145
R1563 VDD.n597 VDD.n592 0.145
R1564 VDD.n601 VDD.n597 0.145
R1565 VDD.n631 VDD.n627 0.145
R1566 VDD.n635 VDD.n631 0.145
R1567 VDD.n639 VDD.n635 0.145
R1568 VDD.n645 VDD.n639 0.145
R1569 VDD.n649 VDD.n645 0.145
R1570 VDD.n659 VDD.n653 0.145
R1571 VDD.n663 VDD.n659 0.145
R1572 VDD.n668 VDD.n663 0.145
R1573 VDD.n672 VDD.n668 0.145
R1574 VDD.n676 VDD.n672 0.145
R1575 VDD.n707 VDD.n702 0.145
R1576 VDD.n711 VDD.n707 0.145
R1577 VDD.n1408 VDD.n1404 0.145
R1578 VDD.n1404 VDD.n1400 0.145
R1579 VDD.n1400 VDD.n1395 0.145
R1580 VDD.n1369 VDD.n1365 0.145
R1581 VDD.n1365 VDD.n1360 0.145
R1582 VDD.n1360 VDD.n1356 0.145
R1583 VDD.n1351 VDD.n1347 0.145
R1584 VDD.n1347 VDD.n1343 0.145
R1585 VDD.n1343 VDD.n1338 0.145
R1586 VDD.n1312 VDD.n1308 0.145
R1587 VDD.n1308 VDD.n1304 0.145
R1588 VDD.n1304 VDD.n1300 0.145
R1589 VDD.n1300 VDD.n1296 0.145
R1590 VDD.n1296 VDD.n1290 0.145
R1591 VDD.n1286 VDD.n1282 0.145
R1592 VDD.n1282 VDD.n1276 0.145
R1593 VDD.n1276 VDD.n1272 0.145
R1594 VDD.n1272 VDD.n1267 0.145
R1595 VDD.n1267 VDD.n1263 0.145
R1596 VDD.n1237 VDD.n1233 0.145
R1597 VDD.n1233 VDD.n1229 0.145
R1598 VDD.n1229 VDD.n1225 0.145
R1599 VDD.n1225 VDD.n1221 0.145
R1600 VDD.n1221 VDD.n1215 0.145
R1601 VDD.n1211 VDD.n1207 0.145
R1602 VDD.n1207 VDD.n1201 0.145
R1603 VDD.n1201 VDD.n1197 0.145
R1604 VDD.n1197 VDD.n1192 0.145
R1605 VDD.n1192 VDD.n1188 0.145
R1606 VDD.n1162 VDD.n1158 0.145
R1607 VDD.n1158 VDD.n1153 0.145
R1608 VDD.n1153 VDD.n1149 0.145
R1609 VDD.n1144 VDD.n1140 0.145
R1610 VDD.n1140 VDD.n1136 0.145
R1611 VDD.n1136 VDD.n1131 0.145
R1612 VDD.n1105 VDD.n1101 0.145
R1613 VDD.n1101 VDD.n1097 0.145
R1614 VDD.n1097 VDD.n1093 0.145
R1615 VDD.n1093 VDD.n1089 0.145
R1616 VDD.n1089 VDD.n1083 0.145
R1617 VDD.n1079 VDD.n1075 0.145
R1618 VDD.n1075 VDD.n1069 0.145
R1619 VDD.n1069 VDD.n1065 0.145
R1620 VDD.n1065 VDD.n1060 0.145
R1621 VDD.n1060 VDD.n1056 0.145
R1622 VDD.n1030 VDD.n1026 0.145
R1623 VDD.n1026 VDD.n1021 0.145
R1624 VDD.n1021 VDD.n1017 0.145
R1625 VDD.n1012 VDD.n1008 0.145
R1626 VDD.n1008 VDD.n1004 0.145
R1627 VDD.n1004 VDD.n999 0.145
R1628 VDD.n973 VDD.n969 0.145
R1629 VDD.n969 VDD.n964 0.145
R1630 VDD.n964 VDD.n960 0.145
R1631 VDD.n955 VDD.n951 0.145
R1632 VDD.n951 VDD.n947 0.145
R1633 VDD.n947 VDD.n942 0.145
R1634 VDD.n916 VDD.n912 0.145
R1635 VDD.n912 VDD.n908 0.145
R1636 VDD.n908 VDD.n904 0.145
R1637 VDD.n904 VDD.n900 0.145
R1638 VDD.n900 VDD.n894 0.145
R1639 VDD.n890 VDD.n886 0.145
R1640 VDD.n886 VDD.n880 0.145
R1641 VDD.n880 VDD.n876 0.145
R1642 VDD.n876 VDD.n871 0.145
R1643 VDD.n871 VDD.n867 0.145
R1644 VDD.n841 VDD.n837 0.145
R1645 VDD.n837 VDD.n833 0.145
R1646 VDD.n833 VDD.n829 0.145
R1647 VDD.n829 VDD.n825 0.145
R1648 VDD.n825 VDD.n819 0.145
R1649 VDD.n815 VDD.n811 0.145
R1650 VDD.n811 VDD.n805 0.145
R1651 VDD.n805 VDD.n801 0.145
R1652 VDD.n801 VDD.n796 0.145
R1653 VDD.n796 VDD.n792 0.145
R1654 VDD.n765 VDD.n761 0.145
R1655 VDD.n761 VDD.n756 0.145
R1656 VDD.n756 VDD.n752 0.145
R1657 VDD.n747 VDD.n743 0.145
R1658 VDD.n743 VDD.n739 0.145
R1659 VDD.n739 VDD.n734 0.145
R1660 VDD VDD.n711 0.086
R1661 VDD VDD.n1413 0.058
R1662 a_6789_1050.n5 a_6789_1050.t9 480.392
R1663 a_6789_1050.n5 a_6789_1050.t8 403.272
R1664 a_6789_1050.n6 a_6789_1050.t7 301.486
R1665 a_6789_1050.n9 a_6789_1050.n7 259.02
R1666 a_6789_1050.n7 a_6789_1050.n4 234.917
R1667 a_6789_1050.n6 a_6789_1050.n5 227.006
R1668 a_6789_1050.n3 a_6789_1050.n2 161.352
R1669 a_6789_1050.n4 a_6789_1050.n0 95.095
R1670 a_6789_1050.n3 a_6789_1050.n1 95.095
R1671 a_6789_1050.n4 a_6789_1050.n3 66.258
R1672 a_6789_1050.n9 a_6789_1050.n8 15.218
R1673 a_6789_1050.n0 a_6789_1050.t2 14.282
R1674 a_6789_1050.n0 a_6789_1050.t1 14.282
R1675 a_6789_1050.n1 a_6789_1050.t6 14.282
R1676 a_6789_1050.n1 a_6789_1050.t5 14.282
R1677 a_6789_1050.n2 a_6789_1050.t0 14.282
R1678 a_6789_1050.n2 a_6789_1050.t4 14.282
R1679 a_6789_1050.n10 a_6789_1050.n9 12.014
R1680 a_6789_1050.n7 a_6789_1050.n6 10.615
R1681 a_7586_101.t0 a_7586_101.n1 93.333
R1682 a_7586_101.n4 a_7586_101.n2 79.092
R1683 a_7586_101.t0 a_7586_101.n0 8.137
R1684 a_7586_101.n4 a_7586_101.n3 4.614
R1685 a_7586_101.t0 a_7586_101.n4 0.111
R1686 GND.n32 GND.n31 237.558
R1687 GND.n64 GND.n63 237.558
R1688 GND.n431 GND.n430 237.558
R1689 GND.n475 GND.n474 237.558
R1690 GND.n519 GND.n518 237.558
R1691 GND.n549 GND.n548 237.558
R1692 GND.n579 GND.n578 237.558
R1693 GND.n624 GND.n623 237.558
R1694 GND.n656 GND.n655 237.558
R1695 GND.n700 GND.n699 237.558
R1696 GND.n744 GND.n743 237.558
R1697 GND.n393 GND.n392 237.558
R1698 GND.n776 GND.n775 237.558
R1699 GND.n348 GND.n347 237.558
R1700 GND.n318 GND.n317 237.558
R1701 GND.n276 GND.n275 237.558
R1702 GND.n232 GND.n231 237.558
R1703 GND.n202 GND.n201 237.558
R1704 GND.n172 GND.n171 237.558
R1705 GND.n130 GND.n129 237.558
R1706 GND.n97 GND.n96 237.558
R1707 GND.n29 GND.n28 210.82
R1708 GND.n61 GND.n60 210.82
R1709 GND.n94 GND.n93 210.82
R1710 GND.n433 GND.n432 210.82
R1711 GND.n477 GND.n476 210.82
R1712 GND.n521 GND.n520 210.82
R1713 GND.n551 GND.n550 210.82
R1714 GND.n581 GND.n580 210.82
R1715 GND.n626 GND.n625 210.82
R1716 GND.n658 GND.n657 210.82
R1717 GND.n702 GND.n701 210.82
R1718 GND.n746 GND.n745 210.82
R1719 GND.n778 GND.n777 210.82
R1720 GND.n390 GND.n389 210.82
R1721 GND.n345 GND.n344 210.82
R1722 GND.n315 GND.n314 210.82
R1723 GND.n273 GND.n272 210.82
R1724 GND.n229 GND.n228 210.82
R1725 GND.n199 GND.n198 210.82
R1726 GND.n169 GND.n168 210.82
R1727 GND.n127 GND.n126 210.82
R1728 GND.n159 GND.n158 173.365
R1729 GND.n305 GND.n304 173.365
R1730 GND.n188 GND.n187 172.612
R1731 GND.n218 GND.n217 172.612
R1732 GND.n334 GND.n333 172.612
R1733 GND.n786 GND.n785 172.612
R1734 GND.n559 GND.n558 172.612
R1735 GND.n529 GND.n528 172.612
R1736 GND.n263 GND.n262 167.358
R1737 GND.n713 GND.n712 167.358
R1738 GND.n669 GND.n668 167.358
R1739 GND.n488 GND.n487 167.358
R1740 GND.n444 GND.n443 167.358
R1741 GND.n756 GND.n755 166.605
R1742 GND.n636 GND.n635 166.605
R1743 GND.n411 GND.n410 166.605
R1744 GND.n50 GND.n49 166.605
R1745 GND.n380 GND.n379 152.358
R1746 GND.n593 GND.n592 152.358
R1747 GND.n83 GND.n82 151.605
R1748 GND.n116 GND.n115 151.605
R1749 GND.n20 GND.n19 37.582
R1750 GND.t28 GND.n17 32.601
R1751 GND.n82 GND.n81 28.421
R1752 GND.n115 GND.n114 28.421
R1753 GND.n379 GND.n378 28.421
R1754 GND.n592 GND.n591 28.421
R1755 GND.n82 GND.n80 25.263
R1756 GND.n115 GND.n113 25.263
R1757 GND.n379 GND.n377 25.263
R1758 GND.n592 GND.n590 25.263
R1759 GND.n80 GND.n79 24.383
R1760 GND.n113 GND.n112 24.383
R1761 GND.n377 GND.n376 24.383
R1762 GND.n590 GND.n589 24.383
R1763 GND.n262 GND.n260 23.03
R1764 GND.n755 GND.n753 23.03
R1765 GND.n712 GND.n710 23.03
R1766 GND.n668 GND.n666 23.03
R1767 GND.n635 GND.n633 23.03
R1768 GND.n487 GND.n485 23.03
R1769 GND.n443 GND.n441 23.03
R1770 GND.n410 GND.n408 23.03
R1771 GND.n49 GND.n47 23.03
R1772 GND.n17 GND.n16 21.734
R1773 GND.n4 GND.n3 20.705
R1774 GND.n10 GND.n9 20.705
R1775 GND.n21 GND.n20 20.705
R1776 GND.n3 GND.n2 19.952
R1777 GND.n30 GND.n29 18.953
R1778 GND.n62 GND.n61 18.953
R1779 GND.n95 GND.n94 18.953
R1780 GND.n434 GND.n433 18.953
R1781 GND.n478 GND.n477 18.953
R1782 GND.n522 GND.n521 18.953
R1783 GND.n552 GND.n551 18.953
R1784 GND.n582 GND.n581 18.953
R1785 GND.n627 GND.n626 18.953
R1786 GND.n659 GND.n658 18.953
R1787 GND.n703 GND.n702 18.953
R1788 GND.n747 GND.n746 18.953
R1789 GND.n779 GND.n778 18.953
R1790 GND.n391 GND.n390 18.953
R1791 GND.n346 GND.n345 18.953
R1792 GND.n316 GND.n315 18.953
R1793 GND.n274 GND.n273 18.953
R1794 GND.n230 GND.n229 18.953
R1795 GND.n200 GND.n199 18.953
R1796 GND.n170 GND.n169 18.953
R1797 GND.n128 GND.n127 18.953
R1798 GND.n19 GND.t28 15.644
R1799 GND.n33 GND.n30 14.864
R1800 GND.n65 GND.n62 14.864
R1801 GND.n98 GND.n95 14.864
R1802 GND.n131 GND.n128 14.864
R1803 GND.n173 GND.n170 14.864
R1804 GND.n203 GND.n200 14.864
R1805 GND.n233 GND.n230 14.864
R1806 GND.n277 GND.n274 14.864
R1807 GND.n319 GND.n316 14.864
R1808 GND.n349 GND.n346 14.864
R1809 GND.n394 GND.n391 14.864
R1810 GND.n780 GND.n779 14.864
R1811 GND.n748 GND.n747 14.864
R1812 GND.n704 GND.n703 14.864
R1813 GND.n660 GND.n659 14.864
R1814 GND.n628 GND.n627 14.864
R1815 GND.n583 GND.n582 14.864
R1816 GND.n553 GND.n552 14.864
R1817 GND.n523 GND.n522 14.864
R1818 GND.n479 GND.n478 14.864
R1819 GND.n435 GND.n434 14.864
R1820 GND.n19 GND.n18 13.541
R1821 GND.n406 GND.n405 9.154
R1822 GND.n413 GND.n412 9.154
R1823 GND.n416 GND.n415 9.154
R1824 GND.n419 GND.n418 9.154
R1825 GND.n422 GND.n421 9.154
R1826 GND.n425 GND.n424 9.154
R1827 GND.n428 GND.n427 9.154
R1828 GND.n435 GND.n431 9.154
R1829 GND.n438 GND.n437 9.154
R1830 GND.n445 GND.n440 9.154
R1831 GND.n448 GND.n447 9.154
R1832 GND.n451 GND.n450 9.154
R1833 GND.n454 GND.n453 9.154
R1834 GND.n457 GND.n456 9.154
R1835 GND.n460 GND.n459 9.154
R1836 GND.n463 GND.n462 9.154
R1837 GND.n466 GND.n465 9.154
R1838 GND.n469 GND.n468 9.154
R1839 GND.n472 GND.n471 9.154
R1840 GND.n479 GND.n475 9.154
R1841 GND.n482 GND.n481 9.154
R1842 GND.n489 GND.n484 9.154
R1843 GND.n492 GND.n491 9.154
R1844 GND.n495 GND.n494 9.154
R1845 GND.n498 GND.n497 9.154
R1846 GND.n501 GND.n500 9.154
R1847 GND.n504 GND.n503 9.154
R1848 GND.n507 GND.n506 9.154
R1849 GND.n510 GND.n509 9.154
R1850 GND.n513 GND.n512 9.154
R1851 GND.n516 GND.n515 9.154
R1852 GND.n523 GND.n519 9.154
R1853 GND.n526 GND.n525 9.154
R1854 GND.n531 GND.n530 9.154
R1855 GND.n534 GND.n533 9.154
R1856 GND.n537 GND.n536 9.154
R1857 GND.n540 GND.n539 9.154
R1858 GND.n543 GND.n542 9.154
R1859 GND.n546 GND.n545 9.154
R1860 GND.n553 GND.n549 9.154
R1861 GND.n556 GND.n555 9.154
R1862 GND.n561 GND.n560 9.154
R1863 GND.n564 GND.n563 9.154
R1864 GND.n567 GND.n566 9.154
R1865 GND.n570 GND.n569 9.154
R1866 GND.n573 GND.n572 9.154
R1867 GND.n576 GND.n575 9.154
R1868 GND.n583 GND.n579 9.154
R1869 GND.n586 GND.n585 9.154
R1870 GND.n594 GND.n588 9.154
R1871 GND.n597 GND.n596 9.154
R1872 GND.n600 GND.n599 9.154
R1873 GND.n603 GND.n602 9.154
R1874 GND.n606 GND.n605 9.154
R1875 GND.n609 GND.n608 9.154
R1876 GND.n612 GND.n611 9.154
R1877 GND.n615 GND.n614 9.154
R1878 GND.n618 GND.n617 9.154
R1879 GND.n621 GND.n620 9.154
R1880 GND.n628 GND.n624 9.154
R1881 GND.n631 GND.n630 9.154
R1882 GND.n638 GND.n637 9.154
R1883 GND.n641 GND.n640 9.154
R1884 GND.n644 GND.n643 9.154
R1885 GND.n647 GND.n646 9.154
R1886 GND.n650 GND.n649 9.154
R1887 GND.n653 GND.n652 9.154
R1888 GND.n660 GND.n656 9.154
R1889 GND.n663 GND.n662 9.154
R1890 GND.n670 GND.n665 9.154
R1891 GND.n673 GND.n672 9.154
R1892 GND.n676 GND.n675 9.154
R1893 GND.n679 GND.n678 9.154
R1894 GND.n682 GND.n681 9.154
R1895 GND.n685 GND.n684 9.154
R1896 GND.n688 GND.n687 9.154
R1897 GND.n691 GND.n690 9.154
R1898 GND.n694 GND.n693 9.154
R1899 GND.n697 GND.n696 9.154
R1900 GND.n704 GND.n700 9.154
R1901 GND.n707 GND.n706 9.154
R1902 GND.n714 GND.n709 9.154
R1903 GND.n717 GND.n716 9.154
R1904 GND.n720 GND.n719 9.154
R1905 GND.n723 GND.n722 9.154
R1906 GND.n726 GND.n725 9.154
R1907 GND.n729 GND.n728 9.154
R1908 GND.n732 GND.n731 9.154
R1909 GND.n735 GND.n734 9.154
R1910 GND.n738 GND.n737 9.154
R1911 GND.n741 GND.n740 9.154
R1912 GND.n748 GND.n744 9.154
R1913 GND.n751 GND.n750 9.154
R1914 GND.n758 GND.n757 9.154
R1915 GND.n761 GND.n760 9.154
R1916 GND.n764 GND.n763 9.154
R1917 GND.n767 GND.n766 9.154
R1918 GND.n770 GND.n769 9.154
R1919 GND.n773 GND.n772 9.154
R1920 GND.n780 GND.n776 9.154
R1921 GND.n783 GND.n782 9.154
R1922 GND.n788 GND.n787 9.154
R1923 GND.n791 GND.n790 9.154
R1924 GND.n794 GND.n793 9.154
R1925 GND.n400 GND.n399 9.154
R1926 GND.n397 GND.n396 9.154
R1927 GND.n394 GND.n393 9.154
R1928 GND.n387 GND.n386 9.154
R1929 GND.n384 GND.n383 9.154
R1930 GND.n381 GND.n375 9.154
R1931 GND.n373 GND.n372 9.154
R1932 GND.n370 GND.n369 9.154
R1933 GND.n367 GND.n366 9.154
R1934 GND.n364 GND.n363 9.154
R1935 GND.n361 GND.n360 9.154
R1936 GND.n358 GND.n357 9.154
R1937 GND.n355 GND.n354 9.154
R1938 GND.n352 GND.n351 9.154
R1939 GND.n349 GND.n348 9.154
R1940 GND.n342 GND.n341 9.154
R1941 GND.n339 GND.n338 9.154
R1942 GND.n336 GND.n335 9.154
R1943 GND.n331 GND.n330 9.154
R1944 GND.n328 GND.n327 9.154
R1945 GND.n325 GND.n324 9.154
R1946 GND.n322 GND.n321 9.154
R1947 GND.n319 GND.n318 9.154
R1948 GND.n312 GND.n311 9.154
R1949 GND.n309 GND.n308 9.154
R1950 GND.n306 GND.n303 9.154
R1951 GND.n301 GND.n300 9.154
R1952 GND.n298 GND.n297 9.154
R1953 GND.n295 GND.n294 9.154
R1954 GND.n292 GND.n291 9.154
R1955 GND.n289 GND.n288 9.154
R1956 GND.n286 GND.n285 9.154
R1957 GND.n283 GND.n282 9.154
R1958 GND.n280 GND.n279 9.154
R1959 GND.n277 GND.n276 9.154
R1960 GND.n270 GND.n269 9.154
R1961 GND.n267 GND.n266 9.154
R1962 GND.n264 GND.n259 9.154
R1963 GND.n257 GND.n256 9.154
R1964 GND.n254 GND.n253 9.154
R1965 GND.n251 GND.n250 9.154
R1966 GND.n248 GND.n247 9.154
R1967 GND.n245 GND.n244 9.154
R1968 GND.n242 GND.n241 9.154
R1969 GND.n239 GND.n238 9.154
R1970 GND.n236 GND.n235 9.154
R1971 GND.n233 GND.n232 9.154
R1972 GND.n226 GND.n225 9.154
R1973 GND.n223 GND.n222 9.154
R1974 GND.n220 GND.n219 9.154
R1975 GND.n215 GND.n214 9.154
R1976 GND.n212 GND.n211 9.154
R1977 GND.n209 GND.n208 9.154
R1978 GND.n206 GND.n205 9.154
R1979 GND.n203 GND.n202 9.154
R1980 GND.n196 GND.n195 9.154
R1981 GND.n193 GND.n192 9.154
R1982 GND.n190 GND.n189 9.154
R1983 GND.n185 GND.n184 9.154
R1984 GND.n182 GND.n181 9.154
R1985 GND.n179 GND.n178 9.154
R1986 GND.n176 GND.n175 9.154
R1987 GND.n173 GND.n172 9.154
R1988 GND.n166 GND.n165 9.154
R1989 GND.n163 GND.n162 9.154
R1990 GND.n160 GND.n157 9.154
R1991 GND.n155 GND.n154 9.154
R1992 GND.n152 GND.n151 9.154
R1993 GND.n149 GND.n148 9.154
R1994 GND.n146 GND.n145 9.154
R1995 GND.n143 GND.n142 9.154
R1996 GND.n140 GND.n139 9.154
R1997 GND.n137 GND.n136 9.154
R1998 GND.n134 GND.n133 9.154
R1999 GND.n131 GND.n130 9.154
R2000 GND.n124 GND.n123 9.154
R2001 GND.n121 GND.n120 9.154
R2002 GND.n118 GND.n117 9.154
R2003 GND.n110 GND.n109 9.154
R2004 GND.n107 GND.n106 9.154
R2005 GND.n104 GND.n103 9.154
R2006 GND.n101 GND.n100 9.154
R2007 GND.n98 GND.n97 9.154
R2008 GND.n91 GND.n90 9.154
R2009 GND.n88 GND.n87 9.154
R2010 GND.n85 GND.n84 9.154
R2011 GND.n77 GND.n76 9.154
R2012 GND.n74 GND.n73 9.154
R2013 GND.n6 GND.n5 9.154
R2014 GND.n12 GND.n11 9.154
R2015 GND.n23 GND.n22 9.154
R2016 GND.n26 GND.n25 9.154
R2017 GND.n33 GND.n32 9.154
R2018 GND.n36 GND.n35 9.154
R2019 GND.n39 GND.n38 9.154
R2020 GND.n42 GND.n41 9.154
R2021 GND.n45 GND.n44 9.154
R2022 GND.n52 GND.n51 9.154
R2023 GND.n55 GND.n54 9.154
R2024 GND.n58 GND.n57 9.154
R2025 GND.n65 GND.n64 9.154
R2026 GND.n68 GND.n67 9.154
R2027 GND.n71 GND.n70 9.154
R2028 GND.n262 GND.n261 8.128
R2029 GND.n755 GND.n754 8.128
R2030 GND.n712 GND.n711 8.128
R2031 GND.n668 GND.n667 8.128
R2032 GND.n635 GND.n634 8.128
R2033 GND.n487 GND.n486 8.128
R2034 GND.n443 GND.n442 8.128
R2035 GND.n410 GND.n409 8.128
R2036 GND.n49 GND.n48 8.128
R2037 GND.n7 GND.n1 4.795
R2038 GND.n404 GND.n403 4.65
R2039 GND.n75 GND.n74 4.65
R2040 GND.n78 GND.n77 4.65
R2041 GND.n86 GND.n85 4.65
R2042 GND.n89 GND.n88 4.65
R2043 GND.n92 GND.n91 4.65
R2044 GND.n99 GND.n98 4.65
R2045 GND.n102 GND.n101 4.65
R2046 GND.n105 GND.n104 4.65
R2047 GND.n108 GND.n107 4.65
R2048 GND.n111 GND.n110 4.65
R2049 GND.n119 GND.n118 4.65
R2050 GND.n122 GND.n121 4.65
R2051 GND.n125 GND.n124 4.65
R2052 GND.n132 GND.n131 4.65
R2053 GND.n135 GND.n134 4.65
R2054 GND.n138 GND.n137 4.65
R2055 GND.n141 GND.n140 4.65
R2056 GND.n144 GND.n143 4.65
R2057 GND.n147 GND.n146 4.65
R2058 GND.n150 GND.n149 4.65
R2059 GND.n153 GND.n152 4.65
R2060 GND.n156 GND.n155 4.65
R2061 GND.n161 GND.n160 4.65
R2062 GND.n164 GND.n163 4.65
R2063 GND.n167 GND.n166 4.65
R2064 GND.n174 GND.n173 4.65
R2065 GND.n177 GND.n176 4.65
R2066 GND.n180 GND.n179 4.65
R2067 GND.n183 GND.n182 4.65
R2068 GND.n186 GND.n185 4.65
R2069 GND.n191 GND.n190 4.65
R2070 GND.n194 GND.n193 4.65
R2071 GND.n197 GND.n196 4.65
R2072 GND.n204 GND.n203 4.65
R2073 GND.n207 GND.n206 4.65
R2074 GND.n210 GND.n209 4.65
R2075 GND.n213 GND.n212 4.65
R2076 GND.n216 GND.n215 4.65
R2077 GND.n221 GND.n220 4.65
R2078 GND.n224 GND.n223 4.65
R2079 GND.n227 GND.n226 4.65
R2080 GND.n234 GND.n233 4.65
R2081 GND.n237 GND.n236 4.65
R2082 GND.n240 GND.n239 4.65
R2083 GND.n243 GND.n242 4.65
R2084 GND.n246 GND.n245 4.65
R2085 GND.n249 GND.n248 4.65
R2086 GND.n252 GND.n251 4.65
R2087 GND.n255 GND.n254 4.65
R2088 GND.n258 GND.n257 4.65
R2089 GND.n265 GND.n264 4.65
R2090 GND.n268 GND.n267 4.65
R2091 GND.n271 GND.n270 4.65
R2092 GND.n278 GND.n277 4.65
R2093 GND.n281 GND.n280 4.65
R2094 GND.n284 GND.n283 4.65
R2095 GND.n287 GND.n286 4.65
R2096 GND.n290 GND.n289 4.65
R2097 GND.n293 GND.n292 4.65
R2098 GND.n296 GND.n295 4.65
R2099 GND.n299 GND.n298 4.65
R2100 GND.n302 GND.n301 4.65
R2101 GND.n307 GND.n306 4.65
R2102 GND.n310 GND.n309 4.65
R2103 GND.n313 GND.n312 4.65
R2104 GND.n320 GND.n319 4.65
R2105 GND.n323 GND.n322 4.65
R2106 GND.n326 GND.n325 4.65
R2107 GND.n329 GND.n328 4.65
R2108 GND.n332 GND.n331 4.65
R2109 GND.n337 GND.n336 4.65
R2110 GND.n340 GND.n339 4.65
R2111 GND.n343 GND.n342 4.65
R2112 GND.n350 GND.n349 4.65
R2113 GND.n353 GND.n352 4.65
R2114 GND.n356 GND.n355 4.65
R2115 GND.n359 GND.n358 4.65
R2116 GND.n362 GND.n361 4.65
R2117 GND.n365 GND.n364 4.65
R2118 GND.n368 GND.n367 4.65
R2119 GND.n371 GND.n370 4.65
R2120 GND.n374 GND.n373 4.65
R2121 GND.n382 GND.n381 4.65
R2122 GND.n385 GND.n384 4.65
R2123 GND.n388 GND.n387 4.65
R2124 GND.n395 GND.n394 4.65
R2125 GND.n398 GND.n397 4.65
R2126 GND.n401 GND.n400 4.65
R2127 GND.n795 GND.n794 4.65
R2128 GND.n792 GND.n791 4.65
R2129 GND.n789 GND.n788 4.65
R2130 GND.n784 GND.n783 4.65
R2131 GND.n781 GND.n780 4.65
R2132 GND.n774 GND.n773 4.65
R2133 GND.n771 GND.n770 4.65
R2134 GND.n768 GND.n767 4.65
R2135 GND.n765 GND.n764 4.65
R2136 GND.n762 GND.n761 4.65
R2137 GND.n759 GND.n758 4.65
R2138 GND.n752 GND.n751 4.65
R2139 GND.n749 GND.n748 4.65
R2140 GND.n742 GND.n741 4.65
R2141 GND.n739 GND.n738 4.65
R2142 GND.n736 GND.n735 4.65
R2143 GND.n733 GND.n732 4.65
R2144 GND.n730 GND.n729 4.65
R2145 GND.n727 GND.n726 4.65
R2146 GND.n724 GND.n723 4.65
R2147 GND.n721 GND.n720 4.65
R2148 GND.n718 GND.n717 4.65
R2149 GND.n715 GND.n714 4.65
R2150 GND.n708 GND.n707 4.65
R2151 GND.n705 GND.n704 4.65
R2152 GND.n698 GND.n697 4.65
R2153 GND.n695 GND.n694 4.65
R2154 GND.n692 GND.n691 4.65
R2155 GND.n689 GND.n688 4.65
R2156 GND.n686 GND.n685 4.65
R2157 GND.n683 GND.n682 4.65
R2158 GND.n680 GND.n679 4.65
R2159 GND.n677 GND.n676 4.65
R2160 GND.n674 GND.n673 4.65
R2161 GND.n671 GND.n670 4.65
R2162 GND.n664 GND.n663 4.65
R2163 GND.n661 GND.n660 4.65
R2164 GND.n654 GND.n653 4.65
R2165 GND.n651 GND.n650 4.65
R2166 GND.n648 GND.n647 4.65
R2167 GND.n645 GND.n644 4.65
R2168 GND.n642 GND.n641 4.65
R2169 GND.n639 GND.n638 4.65
R2170 GND.n632 GND.n631 4.65
R2171 GND.n629 GND.n628 4.65
R2172 GND.n622 GND.n621 4.65
R2173 GND.n619 GND.n618 4.65
R2174 GND.n616 GND.n615 4.65
R2175 GND.n613 GND.n612 4.65
R2176 GND.n610 GND.n609 4.65
R2177 GND.n607 GND.n606 4.65
R2178 GND.n604 GND.n603 4.65
R2179 GND.n601 GND.n600 4.65
R2180 GND.n598 GND.n597 4.65
R2181 GND.n595 GND.n594 4.65
R2182 GND.n587 GND.n586 4.65
R2183 GND.n584 GND.n583 4.65
R2184 GND.n577 GND.n576 4.65
R2185 GND.n574 GND.n573 4.65
R2186 GND.n571 GND.n570 4.65
R2187 GND.n568 GND.n567 4.65
R2188 GND.n565 GND.n564 4.65
R2189 GND.n562 GND.n561 4.65
R2190 GND.n557 GND.n556 4.65
R2191 GND.n554 GND.n553 4.65
R2192 GND.n547 GND.n546 4.65
R2193 GND.n544 GND.n543 4.65
R2194 GND.n541 GND.n540 4.65
R2195 GND.n538 GND.n537 4.65
R2196 GND.n535 GND.n534 4.65
R2197 GND.n532 GND.n531 4.65
R2198 GND.n527 GND.n526 4.65
R2199 GND.n524 GND.n523 4.65
R2200 GND.n517 GND.n516 4.65
R2201 GND.n514 GND.n513 4.65
R2202 GND.n511 GND.n510 4.65
R2203 GND.n508 GND.n507 4.65
R2204 GND.n505 GND.n504 4.65
R2205 GND.n502 GND.n501 4.65
R2206 GND.n499 GND.n498 4.65
R2207 GND.n496 GND.n495 4.65
R2208 GND.n493 GND.n492 4.65
R2209 GND.n490 GND.n489 4.65
R2210 GND.n483 GND.n482 4.65
R2211 GND.n480 GND.n479 4.65
R2212 GND.n473 GND.n472 4.65
R2213 GND.n470 GND.n469 4.65
R2214 GND.n467 GND.n466 4.65
R2215 GND.n464 GND.n463 4.65
R2216 GND.n461 GND.n460 4.65
R2217 GND.n458 GND.n457 4.65
R2218 GND.n455 GND.n454 4.65
R2219 GND.n452 GND.n451 4.65
R2220 GND.n449 GND.n448 4.65
R2221 GND.n446 GND.n445 4.65
R2222 GND.n439 GND.n438 4.65
R2223 GND.n436 GND.n435 4.65
R2224 GND.n429 GND.n428 4.65
R2225 GND.n426 GND.n425 4.65
R2226 GND.n423 GND.n422 4.65
R2227 GND.n420 GND.n419 4.65
R2228 GND.n417 GND.n416 4.65
R2229 GND.n414 GND.n413 4.65
R2230 GND.n407 GND.n406 4.65
R2231 GND.n7 GND.n6 4.65
R2232 GND.n13 GND.n12 4.65
R2233 GND.n24 GND.n23 4.65
R2234 GND.n27 GND.n26 4.65
R2235 GND.n34 GND.n33 4.65
R2236 GND.n37 GND.n36 4.65
R2237 GND.n40 GND.n39 4.65
R2238 GND.n43 GND.n42 4.65
R2239 GND.n46 GND.n45 4.65
R2240 GND.n53 GND.n52 4.65
R2241 GND.n56 GND.n55 4.65
R2242 GND.n59 GND.n58 4.65
R2243 GND.n66 GND.n65 4.65
R2244 GND.n69 GND.n68 4.65
R2245 GND.n72 GND.n71 4.65
R2246 GND.n15 GND.n14 4.504
R2247 GND.n6 GND.n4 4.129
R2248 GND.n52 GND.n50 4.129
R2249 GND.n85 GND.n83 4.129
R2250 GND.n118 GND.n116 4.129
R2251 GND.n190 GND.n188 4.129
R2252 GND.n220 GND.n218 4.129
R2253 GND.n336 GND.n334 4.129
R2254 GND.n788 GND.n786 4.129
R2255 GND.n758 GND.n756 4.129
R2256 GND.n638 GND.n636 4.129
R2257 GND.n561 GND.n559 4.129
R2258 GND.n531 GND.n529 4.129
R2259 GND.n413 GND.n411 4.129
R2260 GND.n23 GND.n21 3.716
R2261 GND.t28 GND.n15 2.452
R2262 GND.n1 GND.n0 0.475
R2263 GND.n403 GND.n402 0.474
R2264 GND.n9 GND.n8 0.376
R2265 GND.n34 GND.n27 0.29
R2266 GND.n66 GND.n59 0.29
R2267 GND.n99 GND.n92 0.29
R2268 GND.n132 GND.n125 0.29
R2269 GND.n174 GND.n167 0.29
R2270 GND.n204 GND.n197 0.29
R2271 GND.n234 GND.n227 0.29
R2272 GND.n278 GND.n271 0.29
R2273 GND.n320 GND.n313 0.29
R2274 GND.n350 GND.n343 0.29
R2275 GND.n395 GND.n388 0.29
R2276 GND.n781 GND.n774 0.29
R2277 GND.n749 GND.n742 0.29
R2278 GND.n705 GND.n698 0.29
R2279 GND.n661 GND.n654 0.29
R2280 GND.n629 GND.n622 0.29
R2281 GND.n584 GND.n577 0.29
R2282 GND.n554 GND.n547 0.29
R2283 GND.n524 GND.n517 0.29
R2284 GND.n480 GND.n473 0.29
R2285 GND.n436 GND.n429 0.29
R2286 GND.n404 GND 0.207
R2287 GND.n12 GND.n10 0.206
R2288 GND.n160 GND.n159 0.206
R2289 GND.n264 GND.n263 0.206
R2290 GND.n306 GND.n305 0.206
R2291 GND.n381 GND.n380 0.206
R2292 GND.n714 GND.n713 0.206
R2293 GND.n670 GND.n669 0.206
R2294 GND.n594 GND.n593 0.206
R2295 GND.n489 GND.n488 0.206
R2296 GND.n445 GND.n444 0.206
R2297 GND.n150 GND.n147 0.197
R2298 GND.n252 GND.n249 0.197
R2299 GND.n296 GND.n293 0.197
R2300 GND.n368 GND.n365 0.197
R2301 GND.n727 GND.n724 0.197
R2302 GND.n683 GND.n680 0.197
R2303 GND.n607 GND.n604 0.197
R2304 GND.n502 GND.n499 0.197
R2305 GND.n458 GND.n455 0.197
R2306 GND.n46 GND.n43 0.181
R2307 GND.n78 GND.n75 0.181
R2308 GND.n111 GND.n108 0.181
R2309 GND.n186 GND.n183 0.181
R2310 GND.n216 GND.n213 0.181
R2311 GND.n332 GND.n329 0.181
R2312 GND.n795 GND.n792 0.181
R2313 GND.n765 GND.n762 0.181
R2314 GND.n645 GND.n642 0.181
R2315 GND.n568 GND.n565 0.181
R2316 GND.n538 GND.n535 0.181
R2317 GND.n420 GND.n417 0.181
R2318 GND.n13 GND.n7 0.157
R2319 GND.n24 GND.n13 0.157
R2320 GND.n27 GND.n24 0.145
R2321 GND.n37 GND.n34 0.145
R2322 GND.n40 GND.n37 0.145
R2323 GND.n43 GND.n40 0.145
R2324 GND.n53 GND.n46 0.145
R2325 GND.n56 GND.n53 0.145
R2326 GND.n59 GND.n56 0.145
R2327 GND.n69 GND.n66 0.145
R2328 GND.n72 GND.n69 0.145
R2329 GND.n75 GND.n72 0.145
R2330 GND.n86 GND.n78 0.145
R2331 GND.n89 GND.n86 0.145
R2332 GND.n92 GND.n89 0.145
R2333 GND.n102 GND.n99 0.145
R2334 GND.n105 GND.n102 0.145
R2335 GND.n108 GND.n105 0.145
R2336 GND.n119 GND.n111 0.145
R2337 GND.n122 GND.n119 0.145
R2338 GND.n125 GND.n122 0.145
R2339 GND.n135 GND.n132 0.145
R2340 GND.n138 GND.n135 0.145
R2341 GND.n141 GND.n138 0.145
R2342 GND.n144 GND.n141 0.145
R2343 GND.n147 GND.n144 0.145
R2344 GND.n153 GND.n150 0.145
R2345 GND.n156 GND.n153 0.145
R2346 GND.n161 GND.n156 0.145
R2347 GND.n164 GND.n161 0.145
R2348 GND.n167 GND.n164 0.145
R2349 GND.n177 GND.n174 0.145
R2350 GND.n180 GND.n177 0.145
R2351 GND.n183 GND.n180 0.145
R2352 GND.n191 GND.n186 0.145
R2353 GND.n194 GND.n191 0.145
R2354 GND.n197 GND.n194 0.145
R2355 GND.n207 GND.n204 0.145
R2356 GND.n210 GND.n207 0.145
R2357 GND.n213 GND.n210 0.145
R2358 GND.n221 GND.n216 0.145
R2359 GND.n224 GND.n221 0.145
R2360 GND.n227 GND.n224 0.145
R2361 GND.n237 GND.n234 0.145
R2362 GND.n240 GND.n237 0.145
R2363 GND.n243 GND.n240 0.145
R2364 GND.n246 GND.n243 0.145
R2365 GND.n249 GND.n246 0.145
R2366 GND.n255 GND.n252 0.145
R2367 GND.n258 GND.n255 0.145
R2368 GND.n265 GND.n258 0.145
R2369 GND.n268 GND.n265 0.145
R2370 GND.n271 GND.n268 0.145
R2371 GND.n281 GND.n278 0.145
R2372 GND.n284 GND.n281 0.145
R2373 GND.n287 GND.n284 0.145
R2374 GND.n290 GND.n287 0.145
R2375 GND.n293 GND.n290 0.145
R2376 GND.n299 GND.n296 0.145
R2377 GND.n302 GND.n299 0.145
R2378 GND.n307 GND.n302 0.145
R2379 GND.n310 GND.n307 0.145
R2380 GND.n313 GND.n310 0.145
R2381 GND.n323 GND.n320 0.145
R2382 GND.n326 GND.n323 0.145
R2383 GND.n329 GND.n326 0.145
R2384 GND.n337 GND.n332 0.145
R2385 GND.n340 GND.n337 0.145
R2386 GND.n343 GND.n340 0.145
R2387 GND.n353 GND.n350 0.145
R2388 GND.n356 GND.n353 0.145
R2389 GND.n359 GND.n356 0.145
R2390 GND.n362 GND.n359 0.145
R2391 GND.n365 GND.n362 0.145
R2392 GND.n371 GND.n368 0.145
R2393 GND.n374 GND.n371 0.145
R2394 GND.n382 GND.n374 0.145
R2395 GND.n385 GND.n382 0.145
R2396 GND.n388 GND.n385 0.145
R2397 GND.n398 GND.n395 0.145
R2398 GND.n401 GND.n398 0.145
R2399 GND.n792 GND.n789 0.145
R2400 GND.n789 GND.n784 0.145
R2401 GND.n784 GND.n781 0.145
R2402 GND.n774 GND.n771 0.145
R2403 GND.n771 GND.n768 0.145
R2404 GND.n768 GND.n765 0.145
R2405 GND.n762 GND.n759 0.145
R2406 GND.n759 GND.n752 0.145
R2407 GND.n752 GND.n749 0.145
R2408 GND.n742 GND.n739 0.145
R2409 GND.n739 GND.n736 0.145
R2410 GND.n736 GND.n733 0.145
R2411 GND.n733 GND.n730 0.145
R2412 GND.n730 GND.n727 0.145
R2413 GND.n724 GND.n721 0.145
R2414 GND.n721 GND.n718 0.145
R2415 GND.n718 GND.n715 0.145
R2416 GND.n715 GND.n708 0.145
R2417 GND.n708 GND.n705 0.145
R2418 GND.n698 GND.n695 0.145
R2419 GND.n695 GND.n692 0.145
R2420 GND.n692 GND.n689 0.145
R2421 GND.n689 GND.n686 0.145
R2422 GND.n686 GND.n683 0.145
R2423 GND.n680 GND.n677 0.145
R2424 GND.n677 GND.n674 0.145
R2425 GND.n674 GND.n671 0.145
R2426 GND.n671 GND.n664 0.145
R2427 GND.n664 GND.n661 0.145
R2428 GND.n654 GND.n651 0.145
R2429 GND.n651 GND.n648 0.145
R2430 GND.n648 GND.n645 0.145
R2431 GND.n642 GND.n639 0.145
R2432 GND.n639 GND.n632 0.145
R2433 GND.n632 GND.n629 0.145
R2434 GND.n622 GND.n619 0.145
R2435 GND.n619 GND.n616 0.145
R2436 GND.n616 GND.n613 0.145
R2437 GND.n613 GND.n610 0.145
R2438 GND.n610 GND.n607 0.145
R2439 GND.n604 GND.n601 0.145
R2440 GND.n601 GND.n598 0.145
R2441 GND.n598 GND.n595 0.145
R2442 GND.n595 GND.n587 0.145
R2443 GND.n587 GND.n584 0.145
R2444 GND.n577 GND.n574 0.145
R2445 GND.n574 GND.n571 0.145
R2446 GND.n571 GND.n568 0.145
R2447 GND.n565 GND.n562 0.145
R2448 GND.n562 GND.n557 0.145
R2449 GND.n557 GND.n554 0.145
R2450 GND.n547 GND.n544 0.145
R2451 GND.n544 GND.n541 0.145
R2452 GND.n541 GND.n538 0.145
R2453 GND.n535 GND.n532 0.145
R2454 GND.n532 GND.n527 0.145
R2455 GND.n527 GND.n524 0.145
R2456 GND.n517 GND.n514 0.145
R2457 GND.n514 GND.n511 0.145
R2458 GND.n511 GND.n508 0.145
R2459 GND.n508 GND.n505 0.145
R2460 GND.n505 GND.n502 0.145
R2461 GND.n499 GND.n496 0.145
R2462 GND.n496 GND.n493 0.145
R2463 GND.n493 GND.n490 0.145
R2464 GND.n490 GND.n483 0.145
R2465 GND.n483 GND.n480 0.145
R2466 GND.n473 GND.n470 0.145
R2467 GND.n470 GND.n467 0.145
R2468 GND.n467 GND.n464 0.145
R2469 GND.n464 GND.n461 0.145
R2470 GND.n461 GND.n458 0.145
R2471 GND.n455 GND.n452 0.145
R2472 GND.n452 GND.n449 0.145
R2473 GND.n449 GND.n446 0.145
R2474 GND.n446 GND.n439 0.145
R2475 GND.n439 GND.n436 0.145
R2476 GND.n429 GND.n426 0.145
R2477 GND.n426 GND.n423 0.145
R2478 GND.n423 GND.n420 0.145
R2479 GND.n417 GND.n414 0.145
R2480 GND.n414 GND.n407 0.145
R2481 GND.n407 GND.n404 0.145
R2482 GND GND.n401 0.086
R2483 GND GND.n795 0.058
R2484 D.n5 D.t1 480.392
R2485 D.n2 D.t0 480.392
R2486 D.n0 D.t5 480.392
R2487 D.n5 D.t4 403.272
R2488 D.n2 D.t7 403.272
R2489 D.n0 D.t8 403.272
R2490 D.n6 D.n5 282.724
R2491 D.n3 D.n2 282.724
R2492 D.n1 D.n0 282.724
R2493 D.n6 D.t3 178.533
R2494 D.n3 D.t2 178.533
R2495 D.n1 D.t6 178.533
R2496 D.n4 D.n1 22.56
R2497 D.n7 D.n4 17.91
R2498 D.n4 D.n3 4.65
R2499 D.n7 D.n6 4.65
R2500 D.n7 D 0.046
R2501 a_5101_1050.n3 a_5101_1050.t6 512.525
R2502 a_5101_1050.n1 a_5101_1050.t5 512.525
R2503 a_5101_1050.n3 a_5101_1050.t9 371.139
R2504 a_5101_1050.n1 a_5101_1050.t7 371.139
R2505 a_5101_1050.n2 a_5101_1050.t10 305.674
R2506 a_5101_1050.n4 a_5101_1050.t8 305.298
R2507 a_5101_1050.n4 a_5101_1050.n3 291.648
R2508 a_5101_1050.n2 a_5101_1050.n1 291.272
R2509 a_5101_1050.n7 a_5101_1050.n6 271.602
R2510 a_5101_1050.n8 a_5101_1050.n7 215.717
R2511 a_5101_1050.n9 a_5101_1050.n8 157.963
R2512 a_5101_1050.n8 a_5101_1050.n0 91.706
R2513 a_5101_1050.n0 a_5101_1050.t2 14.282
R2514 a_5101_1050.n0 a_5101_1050.t1 14.282
R2515 a_5101_1050.t4 a_5101_1050.n9 14.282
R2516 a_5101_1050.n9 a_5101_1050.t3 14.282
R2517 a_5101_1050.n5 a_5101_1050.n2 8.138
R2518 a_5101_1050.n7 a_5101_1050.n5 5.964
R2519 a_5101_1050.n5 a_5101_1050.n4 4.65
R2520 CLK.n15 CLK.t12 472.359
R2521 CLK.n6 CLK.t13 472.359
R2522 CLK.n0 CLK.t17 472.359
R2523 CLK.n20 CLK.t5 459.505
R2524 CLK.n11 CLK.t15 459.505
R2525 CLK.n2 CLK.t11 459.505
R2526 CLK.n21 CLK.t9 399.181
R2527 CLK.n12 CLK.t16 399.181
R2528 CLK.n3 CLK.t4 399.181
R2529 CLK.n1 CLK.t7 398.558
R2530 CLK.n17 CLK.t1 397.101
R2531 CLK.n8 CLK.t6 397.101
R2532 CLK.n20 CLK.t10 384.527
R2533 CLK.n15 CLK.t14 384.527
R2534 CLK.n11 CLK.t0 384.527
R2535 CLK.n6 CLK.t3 384.527
R2536 CLK.n2 CLK.t2 384.527
R2537 CLK.n0 CLK.t8 384.527
R2538 CLK.n21 CLK.n20 33.832
R2539 CLK.n3 CLK.n2 33.832
R2540 CLK.n12 CLK.n11 33.832
R2541 CLK.n1 CLK.n0 32.394
R2542 CLK.n16 CLK.n15 30.822
R2543 CLK.n7 CLK.n6 30.822
R2544 CLK.n5 CLK.n4 11.101
R2545 CLK.n14 CLK.n13 11.101
R2546 CLK.n4 CLK.n1 8.215
R2547 CLK.n13 CLK.n10 6.718
R2548 CLK.n22 CLK.n19 6.718
R2549 CLK.n17 CLK.n16 4.577
R2550 CLK.n8 CLK.n7 4.577
R2551 CLK.n9 CLK.n8 4.282
R2552 CLK.n18 CLK.n17 4.282
R2553 CLK.n4 CLK.n3 2.079
R2554 CLK.n13 CLK.n12 2.079
R2555 CLK.n22 CLK.n21 2.079
R2556 CLK.n22 CLK 0.046
R2557 CLK.n10 CLK.n9 0.038
R2558 CLK.n19 CLK.n18 0.038
R2559 CLK.n9 CLK.n5 0.008
R2560 CLK.n18 CLK.n14 0.008
R2561 a_5227_411.n1 a_5227_411.t8 480.392
R2562 a_5227_411.n3 a_5227_411.t7 472.359
R2563 a_5227_411.n2 a_5227_411.t12 412.921
R2564 a_5227_411.n1 a_5227_411.t11 403.272
R2565 a_5227_411.n3 a_5227_411.t10 384.527
R2566 a_5227_411.n9 a_5227_411.n8 379.101
R2567 a_5227_411.n4 a_5227_411.t9 370.613
R2568 a_5227_411.n12 a_5227_411.n11 161.352
R2569 a_5227_411.n4 a_5227_411.n3 127.096
R2570 a_5227_411.n10 a_5227_411.n9 123.126
R2571 a_5227_411.n2 a_5227_411.n1 115.571
R2572 a_5227_411.n10 a_5227_411.n0 95.095
R2573 a_5227_411.n13 a_5227_411.n12 95.094
R2574 a_5227_411.n12 a_5227_411.n10 66.258
R2575 a_5227_411.n8 a_5227_411.n7 22.578
R2576 a_5227_411.n0 a_5227_411.t2 14.282
R2577 a_5227_411.n0 a_5227_411.t1 14.282
R2578 a_5227_411.n11 a_5227_411.t6 14.282
R2579 a_5227_411.n11 a_5227_411.t5 14.282
R2580 a_5227_411.n13 a_5227_411.t3 14.282
R2581 a_5227_411.t4 a_5227_411.n13 14.282
R2582 a_5227_411.n5 a_5227_411.n2 11.954
R2583 a_5227_411.n5 a_5227_411.n4 8.682
R2584 a_5227_411.n8 a_5227_411.n6 8.58
R2585 a_5227_411.n9 a_5227_411.n5 4.65
R2586 a_3599_411.n7 a_3599_411.t15 512.525
R2587 a_3599_411.n6 a_3599_411.t10 512.525
R2588 a_3599_411.n11 a_3599_411.t13 472.359
R2589 a_3599_411.n11 a_3599_411.t9 384.527
R2590 a_3599_411.n7 a_3599_411.t11 371.139
R2591 a_3599_411.n6 a_3599_411.t7 371.139
R2592 a_3599_411.n8 a_3599_411.n7 343.521
R2593 a_3599_411.n12 a_3599_411.t14 287.037
R2594 a_3599_411.n16 a_3599_411.n14 280.357
R2595 a_3599_411.n10 a_3599_411.n6 259.945
R2596 a_3599_411.n12 a_3599_411.n11 210.673
R2597 a_3599_411.n14 a_3599_411.n5 207.058
R2598 a_3599_411.n8 a_3599_411.t8 172.106
R2599 a_3599_411.n9 a_3599_411.t12 165.68
R2600 a_3599_411.n4 a_3599_411.n3 161.352
R2601 a_3599_411.n5 a_3599_411.n1 95.095
R2602 a_3599_411.n4 a_3599_411.n2 95.095
R2603 a_3599_411.n10 a_3599_411.n9 83.576
R2604 a_3599_411.n5 a_3599_411.n4 66.258
R2605 a_3599_411.n17 a_3599_411.n0 55.263
R2606 a_3599_411.n13 a_3599_411.n10 45.413
R2607 a_3599_411.n16 a_3599_411.n15 30
R2608 a_3599_411.n17 a_3599_411.n16 23.684
R2609 a_3599_411.n1 a_3599_411.t3 14.282
R2610 a_3599_411.n1 a_3599_411.t0 14.282
R2611 a_3599_411.n2 a_3599_411.t5 14.282
R2612 a_3599_411.n2 a_3599_411.t4 14.282
R2613 a_3599_411.n3 a_3599_411.t1 14.282
R2614 a_3599_411.n3 a_3599_411.t6 14.282
R2615 a_3599_411.n9 a_3599_411.n8 10.343
R2616 a_3599_411.n13 a_3599_411.n12 8.685
R2617 a_3599_411.n14 a_3599_411.n13 4.65
R2618 a_15533_1051.t0 a_15533_1051.n5 179.898
R2619 a_15533_1051.n3 a_15533_1051.n2 165.613
R2620 a_15533_1051.n3 a_15533_1051.n1 142.653
R2621 a_15533_1051.n5 a_15533_1051.n4 106.183
R2622 a_15533_1051.n5 a_15533_1051.n0 99.355
R2623 a_15533_1051.n4 a_15533_1051.n3 82.665
R2624 a_15533_1051.n4 a_15533_1051.t6 73.712
R2625 a_15533_1051.n1 a_15533_1051.t7 14.282
R2626 a_15533_1051.n1 a_15533_1051.t4 14.282
R2627 a_15533_1051.n2 a_15533_1051.t1 14.282
R2628 a_15533_1051.n2 a_15533_1051.t2 14.282
R2629 a_15533_1051.n0 a_15533_1051.t3 14.282
R2630 a_15533_1051.n0 a_15533_1051.t5 14.282
R2631 a_14869_1051.n4 a_14869_1051.t5 179.895
R2632 a_14869_1051.n2 a_14869_1051.n1 157.021
R2633 a_14869_1051.n2 a_14869_1051.n0 124.955
R2634 a_14869_1051.n4 a_14869_1051.n3 106.183
R2635 a_14869_1051.n5 a_14869_1051.n4 99.358
R2636 a_14869_1051.n3 a_14869_1051.n2 82.65
R2637 a_14869_1051.n3 a_14869_1051.t0 73.712
R2638 a_14869_1051.n0 a_14869_1051.t6 14.282
R2639 a_14869_1051.n0 a_14869_1051.t7 14.282
R2640 a_14869_1051.n1 a_14869_1051.t2 14.282
R2641 a_14869_1051.n1 a_14869_1051.t3 14.282
R2642 a_14869_1051.n5 a_14869_1051.t4 14.282
R2643 a_14869_1051.t1 a_14869_1051.n5 14.282
R2644 a_217_1050.n3 a_217_1050.t6 512.525
R2645 a_217_1050.n1 a_217_1050.t10 512.525
R2646 a_217_1050.n3 a_217_1050.t9 371.139
R2647 a_217_1050.n1 a_217_1050.t5 371.139
R2648 a_217_1050.n2 a_217_1050.t8 305.674
R2649 a_217_1050.n4 a_217_1050.t7 305.298
R2650 a_217_1050.n4 a_217_1050.n3 291.648
R2651 a_217_1050.n2 a_217_1050.n1 291.272
R2652 a_217_1050.n7 a_217_1050.n6 271.602
R2653 a_217_1050.n8 a_217_1050.n7 215.717
R2654 a_217_1050.n9 a_217_1050.n8 157.963
R2655 a_217_1050.n8 a_217_1050.n0 91.706
R2656 a_217_1050.n0 a_217_1050.t4 14.282
R2657 a_217_1050.n0 a_217_1050.t1 14.282
R2658 a_217_1050.t3 a_217_1050.n9 14.282
R2659 a_217_1050.n9 a_217_1050.t2 14.282
R2660 a_217_1050.n5 a_217_1050.n2 8.138
R2661 a_217_1050.n7 a_217_1050.n5 5.964
R2662 a_217_1050.n5 a_217_1050.n4 4.65
R2663 a_1265_989.n2 a_1265_989.t11 454.685
R2664 a_1265_989.n4 a_1265_989.t13 454.685
R2665 a_1265_989.n0 a_1265_989.t6 454.685
R2666 a_1265_989.n2 a_1265_989.t5 428.979
R2667 a_1265_989.n4 a_1265_989.t10 428.979
R2668 a_1265_989.n0 a_1265_989.t9 428.979
R2669 a_1265_989.n3 a_1265_989.t7 339.542
R2670 a_1265_989.n5 a_1265_989.t8 339.542
R2671 a_1265_989.n1 a_1265_989.t12 339.542
R2672 a_1265_989.n12 a_1265_989.n11 333.44
R2673 a_1265_989.n14 a_1265_989.n13 157.964
R2674 a_1265_989.n3 a_1265_989.n2 143.429
R2675 a_1265_989.n5 a_1265_989.n4 143.429
R2676 a_1265_989.n1 a_1265_989.n0 143.429
R2677 a_1265_989.n14 a_1265_989.n12 132.141
R2678 a_1265_989.n15 a_1265_989.n14 91.705
R2679 a_1265_989.n11 a_1265_989.n10 30
R2680 a_1265_989.n9 a_1265_989.n8 24.383
R2681 a_1265_989.n11 a_1265_989.n9 23.684
R2682 a_1265_989.n13 a_1265_989.t0 14.282
R2683 a_1265_989.n13 a_1265_989.t4 14.282
R2684 a_1265_989.t2 a_1265_989.n15 14.282
R2685 a_1265_989.n15 a_1265_989.t1 14.282
R2686 a_1265_989.n7 a_1265_989.n1 10.046
R2687 a_1265_989.n6 a_1265_989.n5 8.141
R2688 a_1265_989.n6 a_1265_989.n3 4.65
R2689 a_1265_989.n12 a_1265_989.n7 4.65
R2690 a_1265_989.n7 a_1265_989.n6 2.947
R2691 a_1905_1050.n0 a_1905_1050.t7 480.392
R2692 a_1905_1050.n0 a_1905_1050.t9 403.272
R2693 a_1905_1050.n1 a_1905_1050.t8 301.486
R2694 a_1905_1050.n6 a_1905_1050.n5 252.498
R2695 a_1905_1050.n10 a_1905_1050.n6 234.917
R2696 a_1905_1050.n1 a_1905_1050.n0 227.006
R2697 a_1905_1050.n9 a_1905_1050.n8 161.352
R2698 a_1905_1050.n9 a_1905_1050.n7 95.095
R2699 a_1905_1050.n11 a_1905_1050.n10 95.094
R2700 a_1905_1050.n10 a_1905_1050.n9 66.258
R2701 a_1905_1050.n5 a_1905_1050.n4 30
R2702 a_1905_1050.n3 a_1905_1050.n2 24.383
R2703 a_1905_1050.n5 a_1905_1050.n3 23.684
R2704 a_1905_1050.n7 a_1905_1050.t5 14.282
R2705 a_1905_1050.n7 a_1905_1050.t6 14.282
R2706 a_1905_1050.n8 a_1905_1050.t3 14.282
R2707 a_1905_1050.n8 a_1905_1050.t4 14.282
R2708 a_1905_1050.t1 a_1905_1050.n11 14.282
R2709 a_1905_1050.n11 a_1905_1050.t0 14.282
R2710 a_1905_1050.n6 a_1905_1050.n1 10.615
R2711 a_10111_411.n1 a_10111_411.t11 480.392
R2712 a_10111_411.n3 a_10111_411.t9 472.359
R2713 a_10111_411.n2 a_10111_411.t12 412.921
R2714 a_10111_411.n1 a_10111_411.t8 403.272
R2715 a_10111_411.n3 a_10111_411.t7 384.527
R2716 a_10111_411.n9 a_10111_411.n8 379.101
R2717 a_10111_411.n4 a_10111_411.t10 370.613
R2718 a_10111_411.n12 a_10111_411.n11 161.352
R2719 a_10111_411.n4 a_10111_411.n3 127.096
R2720 a_10111_411.n10 a_10111_411.n9 123.126
R2721 a_10111_411.n2 a_10111_411.n1 115.571
R2722 a_10111_411.n10 a_10111_411.n0 95.095
R2723 a_10111_411.n13 a_10111_411.n12 95.094
R2724 a_10111_411.n12 a_10111_411.n10 66.258
R2725 a_10111_411.n8 a_10111_411.n7 22.578
R2726 a_10111_411.n0 a_10111_411.t6 14.282
R2727 a_10111_411.n0 a_10111_411.t4 14.282
R2728 a_10111_411.n11 a_10111_411.t3 14.282
R2729 a_10111_411.n11 a_10111_411.t0 14.282
R2730 a_10111_411.n13 a_10111_411.t1 14.282
R2731 a_10111_411.t2 a_10111_411.n13 14.282
R2732 a_10111_411.n5 a_10111_411.n2 11.954
R2733 a_10111_411.n5 a_10111_411.n4 8.682
R2734 a_10111_411.n8 a_10111_411.n6 8.58
R2735 a_10111_411.n9 a_10111_411.n5 4.65
R2736 a_9985_1050.n3 a_9985_1050.t9 512.525
R2737 a_9985_1050.n1 a_9985_1050.t8 512.525
R2738 a_9985_1050.n3 a_9985_1050.t7 371.139
R2739 a_9985_1050.n1 a_9985_1050.t10 371.139
R2740 a_9985_1050.n2 a_9985_1050.t6 305.674
R2741 a_9985_1050.n4 a_9985_1050.t5 305.298
R2742 a_9985_1050.n4 a_9985_1050.n3 291.648
R2743 a_9985_1050.n2 a_9985_1050.n1 291.272
R2744 a_9985_1050.n10 a_9985_1050.n9 249.863
R2745 a_9985_1050.n11 a_9985_1050.n10 215.717
R2746 a_9985_1050.n12 a_9985_1050.n11 157.963
R2747 a_9985_1050.n11 a_9985_1050.n0 91.706
R2748 a_9985_1050.n9 a_9985_1050.n8 30
R2749 a_9985_1050.n7 a_9985_1050.n6 24.383
R2750 a_9985_1050.n9 a_9985_1050.n7 23.684
R2751 a_9985_1050.n0 a_9985_1050.t2 14.282
R2752 a_9985_1050.n0 a_9985_1050.t3 14.282
R2753 a_9985_1050.t1 a_9985_1050.n12 14.282
R2754 a_9985_1050.n12 a_9985_1050.t0 14.282
R2755 a_9985_1050.n5 a_9985_1050.n2 8.138
R2756 a_9985_1050.n10 a_9985_1050.n5 5.964
R2757 a_9985_1050.n5 a_9985_1050.n4 4.65
R2758 a_10525_103.t0 a_10525_103.n7 59.616
R2759 a_10525_103.n4 a_10525_103.n2 54.496
R2760 a_10525_103.n4 a_10525_103.n3 54.496
R2761 a_10525_103.n1 a_10525_103.n0 24.679
R2762 a_10525_103.n6 a_10525_103.n4 7.859
R2763 a_10525_103.t0 a_10525_103.n1 7.505
R2764 a_10525_103.t0 a_10525_103.n6 3.034
R2765 a_10525_103.n6 a_10525_103.n5 0.443
R2766 a_16096_101.n3 a_16096_101.n1 42.788
R2767 a_16096_101.t0 a_16096_101.n0 8.137
R2768 a_16096_101.n3 a_16096_101.n2 4.665
R2769 a_16096_101.t0 a_16096_101.n3 0.06
R2770 a_4996_101.n3 a_4996_101.n1 42.788
R2771 a_4996_101.t0 a_4996_101.n0 8.137
R2772 a_4996_101.n3 a_4996_101.n2 4.665
R2773 a_4996_101.t0 a_4996_101.n3 0.06
R2774 a_13367_411.n6 a_13367_411.t7 475.572
R2775 a_13367_411.n11 a_13367_411.t14 472.359
R2776 a_13367_411.n8 a_13367_411.t10 469.145
R2777 a_13367_411.n11 a_13367_411.t9 384.527
R2778 a_13367_411.n8 a_13367_411.t13 384.527
R2779 a_13367_411.n6 a_13367_411.t12 384.527
R2780 a_13367_411.n12 a_13367_411.t8 370.613
R2781 a_13367_411.n9 a_13367_411.t15 370.613
R2782 a_13367_411.n7 a_13367_411.t11 370.613
R2783 a_13367_411.n16 a_13367_411.n14 363.934
R2784 a_13367_411.n4 a_13367_411.n3 161.352
R2785 a_13367_411.n7 a_13367_411.n6 128.028
R2786 a_13367_411.n12 a_13367_411.n11 127.096
R2787 a_13367_411.n9 a_13367_411.n8 126.97
R2788 a_13367_411.n14 a_13367_411.n5 123.481
R2789 a_13367_411.n5 a_13367_411.n1 95.095
R2790 a_13367_411.n4 a_13367_411.n2 95.095
R2791 a_13367_411.n5 a_13367_411.n4 66.258
R2792 a_13367_411.n17 a_13367_411.n0 55.263
R2793 a_13367_411.n16 a_13367_411.n15 30
R2794 a_13367_411.n17 a_13367_411.n16 23.684
R2795 a_13367_411.n1 a_13367_411.t0 14.282
R2796 a_13367_411.n1 a_13367_411.t1 14.282
R2797 a_13367_411.n2 a_13367_411.t5 14.282
R2798 a_13367_411.n2 a_13367_411.t2 14.282
R2799 a_13367_411.n3 a_13367_411.t3 14.282
R2800 a_13367_411.n3 a_13367_411.t4 14.282
R2801 a_13367_411.n10 a_13367_411.n7 9.501
R2802 a_13367_411.n13 a_13367_411.n12 8.685
R2803 a_13367_411.n10 a_13367_411.n9 4.65
R2804 a_13367_411.n14 a_13367_411.n13 4.65
R2805 a_13367_411.n13 a_13367_411.n10 1.859
R2806 a_15044_209.n1 a_15044_209.t7 512.525
R2807 a_15044_209.n1 a_15044_209.t9 371.139
R2808 a_15044_209.n2 a_15044_209.t8 338.57
R2809 a_15044_209.n14 a_15044_209.n13 227.387
R2810 a_15044_209.n2 a_15044_209.n1 191.629
R2811 a_15044_209.n16 a_15044_209.n15 165.613
R2812 a_15044_209.n15 a_15044_209.n14 132.893
R2813 a_15044_209.n13 a_15044_209.n12 127.909
R2814 a_15044_209.n11 a_15044_209.n10 112.771
R2815 a_15044_209.n11 a_15044_209.n6 110.702
R2816 a_15044_209.n15 a_15044_209.n0 99.355
R2817 a_15044_209.n6 a_15044_209.n5 30
R2818 a_15044_209.n10 a_15044_209.n9 30
R2819 a_15044_209.n4 a_15044_209.n3 24.383
R2820 a_15044_209.n8 a_15044_209.n7 24.383
R2821 a_15044_209.n6 a_15044_209.n4 23.684
R2822 a_15044_209.n10 a_15044_209.n8 23.684
R2823 a_15044_209.n0 a_15044_209.t4 14.282
R2824 a_15044_209.n0 a_15044_209.t3 14.282
R2825 a_15044_209.n16 a_15044_209.t0 14.282
R2826 a_15044_209.t1 a_15044_209.n16 14.282
R2827 a_15044_209.n14 a_15044_209.n2 10.343
R2828 a_15044_209.n13 a_15044_209.n11 7.053
R2829 a_6149_989.n2 a_6149_989.t5 454.685
R2830 a_6149_989.n4 a_6149_989.t7 454.685
R2831 a_6149_989.n0 a_6149_989.t10 454.685
R2832 a_6149_989.n2 a_6149_989.t12 428.979
R2833 a_6149_989.n4 a_6149_989.t13 428.979
R2834 a_6149_989.n0 a_6149_989.t8 428.979
R2835 a_6149_989.n11 a_6149_989.n10 348.963
R2836 a_6149_989.n3 a_6149_989.t11 339.542
R2837 a_6149_989.n5 a_6149_989.t9 339.542
R2838 a_6149_989.n1 a_6149_989.t6 339.542
R2839 a_6149_989.n13 a_6149_989.n12 157.964
R2840 a_6149_989.n3 a_6149_989.n2 143.429
R2841 a_6149_989.n5 a_6149_989.n4 143.429
R2842 a_6149_989.n1 a_6149_989.n0 143.429
R2843 a_6149_989.n13 a_6149_989.n11 132.141
R2844 a_6149_989.n14 a_6149_989.n13 91.705
R2845 a_6149_989.n10 a_6149_989.n8 22.578
R2846 a_6149_989.n12 a_6149_989.t3 14.282
R2847 a_6149_989.n12 a_6149_989.t4 14.282
R2848 a_6149_989.n14 a_6149_989.t1 14.282
R2849 a_6149_989.t2 a_6149_989.n14 14.282
R2850 a_6149_989.n7 a_6149_989.n1 10.046
R2851 a_6149_989.n10 a_6149_989.n9 8.58
R2852 a_6149_989.n6 a_6149_989.n5 8.141
R2853 a_6149_989.n6 a_6149_989.n3 4.65
R2854 a_6149_989.n11 a_6149_989.n7 4.65
R2855 a_6149_989.n7 a_6149_989.n6 2.947
R2856 a_11033_989.n2 a_11033_989.t6 454.685
R2857 a_11033_989.n4 a_11033_989.t11 454.685
R2858 a_11033_989.n0 a_11033_989.t13 454.685
R2859 a_11033_989.n2 a_11033_989.t5 428.979
R2860 a_11033_989.n4 a_11033_989.t7 428.979
R2861 a_11033_989.n0 a_11033_989.t9 428.979
R2862 a_11033_989.n3 a_11033_989.t12 339.542
R2863 a_11033_989.n5 a_11033_989.t10 339.542
R2864 a_11033_989.n1 a_11033_989.t8 339.542
R2865 a_11033_989.n12 a_11033_989.n11 333.44
R2866 a_11033_989.n14 a_11033_989.n13 157.964
R2867 a_11033_989.n3 a_11033_989.n2 143.429
R2868 a_11033_989.n5 a_11033_989.n4 143.429
R2869 a_11033_989.n1 a_11033_989.n0 143.429
R2870 a_11033_989.n14 a_11033_989.n12 132.141
R2871 a_11033_989.n15 a_11033_989.n14 91.705
R2872 a_11033_989.n11 a_11033_989.n10 30
R2873 a_11033_989.n9 a_11033_989.n8 24.383
R2874 a_11033_989.n11 a_11033_989.n9 23.684
R2875 a_11033_989.n13 a_11033_989.t0 14.282
R2876 a_11033_989.n13 a_11033_989.t1 14.282
R2877 a_11033_989.n15 a_11033_989.t3 14.282
R2878 a_11033_989.t4 a_11033_989.n15 14.282
R2879 a_11033_989.n7 a_11033_989.n1 10.046
R2880 a_11033_989.n6 a_11033_989.n5 8.141
R2881 a_11033_989.n6 a_11033_989.n3 4.65
R2882 a_11033_989.n12 a_11033_989.n7 4.65
R2883 a_11033_989.n7 a_11033_989.n6 2.947
R2884 a_11673_1050.n0 a_11673_1050.t7 480.392
R2885 a_11673_1050.n0 a_11673_1050.t9 403.272
R2886 a_11673_1050.n1 a_11673_1050.t8 301.486
R2887 a_11673_1050.n6 a_11673_1050.n5 252.498
R2888 a_11673_1050.n10 a_11673_1050.n6 234.917
R2889 a_11673_1050.n1 a_11673_1050.n0 227.006
R2890 a_11673_1050.n9 a_11673_1050.n8 161.352
R2891 a_11673_1050.n9 a_11673_1050.n7 95.095
R2892 a_11673_1050.n11 a_11673_1050.n10 95.094
R2893 a_11673_1050.n10 a_11673_1050.n9 66.258
R2894 a_11673_1050.n5 a_11673_1050.n4 30
R2895 a_11673_1050.n3 a_11673_1050.n2 24.383
R2896 a_11673_1050.n5 a_11673_1050.n3 23.684
R2897 a_11673_1050.n7 a_11673_1050.t1 14.282
R2898 a_11673_1050.n7 a_11673_1050.t0 14.282
R2899 a_11673_1050.n8 a_11673_1050.t6 14.282
R2900 a_11673_1050.n8 a_11673_1050.t5 14.282
R2901 a_11673_1050.t4 a_11673_1050.n11 14.282
R2902 a_11673_1050.n11 a_11673_1050.t3 14.282
R2903 a_11673_1050.n6 a_11673_1050.n1 10.615
R2904 a_2702_101.n3 a_2702_101.n1 42.788
R2905 a_2702_101.t0 a_2702_101.n0 8.137
R2906 a_2702_101.n3 a_2702_101.n2 4.665
R2907 a_2702_101.t0 a_2702_101.n3 0.06
R2908 a_9178_210.n10 a_9178_210.n8 171.558
R2909 a_9178_210.n8 a_9178_210.t1 75.764
R2910 a_9178_210.n11 a_9178_210.n0 49.6
R2911 a_9178_210.n3 a_9178_210.n2 27.476
R2912 a_9178_210.n10 a_9178_210.n9 27.2
R2913 a_9178_210.n11 a_9178_210.n10 22.4
R2914 a_9178_210.t1 a_9178_210.n5 20.241
R2915 a_9178_210.n7 a_9178_210.n6 19.952
R2916 a_9178_210.t1 a_9178_210.n3 13.984
R2917 a_9178_210.n5 a_9178_210.n4 13.494
R2918 a_9178_210.t1 a_9178_210.n1 7.04
R2919 a_9178_210.n8 a_9178_210.n7 1.505
R2920 a_8252_101.n3 a_8252_101.n1 42.788
R2921 a_8252_101.t0 a_8252_101.n0 8.137
R2922 a_8252_101.n3 a_8252_101.n2 4.665
R2923 a_8252_101.t0 a_8252_101.n3 0.06
R2924 a_13241_1050.n0 a_13241_1050.t5 512.525
R2925 a_13241_1050.n1 a_13241_1050.t7 445.142
R2926 a_13241_1050.n6 a_13241_1050.n5 389.157
R2927 a_13241_1050.n0 a_13241_1050.t6 371.139
R2928 a_13241_1050.n8 a_13241_1050.n7 157.964
R2929 a_13241_1050.n9 a_13241_1050.n8 91.705
R2930 a_13241_1050.n1 a_13241_1050.n0 85.101
R2931 a_13241_1050.n8 a_13241_1050.n6 76.423
R2932 a_13241_1050.n5 a_13241_1050.n4 30
R2933 a_13241_1050.n3 a_13241_1050.n2 24.383
R2934 a_13241_1050.n5 a_13241_1050.n3 23.684
R2935 a_13241_1050.n7 a_13241_1050.t3 14.282
R2936 a_13241_1050.n7 a_13241_1050.t4 14.282
R2937 a_13241_1050.n9 a_13241_1050.t1 14.282
R2938 a_13241_1050.t2 a_13241_1050.n9 14.282
R2939 a_13241_1050.n6 a_13241_1050.n1 8.044
R2940 SN.n14 SN.t16 479.223
R2941 SN.n11 SN.t7 479.223
R2942 SN.n8 SN.t8 479.223
R2943 SN.n5 SN.t15 479.223
R2944 SN.n2 SN.t4 479.223
R2945 SN.n0 SN.t3 479.223
R2946 SN.n14 SN.t9 375.52
R2947 SN.n11 SN.t17 375.52
R2948 SN.n8 SN.t10 375.52
R2949 SN.n5 SN.t2 375.52
R2950 SN.n2 SN.t13 375.52
R2951 SN.n0 SN.t12 375.52
R2952 SN.n15 SN.n14 252.188
R2953 SN.n12 SN.n11 252.188
R2954 SN.n9 SN.n8 252.188
R2955 SN.n6 SN.n5 252.188
R2956 SN.n3 SN.n2 252.188
R2957 SN.n1 SN.n0 252.188
R2958 SN.n15 SN.t14 231.854
R2959 SN.n12 SN.t1 231.854
R2960 SN.n9 SN.t0 231.854
R2961 SN.n6 SN.t6 231.854
R2962 SN.n3 SN.t5 231.854
R2963 SN.n1 SN.t11 231.854
R2964 SN.n4 SN.n1 13.038
R2965 SN.n7 SN.n4 9.476
R2966 SN.n13 SN.n10 9.476
R2967 SN.n10 SN.n7 8.388
R2968 SN.n16 SN.n13 8.388
R2969 SN.n4 SN.n3 4.65
R2970 SN.n7 SN.n6 4.65
R2971 SN.n10 SN.n9 4.65
R2972 SN.n13 SN.n12 4.65
R2973 SN.n16 SN.n15 4.65
R2974 SN.n16 SN 0.046
R2975 a_6603_103.n5 a_6603_103.n4 66.708
R2976 a_6603_103.n2 a_6603_103.n0 32.662
R2977 a_6603_103.n5 a_6603_103.n3 19.496
R2978 a_6603_103.t0 a_6603_103.n5 13.756
R2979 a_6603_103.t0 a_6603_103.n2 3.034
R2980 a_6603_103.n2 a_6603_103.n1 0.443
R2981 a_6884_210.n10 a_6884_210.n8 171.558
R2982 a_6884_210.n8 a_6884_210.t1 75.764
R2983 a_6884_210.n11 a_6884_210.n0 49.6
R2984 a_6884_210.n3 a_6884_210.n2 27.476
R2985 a_6884_210.n10 a_6884_210.n9 27.2
R2986 a_6884_210.n11 a_6884_210.n10 22.4
R2987 a_6884_210.t1 a_6884_210.n5 20.241
R2988 a_6884_210.n7 a_6884_210.n6 19.952
R2989 a_6884_210.t1 a_6884_210.n3 13.984
R2990 a_6884_210.n5 a_6884_210.n4 13.494
R2991 a_6884_210.t1 a_6884_210.n1 7.04
R2992 a_6884_210.n8 a_6884_210.n7 1.505
R2993 a_13136_101.n3 a_13136_101.n1 42.788
R2994 a_13136_101.t0 a_13136_101.n0 8.137
R2995 a_13136_101.n3 a_13136_101.n2 4.665
R2996 a_13136_101.t0 a_13136_101.n3 0.06
R2997 a_4013_103.t0 a_4013_103.n7 59.616
R2998 a_4013_103.n4 a_4013_103.n2 54.496
R2999 a_4013_103.n4 a_4013_103.n3 54.496
R3000 a_4013_103.n1 a_4013_103.n0 24.679
R3001 a_4013_103.n6 a_4013_103.n4 7.859
R3002 a_4013_103.t0 a_4013_103.n1 7.505
R3003 a_4013_103.t0 a_4013_103.n6 3.034
R3004 a_4013_103.n6 a_4013_103.n5 0.443
R3005 a_4294_210.n8 a_4294_210.n6 185.173
R3006 a_4294_210.t0 a_4294_210.n8 75.765
R3007 a_4294_210.n3 a_4294_210.n1 74.827
R3008 a_4294_210.n3 a_4294_210.n2 27.476
R3009 a_4294_210.n6 a_4294_210.n5 22.349
R3010 a_4294_210.t0 a_4294_210.n10 20.241
R3011 a_4294_210.t0 a_4294_210.n3 13.984
R3012 a_4294_210.n10 a_4294_210.n9 13.494
R3013 a_4294_210.n6 a_4294_210.n4 8.443
R3014 a_4294_210.t0 a_4294_210.n0 8.137
R3015 a_4294_210.n8 a_4294_210.n7 1.505
R3016 a_343_411.n0 a_343_411.t12 480.392
R3017 a_343_411.n2 a_343_411.t7 472.359
R3018 a_343_411.n1 a_343_411.t9 412.921
R3019 a_343_411.n0 a_343_411.t8 403.272
R3020 a_343_411.n2 a_343_411.t10 384.527
R3021 a_343_411.n3 a_343_411.t11 370.613
R3022 a_343_411.n9 a_343_411.n8 363.578
R3023 a_343_411.n12 a_343_411.n11 161.352
R3024 a_343_411.n3 a_343_411.n2 127.096
R3025 a_343_411.n13 a_343_411.n9 123.126
R3026 a_343_411.n1 a_343_411.n0 115.571
R3027 a_343_411.n12 a_343_411.n10 95.095
R3028 a_343_411.n14 a_343_411.n13 95.094
R3029 a_343_411.n13 a_343_411.n12 66.258
R3030 a_343_411.n8 a_343_411.n7 30
R3031 a_343_411.n6 a_343_411.n5 24.383
R3032 a_343_411.n8 a_343_411.n6 23.684
R3033 a_343_411.n10 a_343_411.t6 14.282
R3034 a_343_411.n10 a_343_411.t5 14.282
R3035 a_343_411.n11 a_343_411.t4 14.282
R3036 a_343_411.n11 a_343_411.t3 14.282
R3037 a_343_411.t2 a_343_411.n14 14.282
R3038 a_343_411.n14 a_343_411.t1 14.282
R3039 a_343_411.n4 a_343_411.n1 11.954
R3040 a_343_411.n4 a_343_411.n3 8.682
R3041 a_343_411.n9 a_343_411.n4 4.65
R3042 a_11487_103.t0 a_11487_103.n7 59.616
R3043 a_11487_103.n4 a_11487_103.n2 54.496
R3044 a_11487_103.n4 a_11487_103.n3 54.496
R3045 a_11487_103.n1 a_11487_103.n0 24.679
R3046 a_11487_103.n6 a_11487_103.n4 7.859
R3047 a_11487_103.t0 a_11487_103.n1 7.505
R3048 a_11487_103.t0 a_11487_103.n6 3.034
R3049 a_11487_103.n6 a_11487_103.n5 0.443
R3050 a_3473_1050.n1 a_3473_1050.t5 512.525
R3051 a_3473_1050.n2 a_3473_1050.t7 417.109
R3052 a_3473_1050.n1 a_3473_1050.t6 371.139
R3053 a_3473_1050.n7 a_3473_1050.n6 361.298
R3054 a_3473_1050.n2 a_3473_1050.n1 179.837
R3055 a_3473_1050.n9 a_3473_1050.n8 157.963
R3056 a_3473_1050.n8 a_3473_1050.n7 104.282
R3057 a_3473_1050.n8 a_3473_1050.n0 91.706
R3058 a_3473_1050.n6 a_3473_1050.n5 30
R3059 a_3473_1050.n4 a_3473_1050.n3 24.383
R3060 a_3473_1050.n6 a_3473_1050.n4 23.684
R3061 a_3473_1050.n0 a_3473_1050.t3 14.282
R3062 a_3473_1050.n0 a_3473_1050.t4 14.282
R3063 a_3473_1050.n9 a_3473_1050.t0 14.282
R3064 a_3473_1050.t1 a_3473_1050.n9 14.282
R3065 a_3473_1050.n7 a_3473_1050.n2 10.615
R3066 a_2000_210.n9 a_2000_210.n7 171.558
R3067 a_2000_210.t0 a_2000_210.n9 75.765
R3068 a_2000_210.n3 a_2000_210.n1 74.827
R3069 a_2000_210.n3 a_2000_210.n2 27.476
R3070 a_2000_210.n7 a_2000_210.n6 27.2
R3071 a_2000_210.n5 a_2000_210.n4 23.498
R3072 a_2000_210.n7 a_2000_210.n5 22.4
R3073 a_2000_210.t0 a_2000_210.n11 20.241
R3074 a_2000_210.t0 a_2000_210.n3 13.984
R3075 a_2000_210.n11 a_2000_210.n10 13.494
R3076 a_2000_210.t0 a_2000_210.n0 8.137
R3077 a_2000_210.n9 a_2000_210.n8 1.505
R3078 a_10806_210.n10 a_10806_210.n8 171.558
R3079 a_10806_210.n8 a_10806_210.t1 75.764
R3080 a_10806_210.n11 a_10806_210.n0 49.6
R3081 a_10806_210.n3 a_10806_210.n2 27.476
R3082 a_10806_210.n10 a_10806_210.n9 27.2
R3083 a_10806_210.n11 a_10806_210.n10 22.4
R3084 a_10806_210.t1 a_10806_210.n5 20.241
R3085 a_10806_210.n7 a_10806_210.n6 19.952
R3086 a_10806_210.t1 a_10806_210.n3 13.984
R3087 a_10806_210.n5 a_10806_210.n4 13.494
R3088 a_10806_210.t1 a_10806_210.n1 7.04
R3089 a_10806_210.n8 a_10806_210.n7 1.505
R3090 a_12470_101.n3 a_12470_101.n1 42.788
R3091 a_12470_101.t0 a_12470_101.n0 8.137
R3092 a_12470_101.n3 a_12470_101.n2 4.665
R3093 a_12470_101.t0 a_12470_101.n3 0.06
R3094 a_15430_101.n2 a_15430_101.n0 42.755
R3095 a_15430_101.n2 a_15430_101.n1 2.198
R3096 a_15430_101.t0 a_15430_101.n2 0.106
R3097 a_1038_210.n9 a_1038_210.n7 171.558
R3098 a_1038_210.t0 a_1038_210.n9 75.765
R3099 a_1038_210.n3 a_1038_210.n1 74.827
R3100 a_1038_210.n3 a_1038_210.n2 27.476
R3101 a_1038_210.n7 a_1038_210.n6 27.2
R3102 a_1038_210.n5 a_1038_210.n4 23.498
R3103 a_1038_210.n7 a_1038_210.n5 22.4
R3104 a_1038_210.t0 a_1038_210.n11 20.241
R3105 a_1038_210.t0 a_1038_210.n3 13.984
R3106 a_1038_210.n11 a_1038_210.n10 13.494
R3107 a_1038_210.t0 a_1038_210.n0 8.137
R3108 a_1038_210.n9 a_1038_210.n8 1.505
R3109 a_14062_210.n10 a_14062_210.n8 171.558
R3110 a_14062_210.n8 a_14062_210.t1 75.764
R3111 a_14062_210.n3 a_14062_210.n2 27.476
R3112 a_14062_210.n10 a_14062_210.n9 27.2
R3113 a_14062_210.n11 a_14062_210.n0 23.498
R3114 a_14062_210.n11 a_14062_210.n10 22.4
R3115 a_14062_210.t1 a_14062_210.n5 20.241
R3116 a_14062_210.n7 a_14062_210.n6 19.952
R3117 a_14062_210.t1 a_14062_210.n3 13.984
R3118 a_14062_210.n5 a_14062_210.n4 13.494
R3119 a_14062_210.t1 a_14062_210.n1 7.04
R3120 a_14062_210.n8 a_14062_210.n7 1.505
R3121 a_11768_210.n10 a_11768_210.n8 171.558
R3122 a_11768_210.n8 a_11768_210.t1 75.764
R3123 a_11768_210.n11 a_11768_210.n0 49.6
R3124 a_11768_210.n3 a_11768_210.n2 27.476
R3125 a_11768_210.n10 a_11768_210.n9 27.2
R3126 a_11768_210.n11 a_11768_210.n10 22.4
R3127 a_11768_210.t1 a_11768_210.n5 20.241
R3128 a_11768_210.n7 a_11768_210.n6 19.952
R3129 a_11768_210.t1 a_11768_210.n3 13.984
R3130 a_11768_210.n5 a_11768_210.n4 13.494
R3131 a_11768_210.t1 a_11768_210.n1 7.04
R3132 a_11768_210.n8 a_11768_210.n7 1.505
R3133 a_757_103.n5 a_757_103.n4 66.708
R3134 a_757_103.n2 a_757_103.n0 25.439
R3135 a_757_103.n5 a_757_103.n3 19.496
R3136 a_757_103.t0 a_757_103.n5 13.756
R3137 a_757_103.n2 a_757_103.n1 2.455
R3138 a_757_103.t0 a_757_103.n2 0.246
R3139 a_5922_210.n10 a_5922_210.n8 171.558
R3140 a_5922_210.n8 a_5922_210.t1 75.764
R3141 a_5922_210.n3 a_5922_210.n2 27.476
R3142 a_5922_210.n10 a_5922_210.n9 27.2
R3143 a_5922_210.n11 a_5922_210.n0 23.498
R3144 a_5922_210.n11 a_5922_210.n10 22.4
R3145 a_5922_210.t1 a_5922_210.n5 20.241
R3146 a_5922_210.n7 a_5922_210.n6 19.952
R3147 a_5922_210.t1 a_5922_210.n3 13.984
R3148 a_5922_210.n5 a_5922_210.n4 13.494
R3149 a_5922_210.t1 a_5922_210.n1 7.04
R3150 a_5922_210.n8 a_5922_210.n7 1.505
R3151 a_112_101.n3 a_112_101.n1 42.788
R3152 a_112_101.t0 a_112_101.n0 8.137
R3153 a_112_101.n3 a_112_101.n2 4.665
R3154 a_112_101.t0 a_112_101.n3 0.06
R3155 Q.n2 Q.n1 349.908
R3156 Q.n2 Q.n0 215.564
R3157 Q.n0 Q.t2 14.282
R3158 Q.n0 Q.t1 14.282
R3159 Q.n3 Q.n2 4.65
R3160 Q.n3 Q 0.046
R3161 a_8897_103.n5 a_8897_103.n4 66.708
R3162 a_8897_103.n2 a_8897_103.n0 25.439
R3163 a_8897_103.n5 a_8897_103.n3 19.496
R3164 a_8897_103.t0 a_8897_103.n5 13.756
R3165 a_8897_103.n2 a_8897_103.n1 2.455
R3166 a_8897_103.t0 a_8897_103.n2 0.246
R3167 a_3368_101.n11 a_3368_101.n10 68.43
R3168 a_3368_101.n3 a_3368_101.n2 62.817
R3169 a_3368_101.n7 a_3368_101.n6 38.626
R3170 a_3368_101.n6 a_3368_101.n5 35.955
R3171 a_3368_101.n3 a_3368_101.n1 26.202
R3172 a_3368_101.t0 a_3368_101.n3 19.737
R3173 a_3368_101.t1 a_3368_101.n8 8.137
R3174 a_3368_101.t0 a_3368_101.n4 7.273
R3175 a_3368_101.t0 a_3368_101.n0 6.109
R3176 a_3368_101.t1 a_3368_101.n7 4.864
R3177 a_3368_101.t0 a_3368_101.n12 2.074
R3178 a_3368_101.n12 a_3368_101.t1 0.937
R3179 a_3368_101.t1 a_3368_101.n11 0.763
R3180 a_3368_101.n11 a_3368_101.n9 0.185
R3181 a_9880_101.n11 a_9880_101.n10 68.43
R3182 a_9880_101.n3 a_9880_101.n2 62.817
R3183 a_9880_101.n7 a_9880_101.n6 38.626
R3184 a_9880_101.n6 a_9880_101.n5 35.955
R3185 a_9880_101.n3 a_9880_101.n1 26.202
R3186 a_9880_101.t0 a_9880_101.n3 19.737
R3187 a_9880_101.t1 a_9880_101.n8 8.137
R3188 a_9880_101.t0 a_9880_101.n4 7.273
R3189 a_9880_101.t0 a_9880_101.n0 6.109
R3190 a_9880_101.t1 a_9880_101.n7 4.864
R3191 a_9880_101.t0 a_9880_101.n12 2.074
R3192 a_9880_101.n12 a_9880_101.t1 0.937
R3193 a_9880_101.t1 a_9880_101.n11 0.763
R3194 a_9880_101.n11 a_9880_101.n9 0.185
R3195 a_1719_103.n5 a_1719_103.n4 66.708
R3196 a_1719_103.n2 a_1719_103.n0 25.439
R3197 a_1719_103.n5 a_1719_103.n3 19.496
R3198 a_1719_103.t0 a_1719_103.n5 13.756
R3199 a_1719_103.n2 a_1719_103.n1 2.455
R3200 a_1719_103.t0 a_1719_103.n2 0.246
R3201 a_13781_103.n5 a_13781_103.n4 66.708
R3202 a_13781_103.n2 a_13781_103.n0 25.439
R3203 a_13781_103.n5 a_13781_103.n3 19.496
R3204 a_13781_103.t0 a_13781_103.n5 13.756
R3205 a_13781_103.n2 a_13781_103.n1 2.455
R3206 a_13781_103.t0 a_13781_103.n2 0.246
R3207 a_5641_103.t0 a_5641_103.n7 59.616
R3208 a_5641_103.n4 a_5641_103.n2 54.496
R3209 a_5641_103.n4 a_5641_103.n3 54.496
R3210 a_5641_103.n1 a_5641_103.n0 24.679
R3211 a_5641_103.t0 a_5641_103.n1 7.505
R3212 a_5641_103.n6 a_5641_103.n5 2.455
R3213 a_5641_103.n6 a_5641_103.n4 0.636
R3214 a_5641_103.t0 a_5641_103.n6 0.246
R3215 a_14764_101.n3 a_14764_101.n2 62.817
R3216 a_14764_101.n11 a_14764_101.n10 46.054
R3217 a_14764_101.n7 a_14764_101.n6 38.626
R3218 a_14764_101.n6 a_14764_101.n5 35.955
R3219 a_14764_101.n12 a_14764_101.n11 27.923
R3220 a_14764_101.n3 a_14764_101.n1 26.202
R3221 a_14764_101.t0 a_14764_101.n3 19.737
R3222 a_14764_101.t0 a_14764_101.n4 7.273
R3223 a_14764_101.n9 a_14764_101.n8 6.883
R3224 a_14764_101.t0 a_14764_101.n0 6.109
R3225 a_14764_101.t1 a_14764_101.n7 4.864
R3226 a_14764_101.t0 a_14764_101.n13 2.074
R3227 a_14764_101.t1 a_14764_101.n9 1.179
R3228 a_14764_101.t1 a_14764_101.n12 0.958
R3229 a_14764_101.n13 a_14764_101.t1 0.937
C7 SN GND 6.35fF
C8 VDD GND 27.71fF
C9 a_14764_101.n0 GND 0.02fF
C10 a_14764_101.n1 GND 0.09fF
C11 a_14764_101.n2 GND 0.07fF
C12 a_14764_101.n3 GND 0.03fF
C13 a_14764_101.n4 GND 0.01fF
C14 a_14764_101.n5 GND 0.03fF
C15 a_14764_101.n6 GND 0.04fF
C16 a_14764_101.n7 GND 0.02fF
C17 a_14764_101.n8 GND 0.04fF
C18 a_14764_101.n9 GND 0.08fF
C19 a_14764_101.n10 GND 0.04fF
C20 a_14764_101.n11 GND 0.12fF
C21 a_14764_101.n12 GND 0.14fF
C22 a_14764_101.t1 GND 0.16fF
C23 a_14764_101.n13 GND 0.01fF
C24 a_5641_103.n0 GND 0.08fF
C25 a_5641_103.n1 GND 0.07fF
C26 a_5641_103.n2 GND 0.04fF
C27 a_5641_103.n3 GND 0.06fF
C28 a_5641_103.n4 GND 0.03fF
C29 a_5641_103.n5 GND 0.04fF
C30 a_5641_103.n7 GND 0.08fF
C31 a_13781_103.n0 GND 0.11fF
C32 a_13781_103.n1 GND 0.04fF
C33 a_13781_103.n2 GND 0.03fF
C34 a_13781_103.n3 GND 0.07fF
C35 a_13781_103.n4 GND 0.08fF
C36 a_13781_103.n5 GND 0.03fF
C37 a_1719_103.n0 GND 0.11fF
C38 a_1719_103.n1 GND 0.04fF
C39 a_1719_103.n2 GND 0.03fF
C40 a_1719_103.n3 GND 0.07fF
C41 a_1719_103.n4 GND 0.08fF
C42 a_1719_103.n5 GND 0.03fF
C43 a_9880_101.n0 GND 0.02fF
C44 a_9880_101.n1 GND 0.09fF
C45 a_9880_101.n2 GND 0.08fF
C46 a_9880_101.n3 GND 0.03fF
C47 a_9880_101.n4 GND 0.01fF
C48 a_9880_101.n5 GND 0.04fF
C49 a_9880_101.n6 GND 0.04fF
C50 a_9880_101.n7 GND 0.02fF
C51 a_9880_101.n8 GND 0.05fF
C52 a_9880_101.n9 GND 0.15fF
C53 a_9880_101.n10 GND 0.08fF
C54 a_9880_101.n11 GND 0.08fF
C55 a_9880_101.t1 GND 0.23fF
C56 a_9880_101.n12 GND 0.01fF
C57 a_3368_101.n0 GND 0.02fF
C58 a_3368_101.n1 GND 0.09fF
C59 a_3368_101.n2 GND 0.08fF
C60 a_3368_101.n3 GND 0.03fF
C61 a_3368_101.n4 GND 0.01fF
C62 a_3368_101.n5 GND 0.04fF
C63 a_3368_101.n6 GND 0.04fF
C64 a_3368_101.n7 GND 0.02fF
C65 a_3368_101.n8 GND 0.05fF
C66 a_3368_101.n9 GND 0.15fF
C67 a_3368_101.n10 GND 0.08fF
C68 a_3368_101.n11 GND 0.08fF
C69 a_3368_101.t1 GND 0.23fF
C70 a_3368_101.n12 GND 0.01fF
C71 a_8897_103.n0 GND 0.11fF
C72 a_8897_103.n1 GND 0.04fF
C73 a_8897_103.n2 GND 0.03fF
C74 a_8897_103.n3 GND 0.07fF
C75 a_8897_103.n4 GND 0.08fF
C76 a_8897_103.n5 GND 0.03fF
C77 Q.n0 GND 0.58fF
C78 Q.n1 GND 0.36fF
C79 Q.n2 GND 0.66fF
C80 Q.n3 GND 0.01fF
C81 a_112_101.n0 GND 0.05fF
C82 a_112_101.n1 GND 0.12fF
C83 a_112_101.n2 GND 0.04fF
C84 a_112_101.n3 GND 0.16fF
C85 a_5922_210.n0 GND 0.02fF
C86 a_5922_210.n1 GND 0.09fF
C87 a_5922_210.n2 GND 0.12fF
C88 a_5922_210.n3 GND 0.08fF
C89 a_5922_210.n4 GND 0.08fF
C90 a_5922_210.n5 GND 0.02fF
C91 a_5922_210.t1 GND 0.29fF
C92 a_5922_210.n6 GND 0.09fF
C93 a_5922_210.n7 GND 0.02fF
C94 a_5922_210.n8 GND 0.13fF
C95 a_5922_210.n9 GND 0.02fF
C96 a_5922_210.n10 GND 0.03fF
C97 a_5922_210.n11 GND 0.03fF
C98 a_757_103.n0 GND 0.11fF
C99 a_757_103.n1 GND 0.04fF
C100 a_757_103.n2 GND 0.03fF
C101 a_757_103.n3 GND 0.07fF
C102 a_757_103.n4 GND 0.08fF
C103 a_757_103.n5 GND 0.03fF
C104 a_11768_210.n0 GND 0.02fF
C105 a_11768_210.n1 GND 0.09fF
C106 a_11768_210.n2 GND 0.12fF
C107 a_11768_210.n3 GND 0.08fF
C108 a_11768_210.n4 GND 0.08fF
C109 a_11768_210.n5 GND 0.02fF
C110 a_11768_210.t1 GND 0.29fF
C111 a_11768_210.n6 GND 0.09fF
C112 a_11768_210.n7 GND 0.02fF
C113 a_11768_210.n8 GND 0.13fF
C114 a_11768_210.n9 GND 0.02fF
C115 a_11768_210.n10 GND 0.03fF
C116 a_11768_210.n11 GND 0.02fF
C117 a_14062_210.n0 GND 0.02fF
C118 a_14062_210.n1 GND 0.09fF
C119 a_14062_210.n2 GND 0.12fF
C120 a_14062_210.n3 GND 0.08fF
C121 a_14062_210.n4 GND 0.08fF
C122 a_14062_210.n5 GND 0.02fF
C123 a_14062_210.t1 GND 0.29fF
C124 a_14062_210.n6 GND 0.09fF
C125 a_14062_210.n7 GND 0.02fF
C126 a_14062_210.n8 GND 0.13fF
C127 a_14062_210.n9 GND 0.02fF
C128 a_14062_210.n10 GND 0.03fF
C129 a_14062_210.n11 GND 0.03fF
C130 a_1038_210.n0 GND 0.07fF
C131 a_1038_210.n1 GND 0.09fF
C132 a_1038_210.n2 GND 0.12fF
C133 a_1038_210.n3 GND 0.08fF
C134 a_1038_210.n4 GND 0.02fF
C135 a_1038_210.n5 GND 0.03fF
C136 a_1038_210.n6 GND 0.02fF
C137 a_1038_210.n7 GND 0.03fF
C138 a_1038_210.n8 GND 0.02fF
C139 a_1038_210.n9 GND 0.13fF
C140 a_1038_210.n10 GND 0.08fF
C141 a_1038_210.n11 GND 0.02fF
C142 a_1038_210.t0 GND 0.31fF
C143 a_15430_101.n0 GND 0.13fF
C144 a_15430_101.n1 GND 0.14fF
C145 a_15430_101.n2 GND 0.14fF
C146 a_12470_101.n0 GND 0.05fF
C147 a_12470_101.n1 GND 0.12fF
C148 a_12470_101.n2 GND 0.04fF
C149 a_12470_101.n3 GND 0.17fF
C150 a_10806_210.n0 GND 0.02fF
C151 a_10806_210.n1 GND 0.09fF
C152 a_10806_210.n2 GND 0.12fF
C153 a_10806_210.n3 GND 0.08fF
C154 a_10806_210.n4 GND 0.08fF
C155 a_10806_210.n5 GND 0.02fF
C156 a_10806_210.t1 GND 0.29fF
C157 a_10806_210.n6 GND 0.09fF
C158 a_10806_210.n7 GND 0.02fF
C159 a_10806_210.n8 GND 0.13fF
C160 a_10806_210.n9 GND 0.02fF
C161 a_10806_210.n10 GND 0.03fF
C162 a_10806_210.n11 GND 0.02fF
C163 a_2000_210.n0 GND 0.07fF
C164 a_2000_210.n1 GND 0.09fF
C165 a_2000_210.n2 GND 0.12fF
C166 a_2000_210.n3 GND 0.08fF
C167 a_2000_210.n4 GND 0.02fF
C168 a_2000_210.n5 GND 0.03fF
C169 a_2000_210.n6 GND 0.02fF
C170 a_2000_210.n7 GND 0.03fF
C171 a_2000_210.n8 GND 0.02fF
C172 a_2000_210.n9 GND 0.13fF
C173 a_2000_210.n10 GND 0.08fF
C174 a_2000_210.n11 GND 0.02fF
C175 a_2000_210.t0 GND 0.31fF
C176 a_3473_1050.n0 GND 0.40fF
C177 a_3473_1050.n1 GND 0.29fF
C178 a_3473_1050.n2 GND 0.67fF
C179 a_3473_1050.n3 GND 0.04fF
C180 a_3473_1050.n4 GND 0.06fF
C181 a_3473_1050.n5 GND 0.04fF
C182 a_3473_1050.n6 GND 0.29fF
C183 a_3473_1050.n7 GND 0.70fF
C184 a_3473_1050.n8 GND 0.53fF
C185 a_3473_1050.n9 GND 0.51fF
C186 a_11487_103.n0 GND 0.08fF
C187 a_11487_103.n1 GND 0.07fF
C188 a_11487_103.n2 GND 0.04fF
C189 a_11487_103.n3 GND 0.06fF
C190 a_11487_103.n4 GND 0.11fF
C191 a_11487_103.n5 GND 0.04fF
C192 a_11487_103.n7 GND 0.08fF
C193 a_343_411.n0 GND 0.41fF
C194 a_343_411.n1 GND 1.38fF
C195 a_343_411.n2 GND 0.40fF
C196 a_343_411.t11 GND 0.84fF
C197 a_343_411.n3 GND 0.89fF
C198 a_343_411.n4 GND 2.70fF
C199 a_343_411.n5 GND 0.06fF
C200 a_343_411.n6 GND 0.08fF
C201 a_343_411.n7 GND 0.05fF
C202 a_343_411.n8 GND 0.41fF
C203 a_343_411.n9 GND 0.77fF
C204 a_343_411.n10 GND 0.57fF
C205 a_343_411.n11 GND 0.72fF
C206 a_343_411.n12 GND 0.69fF
C207 a_343_411.n13 GND 0.56fF
C208 a_343_411.n14 GND 0.57fF
C209 a_4294_210.n0 GND 0.07fF
C210 a_4294_210.n1 GND 0.09fF
C211 a_4294_210.n2 GND 0.12fF
C212 a_4294_210.n3 GND 0.08fF
C213 a_4294_210.n4 GND 0.02fF
C214 a_4294_210.n5 GND 0.03fF
C215 a_4294_210.n6 GND 0.05fF
C216 a_4294_210.n7 GND 0.02fF
C217 a_4294_210.n8 GND 0.14fF
C218 a_4294_210.n9 GND 0.08fF
C219 a_4294_210.n10 GND 0.02fF
C220 a_4294_210.t0 GND 0.31fF
C221 a_4013_103.n0 GND 0.08fF
C222 a_4013_103.n1 GND 0.07fF
C223 a_4013_103.n2 GND 0.04fF
C224 a_4013_103.n3 GND 0.06fF
C225 a_4013_103.n4 GND 0.11fF
C226 a_4013_103.n5 GND 0.04fF
C227 a_4013_103.n7 GND 0.08fF
C228 a_13136_101.n0 GND 0.05fF
C229 a_13136_101.n1 GND 0.12fF
C230 a_13136_101.n2 GND 0.04fF
C231 a_13136_101.n3 GND 0.17fF
C232 a_6884_210.n0 GND 0.02fF
C233 a_6884_210.n1 GND 0.09fF
C234 a_6884_210.n2 GND 0.12fF
C235 a_6884_210.n3 GND 0.08fF
C236 a_6884_210.n4 GND 0.08fF
C237 a_6884_210.n5 GND 0.02fF
C238 a_6884_210.t1 GND 0.29fF
C239 a_6884_210.n6 GND 0.09fF
C240 a_6884_210.n7 GND 0.02fF
C241 a_6884_210.n8 GND 0.13fF
C242 a_6884_210.n9 GND 0.02fF
C243 a_6884_210.n10 GND 0.03fF
C244 a_6884_210.n11 GND 0.02fF
C245 a_6603_103.n0 GND 0.13fF
C246 a_6603_103.n1 GND 0.04fF
C247 a_6603_103.n2 GND 0.09fF
C248 a_6603_103.n3 GND 0.07fF
C249 a_6603_103.n4 GND 0.08fF
C250 a_6603_103.n5 GND 0.03fF
C251 SN.n0 GND 0.76fF
C252 SN.t11 GND 0.83fF
C253 SN.n1 GND 1.82fF
C254 SN.n2 GND 0.76fF
C255 SN.t5 GND 0.83fF
C256 SN.n3 GND 0.71fF
C257 SN.n4 GND 4.21fF
C258 SN.n5 GND 0.76fF
C259 SN.t6 GND 0.83fF
C260 SN.n6 GND 0.71fF
C261 SN.n7 GND 3.60fF
C262 SN.n8 GND 0.76fF
C263 SN.t0 GND 0.83fF
C264 SN.n9 GND 0.71fF
C265 SN.n10 GND 3.60fF
C266 SN.n11 GND 0.76fF
C267 SN.t1 GND 0.83fF
C268 SN.n12 GND 0.71fF
C269 SN.n13 GND 3.60fF
C270 SN.n14 GND 0.76fF
C271 SN.t14 GND 0.83fF
C272 SN.n15 GND 0.71fF
C273 SN.n16 GND 1.71fF
C274 a_13241_1050.n0 GND 0.22fF
C275 a_13241_1050.n1 GND 0.70fF
C276 a_13241_1050.n2 GND 0.04fF
C277 a_13241_1050.n3 GND 0.05fF
C278 a_13241_1050.n4 GND 0.03fF
C279 a_13241_1050.n5 GND 0.30fF
C280 a_13241_1050.n6 GND 0.59fF
C281 a_13241_1050.n7 GND 0.47fF
C282 a_13241_1050.n8 GND 0.46fF
C283 a_13241_1050.n9 GND 0.36fF
C284 a_8252_101.n0 GND 0.05fF
C285 a_8252_101.n1 GND 0.12fF
C286 a_8252_101.n2 GND 0.04fF
C287 a_8252_101.n3 GND 0.17fF
C288 a_9178_210.n0 GND 0.02fF
C289 a_9178_210.n1 GND 0.09fF
C290 a_9178_210.n2 GND 0.12fF
C291 a_9178_210.n3 GND 0.08fF
C292 a_9178_210.n4 GND 0.08fF
C293 a_9178_210.n5 GND 0.02fF
C294 a_9178_210.t1 GND 0.29fF
C295 a_9178_210.n6 GND 0.09fF
C296 a_9178_210.n7 GND 0.02fF
C297 a_9178_210.n8 GND 0.13fF
C298 a_9178_210.n9 GND 0.02fF
C299 a_9178_210.n10 GND 0.03fF
C300 a_9178_210.n11 GND 0.02fF
C301 a_2702_101.n0 GND 0.05fF
C302 a_2702_101.n1 GND 0.12fF
C303 a_2702_101.n2 GND 0.04fF
C304 a_2702_101.n3 GND 0.17fF
C305 a_11673_1050.n0 GND 0.38fF
C306 a_11673_1050.n1 GND 0.59fF
C307 a_11673_1050.n2 GND 0.04fF
C308 a_11673_1050.n3 GND 0.05fF
C309 a_11673_1050.n4 GND 0.03fF
C310 a_11673_1050.n5 GND 0.17fF
C311 a_11673_1050.n6 GND 0.69fF
C312 a_11673_1050.n7 GND 0.39fF
C313 a_11673_1050.n8 GND 0.49fF
C314 a_11673_1050.n9 GND 0.47fF
C315 a_11673_1050.n10 GND 0.51fF
C316 a_11673_1050.n11 GND 0.39fF
C317 a_11033_989.n0 GND 0.52fF
C318 a_11033_989.t8 GND 0.94fF
C319 a_11033_989.n1 GND 1.27fF
C320 a_11033_989.n2 GND 0.52fF
C321 a_11033_989.t12 GND 0.93fF
C322 a_11033_989.n3 GND 0.70fF
C323 a_11033_989.n4 GND 0.52fF
C324 a_11033_989.t10 GND 0.94fF
C325 a_11033_989.n5 GND 1.00fF
C326 a_11033_989.n6 GND 1.65fF
C327 a_11033_989.n7 GND 2.09fF
C328 a_11033_989.n8 GND 0.07fF
C329 a_11033_989.n9 GND 0.09fF
C330 a_11033_989.n10 GND 0.06fF
C331 a_11033_989.n11 GND 0.43fF
C332 a_11033_989.n12 GND 0.84fF
C333 a_11033_989.n13 GND 0.84fF
C334 a_11033_989.n14 GND 0.93fF
C335 a_11033_989.n15 GND 0.65fF
C336 a_6149_989.n0 GND 0.46fF
C337 a_6149_989.t6 GND 0.83fF
C338 a_6149_989.n1 GND 1.13fF
C339 a_6149_989.n2 GND 0.46fF
C340 a_6149_989.t11 GND 0.83fF
C341 a_6149_989.n3 GND 0.62fF
C342 a_6149_989.n4 GND 0.46fF
C343 a_6149_989.t9 GND 0.83fF
C344 a_6149_989.n5 GND 0.89fF
C345 a_6149_989.n6 GND 1.46fF
C346 a_6149_989.n7 GND 1.85fF
C347 a_6149_989.n8 GND 0.11fF
C348 a_6149_989.n9 GND 0.04fF
C349 a_6149_989.n10 GND 0.41fF
C350 a_6149_989.n11 GND 0.77fF
C351 a_6149_989.n12 GND 0.74fF
C352 a_6149_989.n13 GND 0.82fF
C353 a_6149_989.n14 GND 0.58fF
C354 a_15044_209.n0 GND 0.26fF
C355 a_15044_209.n1 GND 0.24fF
C356 a_15044_209.n2 GND 0.47fF
C357 a_15044_209.n3 GND 0.03fF
C358 a_15044_209.n4 GND 0.04fF
C359 a_15044_209.n5 GND 0.03fF
C360 a_15044_209.n6 GND 0.03fF
C361 a_15044_209.n7 GND 0.03fF
C362 a_15044_209.n8 GND 0.04fF
C363 a_15044_209.n9 GND 0.03fF
C364 a_15044_209.n10 GND 0.04fF
C365 a_15044_209.n11 GND 0.94fF
C366 a_15044_209.n12 GND 0.12fF
C367 a_15044_209.n13 GND 0.34fF
C368 a_15044_209.n14 GND 0.43fF
C369 a_15044_209.n15 GND 0.41fF
C370 a_15044_209.n16 GND 0.34fF
C371 a_13367_411.n0 GND 0.05fF
C372 a_13367_411.n1 GND 0.45fF
C373 a_13367_411.n2 GND 0.45fF
C374 a_13367_411.n3 GND 0.57fF
C375 a_13367_411.n4 GND 0.54fF
C376 a_13367_411.n5 GND 0.44fF
C377 a_13367_411.n6 GND 0.33fF
C378 a_13367_411.t11 GND 0.66fF
C379 a_13367_411.n7 GND 0.82fF
C380 a_13367_411.n8 GND 0.32fF
C381 a_13367_411.t15 GND 0.66fF
C382 a_13367_411.n9 GND 0.44fF
C383 a_13367_411.n10 GND 1.19fF
C384 a_13367_411.n11 GND 0.32fF
C385 a_13367_411.t8 GND 0.66fF
C386 a_13367_411.n12 GND 0.70fF
C387 a_13367_411.n13 GND 1.06fF
C388 a_13367_411.n14 GND 0.60fF
C389 a_13367_411.n15 GND 0.05fF
C390 a_13367_411.n16 GND 0.33fF
C391 a_13367_411.n17 GND 0.05fF
C392 a_4996_101.n0 GND 0.05fF
C393 a_4996_101.n1 GND 0.12fF
C394 a_4996_101.n2 GND 0.04fF
C395 a_4996_101.n3 GND 0.17fF
C396 a_16096_101.n0 GND 0.06fF
C397 a_16096_101.n1 GND 0.13fF
C398 a_16096_101.n2 GND 0.04fF
C399 a_16096_101.n3 GND 0.19fF
C400 a_10525_103.n0 GND 0.08fF
C401 a_10525_103.n1 GND 0.07fF
C402 a_10525_103.n2 GND 0.04fF
C403 a_10525_103.n3 GND 0.06fF
C404 a_10525_103.n4 GND 0.11fF
C405 a_10525_103.n5 GND 0.04fF
C406 a_10525_103.n7 GND 0.08fF
C407 a_9985_1050.n0 GND 0.50fF
C408 a_9985_1050.n1 GND 0.49fF
C409 a_9985_1050.n2 GND 0.84fF
C410 a_9985_1050.n3 GND 0.49fF
C411 a_9985_1050.n4 GND 0.61fF
C412 a_9985_1050.n5 GND 1.21fF
C413 a_9985_1050.n6 GND 0.05fF
C414 a_9985_1050.n7 GND 0.07fF
C415 a_9985_1050.n8 GND 0.04fF
C416 a_9985_1050.n9 GND 0.22fF
C417 a_9985_1050.n10 GND 0.69fF
C418 a_9985_1050.n11 GND 0.83fF
C419 a_9985_1050.n12 GND 0.64fF
C420 a_10111_411.n0 GND 0.67fF
C421 a_10111_411.n1 GND 0.48fF
C422 a_10111_411.n2 GND 1.62fF
C423 a_10111_411.n3 GND 0.48fF
C424 a_10111_411.t10 GND 0.99fF
C425 a_10111_411.n4 GND 1.05fF
C426 a_10111_411.n5 GND 3.19fF
C427 a_10111_411.n6 GND 0.07fF
C428 a_10111_411.n7 GND 0.09fF
C429 a_10111_411.n8 GND 0.52fF
C430 a_10111_411.n9 GND 0.93fF
C431 a_10111_411.n10 GND 0.66fF
C432 a_10111_411.n11 GND 0.85fF
C433 a_10111_411.n12 GND 0.81fF
C434 a_10111_411.n13 GND 0.67fF
C435 a_1905_1050.n0 GND 0.35fF
C436 a_1905_1050.n1 GND 0.54fF
C437 a_1905_1050.n2 GND 0.04fF
C438 a_1905_1050.n3 GND 0.05fF
C439 a_1905_1050.n4 GND 0.03fF
C440 a_1905_1050.n5 GND 0.15fF
C441 a_1905_1050.n6 GND 0.63fF
C442 a_1905_1050.n7 GND 0.35fF
C443 a_1905_1050.n8 GND 0.45fF
C444 a_1905_1050.n9 GND 0.43fF
C445 a_1905_1050.n10 GND 0.46fF
C446 a_1905_1050.n11 GND 0.35fF
C447 a_1265_989.n0 GND 0.39fF
C448 a_1265_989.t12 GND 0.71fF
C449 a_1265_989.n1 GND 0.96fF
C450 a_1265_989.n2 GND 0.39fF
C451 a_1265_989.t7 GND 0.70fF
C452 a_1265_989.n3 GND 0.53fF
C453 a_1265_989.n4 GND 0.39fF
C454 a_1265_989.t8 GND 0.71fF
C455 a_1265_989.n5 GND 0.76fF
C456 a_1265_989.n6 GND 1.24fF
C457 a_1265_989.n7 GND 1.58fF
C458 a_1265_989.n8 GND 0.05fF
C459 a_1265_989.n9 GND 0.07fF
C460 a_1265_989.n10 GND 0.04fF
C461 a_1265_989.n11 GND 0.32fF
C462 a_1265_989.n12 GND 0.64fF
C463 a_1265_989.n13 GND 0.63fF
C464 a_1265_989.n14 GND 0.70fF
C465 a_1265_989.n15 GND 0.49fF
C466 a_217_1050.n0 GND 0.32fF
C467 a_217_1050.n1 GND 0.32fF
C468 a_217_1050.n2 GND 0.55fF
C469 a_217_1050.n3 GND 0.32fF
C470 a_217_1050.n4 GND 0.39fF
C471 a_217_1050.n5 GND 0.79fF
C472 a_217_1050.n6 GND 0.23fF
C473 a_217_1050.n7 GND 0.46fF
C474 a_217_1050.n8 GND 0.54fF
C475 a_217_1050.n9 GND 0.42fF
C476 a_14869_1051.n0 GND 0.36fF
C477 a_14869_1051.n1 GND 0.43fF
C478 a_14869_1051.n2 GND 0.80fF
C479 a_14869_1051.n3 GND 0.30fF
C480 a_14869_1051.n4 GND 0.52fF
C481 a_14869_1051.n5 GND 0.32fF
C482 a_15533_1051.n0 GND 0.29fF
C483 a_15533_1051.n1 GND 0.28fF
C484 a_15533_1051.n2 GND 0.37fF
C485 a_15533_1051.n3 GND 0.71fF
C486 a_15533_1051.n4 GND 0.27fF
C487 a_15533_1051.n5 GND 0.46fF
C488 a_3599_411.n0 GND 0.08fF
C489 a_3599_411.n1 GND 0.75fF
C490 a_3599_411.n2 GND 0.75fF
C491 a_3599_411.n3 GND 0.96fF
C492 a_3599_411.n4 GND 0.91fF
C493 a_3599_411.n5 GND 0.92fF
C494 a_3599_411.n6 GND 0.70fF
C495 a_3599_411.n7 GND 0.85fF
C496 a_3599_411.n8 GND 1.18fF
C497 a_3599_411.t12 GND 0.84fF
C498 a_3599_411.n9 GND 0.70fF
C499 a_3599_411.n10 GND 8.46fF
C500 a_3599_411.n11 GND 0.65fF
C501 a_3599_411.t14 GND 0.98fF
C502 a_3599_411.n12 GND 1.19fF
C503 a_3599_411.n13 GND 10.95fF
C504 a_3599_411.n14 GND 1.00fF
C505 a_3599_411.n15 GND 0.08fF
C506 a_3599_411.n16 GND 0.38fF
C507 a_3599_411.n17 GND 0.09fF
C508 a_5227_411.n0 GND 0.65fF
C509 a_5227_411.n1 GND 0.47fF
C510 a_5227_411.n2 GND 1.57fF
C511 a_5227_411.n3 GND 0.46fF
C512 a_5227_411.t9 GND 0.96fF
C513 a_5227_411.n4 GND 1.02fF
C514 a_5227_411.n5 GND 3.09fF
C515 a_5227_411.n6 GND 0.07fF
C516 a_5227_411.n7 GND 0.09fF
C517 a_5227_411.n8 GND 0.50fF
C518 a_5227_411.n9 GND 0.90fF
C519 a_5227_411.n10 GND 0.64fF
C520 a_5227_411.n11 GND 0.83fF
C521 a_5227_411.n12 GND 0.78fF
C522 a_5227_411.n13 GND 0.65fF
C523 a_5101_1050.n0 GND 0.51fF
C524 a_5101_1050.n1 GND 0.49fF
C525 a_5101_1050.n2 GND 0.85fF
C526 a_5101_1050.n3 GND 0.49fF
C527 a_5101_1050.n4 GND 0.62fF
C528 a_5101_1050.n5 GND 1.22fF
C529 a_5101_1050.n6 GND 0.36fF
C530 a_5101_1050.n7 GND 0.72fF
C531 a_5101_1050.n8 GND 0.84fF
C532 a_5101_1050.n9 GND 0.65fF
C533 a_7586_101.n0 GND 0.05fF
C534 a_7586_101.n1 GND 0.02fF
C535 a_7586_101.n2 GND 0.12fF
C536 a_7586_101.n3 GND 0.04fF
C537 a_7586_101.n4 GND 0.17fF
C538 a_6789_1050.n0 GND 0.39fF
C539 a_6789_1050.n1 GND 0.39fF
C540 a_6789_1050.n2 GND 0.50fF
C541 a_6789_1050.n3 GND 0.47fF
C542 a_6789_1050.n4 GND 0.51fF
C543 a_6789_1050.n5 GND 0.38fF
C544 a_6789_1050.n6 GND 0.59fF
C545 a_6789_1050.n7 GND 0.70fF
C546 a_6789_1050.n8 GND 0.08fF
C547 a_6789_1050.n9 GND 0.16fF
C548 a_6789_1050.n10 GND 0.05fF
C549 VDD.n1 GND 0.03fF
C550 VDD.n2 GND 0.10fF
C551 VDD.n3 GND 0.03fF
C552 VDD.n4 GND 0.02fF
C553 VDD.n5 GND 0.06fF
C554 VDD.n6 GND 0.02fF
C555 VDD.n7 GND 0.02fF
C556 VDD.n8 GND 0.02fF
C557 VDD.n9 GND 0.02fF
C558 VDD.n10 GND 0.02fF
C559 VDD.n11 GND 0.02fF
C560 VDD.n12 GND 0.02fF
C561 VDD.n13 GND 0.02fF
C562 VDD.n14 GND 0.04fF
C563 VDD.n15 GND 0.01fF
C564 VDD.n20 GND 0.47fF
C565 VDD.n21 GND 0.28fF
C566 VDD.n22 GND 0.02fF
C567 VDD.n23 GND 0.03fF
C568 VDD.n24 GND 0.06fF
C569 VDD.n25 GND 0.21fF
C570 VDD.n26 GND 0.01fF
C571 VDD.n27 GND 0.01fF
C572 VDD.n28 GND 0.07fF
C573 VDD.n29 GND 0.17fF
C574 VDD.n30 GND 0.01fF
C575 VDD.n31 GND 0.03fF
C576 VDD.n32 GND 0.03fF
C577 VDD.n33 GND 0.21fF
C578 VDD.n34 GND 0.01fF
C579 VDD.n35 GND 0.07fF
C580 VDD.n36 GND 0.01fF
C581 VDD.n37 GND 0.02fF
C582 VDD.n38 GND 0.28fF
C583 VDD.n39 GND 0.01fF
C584 VDD.n40 GND 0.02fF
C585 VDD.n41 GND 0.04fF
C586 VDD.n42 GND 0.06fF
C587 VDD.n43 GND 0.02fF
C588 VDD.n44 GND 0.02fF
C589 VDD.n45 GND 0.02fF
C590 VDD.n46 GND 0.02fF
C591 VDD.n47 GND 0.02fF
C592 VDD.n48 GND 0.02fF
C593 VDD.n49 GND 0.02fF
C594 VDD.n50 GND 0.02fF
C595 VDD.n51 GND 0.02fF
C596 VDD.n52 GND 0.02fF
C597 VDD.n53 GND 0.02fF
C598 VDD.n54 GND 0.03fF
C599 VDD.n55 GND 0.02fF
C600 VDD.n56 GND 0.19fF
C601 VDD.n57 GND 0.02fF
C602 VDD.n58 GND 0.02fF
C603 VDD.n60 GND 0.02fF
C604 VDD.n64 GND 0.28fF
C605 VDD.n65 GND 0.28fF
C606 VDD.n66 GND 0.01fF
C607 VDD.n67 GND 0.02fF
C608 VDD.n68 GND 0.04fF
C609 VDD.n69 GND 0.25fF
C610 VDD.n70 GND 0.01fF
C611 VDD.n71 GND 0.02fF
C612 VDD.n72 GND 0.02fF
C613 VDD.n73 GND 0.17fF
C614 VDD.n74 GND 0.01fF
C615 VDD.n75 GND 0.02fF
C616 VDD.n76 GND 0.02fF
C617 VDD.n77 GND 0.01fF
C618 VDD.n78 GND 0.03fF
C619 VDD.n79 GND 0.03fF
C620 VDD.n80 GND 0.15fF
C621 VDD.n81 GND 0.01fF
C622 VDD.n82 GND 0.03fF
C623 VDD.n83 GND 0.03fF
C624 VDD.n84 GND 0.17fF
C625 VDD.n85 GND 0.01fF
C626 VDD.n86 GND 0.02fF
C627 VDD.n87 GND 0.02fF
C628 VDD.n88 GND 0.26fF
C629 VDD.n89 GND 0.01fF
C630 VDD.n90 GND 0.02fF
C631 VDD.n91 GND 0.02fF
C632 VDD.n92 GND 0.28fF
C633 VDD.n93 GND 0.01fF
C634 VDD.n94 GND 0.02fF
C635 VDD.n95 GND 0.04fF
C636 VDD.n96 GND 0.22fF
C637 VDD.n97 GND 0.02fF
C638 VDD.n98 GND 0.02fF
C639 VDD.n99 GND 0.02fF
C640 VDD.n100 GND 0.06fF
C641 VDD.n101 GND 0.02fF
C642 VDD.n102 GND 0.02fF
C643 VDD.n103 GND 0.02fF
C644 VDD.n104 GND 0.02fF
C645 VDD.n105 GND 0.02fF
C646 VDD.n106 GND 0.02fF
C647 VDD.n107 GND 0.02fF
C648 VDD.n108 GND 0.02fF
C649 VDD.n109 GND 0.02fF
C650 VDD.n110 GND 0.02fF
C651 VDD.n111 GND 0.03fF
C652 VDD.n112 GND 0.02fF
C653 VDD.n113 GND 0.02fF
C654 VDD.n117 GND 0.28fF
C655 VDD.n118 GND 0.28fF
C656 VDD.n119 GND 0.01fF
C657 VDD.n120 GND 0.02fF
C658 VDD.n121 GND 0.04fF
C659 VDD.n122 GND 0.26fF
C660 VDD.n123 GND 0.01fF
C661 VDD.n124 GND 0.02fF
C662 VDD.n125 GND 0.02fF
C663 VDD.n126 GND 0.17fF
C664 VDD.n127 GND 0.01fF
C665 VDD.n128 GND 0.02fF
C666 VDD.n129 GND 0.02fF
C667 VDD.n130 GND 0.15fF
C668 VDD.n131 GND 0.01fF
C669 VDD.n132 GND 0.03fF
C670 VDD.n133 GND 0.03fF
C671 VDD.n134 GND 0.01fF
C672 VDD.n135 GND 0.03fF
C673 VDD.n136 GND 0.03fF
C674 VDD.n137 GND 0.17fF
C675 VDD.n138 GND 0.01fF
C676 VDD.n139 GND 0.02fF
C677 VDD.n140 GND 0.02fF
C678 VDD.n141 GND 0.25fF
C679 VDD.n142 GND 0.01fF
C680 VDD.n143 GND 0.02fF
C681 VDD.n144 GND 0.02fF
C682 VDD.n145 GND 0.28fF
C683 VDD.n146 GND 0.01fF
C684 VDD.n147 GND 0.02fF
C685 VDD.n148 GND 0.04fF
C686 VDD.n149 GND 0.22fF
C687 VDD.n150 GND 0.02fF
C688 VDD.n151 GND 0.02fF
C689 VDD.n152 GND 0.02fF
C690 VDD.n153 GND 0.06fF
C691 VDD.n154 GND 0.02fF
C692 VDD.n155 GND 0.02fF
C693 VDD.n156 GND 0.02fF
C694 VDD.n157 GND 0.02fF
C695 VDD.n158 GND 0.02fF
C696 VDD.n159 GND 0.02fF
C697 VDD.n160 GND 0.02fF
C698 VDD.n161 GND 0.02fF
C699 VDD.n162 GND 0.02fF
C700 VDD.n163 GND 0.02fF
C701 VDD.n164 GND 0.03fF
C702 VDD.n165 GND 0.02fF
C703 VDD.n166 GND 0.02fF
C704 VDD.n170 GND 0.28fF
C705 VDD.n171 GND 0.28fF
C706 VDD.n172 GND 0.01fF
C707 VDD.n173 GND 0.02fF
C708 VDD.n174 GND 0.04fF
C709 VDD.n175 GND 0.07fF
C710 VDD.n176 GND 0.25fF
C711 VDD.n177 GND 0.01fF
C712 VDD.n178 GND 0.01fF
C713 VDD.n179 GND 0.02fF
C714 VDD.n180 GND 0.17fF
C715 VDD.n181 GND 0.01fF
C716 VDD.n182 GND 0.02fF
C717 VDD.n183 GND 0.02fF
C718 VDD.n184 GND 0.08fF
C719 VDD.n185 GND 0.05fF
C720 VDD.n186 GND 0.01fF
C721 VDD.n187 GND 0.02fF
C722 VDD.n188 GND 0.03fF
C723 VDD.n189 GND 0.15fF
C724 VDD.n190 GND 0.01fF
C725 VDD.n191 GND 0.02fF
C726 VDD.n192 GND 0.03fF
C727 VDD.n193 GND 0.17fF
C728 VDD.n194 GND 0.01fF
C729 VDD.n195 GND 0.02fF
C730 VDD.n196 GND 0.02fF
C731 VDD.n197 GND 0.07fF
C732 VDD.n198 GND 0.26fF
C733 VDD.n199 GND 0.01fF
C734 VDD.n200 GND 0.01fF
C735 VDD.n201 GND 0.02fF
C736 VDD.n202 GND 0.28fF
C737 VDD.n203 GND 0.01fF
C738 VDD.n204 GND 0.02fF
C739 VDD.n205 GND 0.04fF
C740 VDD.n206 GND 0.27fF
C741 VDD.n207 GND 0.02fF
C742 VDD.n208 GND 0.02fF
C743 VDD.n209 GND 0.02fF
C744 VDD.n210 GND 0.06fF
C745 VDD.n211 GND 0.02fF
C746 VDD.n212 GND 0.02fF
C747 VDD.n213 GND 0.02fF
C748 VDD.n214 GND 0.02fF
C749 VDD.n215 GND 0.02fF
C750 VDD.n216 GND 0.02fF
C751 VDD.n217 GND 0.02fF
C752 VDD.n218 GND 0.02fF
C753 VDD.n219 GND 0.02fF
C754 VDD.n220 GND 0.02fF
C755 VDD.n221 GND 0.03fF
C756 VDD.n222 GND 0.02fF
C757 VDD.n223 GND 0.02fF
C758 VDD.n227 GND 0.28fF
C759 VDD.n228 GND 0.28fF
C760 VDD.n229 GND 0.01fF
C761 VDD.n230 GND 0.02fF
C762 VDD.n231 GND 0.04fF
C763 VDD.n232 GND 0.28fF
C764 VDD.n233 GND 0.01fF
C765 VDD.n234 GND 0.02fF
C766 VDD.n235 GND 0.02fF
C767 VDD.n236 GND 0.23fF
C768 VDD.n237 GND 0.01fF
C769 VDD.n238 GND 0.07fF
C770 VDD.n239 GND 0.02fF
C771 VDD.n240 GND 0.17fF
C772 VDD.n241 GND 0.01fF
C773 VDD.n242 GND 0.02fF
C774 VDD.n243 GND 0.02fF
C775 VDD.n244 GND 0.17fF
C776 VDD.n245 GND 0.01fF
C777 VDD.n246 GND 0.08fF
C778 VDD.n247 GND 0.05fF
C779 VDD.n248 GND 0.02fF
C780 VDD.n249 GND 0.02fF
C781 VDD.n250 GND 0.15fF
C782 VDD.n251 GND 0.02fF
C783 VDD.n252 GND 0.02fF
C784 VDD.n253 GND 0.03fF
C785 VDD.n254 GND 0.15fF
C786 VDD.n255 GND 0.02fF
C787 VDD.n256 GND 0.02fF
C788 VDD.n257 GND 0.03fF
C789 VDD.n258 GND 0.08fF
C790 VDD.n259 GND 0.05fF
C791 VDD.n260 GND 0.16fF
C792 VDD.n261 GND 0.01fF
C793 VDD.n262 GND 0.02fF
C794 VDD.n263 GND 0.02fF
C795 VDD.n264 GND 0.17fF
C796 VDD.n265 GND 0.01fF
C797 VDD.n266 GND 0.02fF
C798 VDD.n267 GND 0.02fF
C799 VDD.n268 GND 0.06fF
C800 VDD.n269 GND 0.23fF
C801 VDD.n270 GND 0.01fF
C802 VDD.n271 GND 0.01fF
C803 VDD.n272 GND 0.02fF
C804 VDD.n273 GND 0.28fF
C805 VDD.n274 GND 0.01fF
C806 VDD.n275 GND 0.02fF
C807 VDD.n276 GND 0.02fF
C808 VDD.n277 GND 0.28fF
C809 VDD.n278 GND 0.01fF
C810 VDD.n279 GND 0.02fF
C811 VDD.n280 GND 0.04fF
C812 VDD.n281 GND 0.27fF
C813 VDD.n282 GND 0.02fF
C814 VDD.n283 GND 0.02fF
C815 VDD.n284 GND 0.02fF
C816 VDD.n285 GND 0.06fF
C817 VDD.n286 GND 0.02fF
C818 VDD.n287 GND 0.02fF
C819 VDD.n288 GND 0.02fF
C820 VDD.n289 GND 0.02fF
C821 VDD.n290 GND 0.02fF
C822 VDD.n291 GND 0.02fF
C823 VDD.n292 GND 0.02fF
C824 VDD.n293 GND 0.02fF
C825 VDD.n294 GND 0.02fF
C826 VDD.n295 GND 0.02fF
C827 VDD.n296 GND 0.03fF
C828 VDD.n297 GND 0.02fF
C829 VDD.n298 GND 0.02fF
C830 VDD.n302 GND 0.28fF
C831 VDD.n303 GND 0.28fF
C832 VDD.n304 GND 0.01fF
C833 VDD.n305 GND 0.02fF
C834 VDD.n306 GND 0.04fF
C835 VDD.n307 GND 0.06fF
C836 VDD.n308 GND 0.25fF
C837 VDD.n309 GND 0.01fF
C838 VDD.n310 GND 0.01fF
C839 VDD.n311 GND 0.02fF
C840 VDD.n312 GND 0.17fF
C841 VDD.n313 GND 0.01fF
C842 VDD.n314 GND 0.02fF
C843 VDD.n315 GND 0.02fF
C844 VDD.n316 GND 0.08fF
C845 VDD.n317 GND 0.05fF
C846 VDD.n318 GND 0.01fF
C847 VDD.n319 GND 0.02fF
C848 VDD.n320 GND 0.03fF
C849 VDD.n321 GND 0.15fF
C850 VDD.n322 GND 0.01fF
C851 VDD.n323 GND 0.02fF
C852 VDD.n324 GND 0.03fF
C853 VDD.n325 GND 0.17fF
C854 VDD.n326 GND 0.01fF
C855 VDD.n327 GND 0.02fF
C856 VDD.n328 GND 0.02fF
C857 VDD.n329 GND 0.07fF
C858 VDD.n330 GND 0.26fF
C859 VDD.n331 GND 0.01fF
C860 VDD.n332 GND 0.01fF
C861 VDD.n333 GND 0.02fF
C862 VDD.n334 GND 0.28fF
C863 VDD.n335 GND 0.01fF
C864 VDD.n336 GND 0.02fF
C865 VDD.n337 GND 0.04fF
C866 VDD.n338 GND 0.22fF
C867 VDD.n339 GND 0.02fF
C868 VDD.n340 GND 0.02fF
C869 VDD.n341 GND 0.02fF
C870 VDD.n342 GND 0.06fF
C871 VDD.n343 GND 0.02fF
C872 VDD.n344 GND 0.02fF
C873 VDD.n345 GND 0.02fF
C874 VDD.n346 GND 0.02fF
C875 VDD.n347 GND 0.02fF
C876 VDD.n348 GND 0.02fF
C877 VDD.n349 GND 0.02fF
C878 VDD.n350 GND 0.02fF
C879 VDD.n351 GND 0.02fF
C880 VDD.n352 GND 0.02fF
C881 VDD.n353 GND 0.03fF
C882 VDD.n354 GND 0.02fF
C883 VDD.n355 GND 0.02fF
C884 VDD.n359 GND 0.28fF
C885 VDD.n360 GND 0.28fF
C886 VDD.n361 GND 0.01fF
C887 VDD.n362 GND 0.02fF
C888 VDD.n363 GND 0.04fF
C889 VDD.n364 GND 0.06fF
C890 VDD.n365 GND 0.25fF
C891 VDD.n366 GND 0.01fF
C892 VDD.n367 GND 0.01fF
C893 VDD.n368 GND 0.02fF
C894 VDD.n369 GND 0.17fF
C895 VDD.n370 GND 0.01fF
C896 VDD.n371 GND 0.02fF
C897 VDD.n372 GND 0.02fF
C898 VDD.n373 GND 0.08fF
C899 VDD.n374 GND 0.05fF
C900 VDD.n375 GND 0.01fF
C901 VDD.n376 GND 0.02fF
C902 VDD.n377 GND 0.03fF
C903 VDD.n378 GND 0.15fF
C904 VDD.n379 GND 0.01fF
C905 VDD.n380 GND 0.02fF
C906 VDD.n381 GND 0.03fF
C907 VDD.n382 GND 0.17fF
C908 VDD.n383 GND 0.01fF
C909 VDD.n384 GND 0.02fF
C910 VDD.n385 GND 0.02fF
C911 VDD.n386 GND 0.07fF
C912 VDD.n387 GND 0.26fF
C913 VDD.n388 GND 0.01fF
C914 VDD.n389 GND 0.01fF
C915 VDD.n390 GND 0.02fF
C916 VDD.n391 GND 0.28fF
C917 VDD.n392 GND 0.01fF
C918 VDD.n393 GND 0.02fF
C919 VDD.n394 GND 0.04fF
C920 VDD.n395 GND 0.27fF
C921 VDD.n396 GND 0.02fF
C922 VDD.n397 GND 0.02fF
C923 VDD.n398 GND 0.02fF
C924 VDD.n399 GND 0.06fF
C925 VDD.n400 GND 0.02fF
C926 VDD.n401 GND 0.02fF
C927 VDD.n402 GND 0.02fF
C928 VDD.n403 GND 0.02fF
C929 VDD.n404 GND 0.02fF
C930 VDD.n405 GND 0.02fF
C931 VDD.n406 GND 0.02fF
C932 VDD.n407 GND 0.02fF
C933 VDD.n408 GND 0.02fF
C934 VDD.n409 GND 0.02fF
C935 VDD.n410 GND 0.03fF
C936 VDD.n411 GND 0.02fF
C937 VDD.n412 GND 0.02fF
C938 VDD.n416 GND 0.28fF
C939 VDD.n417 GND 0.28fF
C940 VDD.n418 GND 0.01fF
C941 VDD.n419 GND 0.02fF
C942 VDD.n420 GND 0.04fF
C943 VDD.n421 GND 0.28fF
C944 VDD.n422 GND 0.01fF
C945 VDD.n423 GND 0.02fF
C946 VDD.n424 GND 0.02fF
C947 VDD.n425 GND 0.23fF
C948 VDD.n426 GND 0.01fF
C949 VDD.n427 GND 0.07fF
C950 VDD.n428 GND 0.02fF
C951 VDD.n429 GND 0.17fF
C952 VDD.n430 GND 0.01fF
C953 VDD.n431 GND 0.02fF
C954 VDD.n432 GND 0.02fF
C955 VDD.n433 GND 0.17fF
C956 VDD.n434 GND 0.01fF
C957 VDD.n435 GND 0.08fF
C958 VDD.n436 GND 0.05fF
C959 VDD.n437 GND 0.02fF
C960 VDD.n438 GND 0.02fF
C961 VDD.n439 GND 0.15fF
C962 VDD.n440 GND 0.02fF
C963 VDD.n441 GND 0.02fF
C964 VDD.n442 GND 0.03fF
C965 VDD.n443 GND 0.15fF
C966 VDD.n444 GND 0.02fF
C967 VDD.n445 GND 0.02fF
C968 VDD.n446 GND 0.03fF
C969 VDD.n447 GND 0.08fF
C970 VDD.n448 GND 0.05fF
C971 VDD.n449 GND 0.16fF
C972 VDD.n450 GND 0.01fF
C973 VDD.n451 GND 0.02fF
C974 VDD.n452 GND 0.02fF
C975 VDD.n453 GND 0.17fF
C976 VDD.n454 GND 0.01fF
C977 VDD.n455 GND 0.02fF
C978 VDD.n456 GND 0.02fF
C979 VDD.n457 GND 0.06fF
C980 VDD.n458 GND 0.23fF
C981 VDD.n459 GND 0.01fF
C982 VDD.n460 GND 0.01fF
C983 VDD.n461 GND 0.02fF
C984 VDD.n462 GND 0.28fF
C985 VDD.n463 GND 0.01fF
C986 VDD.n464 GND 0.02fF
C987 VDD.n465 GND 0.02fF
C988 VDD.n466 GND 0.28fF
C989 VDD.n467 GND 0.01fF
C990 VDD.n468 GND 0.02fF
C991 VDD.n469 GND 0.04fF
C992 VDD.n470 GND 0.32fF
C993 VDD.n471 GND 0.02fF
C994 VDD.n472 GND 0.02fF
C995 VDD.n473 GND 0.02fF
C996 VDD.n474 GND 0.06fF
C997 VDD.n475 GND 0.02fF
C998 VDD.n476 GND 0.02fF
C999 VDD.n477 GND 0.02fF
C1000 VDD.n478 GND 0.02fF
C1001 VDD.n479 GND 0.02fF
C1002 VDD.n480 GND 0.02fF
C1003 VDD.n481 GND 0.02fF
C1004 VDD.n482 GND 0.02fF
C1005 VDD.n483 GND 0.02fF
C1006 VDD.n484 GND 0.02fF
C1007 VDD.n485 GND 0.03fF
C1008 VDD.n486 GND 0.02fF
C1009 VDD.n487 GND 0.02fF
C1010 VDD.n491 GND 0.28fF
C1011 VDD.n492 GND 0.28fF
C1012 VDD.n493 GND 0.01fF
C1013 VDD.n494 GND 0.02fF
C1014 VDD.n495 GND 0.04fF
C1015 VDD.n496 GND 0.28fF
C1016 VDD.n497 GND 0.01fF
C1017 VDD.n498 GND 0.02fF
C1018 VDD.n499 GND 0.02fF
C1019 VDD.n500 GND 0.23fF
C1020 VDD.n501 GND 0.01fF
C1021 VDD.n502 GND 0.07fF
C1022 VDD.n503 GND 0.02fF
C1023 VDD.n504 GND 0.17fF
C1024 VDD.n505 GND 0.01fF
C1025 VDD.n506 GND 0.02fF
C1026 VDD.n507 GND 0.02fF
C1027 VDD.n508 GND 0.17fF
C1028 VDD.n509 GND 0.01fF
C1029 VDD.n510 GND 0.08fF
C1030 VDD.n511 GND 0.05fF
C1031 VDD.n512 GND 0.02fF
C1032 VDD.n513 GND 0.02fF
C1033 VDD.n514 GND 0.15fF
C1034 VDD.n515 GND 0.02fF
C1035 VDD.n516 GND 0.02fF
C1036 VDD.n517 GND 0.03fF
C1037 VDD.n518 GND 0.15fF
C1038 VDD.n519 GND 0.02fF
C1039 VDD.n520 GND 0.02fF
C1040 VDD.n521 GND 0.03fF
C1041 VDD.n522 GND 0.08fF
C1042 VDD.n523 GND 0.05fF
C1043 VDD.n524 GND 0.16fF
C1044 VDD.n525 GND 0.01fF
C1045 VDD.n526 GND 0.02fF
C1046 VDD.n527 GND 0.02fF
C1047 VDD.n528 GND 0.17fF
C1048 VDD.n529 GND 0.01fF
C1049 VDD.n530 GND 0.02fF
C1050 VDD.n531 GND 0.02fF
C1051 VDD.n532 GND 0.06fF
C1052 VDD.n533 GND 0.23fF
C1053 VDD.n534 GND 0.01fF
C1054 VDD.n535 GND 0.01fF
C1055 VDD.n536 GND 0.02fF
C1056 VDD.n537 GND 0.28fF
C1057 VDD.n538 GND 0.01fF
C1058 VDD.n539 GND 0.02fF
C1059 VDD.n540 GND 0.02fF
C1060 VDD.n541 GND 0.28fF
C1061 VDD.n542 GND 0.01fF
C1062 VDD.n543 GND 0.02fF
C1063 VDD.n544 GND 0.04fF
C1064 VDD.n545 GND 0.27fF
C1065 VDD.n546 GND 0.02fF
C1066 VDD.n547 GND 0.02fF
C1067 VDD.n548 GND 0.02fF
C1068 VDD.n549 GND 0.06fF
C1069 VDD.n550 GND 0.02fF
C1070 VDD.n551 GND 0.02fF
C1071 VDD.n552 GND 0.02fF
C1072 VDD.n553 GND 0.02fF
C1073 VDD.n554 GND 0.02fF
C1074 VDD.n555 GND 0.02fF
C1075 VDD.n556 GND 0.02fF
C1076 VDD.n557 GND 0.02fF
C1077 VDD.n558 GND 0.02fF
C1078 VDD.n559 GND 0.02fF
C1079 VDD.n560 GND 0.03fF
C1080 VDD.n561 GND 0.02fF
C1081 VDD.n562 GND 0.02fF
C1082 VDD.n566 GND 0.28fF
C1083 VDD.n567 GND 0.28fF
C1084 VDD.n568 GND 0.01fF
C1085 VDD.n569 GND 0.02fF
C1086 VDD.n570 GND 0.04fF
C1087 VDD.n571 GND 0.06fF
C1088 VDD.n572 GND 0.25fF
C1089 VDD.n573 GND 0.01fF
C1090 VDD.n574 GND 0.01fF
C1091 VDD.n575 GND 0.02fF
C1092 VDD.n576 GND 0.17fF
C1093 VDD.n577 GND 0.01fF
C1094 VDD.n578 GND 0.02fF
C1095 VDD.n579 GND 0.02fF
C1096 VDD.n580 GND 0.08fF
C1097 VDD.n581 GND 0.05fF
C1098 VDD.n582 GND 0.01fF
C1099 VDD.n583 GND 0.02fF
C1100 VDD.n584 GND 0.03fF
C1101 VDD.n585 GND 0.15fF
C1102 VDD.n586 GND 0.01fF
C1103 VDD.n587 GND 0.02fF
C1104 VDD.n588 GND 0.03fF
C1105 VDD.n589 GND 0.17fF
C1106 VDD.n590 GND 0.01fF
C1107 VDD.n591 GND 0.02fF
C1108 VDD.n592 GND 0.02fF
C1109 VDD.n593 GND 0.07fF
C1110 VDD.n594 GND 0.26fF
C1111 VDD.n595 GND 0.01fF
C1112 VDD.n596 GND 0.01fF
C1113 VDD.n597 GND 0.02fF
C1114 VDD.n598 GND 0.28fF
C1115 VDD.n599 GND 0.01fF
C1116 VDD.n600 GND 0.02fF
C1117 VDD.n601 GND 0.04fF
C1118 VDD.n602 GND 0.27fF
C1119 VDD.n603 GND 0.02fF
C1120 VDD.n604 GND 0.02fF
C1121 VDD.n605 GND 0.02fF
C1122 VDD.n606 GND 0.06fF
C1123 VDD.n607 GND 0.02fF
C1124 VDD.n608 GND 0.02fF
C1125 VDD.n609 GND 0.02fF
C1126 VDD.n610 GND 0.02fF
C1127 VDD.n611 GND 0.02fF
C1128 VDD.n612 GND 0.02fF
C1129 VDD.n613 GND 0.02fF
C1130 VDD.n614 GND 0.02fF
C1131 VDD.n615 GND 0.02fF
C1132 VDD.n616 GND 0.02fF
C1133 VDD.n617 GND 0.03fF
C1134 VDD.n618 GND 0.02fF
C1135 VDD.n619 GND 0.02fF
C1136 VDD.n623 GND 0.28fF
C1137 VDD.n624 GND 0.28fF
C1138 VDD.n625 GND 0.01fF
C1139 VDD.n626 GND 0.02fF
C1140 VDD.n627 GND 0.04fF
C1141 VDD.n628 GND 0.28fF
C1142 VDD.n629 GND 0.01fF
C1143 VDD.n630 GND 0.02fF
C1144 VDD.n631 GND 0.02fF
C1145 VDD.n632 GND 0.23fF
C1146 VDD.n633 GND 0.01fF
C1147 VDD.n634 GND 0.07fF
C1148 VDD.n635 GND 0.02fF
C1149 VDD.n636 GND 0.17fF
C1150 VDD.n637 GND 0.01fF
C1151 VDD.n638 GND 0.02fF
C1152 VDD.n639 GND 0.02fF
C1153 VDD.n640 GND 0.17fF
C1154 VDD.n641 GND 0.01fF
C1155 VDD.n642 GND 0.08fF
C1156 VDD.n643 GND 0.05fF
C1157 VDD.n644 GND 0.02fF
C1158 VDD.n645 GND 0.02fF
C1159 VDD.n646 GND 0.15fF
C1160 VDD.n647 GND 0.02fF
C1161 VDD.n648 GND 0.02fF
C1162 VDD.n649 GND 0.03fF
C1163 VDD.n650 GND 0.15fF
C1164 VDD.n651 GND 0.02fF
C1165 VDD.n652 GND 0.02fF
C1166 VDD.n653 GND 0.03fF
C1167 VDD.n654 GND 0.08fF
C1168 VDD.n655 GND 0.05fF
C1169 VDD.n656 GND 0.16fF
C1170 VDD.n657 GND 0.01fF
C1171 VDD.n658 GND 0.02fF
C1172 VDD.n659 GND 0.02fF
C1173 VDD.n660 GND 0.17fF
C1174 VDD.n661 GND 0.01fF
C1175 VDD.n662 GND 0.02fF
C1176 VDD.n663 GND 0.02fF
C1177 VDD.n664 GND 0.06fF
C1178 VDD.n665 GND 0.23fF
C1179 VDD.n666 GND 0.01fF
C1180 VDD.n667 GND 0.01fF
C1181 VDD.n668 GND 0.02fF
C1182 VDD.n669 GND 0.28fF
C1183 VDD.n670 GND 0.01fF
C1184 VDD.n671 GND 0.02fF
C1185 VDD.n672 GND 0.02fF
C1186 VDD.n673 GND 0.28fF
C1187 VDD.n674 GND 0.01fF
C1188 VDD.n675 GND 0.02fF
C1189 VDD.n676 GND 0.04fF
C1190 VDD.n677 GND 0.27fF
C1191 VDD.n678 GND 0.02fF
C1192 VDD.n679 GND 0.02fF
C1193 VDD.n680 GND 0.02fF
C1194 VDD.n681 GND 0.06fF
C1195 VDD.n682 GND 0.02fF
C1196 VDD.n683 GND 0.02fF
C1197 VDD.n684 GND 0.02fF
C1198 VDD.n685 GND 0.02fF
C1199 VDD.n686 GND 0.02fF
C1200 VDD.n687 GND 0.02fF
C1201 VDD.n688 GND 0.02fF
C1202 VDD.n689 GND 0.02fF
C1203 VDD.n690 GND 0.02fF
C1204 VDD.n691 GND 0.02fF
C1205 VDD.n692 GND 0.03fF
C1206 VDD.n693 GND 0.02fF
C1207 VDD.n694 GND 0.02fF
C1208 VDD.n698 GND 0.28fF
C1209 VDD.n699 GND 0.28fF
C1210 VDD.n700 GND 0.01fF
C1211 VDD.n701 GND 0.02fF
C1212 VDD.n702 GND 0.04fF
C1213 VDD.n703 GND 0.06fF
C1214 VDD.n704 GND 0.25fF
C1215 VDD.n705 GND 0.01fF
C1216 VDD.n706 GND 0.01fF
C1217 VDD.n707 GND 0.02fF
C1218 VDD.n708 GND 0.17fF
C1219 VDD.n709 GND 0.01fF
C1220 VDD.n710 GND 0.02fF
C1221 VDD.n711 GND 0.02fF
C1222 VDD.n712 GND 0.14fF
C1223 VDD.n713 GND 0.02fF
C1224 VDD.n714 GND 0.02fF
C1225 VDD.n715 GND 0.06fF
C1226 VDD.n716 GND 0.02fF
C1227 VDD.n717 GND 0.02fF
C1228 VDD.n718 GND 0.02fF
C1229 VDD.n719 GND 0.02fF
C1230 VDD.n720 GND 0.02fF
C1231 VDD.n721 GND 0.02fF
C1232 VDD.n722 GND 0.02fF
C1233 VDD.n723 GND 0.02fF
C1234 VDD.n724 GND 0.03fF
C1235 VDD.n725 GND 0.04fF
C1236 VDD.n726 GND 0.02fF
C1237 VDD.n730 GND 0.47fF
C1238 VDD.n731 GND 0.28fF
C1239 VDD.n732 GND 0.02fF
C1240 VDD.n733 GND 0.03fF
C1241 VDD.n734 GND 0.03fF
C1242 VDD.n735 GND 0.07fF
C1243 VDD.n736 GND 0.26fF
C1244 VDD.n737 GND 0.01fF
C1245 VDD.n738 GND 0.01fF
C1246 VDD.n739 GND 0.02fF
C1247 VDD.n740 GND 0.17fF
C1248 VDD.n741 GND 0.01fF
C1249 VDD.n742 GND 0.02fF
C1250 VDD.n743 GND 0.02fF
C1251 VDD.n744 GND 0.15fF
C1252 VDD.n745 GND 0.01fF
C1253 VDD.n746 GND 0.02fF
C1254 VDD.n747 GND 0.03fF
C1255 VDD.n748 GND 0.08fF
C1256 VDD.n749 GND 0.05fF
C1257 VDD.n750 GND 0.01fF
C1258 VDD.n751 GND 0.02fF
C1259 VDD.n752 GND 0.03fF
C1260 VDD.n753 GND 0.17fF
C1261 VDD.n754 GND 0.01fF
C1262 VDD.n755 GND 0.02fF
C1263 VDD.n756 GND 0.02fF
C1264 VDD.n757 GND 0.06fF
C1265 VDD.n758 GND 0.25fF
C1266 VDD.n759 GND 0.01fF
C1267 VDD.n760 GND 0.01fF
C1268 VDD.n761 GND 0.02fF
C1269 VDD.n762 GND 0.28fF
C1270 VDD.n763 GND 0.01fF
C1271 VDD.n764 GND 0.02fF
C1272 VDD.n765 GND 0.04fF
C1273 VDD.n766 GND 0.06fF
C1274 VDD.n767 GND 0.02fF
C1275 VDD.n768 GND 0.02fF
C1276 VDD.n769 GND 0.02fF
C1277 VDD.n770 GND 0.02fF
C1278 VDD.n771 GND 0.02fF
C1279 VDD.n772 GND 0.02fF
C1280 VDD.n773 GND 0.02fF
C1281 VDD.n774 GND 0.02fF
C1282 VDD.n775 GND 0.02fF
C1283 VDD.n776 GND 0.02fF
C1284 VDD.n777 GND 0.02fF
C1285 VDD.n778 GND 0.03fF
C1286 VDD.n779 GND 0.02fF
C1287 VDD.n782 GND 0.02fF
C1288 VDD.n784 GND 0.02fF
C1289 VDD.n785 GND 0.27fF
C1290 VDD.n786 GND 0.02fF
C1291 VDD.n788 GND 0.28fF
C1292 VDD.n789 GND 0.28fF
C1293 VDD.n790 GND 0.01fF
C1294 VDD.n791 GND 0.02fF
C1295 VDD.n792 GND 0.04fF
C1296 VDD.n793 GND 0.28fF
C1297 VDD.n794 GND 0.01fF
C1298 VDD.n795 GND 0.02fF
C1299 VDD.n796 GND 0.02fF
C1300 VDD.n797 GND 0.06fF
C1301 VDD.n798 GND 0.23fF
C1302 VDD.n799 GND 0.01fF
C1303 VDD.n800 GND 0.01fF
C1304 VDD.n801 GND 0.02fF
C1305 VDD.n802 GND 0.17fF
C1306 VDD.n803 GND 0.01fF
C1307 VDD.n804 GND 0.02fF
C1308 VDD.n805 GND 0.02fF
C1309 VDD.n806 GND 0.08fF
C1310 VDD.n807 GND 0.05fF
C1311 VDD.n808 GND 0.16fF
C1312 VDD.n809 GND 0.01fF
C1313 VDD.n810 GND 0.02fF
C1314 VDD.n811 GND 0.02fF
C1315 VDD.n812 GND 0.15fF
C1316 VDD.n813 GND 0.02fF
C1317 VDD.n814 GND 0.02fF
C1318 VDD.n815 GND 0.03fF
C1319 VDD.n816 GND 0.15fF
C1320 VDD.n817 GND 0.02fF
C1321 VDD.n818 GND 0.02fF
C1322 VDD.n819 GND 0.03fF
C1323 VDD.n820 GND 0.17fF
C1324 VDD.n821 GND 0.01fF
C1325 VDD.n822 GND 0.08fF
C1326 VDD.n823 GND 0.05fF
C1327 VDD.n824 GND 0.02fF
C1328 VDD.n825 GND 0.02fF
C1329 VDD.n826 GND 0.17fF
C1330 VDD.n827 GND 0.01fF
C1331 VDD.n828 GND 0.02fF
C1332 VDD.n829 GND 0.02fF
C1333 VDD.n830 GND 0.23fF
C1334 VDD.n831 GND 0.01fF
C1335 VDD.n832 GND 0.07fF
C1336 VDD.n833 GND 0.02fF
C1337 VDD.n834 GND 0.28fF
C1338 VDD.n835 GND 0.01fF
C1339 VDD.n836 GND 0.02fF
C1340 VDD.n837 GND 0.02fF
C1341 VDD.n838 GND 0.28fF
C1342 VDD.n839 GND 0.01fF
C1343 VDD.n840 GND 0.02fF
C1344 VDD.n841 GND 0.04fF
C1345 VDD.n842 GND 0.32fF
C1346 VDD.n843 GND 0.02fF
C1347 VDD.n844 GND 0.02fF
C1348 VDD.n845 GND 0.02fF
C1349 VDD.n846 GND 0.06fF
C1350 VDD.n847 GND 0.02fF
C1351 VDD.n848 GND 0.02fF
C1352 VDD.n849 GND 0.02fF
C1353 VDD.n850 GND 0.02fF
C1354 VDD.n851 GND 0.02fF
C1355 VDD.n852 GND 0.02fF
C1356 VDD.n853 GND 0.02fF
C1357 VDD.n854 GND 0.02fF
C1358 VDD.n855 GND 0.02fF
C1359 VDD.n856 GND 0.02fF
C1360 VDD.n857 GND 0.03fF
C1361 VDD.n858 GND 0.02fF
C1362 VDD.n859 GND 0.02fF
C1363 VDD.n863 GND 0.28fF
C1364 VDD.n864 GND 0.28fF
C1365 VDD.n865 GND 0.01fF
C1366 VDD.n866 GND 0.02fF
C1367 VDD.n867 GND 0.04fF
C1368 VDD.n868 GND 0.28fF
C1369 VDD.n869 GND 0.01fF
C1370 VDD.n870 GND 0.02fF
C1371 VDD.n871 GND 0.02fF
C1372 VDD.n872 GND 0.06fF
C1373 VDD.n873 GND 0.23fF
C1374 VDD.n874 GND 0.01fF
C1375 VDD.n875 GND 0.01fF
C1376 VDD.n876 GND 0.02fF
C1377 VDD.n877 GND 0.17fF
C1378 VDD.n878 GND 0.01fF
C1379 VDD.n879 GND 0.02fF
C1380 VDD.n880 GND 0.02fF
C1381 VDD.n881 GND 0.08fF
C1382 VDD.n882 GND 0.05fF
C1383 VDD.n883 GND 0.16fF
C1384 VDD.n884 GND 0.01fF
C1385 VDD.n885 GND 0.02fF
C1386 VDD.n886 GND 0.02fF
C1387 VDD.n887 GND 0.15fF
C1388 VDD.n888 GND 0.02fF
C1389 VDD.n889 GND 0.02fF
C1390 VDD.n890 GND 0.03fF
C1391 VDD.n891 GND 0.15fF
C1392 VDD.n892 GND 0.02fF
C1393 VDD.n893 GND 0.02fF
C1394 VDD.n894 GND 0.03fF
C1395 VDD.n895 GND 0.17fF
C1396 VDD.n896 GND 0.01fF
C1397 VDD.n897 GND 0.08fF
C1398 VDD.n898 GND 0.05fF
C1399 VDD.n899 GND 0.02fF
C1400 VDD.n900 GND 0.02fF
C1401 VDD.n901 GND 0.17fF
C1402 VDD.n902 GND 0.01fF
C1403 VDD.n903 GND 0.02fF
C1404 VDD.n904 GND 0.02fF
C1405 VDD.n905 GND 0.23fF
C1406 VDD.n906 GND 0.01fF
C1407 VDD.n907 GND 0.07fF
C1408 VDD.n908 GND 0.02fF
C1409 VDD.n909 GND 0.28fF
C1410 VDD.n910 GND 0.01fF
C1411 VDD.n911 GND 0.02fF
C1412 VDD.n912 GND 0.02fF
C1413 VDD.n913 GND 0.28fF
C1414 VDD.n914 GND 0.01fF
C1415 VDD.n915 GND 0.02fF
C1416 VDD.n916 GND 0.04fF
C1417 VDD.n917 GND 0.27fF
C1418 VDD.n918 GND 0.02fF
C1419 VDD.n919 GND 0.02fF
C1420 VDD.n920 GND 0.02fF
C1421 VDD.n921 GND 0.06fF
C1422 VDD.n922 GND 0.02fF
C1423 VDD.n923 GND 0.02fF
C1424 VDD.n924 GND 0.02fF
C1425 VDD.n925 GND 0.02fF
C1426 VDD.n926 GND 0.02fF
C1427 VDD.n927 GND 0.02fF
C1428 VDD.n928 GND 0.02fF
C1429 VDD.n929 GND 0.02fF
C1430 VDD.n930 GND 0.02fF
C1431 VDD.n931 GND 0.02fF
C1432 VDD.n932 GND 0.03fF
C1433 VDD.n933 GND 0.02fF
C1434 VDD.n934 GND 0.02fF
C1435 VDD.n938 GND 0.28fF
C1436 VDD.n939 GND 0.28fF
C1437 VDD.n940 GND 0.01fF
C1438 VDD.n941 GND 0.02fF
C1439 VDD.n942 GND 0.04fF
C1440 VDD.n943 GND 0.07fF
C1441 VDD.n944 GND 0.26fF
C1442 VDD.n945 GND 0.01fF
C1443 VDD.n946 GND 0.01fF
C1444 VDD.n947 GND 0.02fF
C1445 VDD.n948 GND 0.17fF
C1446 VDD.n949 GND 0.01fF
C1447 VDD.n950 GND 0.02fF
C1448 VDD.n951 GND 0.02fF
C1449 VDD.n952 GND 0.15fF
C1450 VDD.n953 GND 0.01fF
C1451 VDD.n954 GND 0.02fF
C1452 VDD.n955 GND 0.03fF
C1453 VDD.n956 GND 0.08fF
C1454 VDD.n957 GND 0.05fF
C1455 VDD.n958 GND 0.01fF
C1456 VDD.n959 GND 0.02fF
C1457 VDD.n960 GND 0.03fF
C1458 VDD.n961 GND 0.17fF
C1459 VDD.n962 GND 0.01fF
C1460 VDD.n963 GND 0.02fF
C1461 VDD.n964 GND 0.02fF
C1462 VDD.n965 GND 0.06fF
C1463 VDD.n966 GND 0.25fF
C1464 VDD.n967 GND 0.01fF
C1465 VDD.n968 GND 0.01fF
C1466 VDD.n969 GND 0.02fF
C1467 VDD.n970 GND 0.28fF
C1468 VDD.n971 GND 0.01fF
C1469 VDD.n972 GND 0.02fF
C1470 VDD.n973 GND 0.04fF
C1471 VDD.n974 GND 0.22fF
C1472 VDD.n975 GND 0.02fF
C1473 VDD.n976 GND 0.02fF
C1474 VDD.n977 GND 0.02fF
C1475 VDD.n978 GND 0.06fF
C1476 VDD.n979 GND 0.02fF
C1477 VDD.n980 GND 0.02fF
C1478 VDD.n981 GND 0.02fF
C1479 VDD.n982 GND 0.02fF
C1480 VDD.n983 GND 0.02fF
C1481 VDD.n984 GND 0.02fF
C1482 VDD.n985 GND 0.02fF
C1483 VDD.n986 GND 0.02fF
C1484 VDD.n987 GND 0.02fF
C1485 VDD.n988 GND 0.02fF
C1486 VDD.n989 GND 0.03fF
C1487 VDD.n990 GND 0.02fF
C1488 VDD.n991 GND 0.02fF
C1489 VDD.n995 GND 0.28fF
C1490 VDD.n996 GND 0.28fF
C1491 VDD.n997 GND 0.01fF
C1492 VDD.n998 GND 0.02fF
C1493 VDD.n999 GND 0.04fF
C1494 VDD.n1000 GND 0.07fF
C1495 VDD.n1001 GND 0.26fF
C1496 VDD.n1002 GND 0.01fF
C1497 VDD.n1003 GND 0.01fF
C1498 VDD.n1004 GND 0.02fF
C1499 VDD.n1005 GND 0.17fF
C1500 VDD.n1006 GND 0.01fF
C1501 VDD.n1007 GND 0.02fF
C1502 VDD.n1008 GND 0.02fF
C1503 VDD.n1009 GND 0.15fF
C1504 VDD.n1010 GND 0.01fF
C1505 VDD.n1011 GND 0.02fF
C1506 VDD.n1012 GND 0.03fF
C1507 VDD.n1013 GND 0.08fF
C1508 VDD.n1014 GND 0.05fF
C1509 VDD.n1015 GND 0.01fF
C1510 VDD.n1016 GND 0.02fF
C1511 VDD.n1017 GND 0.03fF
C1512 VDD.n1018 GND 0.17fF
C1513 VDD.n1019 GND 0.01fF
C1514 VDD.n1020 GND 0.02fF
C1515 VDD.n1021 GND 0.02fF
C1516 VDD.n1022 GND 0.06fF
C1517 VDD.n1023 GND 0.25fF
C1518 VDD.n1024 GND 0.01fF
C1519 VDD.n1025 GND 0.01fF
C1520 VDD.n1026 GND 0.02fF
C1521 VDD.n1027 GND 0.28fF
C1522 VDD.n1028 GND 0.01fF
C1523 VDD.n1029 GND 0.02fF
C1524 VDD.n1030 GND 0.04fF
C1525 VDD.n1031 GND 0.27fF
C1526 VDD.n1032 GND 0.02fF
C1527 VDD.n1033 GND 0.02fF
C1528 VDD.n1034 GND 0.02fF
C1529 VDD.n1035 GND 0.06fF
C1530 VDD.n1036 GND 0.02fF
C1531 VDD.n1037 GND 0.02fF
C1532 VDD.n1038 GND 0.02fF
C1533 VDD.n1039 GND 0.02fF
C1534 VDD.n1040 GND 0.02fF
C1535 VDD.n1041 GND 0.02fF
C1536 VDD.n1042 GND 0.02fF
C1537 VDD.n1043 GND 0.02fF
C1538 VDD.n1044 GND 0.02fF
C1539 VDD.n1045 GND 0.02fF
C1540 VDD.n1046 GND 0.03fF
C1541 VDD.n1047 GND 0.02fF
C1542 VDD.n1048 GND 0.02fF
C1543 VDD.n1052 GND 0.28fF
C1544 VDD.n1053 GND 0.28fF
C1545 VDD.n1054 GND 0.01fF
C1546 VDD.n1055 GND 0.02fF
C1547 VDD.n1056 GND 0.04fF
C1548 VDD.n1057 GND 0.28fF
C1549 VDD.n1058 GND 0.01fF
C1550 VDD.n1059 GND 0.02fF
C1551 VDD.n1060 GND 0.02fF
C1552 VDD.n1061 GND 0.06fF
C1553 VDD.n1062 GND 0.23fF
C1554 VDD.n1063 GND 0.01fF
C1555 VDD.n1064 GND 0.01fF
C1556 VDD.n1065 GND 0.02fF
C1557 VDD.n1066 GND 0.17fF
C1558 VDD.n1067 GND 0.01fF
C1559 VDD.n1068 GND 0.02fF
C1560 VDD.n1069 GND 0.02fF
C1561 VDD.n1070 GND 0.08fF
C1562 VDD.n1071 GND 0.05fF
C1563 VDD.n1072 GND 0.16fF
C1564 VDD.n1073 GND 0.01fF
C1565 VDD.n1074 GND 0.02fF
C1566 VDD.n1075 GND 0.02fF
C1567 VDD.n1076 GND 0.15fF
C1568 VDD.n1077 GND 0.02fF
C1569 VDD.n1078 GND 0.02fF
C1570 VDD.n1079 GND 0.03fF
C1571 VDD.n1080 GND 0.15fF
C1572 VDD.n1081 GND 0.02fF
C1573 VDD.n1082 GND 0.02fF
C1574 VDD.n1083 GND 0.03fF
C1575 VDD.n1084 GND 0.17fF
C1576 VDD.n1085 GND 0.01fF
C1577 VDD.n1086 GND 0.08fF
C1578 VDD.n1087 GND 0.05fF
C1579 VDD.n1088 GND 0.02fF
C1580 VDD.n1089 GND 0.02fF
C1581 VDD.n1090 GND 0.17fF
C1582 VDD.n1091 GND 0.01fF
C1583 VDD.n1092 GND 0.02fF
C1584 VDD.n1093 GND 0.02fF
C1585 VDD.n1094 GND 0.23fF
C1586 VDD.n1095 GND 0.01fF
C1587 VDD.n1096 GND 0.07fF
C1588 VDD.n1097 GND 0.02fF
C1589 VDD.n1098 GND 0.28fF
C1590 VDD.n1099 GND 0.01fF
C1591 VDD.n1100 GND 0.02fF
C1592 VDD.n1101 GND 0.02fF
C1593 VDD.n1102 GND 0.28fF
C1594 VDD.n1103 GND 0.01fF
C1595 VDD.n1104 GND 0.02fF
C1596 VDD.n1105 GND 0.04fF
C1597 VDD.n1106 GND 0.27fF
C1598 VDD.n1107 GND 0.02fF
C1599 VDD.n1108 GND 0.02fF
C1600 VDD.n1109 GND 0.02fF
C1601 VDD.n1110 GND 0.06fF
C1602 VDD.n1111 GND 0.02fF
C1603 VDD.n1112 GND 0.02fF
C1604 VDD.n1113 GND 0.02fF
C1605 VDD.n1114 GND 0.02fF
C1606 VDD.n1115 GND 0.02fF
C1607 VDD.n1116 GND 0.02fF
C1608 VDD.n1117 GND 0.02fF
C1609 VDD.n1118 GND 0.02fF
C1610 VDD.n1119 GND 0.02fF
C1611 VDD.n1120 GND 0.02fF
C1612 VDD.n1121 GND 0.03fF
C1613 VDD.n1122 GND 0.02fF
C1614 VDD.n1123 GND 0.02fF
C1615 VDD.n1127 GND 0.28fF
C1616 VDD.n1128 GND 0.28fF
C1617 VDD.n1129 GND 0.01fF
C1618 VDD.n1130 GND 0.02fF
C1619 VDD.n1131 GND 0.04fF
C1620 VDD.n1132 GND 0.07fF
C1621 VDD.n1133 GND 0.26fF
C1622 VDD.n1134 GND 0.01fF
C1623 VDD.n1135 GND 0.01fF
C1624 VDD.n1136 GND 0.02fF
C1625 VDD.n1137 GND 0.17fF
C1626 VDD.n1138 GND 0.01fF
C1627 VDD.n1139 GND 0.02fF
C1628 VDD.n1140 GND 0.02fF
C1629 VDD.n1141 GND 0.15fF
C1630 VDD.n1142 GND 0.01fF
C1631 VDD.n1143 GND 0.02fF
C1632 VDD.n1144 GND 0.03fF
C1633 VDD.n1145 GND 0.08fF
C1634 VDD.n1146 GND 0.05fF
C1635 VDD.n1147 GND 0.01fF
C1636 VDD.n1148 GND 0.02fF
C1637 VDD.n1149 GND 0.03fF
C1638 VDD.n1150 GND 0.17fF
C1639 VDD.n1151 GND 0.01fF
C1640 VDD.n1152 GND 0.02fF
C1641 VDD.n1153 GND 0.02fF
C1642 VDD.n1154 GND 0.06fF
C1643 VDD.n1155 GND 0.25fF
C1644 VDD.n1156 GND 0.01fF
C1645 VDD.n1157 GND 0.01fF
C1646 VDD.n1158 GND 0.02fF
C1647 VDD.n1159 GND 0.28fF
C1648 VDD.n1160 GND 0.01fF
C1649 VDD.n1161 GND 0.02fF
C1650 VDD.n1162 GND 0.04fF
C1651 VDD.n1163 GND 0.27fF
C1652 VDD.n1164 GND 0.02fF
C1653 VDD.n1165 GND 0.02fF
C1654 VDD.n1166 GND 0.02fF
C1655 VDD.n1167 GND 0.06fF
C1656 VDD.n1168 GND 0.02fF
C1657 VDD.n1169 GND 0.02fF
C1658 VDD.n1170 GND 0.02fF
C1659 VDD.n1171 GND 0.02fF
C1660 VDD.n1172 GND 0.02fF
C1661 VDD.n1173 GND 0.02fF
C1662 VDD.n1174 GND 0.02fF
C1663 VDD.n1175 GND 0.02fF
C1664 VDD.n1176 GND 0.02fF
C1665 VDD.n1177 GND 0.02fF
C1666 VDD.n1178 GND 0.03fF
C1667 VDD.n1179 GND 0.02fF
C1668 VDD.n1180 GND 0.02fF
C1669 VDD.n1184 GND 0.28fF
C1670 VDD.n1185 GND 0.28fF
C1671 VDD.n1186 GND 0.01fF
C1672 VDD.n1187 GND 0.02fF
C1673 VDD.n1188 GND 0.04fF
C1674 VDD.n1189 GND 0.28fF
C1675 VDD.n1190 GND 0.01fF
C1676 VDD.n1191 GND 0.02fF
C1677 VDD.n1192 GND 0.02fF
C1678 VDD.n1193 GND 0.06fF
C1679 VDD.n1194 GND 0.23fF
C1680 VDD.n1195 GND 0.01fF
C1681 VDD.n1196 GND 0.01fF
C1682 VDD.n1197 GND 0.02fF
C1683 VDD.n1198 GND 0.17fF
C1684 VDD.n1199 GND 0.01fF
C1685 VDD.n1200 GND 0.02fF
C1686 VDD.n1201 GND 0.02fF
C1687 VDD.n1202 GND 0.08fF
C1688 VDD.n1203 GND 0.05fF
C1689 VDD.n1204 GND 0.16fF
C1690 VDD.n1205 GND 0.01fF
C1691 VDD.n1206 GND 0.02fF
C1692 VDD.n1207 GND 0.02fF
C1693 VDD.n1208 GND 0.15fF
C1694 VDD.n1209 GND 0.02fF
C1695 VDD.n1210 GND 0.02fF
C1696 VDD.n1211 GND 0.03fF
C1697 VDD.n1212 GND 0.15fF
C1698 VDD.n1213 GND 0.02fF
C1699 VDD.n1214 GND 0.02fF
C1700 VDD.n1215 GND 0.03fF
C1701 VDD.n1216 GND 0.17fF
C1702 VDD.n1217 GND 0.01fF
C1703 VDD.n1218 GND 0.08fF
C1704 VDD.n1219 GND 0.05fF
C1705 VDD.n1220 GND 0.02fF
C1706 VDD.n1221 GND 0.02fF
C1707 VDD.n1222 GND 0.17fF
C1708 VDD.n1223 GND 0.01fF
C1709 VDD.n1224 GND 0.02fF
C1710 VDD.n1225 GND 0.02fF
C1711 VDD.n1226 GND 0.23fF
C1712 VDD.n1227 GND 0.01fF
C1713 VDD.n1228 GND 0.07fF
C1714 VDD.n1229 GND 0.02fF
C1715 VDD.n1230 GND 0.28fF
C1716 VDD.n1231 GND 0.01fF
C1717 VDD.n1232 GND 0.02fF
C1718 VDD.n1233 GND 0.02fF
C1719 VDD.n1234 GND 0.28fF
C1720 VDD.n1235 GND 0.01fF
C1721 VDD.n1236 GND 0.02fF
C1722 VDD.n1237 GND 0.04fF
C1723 VDD.n1238 GND 0.32fF
C1724 VDD.n1239 GND 0.02fF
C1725 VDD.n1240 GND 0.02fF
C1726 VDD.n1241 GND 0.02fF
C1727 VDD.n1242 GND 0.06fF
C1728 VDD.n1243 GND 0.02fF
C1729 VDD.n1244 GND 0.02fF
C1730 VDD.n1245 GND 0.02fF
C1731 VDD.n1246 GND 0.02fF
C1732 VDD.n1247 GND 0.02fF
C1733 VDD.n1248 GND 0.02fF
C1734 VDD.n1249 GND 0.02fF
C1735 VDD.n1250 GND 0.02fF
C1736 VDD.n1251 GND 0.02fF
C1737 VDD.n1252 GND 0.02fF
C1738 VDD.n1253 GND 0.03fF
C1739 VDD.n1254 GND 0.02fF
C1740 VDD.n1255 GND 0.02fF
C1741 VDD.n1259 GND 0.28fF
C1742 VDD.n1260 GND 0.28fF
C1743 VDD.n1261 GND 0.01fF
C1744 VDD.n1262 GND 0.02fF
C1745 VDD.n1263 GND 0.04fF
C1746 VDD.n1264 GND 0.28fF
C1747 VDD.n1265 GND 0.01fF
C1748 VDD.n1266 GND 0.02fF
C1749 VDD.n1267 GND 0.02fF
C1750 VDD.n1268 GND 0.06fF
C1751 VDD.n1269 GND 0.23fF
C1752 VDD.n1270 GND 0.01fF
C1753 VDD.n1271 GND 0.01fF
C1754 VDD.n1272 GND 0.02fF
C1755 VDD.n1273 GND 0.17fF
C1756 VDD.n1274 GND 0.01fF
C1757 VDD.n1275 GND 0.02fF
C1758 VDD.n1276 GND 0.02fF
C1759 VDD.n1277 GND 0.08fF
C1760 VDD.n1278 GND 0.05fF
C1761 VDD.n1279 GND 0.16fF
C1762 VDD.n1280 GND 0.01fF
C1763 VDD.n1281 GND 0.02fF
C1764 VDD.n1282 GND 0.02fF
C1765 VDD.n1283 GND 0.15fF
C1766 VDD.n1284 GND 0.02fF
C1767 VDD.n1285 GND 0.02fF
C1768 VDD.n1286 GND 0.03fF
C1769 VDD.n1287 GND 0.15fF
C1770 VDD.n1288 GND 0.02fF
C1771 VDD.n1289 GND 0.02fF
C1772 VDD.n1290 GND 0.03fF
C1773 VDD.n1291 GND 0.17fF
C1774 VDD.n1292 GND 0.01fF
C1775 VDD.n1293 GND 0.08fF
C1776 VDD.n1294 GND 0.05fF
C1777 VDD.n1295 GND 0.02fF
C1778 VDD.n1296 GND 0.02fF
C1779 VDD.n1297 GND 0.17fF
C1780 VDD.n1298 GND 0.01fF
C1781 VDD.n1299 GND 0.02fF
C1782 VDD.n1300 GND 0.02fF
C1783 VDD.n1301 GND 0.23fF
C1784 VDD.n1302 GND 0.01fF
C1785 VDD.n1303 GND 0.07fF
C1786 VDD.n1304 GND 0.02fF
C1787 VDD.n1305 GND 0.28fF
C1788 VDD.n1306 GND 0.01fF
C1789 VDD.n1307 GND 0.02fF
C1790 VDD.n1308 GND 0.02fF
C1791 VDD.n1309 GND 0.28fF
C1792 VDD.n1310 GND 0.01fF
C1793 VDD.n1311 GND 0.02fF
C1794 VDD.n1312 GND 0.04fF
C1795 VDD.n1313 GND 0.27fF
C1796 VDD.n1314 GND 0.02fF
C1797 VDD.n1315 GND 0.02fF
C1798 VDD.n1316 GND 0.02fF
C1799 VDD.n1317 GND 0.06fF
C1800 VDD.n1318 GND 0.02fF
C1801 VDD.n1319 GND 0.02fF
C1802 VDD.n1320 GND 0.02fF
C1803 VDD.n1321 GND 0.02fF
C1804 VDD.n1322 GND 0.02fF
C1805 VDD.n1323 GND 0.02fF
C1806 VDD.n1324 GND 0.02fF
C1807 VDD.n1325 GND 0.02fF
C1808 VDD.n1326 GND 0.02fF
C1809 VDD.n1327 GND 0.02fF
C1810 VDD.n1328 GND 0.03fF
C1811 VDD.n1329 GND 0.02fF
C1812 VDD.n1330 GND 0.02fF
C1813 VDD.n1334 GND 0.28fF
C1814 VDD.n1335 GND 0.28fF
C1815 VDD.n1336 GND 0.01fF
C1816 VDD.n1337 GND 0.02fF
C1817 VDD.n1338 GND 0.04fF
C1818 VDD.n1339 GND 0.07fF
C1819 VDD.n1340 GND 0.26fF
C1820 VDD.n1341 GND 0.01fF
C1821 VDD.n1342 GND 0.01fF
C1822 VDD.n1343 GND 0.02fF
C1823 VDD.n1344 GND 0.17fF
C1824 VDD.n1345 GND 0.01fF
C1825 VDD.n1346 GND 0.02fF
C1826 VDD.n1347 GND 0.02fF
C1827 VDD.n1348 GND 0.15fF
C1828 VDD.n1349 GND 0.01fF
C1829 VDD.n1350 GND 0.02fF
C1830 VDD.n1351 GND 0.03fF
C1831 VDD.n1352 GND 0.08fF
C1832 VDD.n1353 GND 0.05fF
C1833 VDD.n1354 GND 0.01fF
C1834 VDD.n1355 GND 0.02fF
C1835 VDD.n1356 GND 0.03fF
C1836 VDD.n1357 GND 0.17fF
C1837 VDD.n1358 GND 0.01fF
C1838 VDD.n1359 GND 0.02fF
C1839 VDD.n1360 GND 0.02fF
C1840 VDD.n1361 GND 0.06fF
C1841 VDD.n1362 GND 0.25fF
C1842 VDD.n1363 GND 0.01fF
C1843 VDD.n1364 GND 0.01