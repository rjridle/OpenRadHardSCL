magic
tech sky130
magscale 1 2
timestamp 1645232802
<< nmos >>
rect 160 222 190 276
rect 54 192 190 222
rect 54 92 84 192
rect 160 92 190 192
rect 54 62 190 92
<< ndiff >>
rect -1 260 160 276
rect -1 226 9 260
rect 43 226 160 260
rect -1 222 160 226
rect 190 260 246 276
rect 190 226 202 260
rect 236 226 246 260
rect -1 189 54 222
rect -1 155 9 189
rect 43 155 54 189
rect -1 121 54 155
rect -1 87 9 121
rect 43 87 54 121
rect 84 156 160 192
rect 84 122 107 156
rect 141 122 160 156
rect 84 92 160 122
rect 190 189 246 226
rect 190 155 202 189
rect 236 155 246 189
rect 190 121 246 155
rect -1 62 54 87
rect 190 87 202 121
rect 236 87 246 121
rect 190 62 246 87
rect -1 50 246 62
rect -1 16 9 50
rect 43 16 110 50
rect 144 16 202 50
rect 236 16 246 50
rect -1 0 246 16
<< ndiffc >>
rect 9 226 43 260
rect 202 226 236 260
rect 9 155 43 189
rect 9 87 43 121
rect 107 122 141 156
rect 202 155 236 189
rect 202 87 236 121
rect 9 16 43 50
rect 110 16 144 50
rect 202 16 236 50
<< poly >>
rect 160 276 190 309
<< locali >>
rect 9 260 43 276
rect 9 189 43 226
rect 202 260 236 276
rect 202 189 236 226
rect 9 121 43 155
rect 107 156 141 172
rect 107 106 141 122
rect 202 121 236 155
rect 9 50 43 87
rect 202 50 236 87
rect 43 16 110 50
rect 144 16 202 50
rect 9 0 43 16
rect 202 0 236 16
<< end >>
