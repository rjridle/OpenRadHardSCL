* HSPICE file created from tmp.ext - technology: sky130A

.option scale=5000u

.subckt tmp Y A B VDD VSS
X0 VDD A a_217_1051 VDD sky130_fd_pr__pfet_01v8 ad=55600 pd=2278 as=0 ps=0 w=400 l=30 M=2
X1 Y a_217_1051 VDD VDD sky130_fd_pr__pfet_01v8 ad=11600 pd=458 as=0 ps=0 w=400 l=30 M=2
X2 VDD B a_217_1051 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=400 l=30 M=2
X3 VSS A a_112_101 VSS sky130_fd_pr__nfet_01v8 ad=53378 pd=1936 as=0 ps=0 w=598 l=30
X4 a_217_1051 B a_112_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=598 l=30
X5 Y a_217_1051 VSS VSS sky130_fd_pr__nfet_01v8 ad=7088 pd=312 as=0 ps=0 w=598 l=30
C0 VDD a_217_1051 2.25fF
.ends

** hspice subcircuit dictionary
