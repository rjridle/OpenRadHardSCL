* SPICE3 file created from AND2X1.ext - technology: sky130A

.subckt AND2X1 Y A B VDD VSS
X0 VDD A a_217_1050# VDD sky130_fd_pr__pfet_01v8 ad=2.78p pd=2.278u as=0p ps=0u w=2u l=0.15u M=2
X1 Y a_217_1050# VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8p pd=4.58u as=0p ps=0u w=2u l=0.15u M=2
X2 Y a_217_1050# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=1.3199p ps=9.67u w=3u l=0.15u
X3 VDD B a_217_1050# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X4 VSS A a_112_101# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X5 a_217_1050# B a_112_101# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
C0 a_217_1050# VDD 2.24fF
.ends
