magic
tech sky130A
magscale 1 2
timestamp 1647328314
<< nwell >>
rect 55 1505 89 1539
<< psubdiffcont >>
rect 55 13 89 47
<< nsubdiffcont >>
rect 55 1505 89 1539
<< viali >>
rect 55 1505 89 1539
rect 55 13 89 47
<< metal1 >>
rect 547 649 761 683
use invx1_pcell  invx1_pcell_0
timestamp 1647328248
transform 1 0 666 0 1 0
box -84 0 528 1575
use li1_M1_contact  li1_M1_contact_0
timestamp 1646004885
transform -1 0 518 0 -1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_1
timestamp 1646004885
transform 1 0 814 0 1 666
box -53 -33 29 33
use nor2x1_pcell  nor2x1_pcell_0
timestamp 1647327768
transform 1 0 0 0 1 0
box -84 0 750 1575
<< labels >>
rlabel metal1 72 30 72 30 1 VSS
port 1 n
rlabel metal1 72 1522 72 1522 1 VDD
port 2 n
<< end >>
