* SPICE3 file created from DFFSNQX1.ext - technology: sky130A

.subckt DFFSNQX1 Q D CLK SN VDD GND
X0 VDD.t17 D.t0 a_217_1050.t2 �A�U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X1 VDD.t57 a_1265_989.t5 a_1905_1050.t2 @�[�U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X2 Q.t4 a_1265_989.t6 VDD.t5 ����U sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X3 a_1905_1050.t5 a_217_1050.t5 VDD.t37  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X4 VDD.t43 a_343_411.t7 a_217_1050.t4 VDD.t42 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X5 VDD.t35 a_217_1050.t6 a_343_411.t6 쒤[ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X6 a_3473_1050.t1 Q.t7 VDD.t11 쒤[ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X7 GND a_217_1050.t7 a_757_103.t0 GND sky130_fd_pr__nfet_01v8 ad=1.0746p pd=9.42u as=0p ps=0u w=0u l=0u
X8 GND D.t1 a_112_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X9 VDD.t39 CLK.t1 a_343_411.t1  쒤[ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X10 a_3473_1050.t4 a_343_411.t8 VDD.t1 �뒤[ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X11 GND a_343_411.t9 a_3368_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X12 VDD.t41 a_1905_1050.t7 a_1265_989.t3  쒤[ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X13 VDD.t49 a_3473_1050.t5 Q.t6 �뒤[ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X14 VDD.t51 a_1265_989.t9 Q.t3  쒤[ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X15 VDD.t55 a_1265_989.t10 a_343_411.t3 �뒤[ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X16 a_217_1050.t1 D.t2 VDD.t15  쒤[ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X17 a_1905_1050.t1 a_1265_989.t11 VDD.t53 �뒤[ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X18 GND a_217_1050.t8 a_1719_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X19 VDD.t19 SN.t1 Q.t0  쒤[ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X20 a_1905_1050.t6 SN.t2 VDD.t45 �뒤[ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X21 GND a_1905_1050.t8 a_2702_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X22 a_217_1050.t3 a_343_411.t10 VDD.t27  쒤[ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X23 a_343_411.t5 a_217_1050.t9 VDD.t33 �뒤[ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X24 Q a_1265_989.t12 a_4294_210.t0 GND sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=0p ps=0u w=0u l=0u
X25 VDD.t31 a_217_1050.t10 a_1905_1050.t4  쒤[ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X26 a_343_411.t0 CLK.t3 VDD.t9 �뒤[ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X27 a_1265_989.t4 a_1905_1050.t9 VDD.t59  쒤[ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X28 VDD.t13 Q.t8 a_3473_1050.t0 �뒤[ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X29 VDD.t3 CLK.t4 a_1265_989.t0  쒤[ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X30 GND a_3473_1050.t7 a_4013_103.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X31 Q.t5 a_3473_1050.t6 VDD.t47 �뒤[ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X32 a_343_411.t2 a_1265_989.t13 VDD.t7  쒤[ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X33 VDD.t23 SN.t4 a_1905_1050.t0 �뒤[ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X34 a_1265_989.t1 CLK.t5 VDD.t29  쒤[ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X35 VDD.t21 a_343_411.t12 a_3473_1050.t3 �뒤[ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X36 Q.t1 SN.t5 VDD.t25  쒤[ sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
C0 CLK VDD 1.61fF
C1 Q SN 0.39fF
C2 Q VDD 2.82fF
C3 D VDD 0.33fF
C4 SN VDD 0.59fF
C5 SN CLK 0.09fF
R0 D.n0 D.t0 480.392
R1 D.n0 D.t2 403.272
R2 D.n1 D.t1 385.063
R3 D.n1 D.n0 143.429
R4 D.n2 D.n1 4.65
R5 D.n2 D 0.046
R6 a_217_1050.n5 a_217_1050.t6 512.525
R7 a_217_1050.n3 a_217_1050.t10 512.525
R8 a_217_1050.n5 a_217_1050.t9 371.139
R9 a_217_1050.n3 a_217_1050.t5 371.139
R10 a_217_1050.n4 a_217_1050.t8 305.674
R11 a_217_1050.n6 a_217_1050.t7 305.298
R12 a_217_1050.n6 a_217_1050.n5 291.648
R13 a_217_1050.n4 a_217_1050.n3 291.272
R14 a_217_1050.n10 a_217_1050.n8 256.385
R15 a_217_1050.n8 a_217_1050.n2 215.717
R16 a_217_1050.n2 a_217_1050.n1 157.964
R17 a_217_1050.n2 a_217_1050.n0 91.706
R18 a_217_1050.n10 a_217_1050.n9 15.218
R19 a_217_1050.n0 a_217_1050.t4 14.282
R20 a_217_1050.n0 a_217_1050.t3 14.282
R21 a_217_1050.n1 a_217_1050.t2 14.282
R22 a_217_1050.n1 a_217_1050.t1 14.282
R23 a_217_1050.n11 a_217_1050.n10 12.014
R24 a_217_1050.n7 a_217_1050.n4 8.138
R25 a_217_1050.n8 a_217_1050.n7 5.964
R26 a_217_1050.n7 a_217_1050.n6 4.65
R27 VDD.n296 VDD.n285 144.705
R28 VDD.n211 VDD.n204 144.705
R29 VDD.n371 VDD.n364 144.705
R30 VDD.n154 VDD.n147 144.705
R31 VDD.n97 VDD.n86 144.705
R32 VDD.n338 VDD.t55 143.754
R33 VDD.n413 VDD.t57 143.754
R34 VDD.n30 VDD.t51 143.754
R35 VDD.n263 VDD.t43 143.754
R36 VDD.n157 VDD.t3 143.754
R37 VDD.n100 VDD.t13 143.754
R38 VDD.n241 VDD.t15 135.17
R39 VDD.n303 VDD.t33 135.17
R40 VDD.n378 VDD.t37 135.17
R41 VDD.n179 VDD.t59 135.17
R42 VDD.n122 VDD.t1 135.17
R43 VDD.n60 VDD.t47 135.17
R44 VDD.n255 VDD.n254 129.472
R45 VDD.n313 VDD.n312 129.472
R46 VDD.n329 VDD.n328 129.472
R47 VDD.n388 VDD.n387 129.472
R48 VDD.n404 VDD.n403 129.472
R49 VDD.n167 VDD.n166 129.472
R50 VDD.n110 VDD.n109 129.472
R51 VDD.n51 VDD.n50 129.472
R52 VDD.n39 VDD.n38 129.472
R53 VDD.n82 VDD.n81 92.5
R54 VDD.n80 VDD.n79 92.5
R55 VDD.n78 VDD.n77 92.5
R56 VDD.n76 VDD.n75 92.5
R57 VDD.n84 VDD.n83 92.5
R58 VDD.n143 VDD.n142 92.5
R59 VDD.n141 VDD.n140 92.5
R60 VDD.n139 VDD.n138 92.5
R61 VDD.n137 VDD.n136 92.5
R62 VDD.n145 VDD.n144 92.5
R63 VDD.n200 VDD.n199 92.5
R64 VDD.n198 VDD.n197 92.5
R65 VDD.n196 VDD.n195 92.5
R66 VDD.n194 VDD.n193 92.5
R67 VDD.n202 VDD.n201 92.5
R68 VDD.n360 VDD.n359 92.5
R69 VDD.n358 VDD.n357 92.5
R70 VDD.n356 VDD.n355 92.5
R71 VDD.n354 VDD.n353 92.5
R72 VDD.n362 VDD.n361 92.5
R73 VDD.n281 VDD.n280 92.5
R74 VDD.n279 VDD.n278 92.5
R75 VDD.n277 VDD.n276 92.5
R76 VDD.n275 VDD.n274 92.5
R77 VDD.n283 VDD.n282 92.5
R78 VDD.n229 VDD.n228 92.5
R79 VDD.n227 VDD.n226 92.5
R80 VDD.n225 VDD.n224 92.5
R81 VDD.n223 VDD.n222 92.5
R82 VDD.n231 VDD.n230 92.5
R83 VDD.n14 VDD.n1 92.5
R84 VDD.n5 VDD.n4 92.5
R85 VDD.n7 VDD.n6 92.5
R86 VDD.n9 VDD.n8 92.5
R87 VDD.n11 VDD.n10 92.5
R88 VDD.n13 VDD.n12 92.5
R89 VDD.n21 VDD.n20 92.059
R90 VDD.n96 VDD.n95 92.059
R91 VDD.n153 VDD.n152 92.059
R92 VDD.n210 VDD.n209 92.059
R93 VDD.n370 VDD.n369 92.059
R94 VDD.n295 VDD.n294 92.059
R95 VDD.n237 VDD.n236 92.059
R96 VDD.n20 VDD.n16 67.194
R97 VDD.n20 VDD.n17 67.194
R98 VDD.n20 VDD.n18 67.194
R99 VDD.n20 VDD.n19 67.194
R100 VDD.n221 VDD.n220 44.141
R101 VDD.n352 VDD.n351 44.141
R102 VDD.n192 VDD.n191 44.141
R103 VDD.n135 VDD.n134 44.141
R104 VDD.n5 VDD.n3 44.141
R105 VDD.n351 VDD.n349 44.107
R106 VDD.n191 VDD.n189 44.107
R107 VDD.n134 VDD.n132 44.107
R108 VDD.n220 VDD.n218 44.107
R109 VDD.n3 VDD.n2 44.107
R110 VDD.n20 VDD.n15 41.052
R111 VDD.n90 VDD.n88 39.742
R112 VDD.n90 VDD.n89 39.742
R113 VDD.n92 VDD.n91 39.742
R114 VDD.n149 VDD.n148 39.742
R115 VDD.n206 VDD.n205 39.742
R116 VDD.n366 VDD.n365 39.742
R117 VDD.n233 VDD.n232 39.742
R118 VDD.n293 VDD.n290 39.742
R119 VDD.n293 VDD.n292 39.742
R120 VDD.n289 VDD.n288 39.742
R121 VDD.n134 VDD.n133 38
R122 VDD.n191 VDD.n190 38
R123 VDD.n351 VDD.n350 38
R124 VDD.n220 VDD.n219 38
R125 VDD.n349 VDD.n348 36.774
R126 VDD.n189 VDD.n188 36.774
R127 VDD.n132 VDD.n131 36.774
R128 VDD.n88 VDD.n87 36.774
R129 VDD.n292 VDD.n291 36.774
R130 VDD.n32  쒤[ 35.8
R131 VDD.n407 @�[�U 35.8
R132 VDD.n332 �뒤[ 35.8
R133 VDD.n56 �뒤[ 33.243
R134 VDD.n383 �r�U 33.243
R135 VDD.n308 �뒤[ 33.243
R136 VDD.n1 VDD.n0 30.923
R137 VDD.n95 VDD.n93 26.38
R138 VDD.n95 VDD.n92 26.38
R139 VDD.n95 VDD.n90 26.38
R140 VDD.n95 VDD.n94 26.38
R141 VDD.n152 VDD.n150 26.38
R142 VDD.n152 VDD.n149 26.38
R143 VDD.n152 VDD.n151 26.38
R144 VDD.n209 VDD.n207 26.38
R145 VDD.n209 VDD.n206 26.38
R146 VDD.n209 VDD.n208 26.38
R147 VDD.n369 VDD.n367 26.38
R148 VDD.n369 VDD.n366 26.38
R149 VDD.n369 VDD.n368 26.38
R150 VDD.n236 VDD.n234 26.38
R151 VDD.n236 VDD.n233 26.38
R152 VDD.n236 VDD.n235 26.38
R153 VDD.n294 VDD.n293 26.38
R154 VDD.n294 VDD.n289 26.38
R155 VDD.n294 VDD.n287 26.38
R156 VDD.n294 VDD.n286 26.38
R157 VDD.n239 VDD.n231 22.915
R158 VDD.n23 VDD.n14 22.915
R159 VDD.n105 �뒤[ 20.457
R160 VDD.n162  쒤[ 20.457
R161 VDD.n259 VDD.t42 20.457
R162 VDD.n118 �뒤[ 17.9
R163 VDD.n175  쒤[ 17.9
R164 VDD.n246  쒤[ 17.9
R165 VDD.n36 ����U 15.343
R166 VDD.n401 �뒤[ 15.343
R167 VDD.n326  쒤[ 15.343
R168 VDD.n231 VDD.n229 14.864
R169 VDD.n229 VDD.n227 14.864
R170 VDD.n227 VDD.n225 14.864
R171 VDD.n225 VDD.n223 14.864
R172 VDD.n223 VDD.n221 14.864
R173 VDD.n362 VDD.n360 14.864
R174 VDD.n360 VDD.n358 14.864
R175 VDD.n358 VDD.n356 14.864
R176 VDD.n356 VDD.n354 14.864
R177 VDD.n354 VDD.n352 14.864
R178 VDD.n202 VDD.n200 14.864
R179 VDD.n200 VDD.n198 14.864
R180 VDD.n198 VDD.n196 14.864
R181 VDD.n196 VDD.n194 14.864
R182 VDD.n194 VDD.n192 14.864
R183 VDD.n145 VDD.n143 14.864
R184 VDD.n143 VDD.n141 14.864
R185 VDD.n141 VDD.n139 14.864
R186 VDD.n139 VDD.n137 14.864
R187 VDD.n137 VDD.n135 14.864
R188 VDD.n84 VDD.n82 14.864
R189 VDD.n82 VDD.n80 14.864
R190 VDD.n80 VDD.n78 14.864
R191 VDD.n78 VDD.n76 14.864
R192 VDD.n76 VDD.n74 14.864
R193 VDD.n74 VDD.n73 14.864
R194 VDD.n283 VDD.n281 14.864
R195 VDD.n281 VDD.n279 14.864
R196 VDD.n279 VDD.n277 14.864
R197 VDD.n277 VDD.n275 14.864
R198 VDD.n275 VDD.n273 14.864
R199 VDD.n273 VDD.n272 14.864
R200 VDD.n14 VDD.n13 14.864
R201 VDD.n13 VDD.n11 14.864
R202 VDD.n11 VDD.n9 14.864
R203 VDD.n9 VDD.n7 14.864
R204 VDD.n7 VDD.n5 14.864
R205 VDD.n98 VDD.n85 14.864
R206 VDD.n155 VDD.n146 14.864
R207 VDD.n212 VDD.n203 14.864
R208 VDD.n372 VDD.n363 14.864
R209 VDD.n297 VDD.n284 14.864
R210 VDD.n254 VDD.t27 14.282
R211 VDD.n254 VDD.t17 14.282
R212 VDD.n312 VDD.t9 14.282
R213 VDD.n312 VDD.t35 14.282
R214 VDD.n328 VDD.t7 14.282
R215 VDD.n328 VDD.t39 14.282
R216 VDD.n387 VDD.t45 14.282
R217 VDD.n387 VDD.t31 14.282
R218 VDD.n403 VDD.t53 14.282
R219 VDD.n403 VDD.t23 14.282
R220 VDD.n166 VDD.t29 14.282
R221 VDD.n166 VDD.t41 14.282
R222 VDD.n109 VDD.t11 14.282
R223 VDD.n109 VDD.t21 14.282
R224 VDD.n50 VDD.t25 14.282
R225 VDD.n50 VDD.t49 14.282
R226 VDD.n38 VDD.t5 14.282
R227 VDD.n38 VDD.t19 14.282
R228 VDD.n52 �뒤[ 12.786
R229 VDD.n389  쒤[ 12.786
R230 VDD.n314 쒤[ 12.786
R231 VDD.n112 VDD.n110 9.083
R232 VDD.n169 VDD.n167 9.083
R233 VDD.n257 VDD.n255 9.083
R234 VDD.n23 VDD.n22 8.855
R235 VDD.n22 VDD.n21 8.855
R236 VDD.n26 VDD.n25 8.855
R237 VDD.n25 VDD.n24 8.855
R238 VDD.n30 VDD.n29 8.855
R239 VDD.n29 VDD.n28 8.855
R240 VDD.n34 VDD.n33 8.855
R241 VDD.n33 VDD.n32 8.855
R242 VDD.n40 VDD.n37 8.855
R243 VDD.n37 VDD.n36 8.855
R244 VDD.n44 VDD.n43 8.855
R245 VDD.n43 VDD.n42 8.855
R246 VDD.n48 VDD.n47 8.855
R247 VDD.n47 VDD.n46 8.855
R248 VDD.n54 VDD.n53 8.855
R249 VDD.n53 VDD.n52 8.855
R250 VDD.n58 VDD.n57 8.855
R251 VDD.n57 VDD.n56 8.855
R252 VDD.n63 VDD.n62 8.855
R253 VDD.n62 VDD.n61 8.855
R254 VDD.n67 VDD.n66 8.855
R255 VDD.n66 VDD.n65 8.855
R256 VDD.n71 VDD.n70 8.855
R257 VDD.n70 VDD.n69 8.855
R258 VDD.n98 VDD.n97 8.855
R259 VDD.n97 VDD.n96 8.855
R260 VDD.n103 VDD.n102 8.855
R261 VDD.n102 VDD.n101 8.855
R262 VDD.n107 VDD.n106 8.855
R263 VDD.n106 VDD.n105 8.855
R264 VDD.n112 VDD.n111 8.855
R265 VDD.n111 쒤[ 8.855
R266 VDD.n116 VDD.n115 8.855
R267 VDD.n115 VDD.n114 8.855
R268 VDD.n120 VDD.n119 8.855
R269 VDD.n119 VDD.n118 8.855
R270 VDD.n125 VDD.n124 8.855
R271 VDD.n124 VDD.n123 8.855
R272 VDD.n129 VDD.n128 8.855
R273 VDD.n128 VDD.n127 8.855
R274 VDD.n155 VDD.n154 8.855
R275 VDD.n154 VDD.n153 8.855
R276 VDD.n160 VDD.n159 8.855
R277 VDD.n159 VDD.n158 8.855
R278 VDD.n164 VDD.n163 8.855
R279 VDD.n163 VDD.n162 8.855
R280 VDD.n169 VDD.n168 8.855
R281 VDD.n168  쒤[ 8.855
R282 VDD.n173 VDD.n172 8.855
R283 VDD.n172 VDD.n171 8.855
R284 VDD.n177 VDD.n176 8.855
R285 VDD.n176 VDD.n175 8.855
R286 VDD.n182 VDD.n181 8.855
R287 VDD.n181 VDD.n180 8.855
R288 VDD.n186 VDD.n185 8.855
R289 VDD.n185 VDD.n184 8.855
R290 VDD.n212 VDD.n211 8.855
R291 VDD.n211 VDD.n210 8.855
R292 VDD.n216 VDD.n215 8.855
R293 VDD.n215 VDD.n214 8.855
R294 VDD.n413 VDD.n412 8.855
R295 VDD.n412 VDD.n411 8.855
R296 VDD.n409 VDD.n408 8.855
R297 VDD.n408 VDD.n407 8.855
R298 VDD.n405 VDD.n402 8.855
R299 VDD.n402 VDD.n401 8.855
R300 VDD.n399 VDD.n398 8.855
R301 VDD.n398 VDD.n397 8.855
R302 VDD.n395 VDD.n394 8.855
R303 VDD.n394 VDD.n393 8.855
R304 VDD.n391 VDD.n390 8.855
R305 VDD.n390 VDD.n389 8.855
R306 VDD.n385 VDD.n384 8.855
R307 VDD.n384 VDD.n383 8.855
R308 VDD.n381 VDD.n380 8.855
R309 VDD.n380 VDD.n379 8.855
R310 VDD.n376 VDD.n375 8.855
R311 VDD.n375 VDD.n374 8.855
R312 VDD.n372 VDD.n371 8.855
R313 VDD.n371 VDD.n370 8.855
R314 VDD.n346 VDD.n345 8.855
R315 VDD.n345 VDD.n344 8.855
R316 VDD.n342 VDD.n341 8.855
R317 VDD.n341 VDD.n340 8.855
R318 VDD.n338 VDD.n337 8.855
R319 VDD.n337 VDD.n336 8.855
R320 VDD.n334 VDD.n333 8.855
R321 VDD.n333 VDD.n332 8.855
R322 VDD.n330 VDD.n327 8.855
R323 VDD.n327 VDD.n326 8.855
R324 VDD.n324 VDD.n323 8.855
R325 VDD.n323 VDD.n322 8.855
R326 VDD.n320 VDD.n319 8.855
R327 VDD.n319 VDD.n318 8.855
R328 VDD.n316 VDD.n315 8.855
R329 VDD.n315 VDD.n314 8.855
R330 VDD.n310 VDD.n309 8.855
R331 VDD.n309 VDD.n308 8.855
R332 VDD.n306 VDD.n305 8.855
R333 VDD.n305 VDD.n304 8.855
R334 VDD.n301 VDD.n300 8.855
R335 VDD.n300 VDD.n299 8.855
R336 VDD.n297 VDD.n296 8.855
R337 VDD.n296 VDD.n295 8.855
R338 VDD.n270 VDD.n269 8.855
R339 VDD.n269 VDD.n268 8.855
R340 VDD.n266 VDD.n265 8.855
R341 VDD.n265 VDD.n264 8.855
R342 VDD.n261 VDD.n260 8.855
R343 VDD.n260 VDD.n259 8.855
R344 VDD.n257 VDD.n256 8.855
R345 VDD.n256  쒤[ 8.855
R346 VDD.n252 VDD.n251 8.855
R347 VDD.n251 VDD.n250 8.855
R348 VDD.n248 VDD.n247 8.855
R349 VDD.n247 VDD.n246 8.855
R350 VDD.n244 VDD.n243 8.855
R351 VDD.n243 VDD.n242 8.855
R352 VDD.n239 VDD.n238 8.855
R353 VDD.n238 VDD.n237 8.855
R354 VDD.n363 VDD.n362 8.051
R355 VDD.n203 VDD.n202 8.051
R356 VDD.n146 VDD.n145 8.051
R357 VDD.n85 VDD.n84 8.051
R358 VDD.n284 VDD.n283 8.051
R359 VDD.n46  쒤[ 7.671
R360 VDD.n393 �뒤[ 7.671
R361 VDD.n318 �뒤[ 7.671
R362 VDD.n54 VDD.n51 7.019
R363 VDD.n391 VDD.n388 7.019
R364 VDD.n316 VDD.n313 7.019
R365 VDD.n40 VDD.n39 6.606
R366 VDD.n405 VDD.n404 6.606
R367 VDD.n330 VDD.n329 6.606
R368 VDD.n42  쒤[ 5.114
R369 VDD.n397 �뒤[ 5.114
R370 VDD.n322  쒤[ 5.114
R371 VDD.n31 VDD.n30 4.65
R372 VDD.n35 VDD.n34 4.65
R373 VDD.n41 VDD.n40 4.65
R374 VDD.n45 VDD.n44 4.65
R375 VDD.n49 VDD.n48 4.65
R376 VDD.n55 VDD.n54 4.65
R377 VDD.n59 VDD.n58 4.65
R378 VDD.n64 VDD.n63 4.65
R379 VDD.n68 VDD.n67 4.65
R380 VDD.n72 VDD.n71 4.65
R381 VDD.n99 VDD.n98 4.65
R382 VDD.n104 VDD.n103 4.65
R383 VDD.n108 VDD.n107 4.65
R384 VDD.n113 VDD.n112 4.65
R385 VDD.n117 VDD.n116 4.65
R386 VDD.n121 VDD.n120 4.65
R387 VDD.n126 VDD.n125 4.65
R388 VDD.n130 VDD.n129 4.65
R389 VDD.n156 VDD.n155 4.65
R390 VDD.n161 VDD.n160 4.65
R391 VDD.n165 VDD.n164 4.65
R392 VDD.n170 VDD.n169 4.65
R393 VDD.n174 VDD.n173 4.65
R394 VDD.n178 VDD.n177 4.65
R395 VDD.n183 VDD.n182 4.65
R396 VDD.n187 VDD.n186 4.65
R397 VDD.n213 VDD.n212 4.65
R398 VDD.n217 VDD.n216 4.65
R399 VDD.n414 VDD.n413 4.65
R400 VDD.n410 VDD.n409 4.65
R401 VDD.n406 VDD.n405 4.65
R402 VDD.n400 VDD.n399 4.65
R403 VDD.n396 VDD.n395 4.65
R404 VDD.n392 VDD.n391 4.65
R405 VDD.n386 VDD.n385 4.65
R406 VDD.n382 VDD.n381 4.65
R407 VDD.n377 VDD.n376 4.65
R408 VDD.n373 VDD.n372 4.65
R409 VDD.n347 VDD.n346 4.65
R410 VDD.n343 VDD.n342 4.65
R411 VDD.n339 VDD.n338 4.65
R412 VDD.n335 VDD.n334 4.65
R413 VDD.n331 VDD.n330 4.65
R414 VDD.n325 VDD.n324 4.65
R415 VDD.n321 VDD.n320 4.65
R416 VDD.n317 VDD.n316 4.65
R417 VDD.n311 VDD.n310 4.65
R418 VDD.n307 VDD.n306 4.65
R419 VDD.n302 VDD.n301 4.65
R420 VDD.n298 VDD.n297 4.65
R421 VDD.n271 VDD.n270 4.65
R422 VDD.n267 VDD.n266 4.65
R423 VDD.n262 VDD.n261 4.65
R424 VDD.n258 VDD.n257 4.65
R425 VDD.n253 VDD.n252 4.65
R426 VDD.n249 VDD.n248 4.65
R427 VDD.n245 VDD.n244 4.65
R428 VDD.n240 VDD.n239 4.65
R429 VDD.n27 VDD.n23 2.933
R430 VDD.n125 VDD.n122 2.89
R431 VDD.n182 VDD.n179 2.89
R432 VDD.n244 VDD.n241 2.89
R433 VDD.n27 VDD.n26 2.844
R434 VDD.n114 �뒤[ 2.557
R435 VDD.n171  쒤[ 2.557
R436 VDD.n250 �A�U 2.557
R437 VDD.n103 VDD.n100 2.477
R438 VDD.n160 VDD.n157 2.477
R439 VDD.n266 VDD.n263 2.477
R440 VDD.n31 VDD.n27 1.063
R441 VDD.n63 VDD.n60 0.412
R442 VDD.n381 VDD.n378 0.412
R443 VDD.n306 VDD.n303 0.412
R444 VDD.n99 VDD.n72 0.29
R445 VDD.n156 VDD.n130 0.29
R446 VDD.n213 VDD.n187 0.29
R447 VDD.n373 VDD.n347 0.29
R448 VDD.n298 VDD.n271 0.29
R449 VDD.n240 VDD 0.207
R450 VDD.n49 VDD.n45 0.197
R451 VDD.n400 VDD.n396 0.197
R452 VDD.n325 VDD.n321 0.197
R453 VDD.n117 VDD.n113 0.181
R454 VDD.n174 VDD.n170 0.181
R455 VDD.n258 VDD.n253 0.181
R456 VDD.n35 VDD.n31 0.145
R457 VDD.n41 VDD.n35 0.145
R458 VDD.n45 VDD.n41 0.145
R459 VDD.n55 VDD.n49 0.145
R460 VDD.n59 VDD.n55 0.145
R461 VDD.n64 VDD.n59 0.145
R462 VDD.n68 VDD.n64 0.145
R463 VDD.n72 VDD.n68 0.145
R464 VDD.n104 VDD.n99 0.145
R465 VDD.n108 VDD.n104 0.145
R466 VDD.n113 VDD.n108 0.145
R467 VDD.n121 VDD.n117 0.145
R468 VDD.n126 VDD.n121 0.145
R469 VDD.n130 VDD.n126 0.145
R470 VDD.n161 VDD.n156 0.145
R471 VDD.n165 VDD.n161 0.145
R472 VDD.n170 VDD.n165 0.145
R473 VDD.n178 VDD.n174 0.145
R474 VDD.n183 VDD.n178 0.145
R475 VDD.n187 VDD.n183 0.145
R476 VDD.n217 VDD.n213 0.145
R477 VDD.n414 VDD.n410 0.145
R478 VDD.n410 VDD.n406 0.145
R479 VDD.n406 VDD.n400 0.145
R480 VDD.n396 VDD.n392 0.145
R481 VDD.n392 VDD.n386 0.145
R482 VDD.n386 VDD.n382 0.145
R483 VDD.n382 VDD.n377 0.145
R484 VDD.n377 VDD.n373 0.145
R485 VDD.n347 VDD.n343 0.145
R486 VDD.n343 VDD.n339 0.145
R487 VDD.n339 VDD.n335 0.145
R488 VDD.n335 VDD.n331 0.145
R489 VDD.n331 VDD.n325 0.145
R490 VDD.n321 VDD.n317 0.145
R491 VDD.n317 VDD.n311 0.145
R492 VDD.n311 VDD.n307 0.145
R493 VDD.n307 VDD.n302 0.145
R494 VDD.n302 VDD.n298 0.145
R495 VDD.n271 VDD.n267 0.145
R496 VDD.n267 VDD.n262 0.145
R497 VDD.n262 VDD.n258 0.145
R498 VDD.n253 VDD.n249 0.145
R499 VDD.n249 VDD.n245 0.145
R500 VDD.n245 VDD.n240 0.145
R501 VDD VDD.n414 0.137
R502 VDD VDD.n217 0.008
R503 a_1265_989.n6 a_1265_989.t11 454.685
R504 a_1265_989.n8 a_1265_989.t13 454.685
R505 a_1265_989.n4 a_1265_989.t6 454.685
R506 a_1265_989.n6 a_1265_989.t5 428.979
R507 a_1265_989.n8 a_1265_989.t10 428.979
R508 a_1265_989.n4 a_1265_989.t9 428.979
R509 a_1265_989.n7 a_1265_989.t7 339.542
R510 a_1265_989.n9 a_1265_989.t8 339.542
R511 a_1265_989.n5 a_1265_989.t12 339.542
R512 a_1265_989.n14 a_1265_989.n12 333.44
R513 a_1265_989.n3 a_1265_989.n2 157.964
R514 a_1265_989.n7 a_1265_989.n6 143.429
R515 a_1265_989.n9 a_1265_989.n8 143.429
R516 a_1265_989.n5 a_1265_989.n4 143.429
R517 a_1265_989.n12 a_1265_989.n3 132.141
R518 a_1265_989.n3 a_1265_989.n1 91.706
R519 a_1265_989.n15 a_1265_989.n0 55.263
R520 a_1265_989.n14 a_1265_989.n13 30
R521 a_1265_989.n15 a_1265_989.n14 23.684
R522 a_1265_989.n1 a_1265_989.t0 14.282
R523 a_1265_989.n1 a_1265_989.t1 14.282
R524 a_1265_989.n2 a_1265_989.t3 14.282
R525 a_1265_989.n2 a_1265_989.t4 14.282
R526 a_1265_989.n11 a_1265_989.n5 10.046
R527 a_1265_989.n10 a_1265_989.n9 8.141
R528 a_1265_989.n10 a_1265_989.n7 4.65
R529 a_1265_989.n12 a_1265_989.n11 4.65
R530 a_1265_989.n11 a_1265_989.n10 2.947
R531 a_1905_1050.n0 a_1905_1050.t7 480.392
R532 a_1905_1050.n0 a_1905_1050.t9 403.272
R533 a_1905_1050.n1 a_1905_1050.t8 301.486
R534 a_1905_1050.n6 a_1905_1050.n5 252.498
R535 a_1905_1050.n10 a_1905_1050.n6 234.917
R536 a_1905_1050.n1 a_1905_1050.n0 227.006
R537 a_1905_1050.n9 a_1905_1050.n8 161.352
R538 a_1905_1050.n9 a_1905_1050.n7 95.095
R539 a_1905_1050.n11 a_1905_1050.n10 95.094
R540 a_1905_1050.n10 a_1905_1050.n9 66.258
R541 a_1905_1050.n5 a_1905_1050.n4 30
R542 a_1905_1050.n3 a_1905_1050.n2 24.383
R543 a_1905_1050.n5 a_1905_1050.n3 23.684
R544 a_1905_1050.n7 a_1905_1050.t0 14.282
R545 a_1905_1050.n7 a_1905_1050.t6 14.282
R546 a_1905_1050.n8 a_1905_1050.t4 14.282
R547 a_1905_1050.n8 a_1905_1050.t5 14.282
R548 a_1905_1050.t2 a_1905_1050.n11 14.282
R549 a_1905_1050.n11 a_1905_1050.t1 14.282
R550 a_1905_1050.n6 a_1905_1050.n1 10.615
R551 Q.n10 Q.t8 472.359
R552 Q.n10 Q.t7 384.527
R553 Q.n11 Q.t9 314.896
R554 Q.n9 Q.n8 308.216
R555 Q.n11 Q.n10 182.814
R556 Q.n9 Q.n4 179.199
R557 Q.n3 Q.n2 161.352
R558 Q.n4 Q.n0 95.095
R559 Q.n3 Q.n1 95.095
R560 Q.n4 Q.n3 66.258
R561 Q.n8 Q.n7 30
R562 Q.n6 Q.n5 24.383
R563 Q.n8 Q.n6 23.684
R564 Q.n0 Q.t3 14.282
R565 Q.n0 Q.t4 14.282
R566 Q.n1 Q.t0 14.282
R567 Q.n1 Q.t1 14.282
R568 Q.n2 Q.t6 14.282
R569 Q.n2 Q.t5 14.282
R570 Q Q.n11 8.639
R571 Q.n12 Q.n9 4.65
R572 Q.n12 Q 0.046
R573 CLK.n0 CLK.t4 472.359
R574 CLK.n2 CLK.t1 459.505
R575 CLK.n3 CLK.t2 399.181
R576 CLK.n1 CLK.t0 398.558
R577 CLK.n2 CLK.t3 384.527
R578 CLK.n0 CLK.t5 384.527
R579 CLK.n3 CLK.n2 33.832
R580 CLK.n1 CLK.n0 32.394
R581 CLK.n4 CLK.n1 8.215
R582 CLK.n4 CLK.n3 2.079
R583 CLK.n4 CLK 0.046
R584 a_2702_101.n10 a_2702_101.n9 93.333
R585 a_2702_101.n12 a_2702_101.n11 68.43
R586 a_2702_101.n3 a_2702_101.n2 51.907
R587 a_2702_101.n3 a_2702_101.n1 51.594
R588 a_2702_101.t0 a_2702_101.n3 38.864
R589 a_2702_101.n7 a_2702_101.n6 38.626
R590 a_2702_101.n6 a_2702_101.n5 35.955
R591 a_2702_101.t1 a_2702_101.n8 8.137
R592 a_2702_101.t0 a_2702_101.n0 6.109
R593 a_2702_101.t1 a_2702_101.n7 4.864
R594 a_2702_101.t0 a_2702_101.n4 3.871
R595 a_2702_101.t0 a_2702_101.n13 2.535
R596 a_2702_101.n13 a_2702_101.t1 1.145
R597 a_2702_101.t1 a_2702_101.n12 0.763
R598 a_2702_101.n12 a_2702_101.n10 0.185
R599 GND.n141 GND.n140 237.558
R600 GND.n105 GND.n104 237.558
R601 GND.n186 GND.n185 237.558
R602 GND.n75 GND.n74 237.558
R603 GND.n43 GND.n42 237.558
R604 GND.n40 GND.n39 210.82
R605 GND.n143 GND.n142 210.82
R606 GND.n188 GND.n187 210.82
R607 GND.n102 GND.n101 210.82
R608 GND.n72 GND.n71 210.82
R609 GND.n91 GND.n90 172.612
R610 GND.n61 GND.n60 166.605
R611 GND.n30 GND.n29 152.358
R612 GND.n200 GND.n199 152.358
R613 GND.n155 GND.n154 152.358
R614 GND.n121 GND.n120 151.605
R615 GND.n29 GND.n28 28.421
R616 GND.n199 GND.n198 28.421
R617 GND.n154 GND.n153 28.421
R618 GND.n120 GND.n119 28.421
R619 GND.n29 GND.n27 25.263
R620 GND.n199 GND.n197 25.263
R621 GND.n154 GND.n152 25.263
R622 GND.n120 GND.n118 25.263
R623 GND.n27 GND.n26 24.383
R624 GND.n197 GND.n196 24.383
R625 GND.n152 GND.n151 24.383
R626 GND.n118 GND.n117 24.383
R627 GND.n60 GND.n58 23.03
R628 GND.n41 GND.n40 18.953
R629 GND.n144 GND.n143 18.953
R630 GND.n189 GND.n188 18.953
R631 GND.n103 GND.n102 18.953
R632 GND.n73 GND.n72 18.953
R633 GND.n44 GND.n41 14.864
R634 GND.n76 GND.n73 14.864
R635 GND.n106 GND.n103 14.864
R636 GND.n190 GND.n189 14.864
R637 GND.n145 GND.n144 14.864
R638 GND.n115 GND.n114 9.154
R639 GND.n123 GND.n122 9.154
R640 GND.n126 GND.n125 9.154
R641 GND.n129 GND.n128 9.154
R642 GND.n132 GND.n131 9.154
R643 GND.n135 GND.n134 9.154
R644 GND.n138 GND.n137 9.154
R645 GND.n145 GND.n141 9.154
R646 GND.n148 GND.n147 9.154
R647 GND.n156 GND.n150 9.154
R648 GND.n159 GND.n158 9.154
R649 GND.n162 GND.n161 9.154
R650 GND.n165 GND.n164 9.154
R651 GND.n168 GND.n167 9.154
R652 GND.n171 GND.n170 9.154
R653 GND.n174 GND.n173 9.154
R654 GND.n177 GND.n176 9.154
R655 GND.n180 GND.n179 9.154
R656 GND.n183 GND.n182 9.154
R657 GND.n190 GND.n186 9.154
R658 GND.n193 GND.n192 9.154
R659 GND.n201 GND.n195 9.154
R660 GND.n204 GND.n203 9.154
R661 GND.n207 GND.n206 9.154
R662 GND.n210 GND.n209 9.154
R663 GND.n213 GND.n212 9.154
R664 GND.n216 GND.n215 9.154
R665 GND.n219 GND.n218 9.154
R666 GND.n222 GND.n221 9.154
R667 GND.n109 GND.n108 9.154
R668 GND.n106 GND.n105 9.154
R669 GND.n99 GND.n98 9.154
R670 GND.n96 GND.n95 9.154
R671 GND.n93 GND.n92 9.154
R672 GND.n88 GND.n87 9.154
R673 GND.n85 GND.n84 9.154
R674 GND.n82 GND.n81 9.154
R675 GND.n79 GND.n78 9.154
R676 GND.n76 GND.n75 9.154
R677 GND.n69 GND.n68 9.154
R678 GND.n66 GND.n65 9.154
R679 GND.n63 GND.n62 9.154
R680 GND.n56 GND.n55 9.154
R681 GND.n53 GND.n52 9.154
R682 GND.n50 GND.n49 9.154
R683 GND.n47 GND.n46 9.154
R684 GND.n44 GND.n43 9.154
R685 GND.n37 GND.n36 9.154
R686 GND.n34 GND.n33 9.154
R687 GND.n31 GND.n25 9.154
R688 GND.n23 GND.n22 9.154
R689 GND.n20 GND.n19 9.154
R690 GND.n17 GND.n16 9.154
R691 GND.n14 GND.n13 9.154
R692 GND.n11 GND.n10 9.154
R693 GND.n8 GND.n7 9.154
R694 GND.n5 GND.n4 9.154
R695 GND.n2 GND.n1 9.154
R696 GND.n60 GND.n59 8.128
R697 GND.n113 GND.n112 4.65
R698 GND.n6 GND.n5 4.65
R699 GND.n9 GND.n8 4.65
R700 GND.n12 GND.n11 4.65
R701 GND.n15 GND.n14 4.65
R702 GND.n18 GND.n17 4.65
R703 GND.n21 GND.n20 4.65
R704 GND.n24 GND.n23 4.65
R705 GND.n32 GND.n31 4.65
R706 GND.n35 GND.n34 4.65
R707 GND.n38 GND.n37 4.65
R708 GND.n45 GND.n44 4.65
R709 GND.n48 GND.n47 4.65
R710 GND.n51 GND.n50 4.65
R711 GND.n54 GND.n53 4.65
R712 GND.n57 GND.n56 4.65
R713 GND.n64 GND.n63 4.65
R714 GND.n67 GND.n66 4.65
R715 GND.n70 GND.n69 4.65
R716 GND.n77 GND.n76 4.65
R717 GND.n80 GND.n79 4.65
R718 GND.n83 GND.n82 4.65
R719 GND.n86 GND.n85 4.65
R720 GND.n89 GND.n88 4.65
R721 GND.n94 GND.n93 4.65
R722 GND.n97 GND.n96 4.65
R723 GND.n100 GND.n99 4.65
R724 GND.n107 GND.n106 4.65
R725 GND.n110 GND.n109 4.65
R726 GND.n223 GND.n222 4.65
R727 GND.n220 GND.n219 4.65
R728 GND.n217 GND.n216 4.65
R729 GND.n214 GND.n213 4.65
R730 GND.n211 GND.n210 4.65
R731 GND.n208 GND.n207 4.65
R732 GND.n205 GND.n204 4.65
R733 GND.n202 GND.n201 4.65
R734 GND.n194 GND.n193 4.65
R735 GND.n191 GND.n190 4.65
R736 GND.n184 GND.n183 4.65
R737 GND.n181 GND.n180 4.65
R738 GND.n178 GND.n177 4.65
R739 GND.n175 GND.n174 4.65
R740 GND.n172 GND.n171 4.65
R741 GND.n169 GND.n168 4.65
R742 GND.n166 GND.n165 4.65
R743 GND.n163 GND.n162 4.65
R744 GND.n160 GND.n159 4.65
R745 GND.n157 GND.n156 4.65
R746 GND.n149 GND.n148 4.65
R747 GND.n146 GND.n145 4.65
R748 GND.n139 GND.n138 4.65
R749 GND.n136 GND.n135 4.65
R750 GND.n133 GND.n132 4.65
R751 GND.n130 GND.n129 4.65
R752 GND.n127 GND.n126 4.65
R753 GND.n124 GND.n123 4.65
R754 GND.n116 GND.n115 4.65
R755 GND.n63 GND.n61 4.129
R756 GND.n93 GND.n91 4.129
R757 GND.n123 GND.n121 4.129
R758 GND.n3 GND.n0 3.407
R759 GND.n3 GND.n2 2.844
R760 GND.n6 GND.n3 1.063
R761 GND.n112 GND.n111 0.474
R762 GND.n45 GND.n38 0.29
R763 GND.n77 GND.n70 0.29
R764 GND.n107 GND.n100 0.29
R765 GND.n191 GND.n184 0.29
R766 GND.n146 GND.n139 0.29
R767 GND.n113 GND 0.207
R768 GND.n31 GND.n30 0.206
R769 GND.n201 GND.n200 0.206
R770 GND.n156 GND.n155 0.206
R771 GND.n18 GND.n15 0.197
R772 GND.n214 GND.n211 0.197
R773 GND.n169 GND.n166 0.197
R774 GND.n57 GND.n54 0.181
R775 GND.n89 GND.n86 0.181
R776 GND.n130 GND.n127 0.181
R777 GND.n9 GND.n6 0.145
R778 GND.n12 GND.n9 0.145
R779 GND.n15 GND.n12 0.145
R780 GND.n21 GND.n18 0.145
R781 GND.n24 GND.n21 0.145
R782 GND.n32 GND.n24 0.145
R783 GND.n35 GND.n32 0.145
R784 GND.n38 GND.n35 0.145
R785 GND.n48 GND.n45 0.145
R786 GND.n51 GND.n48 0.145
R787 GND.n54 GND.n51 0.145
R788 GND.n64 GND.n57 0.145
R789 GND.n67 GND.n64 0.145
R790 GND.n70 GND.n67 0.145
R791 GND.n80 GND.n77 0.145
R792 GND.n83 GND.n80 0.145
R793 GND.n86 GND.n83 0.145
R794 GND.n94 GND.n89 0.145
R795 GND.n97 GND.n94 0.145
R796 GND.n100 GND.n97 0.145
R797 GND.n110 GND.n107 0.145
R798 GND.n223 GND.n220 0.145
R799 GND.n220 GND.n217 0.145
R800 GND.n217 GND.n214 0.145
R801 GND.n211 GND.n208 0.145
R802 GND.n208 GND.n205 0.145
R803 GND.n205 GND.n202 0.145
R804 GND.n202 GND.n194 0.145
R805 GND.n194 GND.n191 0.145
R806 GND.n184 GND.n181 0.145
R807 GND.n181 GND.n178 0.145
R808 GND.n178 GND.n175 0.145
R809 GND.n175 GND.n172 0.145
R810 GND.n172 GND.n169 0.145
R811 GND.n166 GND.n163 0.145
R812 GND.n163 GND.n160 0.145
R813 GND.n160 GND.n157 0.145
R814 GND.n157 GND.n149 0.145
R815 GND.n149 GND.n146 0.145
R816 GND.n139 GND.n136 0.145
R817 GND.n136 GND.n133 0.145
R818 GND.n133 GND.n130 0.145
R819 GND.n127 GND.n124 0.145
R820 GND.n124 GND.n116 0.145
R821 GND.n116 GND.n113 0.145
R822 GND GND.n223 0.137
R823 GND GND.n110 0.008
R824 SN.n2 SN.t4 479.223
R825 SN.n0 SN.t1 479.223
R826 SN.n2 SN.t2 375.52
R827 SN.n0 SN.t5 375.52
R828 SN.n3 SN.n2 252.188
R829 SN.n1 SN.n0 252.188
R830 SN.n3 SN.t3 231.854
R831 SN.n1 SN.t0 231.854
R832 SN.n4 SN.n1 13.038
R833 SN.n4 SN.n3 4.65
R834 SN.n4 SN 0.046
R835 a_4013_103.t0 a_4013_103.n7 59.616
R836 a_4013_103.n4 a_4013_103.n2 54.496
R837 a_4013_103.n4 a_4013_103.n3 54.496
R838 a_4013_103.n1 a_4013_103.n0 24.679
R839 a_4013_103.n6 a_4013_103.n4 7.859
R840 a_4013_103.t0 a_4013_103.n1 7.505
R841 a_4013_103.t0 a_4013_103.n6 3.034
R842 a_4013_103.n6 a_4013_103.n5 0.443
R843 a_4294_210.n8 a_4294_210.n6 185.173
R844 a_4294_210.t0 a_4294_210.n8 75.765
R845 a_4294_210.n3 a_4294_210.n1 74.827
R846 a_4294_210.n3 a_4294_210.n2 27.476
R847 a_4294_210.n6 a_4294_210.n5 22.349
R848 a_4294_210.t0 a_4294_210.n10 20.241
R849 a_4294_210.t0 a_4294_210.n3 13.984
R850 a_4294_210.n10 a_4294_210.n9 13.494
R851 a_4294_210.n6 a_4294_210.n4 8.443
R852 a_4294_210.t0 a_4294_210.n0 8.137
R853 a_4294_210.n8 a_4294_210.n7 1.505
R854 a_343_411.n1 a_343_411.t12 480.392
R855 a_343_411.n3 a_343_411.t7 472.359
R856 a_343_411.n2 a_343_411.t9 412.921
R857 a_343_411.n1 a_343_411.t8 403.272
R858 a_343_411.n3 a_343_411.t10 384.527
R859 a_343_411.n4 a_343_411.t11 370.613
R860 a_343_411.n10 a_343_411.n9 363.578
R861 a_343_411.n13 a_343_411.n12 161.352
R862 a_343_411.n4 a_343_411.n3 127.096
R863 a_343_411.n11 a_343_411.n10 123.126
R864 a_343_411.n2 a_343_411.n1 115.571
R865 a_343_411.n11 a_343_411.n0 95.095
R866 a_343_411.n14 a_343_411.n13 95.094
R867 a_343_411.n13 a_343_411.n11 66.258
R868 a_343_411.n9 a_343_411.n8 30
R869 a_343_411.n7 a_343_411.n6 24.383
R870 a_343_411.n9 a_343_411.n7 23.684
R871 a_343_411.n0 a_343_411.t3 14.282
R872 a_343_411.n0 a_343_411.t2 14.282
R873 a_343_411.n12 a_343_411.t6 14.282
R874 a_343_411.n12 a_343_411.t5 14.282
R875 a_343_411.t1 a_343_411.n14 14.282
R876 a_343_411.n14 a_343_411.t0 14.282
R877 a_343_411.n5 a_343_411.n2 11.954
R878 a_343_411.n5 a_343_411.n4 8.682
R879 a_343_411.n10 a_343_411.n5 4.65
R880 a_3473_1050.n0 a_3473_1050.t5 512.525
R881 a_3473_1050.n0 a_3473_1050.t6 371.139
R882 a_3473_1050.n1 a_3473_1050.t7 333.533
R883 a_3473_1050.n6 a_3473_1050.n5 277.722
R884 a_3473_1050.n1 a_3473_1050.n0 263.413
R885 a_3473_1050.n8 a_3473_1050.n6 187.858
R886 a_3473_1050.n8 a_3473_1050.n7 157.964
R887 a_3473_1050.n9 a_3473_1050.n8 91.705
R888 a_3473_1050.n5 a_3473_1050.n4 30
R889 a_3473_1050.n3 a_3473_1050.n2 24.383
R890 a_3473_1050.n5 a_3473_1050.n3 23.684
R891 a_3473_1050.n7 a_3473_1050.t3 14.282
R892 a_3473_1050.n7 a_3473_1050.t4 14.282
R893 a_3473_1050.n9 a_3473_1050.t0 14.282
R894 a_3473_1050.t1 a_3473_1050.n9 14.282
R895 a_3473_1050.n6 a_3473_1050.n1 10.615
R896 a_2000_210.n9 a_2000_210.n7 171.558
R897 a_2000_210.t0 a_2000_210.n9 75.765
R898 a_2000_210.n3 a_2000_210.n1 74.827
R899 a_2000_210.n3 a_2000_210.n2 27.476
R900 a_2000_210.n7 a_2000_210.n6 27.2
R901 a_2000_210.n5 a_2000_210.n4 23.498
R902 a_2000_210.n7 a_2000_210.n5 22.4
R903 a_2000_210.t0 a_2000_210.n11 20.241
R904 a_2000_210.t0 a_2000_210.n3 13.984
R905 a_2000_210.n11 a_2000_210.n10 13.494
R906 a_2000_210.t0 a_2000_210.n0 8.137
R907 a_2000_210.n9 a_2000_210.n8 1.505
R908 a_1038_210.n10 a_1038_210.n8 171.558
R909 a_1038_210.n8 a_1038_210.t1 75.764
R910 a_1038_210.n3 a_1038_210.n2 27.476
R911 a_1038_210.n10 a_1038_210.n9 27.2
R912 a_1038_210.n11 a_1038_210.n0 23.498
R913 a_1038_210.n11 a_1038_210.n10 22.4
R914 a_1038_210.t1 a_1038_210.n5 20.241
R915 a_1038_210.n7 a_1038_210.n6 19.952
R916 a_1038_210.t1 a_1038_210.n3 13.984
R917 a_1038_210.n5 a_1038_210.n4 13.494
R918 a_1038_210.t1 a_1038_210.n1 7.04
R919 a_1038_210.n8 a_1038_210.n7 1.505
R920 a_757_103.t0 a_757_103.n7 59.616
R921 a_757_103.n4 a_757_103.n2 54.496
R922 a_757_103.n4 a_757_103.n3 54.496
R923 a_757_103.n1 a_757_103.n0 24.679
R924 a_757_103.t0 a_757_103.n1 7.505
R925 a_757_103.n6 a_757_103.n5 2.455
R926 a_757_103.n6 a_757_103.n4 0.636
R927 a_757_103.t0 a_757_103.n6 0.246
R928 a_112_101.n11 a_112_101.n10 68.43
R929 a_112_101.n3 a_112_101.n2 62.817
R930 a_112_101.n7 a_112_101.n6 38.626
R931 a_112_101.n6 a_112_101.n5 35.955
R932 a_112_101.n3 a_112_101.n1 26.202
R933 a_112_101.t0 a_112_101.n3 19.737
R934 a_112_101.t1 a_112_101.n8 8.137
R935 a_112_101.t0 a_112_101.n4 7.273
R936 a_112_101.t0 a_112_101.n0 6.109
R937 a_112_101.t1 a_112_101.n7 4.864
R938 a_112_101.t0 a_112_101.n12 2.074
R939 a_112_101.n12 a_112_101.t1 0.937
R940 a_112_101.t1 a_112_101.n11 0.763
R941 a_112_101.n11 a_112_101.n9 0.185
R942 a_3368_101.n3 a_3368_101.n1 42.788
R943 a_3368_101.t0 a_3368_101.n0 8.137
R944 a_3368_101.n3 a_3368_101.n2 4.665
R945 a_3368_101.t0 a_3368_101.n3 0.06
R946 a_1719_103.n5 a_1719_103.n4 66.708
R947 a_1719_103.n2 a_1719_103.n0 25.439
R948 a_1719_103.n5 a_1719_103.n3 19.496
R949 a_1719_103.t0 a_1719_103.n5 13.756
R950 a_1719_103.n2 a_1719_103.n1 2.455
R951 a_1719_103.t0 a_1719_103.n2 0.246
C6 SN GND 1.44fF
C7 VDD GND 8.00fF
C8 a_1719_103.n0 GND 0.11fF
C9 a_1719_103.n1 GND 0.04fF
C10 a_1719_103.n2 GND 0.03fF
C11 a_1719_103.n3 GND 0.07fF
C12 a_1719_103.n4 GND 0.08fF
C13 a_1719_103.n5 GND 0.03fF
C14 a_3368_101.n0 GND 0.05fF
C15 a_3368_101.n1 GND 0.12fF
C16 a_3368_101.n2 GND 0.04fF
C17 a_3368_101.n3 GND 0.17fF
C18 a_112_101.n0 GND 0.02fF
C19 a_112_101.n1 GND 0.09fF
C20 a_112_101.n2 GND 0.08fF
C21 a_112_101.n3 GND 0.03fF
C22 a_112_101.n4 GND 0.01fF
C23 a_112_101.n5 GND 0.04fF
C24 a_112_101.n6 GND 0.04fF
C25 a_112_101.n7 GND 0.02fF
C26 a_112_101.n8 GND 0.05fF
C27 a_112_101.n9 GND 0.14fF
C28 a_112_101.n10 GND 0.08fF
C29 a_112_101.n11 GND 0.08fF
C30 a_112_101.t1 GND 0.22fF
C31 a_112_101.n12 GND 0.01fF
C32 a_757_103.n0 GND 0.08fF
C33 a_757_103.n1 GND 0.07fF
C34 a_757_103.n2 GND 0.04fF
C35 a_757_103.n3 GND 0.06fF
C36 a_757_103.n4 GND 0.03fF
C37 a_757_103.n5 GND 0.04fF
C38 a_757_103.n7 GND 0.08fF
C39 a_1038_210.n0 GND 0.02fF
C40 a_1038_210.n1 GND 0.09fF
C41 a_1038_210.n2 GND 0.12fF
C42 a_1038_210.n3 GND 0.08fF
C43 a_1038_210.n4 GND 0.08fF
C44 a_1038_210.n5 GND 0.02fF
C45 a_1038_210.t1 GND 0.29fF
C46 a_1038_210.n6 GND 0.09fF
C47 a_1038_210.n7 GND 0.02fF
C48 a_1038_210.n8 GND 0.13fF
C49 a_1038_210.n9 GND 0.02fF
C50 a_1038_210.n10 GND 0.03fF
C51 a_1038_210.n11 GND 0.03fF
C52 a_2000_210.n0 GND 0.07fF
C53 a_2000_210.n1 GND 0.09fF
C54 a_2000_210.n2 GND 0.12fF
C55 a_2000_210.n3 GND 0.08fF
C56 a_2000_210.n4 GND 0.02fF
C57 a_2000_210.n5 GND 0.03fF
C58 a_2000_210.n6 GND 0.02fF
C59 a_2000_210.n7 GND 0.03fF
C60 a_2000_210.n8 GND 0.02fF
C61 a_2000_210.n9 GND 0.13fF
C62 a_2000_210.n10 GND 0.08fF
C63 a_2000_210.n11 GND 0.02fF
C64 a_2000_210.t0 GND 0.31fF
C65 a_3473_1050.n0 GND 0.32fF
C66 a_3473_1050.n1 GND 0.60fF
C67 a_3473_1050.n2 GND 0.04fF
C68 a_3473_1050.n3 GND 0.05fF
C69 a_3473_1050.n4 GND 0.03fF
C70 a_3473_1050.n5 GND 0.18fF
C71 a_3473_1050.n6 GND 0.62fF
C72 a_3473_1050.n7 GND 0.45fF
C73 a_3473_1050.n8 GND 0.56fF
C74 a_3473_1050.n9 GND 0.35fF
C75 a_343_411.n0 GND 0.54fF
C76 a_343_411.n1 GND 0.39fF
C77 a_343_411.n2 GND 1.30fF
C78 a_343_411.n3 GND 0.38fF
C79 a_343_411.t11 GND 0.79fF
C80 a_343_411.n4 GND 0.84fF
C81 a_343_411.n5 GND 2.54fF
C82 a_343_411.n6 GND 0.06fF
C83 a_343_411.n7 GND 0.07fF
C84 a_343_411.n8 GND 0.05fF
C85 a_343_411.n9 GND 0.39fF
C86 a_343_411.n10 GND 0.72fF
C87 a_343_411.n11 GND 0.53fF
C88 a_343_411.n12 GND 0.68fF
C89 a_343_411.n13 GND 0.65fF
C90 a_343_411.n14 GND 0.54fF
C91 a_4294_210.n0 GND 0.06fF
C92 a_4294_210.n1 GND 0.09fF
C93 a_4294_210.n2 GND 0.11fF
C94 a_4294_210.n3 GND 0.08fF
C95 a_4294_210.n4 GND 0.02fF
C96 a_4294_210.n5 GND 0.03fF
C97 a_4294_210.n6 GND 0.04fF
C98 a_4294_210.n7 GND 0.02fF
C99 a_4294_210.n8 GND 0.13fF
C100 a_4294_210.n9 GND 0.08fF
C101 a_4294_210.n10 GND 0.02fF
C102 a_4013_103.n0 GND 0.08fF
C103 a_4013_103.n1 GND 0.07fF
C104 a_4013_103.n2 GND 0.04fF
C105 a_4013_103.n3 GND 0.06fF
C106 a_4013_103.n4 GND 0.11fF
C107 a_4013_103.n5 GND 0.04fF
C108 a_4013_103.n7 GND 0.08fF
C109 SN.n0 GND 0.41fF
C110 SN.t0 GND 0.44fF
C111 SN.n1 GND 0.97fF
C112 SN.n2 GND 0.41fF
C113 SN.t3 GND 0.44fF
C114 SN.n3 GND 0.38fF
C115 SN.n4 GND 1.24fF
C116 a_2702_101.n0 GND 0.02fF
C117 a_2702_101.n1 GND 0.09fF
C118 a_2702_101.n2 GND 0.07fF
C119 a_2702_101.n3 GND 0.04fF
C120 a_2702_101.n4 GND 0.01fF
C121 a_2702_101.n5 GND 0.04fF
C122 a_2702_101.n6 GND 0.04fF
C123 a_2702_101.n7 GND 0.02fF
C124 a_2702_101.n8 GND 0.05fF
C125 a_2702_101.n9 GND 0.02fF
C126 a_2702_101.n10 GND 0.15fF
C127 a_2702_101.n11 GND 0.08fF
C128 a_2702_101.n12 GND 0.08fF
C129 a_2702_101.t1 GND 0.23fF
C130 a_2702_101.n13 GND 0.01fF
C131 Q.n0 GND 0.39fF
C132 Q.n1 GND 0.39fF
C133 Q.n2 GND 0.50fF
C134 Q.n3 GND 0.47fF
C135 Q.n4 GND 0.45fF
C136 Q.n5 GND 0.04fF
C137 Q.n6 GND 0.05fF
C138 Q.n7 GND 0.03fF
C139 Q.n8 GND 0.22fF
C140 Q.n9 GND 0.52fF
C141 Q.n10 GND 0.31fF
C142 Q.t9 GND 0.53fF
C143 Q.n11 GND 0.61fF
C144 Q.n12 GND 0.03fF
C145 a_1905_1050.n0 GND 0.33fF
C146 a_1905_1050.n1 GND 0.51fF
C147 a_1905_1050.n2 GND 0.03fF
C148 a_1905_1050.n3 GND 0.05fF
C149 a_1905_1050.n4 GND 0.03fF
C150 a_1905_1050.n5 GND 0.14fF
C151 a_1905_1050.n6 GND 0.60fF
C152 a_1905_1050.n7 GND 0.34fF
C153 a_1905_1050.n8 GND 0.43fF
C154 a_1905_1050.n9 GND 0.40fF
C155 a_1905_1050.n10 GND 0.44fF
C156 a_1905_1050.n11 GND 0.34fF
C157 a_1265_989.n0 GND 0.07fF
C158 a_1265_989.n1 GND 0.45fF
C159 a_1265_989.n2 GND 0.58fF
C160 a_1265_989.n3 GND 0.65fF
C161 a_1265_989.n4 GND 0.36fF
C162 a_1265_989.n5 GND 0.89fF
C163 a_1265_989.n6 GND 0.36fF
C164 a_1265_989.t7 GND 0.65fF
C165 a_1265_989.n7 GND 0.49fF
C166 a_1265_989.n8 GND 0.36fF
C167 a_1265_989.t8 GND 0.65fF
C168 a_1265_989.n9 GND 0.70fF
C169 a_1265_989.n10 GND 1.15fF
C170 a_1265_989.n11 GND 1.46fF
C171 a_1265_989.n12 GND 0.59fF
C172 a_1265_989.n13 GND 0.03fF
C173 a_1265_989.n14 GND 0.30fF
C174 a_1265_989.n15 GND 0.05fF
C175 VDD.n1 GND 0.03fF
C176 VDD.n2 GND 0.17fF
C177 VDD.n3 GND 0.03fF
C178 VDD.n4 GND 0.02fF
C179 VDD.n5 GND 0.06fF
C180 VDD.n6 GND 0.02fF
C181 VDD.n7 GND 0.02fF
C182 VDD.n8 GND 0.02fF
C183 VDD.n9 GND 0.02fF
C184 VDD.n10 GND 0.02fF
C185 VDD.n11 GND 0.02fF
C186 VDD.n12 GND 0.02fF
C187 VDD.n13 GND 0.02fF
C188 VDD.n14 GND 0.03fF
C189 VDD.n15 GND 0.01fF
C190 VDD.n20 GND 0.43fF
C191 VDD.n21 GND 0.26fF
C192 VDD.n22 GND 0.02fF
C193 VDD.n23 GND 0.03fF
C194 VDD.n24 GND 0.26fF
C195 VDD.n25 GND 0.01fF
C196 VDD.n26 GND 0.02fF
C197 VDD.n27 GND 0.01fF
C198 VDD.n28 GND 0.21fF
C199 VDD.n29 GND 0.01fF
C200 VDD.n30 GND 0.07fF
C201 VDD.n31 GND 0.08fF
C202 VDD.n32 GND 0.16fF
C203 VDD.n33 GND 0.01fF
C204 VDD.n34 GND 0.02fF
C205 VDD.n35 GND 0.02fF
C206 VDD.n36 GND 0.15fF
C207 VDD.n37 GND 0.01fF
C208 VDD.n38 GND 0.08fF
C209 VDD.n39 GND 0.05fF
C210 VDD.n40 GND 0.02fF
C211 VDD.n41 GND 0.02fF
C212 VDD.n42 GND 0.14fF
C213 VDD.n43 GND 0.01fF
C214 VDD.n44 GND 0.02fF
C215 VDD.n45 GND 0.03fF
C216 VDD.n46 GND 0.14fF
C217 VDD.n47 GND 0.01fF
C218 VDD.n48 GND 0.02fF
C219 VDD.n49 GND 0.03fF
C220 VDD.n50 GND 0.08fF
C221 VDD.n51 GND 0.05fF
C222 VDD.n52 GND 0.15fF
C223 VDD.n53 GND 0.01fF
C224 VDD.n54 GND 0.02fF
C225 VDD.n55 GND 0.02fF
C226 VDD.n56 GND 0.16fF
C227 VDD.n57 GND 0.01fF
C228 VDD.n58 GND 0.02fF
C229 VDD.n59 GND 0.02fF
C230 VDD.n60 GND 0.06fF
C231 VDD.n61 GND 0.21fF
C232 VDD.n62 GND 0.01fF
C233 VDD.n63 GND 0.01fF
C234 VDD.n64 GND 0.02fF
C235 VDD.n65 GND 0.26fF
C236 VDD.n66 GND 0.01fF
C237 VDD.n67 GND 0.02fF
C238 VDD.n68 GND 0.02fF
C239 VDD.n69 GND 0.26fF
C240 VDD.n70 GND 0.01fF
C241 VDD.n71 GND 0.02fF
C242 VDD.n72 GND 0.03fF
C243 VDD.n73 GND 0.05fF
C244 VDD.n74 GND 0.02fF
C245 VDD.n75 GND 0.02fF
C246 VDD.n76 GND 0.02fF
C247 VDD.n77 GND 0.02fF
C248 VDD.n78 GND 0.02fF
C249 VDD.n79 GND 0.02fF
C250 VDD.n80 GND 0.02fF
C251 VDD.n81 GND 0.02fF
C252 VDD.n82 GND 0.02fF
C253 VDD.n83 GND 0.02fF
C254 VDD.n84 GND 0.02fF
C255 VDD.n85 GND 0.03fF
C256 VDD.n86 GND 0.02fF
C257 VDD.n87 GND 0.25fF
C258 VDD.n88 GND 0.02fF
C259 VDD.n89 GND 0.02fF
C260 VDD.n91 GND 0.02fF
C261 VDD.n95 GND 0.26fF
C262 VDD.n96 GND 0.26fF
C263 VDD.n97 GND 0.01fF
C264 VDD.n98 GND 0.02fF
C265 VDD.n99 GND 0.03fF
C266 VDD.n100 GND 0.06fF
C267 VDD.n101 GND 0.23fF
C268 VDD.n102 GND 0.01fF
C269 VDD.n103 GND 0.01fF
C270 VDD.n104 GND 0.02fF
C271 VDD.n105 GND 0.16fF
C272 VDD.n106 GND 0.01fF
C273 VDD.n107 GND 0.02fF
C274 VDD.n108 GND 0.02fF
C275 VDD.n109 GND 0.08fF
C276 VDD.n110 GND 0.05fF
C277 VDD.n111 GND 0.01fF
C278 VDD.n112 GND 0.02fF
C279 VDD.n113 GND 0.02fF
C280 VDD.n114 GND 0.13fF
C281 VDD.n115 GND 0.01fF
C282 VDD.n116 GND 0.02fF
C283 VDD.n117 GND 0.02fF
C284 VDD.n118 GND 0.16fF
C285 VDD.n119 GND 0.01fF
C286 VDD.n120 GND 0.02fF
C287 VDD.n121 GND 0.02fF
C288 VDD.n122 GND 0.06fF
C289 VDD.n123 GND 0.24fF
C290 VDD.n124 GND 0.01fF
C291 VDD.n125 GND 0.01fF
C292 VDD.n126 GND 0.02fF
C293 VDD.n127 GND 0.26fF
C294 VDD.n128 GND 0.01fF
C295 VDD.n129 GND 0.02fF
C296 VDD.n130 GND 0.03fF
C297 VDD.n131 GND 0.20fF
C298 VDD.n132 GND 0.02fF
C299 VDD.n133 GND 0.02fF
C300 VDD.n134 GND 0.02fF
C301 VDD.n135 GND 0.06fF
C302 VDD.n136 GND 0.02fF
C303 VDD.n137 GND 0.02fF
C304 VDD.n138 GND 0.02fF
C305 VDD.n139 GND 0.02fF
C306 VDD.n140 GND 0.02fF
C307 VDD.n141 GND 0.02fF
C308 VDD.n142 GND 0.02fF
C309 VDD.n143 GND 0.02fF
C310 VDD.n144 GND 0.02fF
C311 VDD.n145 GND 0.02fF
C312 VDD.n146 GND 0.03fF
C313 VDD.n147 GND 0.02fF
C314 VDD.n148 GND 0.02fF
C315 VDD.n152 GND 0.26fF
C316 VDD.n153 GND 0.26fF
C317 VDD.n154 GND 0.01fF
C318 VDD.n155 GND 0.02fF
C319 VDD.n156 GND 0.03fF
C320 VDD.n157 GND 0.06fF
C321 VDD.n158 GND 0.23fF
C322 VDD.n159 GND 0.01fF
C323 VDD.n160 GND 0.01fF
C324 VDD.n161 GND 0.02fF
C325 VDD.n162 GND 0.16fF
C326 VDD.n163 GND 0.01fF
C327 VDD.n164 GND 0.02fF
C328 VDD.n165 GND 0.02fF
C329 VDD.n166 GND 0.08fF
C330 VDD.n167 GND 0.05fF
C331 VDD.n168 GND 0.01fF
C332 VDD.n169 GND 0.02fF
C333 VDD.n170 GND 0.02fF
C334 VDD.n171 GND 0.13fF
C335 VDD.n172 GND 0.01fF
C336 VDD.n173 GND 0.02fF
C337 VDD.n174 GND 0.02fF
C338 VDD.n175 GND 0.16fF
C339 VDD.n176 GND 0.01fF
C340 VDD.n177 GND 0.02fF
C341 VDD.n178 GND 0.02fF
C342 VDD.n179 GND 0.06fF
C343 VDD.n180 GND 0.24fF
C344 VDD.n181 GND 0.01fF
C345 VDD.n182 GND 0.01fF
C346 VDD.n183 GND 0.02fF
C347 VDD.n184 GND 0.26fF
C348 VDD.n185 GND 0.01fF
C349 VDD.n186 GND 0.02fF
C350 VDD.n187 GND 0.03fF
C351 VDD.n188 GND 0.25fF
C352 VDD.n189 GND 0.02fF
C353 VDD.n190 GND 0.02fF
C354 VDD.n191 GND 0.02fF
C355 VDD.n192 GND 0.06fF
C356 VDD.n193 GND 0.02fF
C357 VDD.n194 GND 0.02fF
C358 VDD.n195 GND 0.02fF
C359 VDD.n196 GND 0.02fF
C360 VDD.n197 GND 0.02fF
C361 VDD.n198 GND 0.02fF
C362 VDD.n199 GND 0.02fF
C363 VDD.n200 GND 0.02fF
C364 VDD.n201 GND 0.02fF
C365 VDD.n202 GND 0.02fF
C366 VDD.n203 GND 0.03fF
C367 VDD.n204 GND 0.02fF
C368 VDD.n205 GND 0.02fF
C369 VDD.n209 GND 0.26fF
C370 VDD.n210 GND 0.26fF
C371 VDD.n211 GND 0.01fF
C372 VDD.n212 GND 0.02fF
C373 VDD.n213 GND 0.03fF
C374 VDD.n214 GND 0.26fF
C375 VDD.n215 GND 0.01fF
C376 VDD.n216 GND 0.02fF
C377 VDD.n217 GND 0.01fF
C378 VDD.n218 GND 0.13fF
C379 VDD.n219 GND 0.02fF
C380 VDD.n220 GND 0.02fF
C381 VDD.n221 GND 0.06fF
C382 VDD.n222 GND 0.02fF
C383 VDD.n223 GND 0.02fF
C384 VDD.n224 GND 0.02fF
C385 VDD.n225 GND 0.02fF
C386 VDD.n226 GND 0.02fF
C387 VDD.n227 GND 0.02fF
C388 VDD.n228 GND 0.02fF
C389 VDD.n229 GND 0.02fF
C390 VDD.n230 GND 0.03fF
C391 VDD.n231 GND 0.03fF
C392 VDD.n232 GND 0.02fF
C393 VDD.n236 GND 0.43fF
C394 VDD.n237 GND 0.26fF
C395 VDD.n238 GND 0.02fF
C396 VDD.n239 GND 0.03fF
C397 VDD.n240 GND 0.03fF
C398 VDD.n241 GND 0.06fF
C399 VDD.n242 GND 0.24fF
C400 VDD.n243 GND 0.01fF
C401 VDD.n244 GND 0.01fF
C402 VDD.n245 GND 0.02fF
C403 VDD.n246 GND 0.16fF
C404 VDD.n247 GND 0.01fF
C405 VDD.n248 GND 0.02fF
C406 VDD.n249 GND 0.02fF
C407 VDD.n250 GND 0.13fF
C408 VDD.n251 GND 0.01fF
C409 VDD.n252 GND 0.02fF
C410 VDD.n253 GND 0.02fF
C411 VDD.n254 GND 0.08fF
C412 VDD.n255 GND 0.05fF
C413 VDD.n256 GND 0.01fF
C414 VDD.n257 GND 0.02fF
C415 VDD.n258 GND 0.02fF
C416 VDD.n259 GND 0.16fF
C417 VDD.n260 GND 0.01fF
C418 VDD.n261 GND 0.02fF
C419 VDD.n262 GND 0.02fF
C420 VDD.n263 GND 0.06fF
C421 VDD.n264 GND 0.23fF
C422 VDD.n265 GND 0.01fF
C423 VDD.n266 GND 0.01fF
C424 VDD.n267 GND 0.02fF
C425 VDD.n268 GND 0.26fF
C426 VDD.n269 GND 0.01fF
C427 VDD.n270 GND 0.02fF
C428 VDD.n271 GND 0.03fF
C429 VDD.n272 GND 0.05fF
C430 VDD.n273 GND 0.02fF
C431 VDD.n274 GND 0.02fF
C432 VDD.n275 GND 0.02fF
C433 VDD.n276 GND 0.02fF
C434 VDD.n277 GND 0.02fF
C435 VDD.n278 GND 0.02fF
C436 VDD.n279 GND 0.02fF
C437 VDD.n280 GND 0.02fF
C438 VDD.n281 GND 0.02fF
C439 VDD.n282 GND 0.02fF
C440 VDD.n283 GND 0.02fF
C441 VDD.n284 GND 0.03fF
C442 VDD.n285 GND 0.02fF
C443 VDD.n288 GND 0.02fF
C444 VDD.n290 GND 0.02fF
C445 VDD.n291 GND 0.25fF
C446 VDD.n292 GND 0.02fF
C447 VDD.n294 GND 0.26fF
C448 VDD.n295 GND 0.26fF
C449 VDD.n296 GND 0.01fF
C450 VDD.n297 GND 0.02fF
C451 VDD.n298 GND 0.03fF
C452 VDD.n299 GND 0.26fF
C453 VDD.n300 GND 0.01fF
C454 VDD.n301 GND 0.02fF
C455 VDD.n302 GND 0.02fF
C456 VDD.n303 GND 0.06fF
C457 VDD.n304 GND 0.21fF
C458 VDD.n305 GND 0.01fF
C459 VDD.n306 GND 0.01fF
C460 VDD.n307 GND 0.02fF
C461 VDD.n308 GND 0.16fF
C462 VDD.n309 GND 0.01fF
C463 VDD.n310 GND 0.02fF
C464 VDD.n311 GND 0.02fF
C465 VDD.n312 GND 0.08fF
C466 VDD.n313 GND 0.05fF
C467 VD