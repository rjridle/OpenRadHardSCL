magic
tech sky130A
magscale 1 2
timestamp 1649530829
<< nwell >>
rect -84 832 19398 1575
<< nmos >>
rect 147 318 177 379
tri 177 318 193 334 sw
rect 447 318 477 379
rect 147 288 253 318
tri 253 288 283 318 sw
rect 147 187 177 288
tri 177 272 193 288 nw
tri 237 272 253 288 ne
tri 177 187 193 203 sw
tri 237 187 253 203 se
rect 253 187 283 288
tri 342 288 372 318 se
rect 372 288 477 318
rect 342 194 372 288
tri 372 272 388 288 nw
tri 431 272 447 288 ne
tri 372 194 388 210 sw
tri 431 194 447 210 se
rect 447 194 477 288
tri 147 157 177 187 ne
rect 177 157 253 187
tri 253 157 283 187 nw
tri 342 164 372 194 ne
rect 372 164 447 194
tri 447 164 477 194 nw
rect 649 326 679 379
tri 679 326 695 342 sw
rect 649 296 755 326
tri 755 296 785 326 sw
rect 649 195 679 296
tri 679 280 695 296 nw
tri 739 280 755 296 ne
tri 679 195 695 211 sw
tri 739 195 755 211 se
rect 755 195 785 296
tri 649 165 679 195 ne
rect 679 165 755 195
tri 755 165 785 195 nw
rect 1109 318 1139 379
tri 1139 318 1155 334 sw
rect 1409 318 1439 379
rect 1109 288 1215 318
tri 1215 288 1245 318 sw
rect 1109 187 1139 288
tri 1139 272 1155 288 nw
tri 1199 272 1215 288 ne
tri 1139 187 1155 203 sw
tri 1199 187 1215 203 se
rect 1215 187 1245 288
tri 1304 288 1334 318 se
rect 1334 288 1439 318
rect 1304 194 1334 288
tri 1334 272 1350 288 nw
tri 1393 272 1409 288 ne
tri 1334 194 1350 210 sw
tri 1393 194 1409 210 se
rect 1409 194 1439 288
tri 1109 157 1139 187 ne
rect 1139 157 1215 187
tri 1215 157 1245 187 nw
tri 1304 164 1334 194 ne
rect 1334 164 1409 194
tri 1409 164 1439 194 nw
rect 1611 326 1641 379
tri 1641 326 1657 342 sw
rect 1611 296 1717 326
tri 1717 296 1747 326 sw
rect 1611 195 1641 296
tri 1641 280 1657 296 nw
tri 1701 280 1717 296 ne
tri 1641 195 1657 211 sw
tri 1701 195 1717 211 se
rect 1717 195 1747 296
tri 1611 165 1641 195 ne
rect 1641 165 1717 195
tri 1717 165 1747 195 nw
rect 2071 318 2101 379
tri 2101 318 2117 334 sw
rect 2371 318 2401 379
rect 2071 288 2177 318
tri 2177 288 2207 318 sw
rect 2071 187 2101 288
tri 2101 272 2117 288 nw
tri 2161 272 2177 288 ne
tri 2101 187 2117 203 sw
tri 2161 187 2177 203 se
rect 2177 187 2207 288
tri 2266 288 2296 318 se
rect 2296 288 2401 318
rect 2266 194 2296 288
tri 2296 272 2312 288 nw
tri 2355 272 2371 288 ne
tri 2296 194 2312 210 sw
tri 2355 194 2371 210 se
rect 2371 194 2401 288
tri 2071 157 2101 187 ne
rect 2101 157 2177 187
tri 2177 157 2207 187 nw
tri 2266 164 2296 194 ne
rect 2296 164 2371 194
tri 2371 164 2401 194 nw
rect 2573 326 2603 379
tri 2603 326 2619 342 sw
rect 2573 296 2679 326
tri 2679 296 2709 326 sw
rect 2573 195 2603 296
tri 2603 280 2619 296 nw
tri 2663 280 2679 296 ne
tri 2603 195 2619 211 sw
tri 2663 195 2679 211 se
rect 2679 195 2709 296
tri 2573 165 2603 195 ne
rect 2603 165 2679 195
tri 2679 165 2709 195 nw
rect 3033 318 3063 379
tri 3063 318 3079 334 sw
rect 3333 318 3363 379
rect 3033 288 3139 318
tri 3139 288 3169 318 sw
rect 3033 187 3063 288
tri 3063 272 3079 288 nw
tri 3123 272 3139 288 ne
tri 3063 187 3079 203 sw
tri 3123 187 3139 203 se
rect 3139 187 3169 288
tri 3228 288 3258 318 se
rect 3258 288 3363 318
rect 3228 194 3258 288
tri 3258 272 3274 288 nw
tri 3317 272 3333 288 ne
tri 3258 194 3274 210 sw
tri 3317 194 3333 210 se
rect 3333 194 3363 288
tri 3033 157 3063 187 ne
rect 3063 157 3139 187
tri 3139 157 3169 187 nw
tri 3228 164 3258 194 ne
rect 3258 164 3333 194
tri 3333 164 3363 194 nw
rect 3535 326 3565 379
tri 3565 326 3581 342 sw
rect 3535 296 3641 326
tri 3641 296 3671 326 sw
rect 3535 195 3565 296
tri 3565 280 3581 296 nw
tri 3625 280 3641 296 ne
tri 3565 195 3581 211 sw
tri 3625 195 3641 211 se
rect 3641 195 3671 296
tri 3535 165 3565 195 ne
rect 3565 165 3641 195
tri 3641 165 3671 195 nw
rect 3995 318 4025 379
tri 4025 318 4041 334 sw
rect 4295 318 4325 379
rect 3995 288 4101 318
tri 4101 288 4131 318 sw
rect 3995 187 4025 288
tri 4025 272 4041 288 nw
tri 4085 272 4101 288 ne
tri 4025 187 4041 203 sw
tri 4085 187 4101 203 se
rect 4101 187 4131 288
tri 4190 288 4220 318 se
rect 4220 288 4325 318
rect 4190 194 4220 288
tri 4220 272 4236 288 nw
tri 4279 272 4295 288 ne
tri 4220 194 4236 210 sw
tri 4279 194 4295 210 se
rect 4295 194 4325 288
tri 3995 157 4025 187 ne
rect 4025 157 4101 187
tri 4101 157 4131 187 nw
tri 4190 164 4220 194 ne
rect 4220 164 4295 194
tri 4295 164 4325 194 nw
rect 4497 326 4527 379
tri 4527 326 4543 342 sw
rect 4497 296 4603 326
tri 4603 296 4633 326 sw
rect 4497 195 4527 296
tri 4527 280 4543 296 nw
tri 4587 280 4603 296 ne
tri 4527 195 4543 211 sw
tri 4587 195 4603 211 se
rect 4603 195 4633 296
tri 4497 165 4527 195 ne
rect 4527 165 4603 195
tri 4603 165 4633 195 nw
rect 4957 318 4987 379
tri 4987 318 5003 334 sw
rect 5257 318 5287 379
rect 4957 288 5063 318
tri 5063 288 5093 318 sw
rect 4957 187 4987 288
tri 4987 272 5003 288 nw
tri 5047 272 5063 288 ne
tri 4987 187 5003 203 sw
tri 5047 187 5063 203 se
rect 5063 187 5093 288
tri 5152 288 5182 318 se
rect 5182 288 5287 318
rect 5152 194 5182 288
tri 5182 272 5198 288 nw
tri 5241 272 5257 288 ne
tri 5182 194 5198 210 sw
tri 5241 194 5257 210 se
rect 5257 194 5287 288
tri 4957 157 4987 187 ne
rect 4987 157 5063 187
tri 5063 157 5093 187 nw
tri 5152 164 5182 194 ne
rect 5182 164 5257 194
tri 5257 164 5287 194 nw
rect 5459 326 5489 379
tri 5489 326 5505 342 sw
rect 5459 296 5565 326
tri 5565 296 5595 326 sw
rect 5459 195 5489 296
tri 5489 280 5505 296 nw
tri 5549 280 5565 296 ne
tri 5489 195 5505 211 sw
tri 5549 195 5565 211 se
rect 5565 195 5595 296
tri 5459 165 5489 195 ne
rect 5489 165 5565 195
tri 5565 165 5595 195 nw
rect 5919 318 5949 379
tri 5949 318 5965 334 sw
rect 6219 318 6249 379
rect 5919 288 6025 318
tri 6025 288 6055 318 sw
rect 5919 187 5949 288
tri 5949 272 5965 288 nw
tri 6009 272 6025 288 ne
tri 5949 187 5965 203 sw
tri 6009 187 6025 203 se
rect 6025 187 6055 288
tri 6114 288 6144 318 se
rect 6144 288 6249 318
rect 6114 194 6144 288
tri 6144 272 6160 288 nw
tri 6203 272 6219 288 ne
tri 6144 194 6160 210 sw
tri 6203 194 6219 210 se
rect 6219 194 6249 288
tri 5919 157 5949 187 ne
rect 5949 157 6025 187
tri 6025 157 6055 187 nw
tri 6114 164 6144 194 ne
rect 6144 164 6219 194
tri 6219 164 6249 194 nw
rect 6421 326 6451 379
tri 6451 326 6467 342 sw
rect 6421 296 6527 326
tri 6527 296 6557 326 sw
rect 6421 195 6451 296
tri 6451 280 6467 296 nw
tri 6511 280 6527 296 ne
tri 6451 195 6467 211 sw
tri 6511 195 6527 211 se
rect 6527 195 6557 296
tri 6421 165 6451 195 ne
rect 6451 165 6527 195
tri 6527 165 6557 195 nw
rect 6881 318 6911 379
tri 6911 318 6927 334 sw
rect 7181 318 7211 379
rect 6881 288 6987 318
tri 6987 288 7017 318 sw
rect 6881 187 6911 288
tri 6911 272 6927 288 nw
tri 6971 272 6987 288 ne
tri 6911 187 6927 203 sw
tri 6971 187 6987 203 se
rect 6987 187 7017 288
tri 7076 288 7106 318 se
rect 7106 288 7211 318
rect 7076 194 7106 288
tri 7106 272 7122 288 nw
tri 7165 272 7181 288 ne
tri 7106 194 7122 210 sw
tri 7165 194 7181 210 se
rect 7181 194 7211 288
tri 6881 157 6911 187 ne
rect 6911 157 6987 187
tri 6987 157 7017 187 nw
tri 7076 164 7106 194 ne
rect 7106 164 7181 194
tri 7181 164 7211 194 nw
rect 7383 326 7413 379
tri 7413 326 7429 342 sw
rect 7383 296 7489 326
tri 7489 296 7519 326 sw
rect 7383 195 7413 296
tri 7413 280 7429 296 nw
tri 7473 280 7489 296 ne
tri 7413 195 7429 211 sw
tri 7473 195 7489 211 se
rect 7489 195 7519 296
tri 7383 165 7413 195 ne
rect 7413 165 7489 195
tri 7489 165 7519 195 nw
rect 7843 318 7873 379
tri 7873 318 7889 334 sw
rect 8143 318 8173 379
rect 7843 288 7949 318
tri 7949 288 7979 318 sw
rect 7843 187 7873 288
tri 7873 272 7889 288 nw
tri 7933 272 7949 288 ne
tri 7873 187 7889 203 sw
tri 7933 187 7949 203 se
rect 7949 187 7979 288
tri 8038 288 8068 318 se
rect 8068 288 8173 318
rect 8038 194 8068 288
tri 8068 272 8084 288 nw
tri 8127 272 8143 288 ne
tri 8068 194 8084 210 sw
tri 8127 194 8143 210 se
rect 8143 194 8173 288
tri 7843 157 7873 187 ne
rect 7873 157 7949 187
tri 7949 157 7979 187 nw
tri 8038 164 8068 194 ne
rect 8068 164 8143 194
tri 8143 164 8173 194 nw
rect 8345 326 8375 379
tri 8375 326 8391 342 sw
rect 8345 296 8451 326
tri 8451 296 8481 326 sw
rect 8345 195 8375 296
tri 8375 280 8391 296 nw
tri 8435 280 8451 296 ne
tri 8375 195 8391 211 sw
tri 8435 195 8451 211 se
rect 8451 195 8481 296
tri 8345 165 8375 195 ne
rect 8375 165 8451 195
tri 8451 165 8481 195 nw
rect 8805 318 8835 379
tri 8835 318 8851 334 sw
rect 9105 318 9135 379
rect 8805 288 8911 318
tri 8911 288 8941 318 sw
rect 8805 187 8835 288
tri 8835 272 8851 288 nw
tri 8895 272 8911 288 ne
tri 8835 187 8851 203 sw
tri 8895 187 8911 203 se
rect 8911 187 8941 288
tri 9000 288 9030 318 se
rect 9030 288 9135 318
rect 9000 194 9030 288
tri 9030 272 9046 288 nw
tri 9089 272 9105 288 ne
tri 9030 194 9046 210 sw
tri 9089 194 9105 210 se
rect 9105 194 9135 288
tri 8805 157 8835 187 ne
rect 8835 157 8911 187
tri 8911 157 8941 187 nw
tri 9000 164 9030 194 ne
rect 9030 164 9105 194
tri 9105 164 9135 194 nw
rect 9307 326 9337 379
tri 9337 326 9353 342 sw
rect 9307 296 9413 326
tri 9413 296 9443 326 sw
rect 9307 195 9337 296
tri 9337 280 9353 296 nw
tri 9397 280 9413 296 ne
tri 9337 195 9353 211 sw
tri 9397 195 9413 211 se
rect 9413 195 9443 296
tri 9307 165 9337 195 ne
rect 9337 165 9413 195
tri 9413 165 9443 195 nw
rect 9767 318 9797 379
tri 9797 318 9813 334 sw
rect 10067 318 10097 379
rect 9767 288 9873 318
tri 9873 288 9903 318 sw
rect 9767 187 9797 288
tri 9797 272 9813 288 nw
tri 9857 272 9873 288 ne
tri 9797 187 9813 203 sw
tri 9857 187 9873 203 se
rect 9873 187 9903 288
tri 9962 288 9992 318 se
rect 9992 288 10097 318
rect 9962 194 9992 288
tri 9992 272 10008 288 nw
tri 10051 272 10067 288 ne
tri 9992 194 10008 210 sw
tri 10051 194 10067 210 se
rect 10067 194 10097 288
tri 9767 157 9797 187 ne
rect 9797 157 9873 187
tri 9873 157 9903 187 nw
tri 9962 164 9992 194 ne
rect 9992 164 10067 194
tri 10067 164 10097 194 nw
rect 10269 326 10299 379
tri 10299 326 10315 342 sw
rect 10269 296 10375 326
tri 10375 296 10405 326 sw
rect 10269 195 10299 296
tri 10299 280 10315 296 nw
tri 10359 280 10375 296 ne
tri 10299 195 10315 211 sw
tri 10359 195 10375 211 se
rect 10375 195 10405 296
tri 10269 165 10299 195 ne
rect 10299 165 10375 195
tri 10375 165 10405 195 nw
rect 10729 318 10759 379
tri 10759 318 10775 334 sw
rect 11029 318 11059 379
rect 10729 288 10835 318
tri 10835 288 10865 318 sw
rect 10729 187 10759 288
tri 10759 272 10775 288 nw
tri 10819 272 10835 288 ne
tri 10759 187 10775 203 sw
tri 10819 187 10835 203 se
rect 10835 187 10865 288
tri 10924 288 10954 318 se
rect 10954 288 11059 318
rect 10924 194 10954 288
tri 10954 272 10970 288 nw
tri 11013 272 11029 288 ne
tri 10954 194 10970 210 sw
tri 11013 194 11029 210 se
rect 11029 194 11059 288
tri 10729 157 10759 187 ne
rect 10759 157 10835 187
tri 10835 157 10865 187 nw
tri 10924 164 10954 194 ne
rect 10954 164 11029 194
tri 11029 164 11059 194 nw
rect 11231 326 11261 379
tri 11261 326 11277 342 sw
rect 11231 296 11337 326
tri 11337 296 11367 326 sw
rect 11231 195 11261 296
tri 11261 280 11277 296 nw
tri 11321 280 11337 296 ne
tri 11261 195 11277 211 sw
tri 11321 195 11337 211 se
rect 11337 195 11367 296
tri 11231 165 11261 195 ne
rect 11261 165 11337 195
tri 11337 165 11367 195 nw
rect 11691 318 11721 379
tri 11721 318 11737 334 sw
rect 11991 318 12021 379
rect 11691 288 11797 318
tri 11797 288 11827 318 sw
rect 11691 187 11721 288
tri 11721 272 11737 288 nw
tri 11781 272 11797 288 ne
tri 11721 187 11737 203 sw
tri 11781 187 11797 203 se
rect 11797 187 11827 288
tri 11886 288 11916 318 se
rect 11916 288 12021 318
rect 11886 194 11916 288
tri 11916 272 11932 288 nw
tri 11975 272 11991 288 ne
tri 11916 194 11932 210 sw
tri 11975 194 11991 210 se
rect 11991 194 12021 288
tri 11691 157 11721 187 ne
rect 11721 157 11797 187
tri 11797 157 11827 187 nw
tri 11886 164 11916 194 ne
rect 11916 164 11991 194
tri 11991 164 12021 194 nw
rect 12193 326 12223 379
tri 12223 326 12239 342 sw
rect 12193 296 12299 326
tri 12299 296 12329 326 sw
rect 12193 195 12223 296
tri 12223 280 12239 296 nw
tri 12283 280 12299 296 ne
tri 12223 195 12239 211 sw
tri 12283 195 12299 211 se
rect 12299 195 12329 296
tri 12193 165 12223 195 ne
rect 12223 165 12299 195
tri 12299 165 12329 195 nw
rect 12653 318 12683 379
tri 12683 318 12699 334 sw
rect 12953 318 12983 379
rect 12653 288 12759 318
tri 12759 288 12789 318 sw
rect 12653 187 12683 288
tri 12683 272 12699 288 nw
tri 12743 272 12759 288 ne
tri 12683 187 12699 203 sw
tri 12743 187 12759 203 se
rect 12759 187 12789 288
tri 12848 288 12878 318 se
rect 12878 288 12983 318
rect 12848 194 12878 288
tri 12878 272 12894 288 nw
tri 12937 272 12953 288 ne
tri 12878 194 12894 210 sw
tri 12937 194 12953 210 se
rect 12953 194 12983 288
tri 12653 157 12683 187 ne
rect 12683 157 12759 187
tri 12759 157 12789 187 nw
tri 12848 164 12878 194 ne
rect 12878 164 12953 194
tri 12953 164 12983 194 nw
rect 13155 326 13185 379
tri 13185 326 13201 342 sw
rect 13155 296 13261 326
tri 13261 296 13291 326 sw
rect 13155 195 13185 296
tri 13185 280 13201 296 nw
tri 13245 280 13261 296 ne
tri 13185 195 13201 211 sw
tri 13245 195 13261 211 se
rect 13261 195 13291 296
tri 13155 165 13185 195 ne
rect 13185 165 13261 195
tri 13261 165 13291 195 nw
rect 13615 318 13645 379
tri 13645 318 13661 334 sw
rect 13915 318 13945 379
rect 13615 288 13721 318
tri 13721 288 13751 318 sw
rect 13615 187 13645 288
tri 13645 272 13661 288 nw
tri 13705 272 13721 288 ne
tri 13645 187 13661 203 sw
tri 13705 187 13721 203 se
rect 13721 187 13751 288
tri 13810 288 13840 318 se
rect 13840 288 13945 318
rect 13810 194 13840 288
tri 13840 272 13856 288 nw
tri 13899 272 13915 288 ne
tri 13840 194 13856 210 sw
tri 13899 194 13915 210 se
rect 13915 194 13945 288
tri 13615 157 13645 187 ne
rect 13645 157 13721 187
tri 13721 157 13751 187 nw
tri 13810 164 13840 194 ne
rect 13840 164 13915 194
tri 13915 164 13945 194 nw
rect 14117 326 14147 379
tri 14147 326 14163 342 sw
rect 14117 296 14223 326
tri 14223 296 14253 326 sw
rect 14117 195 14147 296
tri 14147 280 14163 296 nw
tri 14207 280 14223 296 ne
tri 14147 195 14163 211 sw
tri 14207 195 14223 211 se
rect 14223 195 14253 296
tri 14117 165 14147 195 ne
rect 14147 165 14223 195
tri 14223 165 14253 195 nw
rect 14577 318 14607 379
tri 14607 318 14623 334 sw
rect 14877 318 14907 379
rect 14577 288 14683 318
tri 14683 288 14713 318 sw
rect 14577 187 14607 288
tri 14607 272 14623 288 nw
tri 14667 272 14683 288 ne
tri 14607 187 14623 203 sw
tri 14667 187 14683 203 se
rect 14683 187 14713 288
tri 14772 288 14802 318 se
rect 14802 288 14907 318
rect 14772 194 14802 288
tri 14802 272 14818 288 nw
tri 14861 272 14877 288 ne
tri 14802 194 14818 210 sw
tri 14861 194 14877 210 se
rect 14877 194 14907 288
tri 14577 157 14607 187 ne
rect 14607 157 14683 187
tri 14683 157 14713 187 nw
tri 14772 164 14802 194 ne
rect 14802 164 14877 194
tri 14877 164 14907 194 nw
rect 15079 326 15109 379
tri 15109 326 15125 342 sw
rect 15079 296 15185 326
tri 15185 296 15215 326 sw
rect 15079 195 15109 296
tri 15109 280 15125 296 nw
tri 15169 280 15185 296 ne
tri 15109 195 15125 211 sw
tri 15169 195 15185 211 se
rect 15185 195 15215 296
tri 15079 165 15109 195 ne
rect 15109 165 15185 195
tri 15185 165 15215 195 nw
rect 15539 318 15569 379
tri 15569 318 15585 334 sw
rect 15839 318 15869 379
rect 15539 288 15645 318
tri 15645 288 15675 318 sw
rect 15539 187 15569 288
tri 15569 272 15585 288 nw
tri 15629 272 15645 288 ne
tri 15569 187 15585 203 sw
tri 15629 187 15645 203 se
rect 15645 187 15675 288
tri 15734 288 15764 318 se
rect 15764 288 15869 318
rect 15734 194 15764 288
tri 15764 272 15780 288 nw
tri 15823 272 15839 288 ne
tri 15764 194 15780 210 sw
tri 15823 194 15839 210 se
rect 15839 194 15869 288
tri 15539 157 15569 187 ne
rect 15569 157 15645 187
tri 15645 157 15675 187 nw
tri 15734 164 15764 194 ne
rect 15764 164 15839 194
tri 15839 164 15869 194 nw
rect 16041 326 16071 379
tri 16071 326 16087 342 sw
rect 16041 296 16147 326
tri 16147 296 16177 326 sw
rect 16041 195 16071 296
tri 16071 280 16087 296 nw
tri 16131 280 16147 296 ne
tri 16071 195 16087 211 sw
tri 16131 195 16147 211 se
rect 16147 195 16177 296
tri 16041 165 16071 195 ne
rect 16071 165 16147 195
tri 16147 165 16177 195 nw
rect 16501 318 16531 379
tri 16531 318 16547 334 sw
rect 16801 318 16831 379
rect 16501 288 16607 318
tri 16607 288 16637 318 sw
rect 16501 187 16531 288
tri 16531 272 16547 288 nw
tri 16591 272 16607 288 ne
tri 16531 187 16547 203 sw
tri 16591 187 16607 203 se
rect 16607 187 16637 288
tri 16696 288 16726 318 se
rect 16726 288 16831 318
rect 16696 194 16726 288
tri 16726 272 16742 288 nw
tri 16785 272 16801 288 ne
tri 16726 194 16742 210 sw
tri 16785 194 16801 210 se
rect 16801 194 16831 288
tri 16501 157 16531 187 ne
rect 16531 157 16607 187
tri 16607 157 16637 187 nw
tri 16696 164 16726 194 ne
rect 16726 164 16801 194
tri 16801 164 16831 194 nw
rect 17003 326 17033 379
tri 17033 326 17049 342 sw
rect 17003 296 17109 326
tri 17109 296 17139 326 sw
rect 17003 195 17033 296
tri 17033 280 17049 296 nw
tri 17093 280 17109 296 ne
tri 17033 195 17049 211 sw
tri 17093 195 17109 211 se
rect 17109 195 17139 296
tri 17003 165 17033 195 ne
rect 17033 165 17109 195
tri 17109 165 17139 195 nw
rect 17484 316 17514 377
tri 17514 316 17530 332 sw
rect 17678 324 17708 377
tri 17708 324 17724 340 sw
rect 17484 286 17590 316
tri 17590 286 17620 316 sw
rect 17678 294 17784 324
tri 17784 294 17814 324 sw
rect 17484 185 17514 286
tri 17514 270 17530 286 nw
tri 17574 270 17590 286 ne
tri 17514 185 17530 201 sw
tri 17574 185 17590 201 se
rect 17590 185 17620 286
rect 17678 193 17708 294
tri 17708 278 17724 294 nw
tri 17768 278 17784 294 ne
tri 17708 193 17724 209 sw
tri 17768 193 17784 209 se
rect 17784 193 17814 294
tri 17484 155 17514 185 ne
rect 17514 155 17590 185
tri 17590 155 17620 185 nw
tri 17678 163 17708 193 ne
rect 17708 163 17784 193
tri 17784 163 17814 193 nw
rect 18150 316 18180 377
tri 18180 316 18196 332 sw
tri 18434 324 18450 340 se
rect 18450 324 18480 377
rect 18150 286 18256 316
tri 18256 286 18286 316 sw
tri 18344 294 18374 324 se
rect 18374 294 18480 324
rect 18150 185 18180 286
tri 18180 270 18196 286 nw
tri 18240 270 18256 286 ne
tri 18180 185 18196 201 sw
tri 18240 185 18256 201 se
rect 18256 185 18286 286
rect 18344 193 18374 294
tri 18374 278 18390 294 nw
tri 18434 278 18450 294 ne
tri 18374 193 18390 209 sw
tri 18434 193 18450 209 se
rect 18450 193 18480 294
tri 18150 155 18180 185 ne
rect 18180 155 18256 185
tri 18256 155 18286 185 nw
tri 18344 163 18374 193 ne
rect 18374 163 18450 193
tri 18450 163 18480 193 nw
rect 18816 316 18846 377
tri 18846 316 18862 332 sw
rect 19010 324 19040 377
tri 19040 324 19056 340 sw
rect 18816 286 18922 316
tri 18922 286 18952 316 sw
rect 19010 294 19116 324
tri 19116 294 19146 324 sw
rect 18816 185 18846 286
tri 18846 270 18862 286 nw
tri 18906 270 18922 286 ne
tri 18846 185 18862 201 sw
tri 18906 185 18922 201 se
rect 18922 185 18952 286
rect 19010 279 19041 294
tri 19041 279 19056 294 nw
tri 19100 279 19115 294 ne
rect 19115 279 19146 294
rect 19010 193 19040 279
tri 19040 193 19056 209 sw
tri 19100 193 19116 209 se
rect 19116 193 19146 279
tri 18816 155 18846 185 ne
rect 18846 155 18922 185
tri 18922 155 18952 185 nw
tri 19010 163 19040 193 ne
rect 19040 163 19116 193
tri 19116 163 19146 193 nw
<< pmos >>
rect 247 1050 277 1450
rect 335 1050 365 1450
rect 423 1050 453 1450
rect 511 1050 541 1450
rect 599 1050 629 1450
rect 687 1050 717 1450
rect 1209 1050 1239 1450
rect 1297 1050 1327 1450
rect 1385 1050 1415 1450
rect 1473 1050 1503 1450
rect 1561 1050 1591 1450
rect 1649 1050 1679 1450
rect 2171 1050 2201 1450
rect 2259 1050 2289 1450
rect 2347 1050 2377 1450
rect 2435 1050 2465 1450
rect 2523 1050 2553 1450
rect 2611 1050 2641 1450
rect 3133 1050 3163 1450
rect 3221 1050 3251 1450
rect 3309 1050 3339 1450
rect 3397 1050 3427 1450
rect 3485 1050 3515 1450
rect 3573 1050 3603 1450
rect 4095 1050 4125 1450
rect 4183 1050 4213 1450
rect 4271 1050 4301 1450
rect 4359 1050 4389 1450
rect 4447 1050 4477 1450
rect 4535 1050 4565 1450
rect 5057 1050 5087 1450
rect 5145 1050 5175 1450
rect 5233 1050 5263 1450
rect 5321 1050 5351 1450
rect 5409 1050 5439 1450
rect 5497 1050 5527 1450
rect 6019 1050 6049 1450
rect 6107 1050 6137 1450
rect 6195 1050 6225 1450
rect 6283 1050 6313 1450
rect 6371 1050 6401 1450
rect 6459 1050 6489 1450
rect 6981 1050 7011 1450
rect 7069 1050 7099 1450
rect 7157 1050 7187 1450
rect 7245 1050 7275 1450
rect 7333 1050 7363 1450
rect 7421 1050 7451 1450
rect 7943 1050 7973 1450
rect 8031 1050 8061 1450
rect 8119 1050 8149 1450
rect 8207 1050 8237 1450
rect 8295 1050 8325 1450
rect 8383 1050 8413 1450
rect 8905 1050 8935 1450
rect 8993 1050 9023 1450
rect 9081 1050 9111 1450
rect 9169 1050 9199 1450
rect 9257 1050 9287 1450
rect 9345 1050 9375 1450
rect 9867 1050 9897 1450
rect 9955 1050 9985 1450
rect 10043 1050 10073 1450
rect 10131 1050 10161 1450
rect 10219 1050 10249 1450
rect 10307 1050 10337 1450
rect 10829 1050 10859 1450
rect 10917 1050 10947 1450
rect 11005 1050 11035 1450
rect 11093 1050 11123 1450
rect 11181 1050 11211 1450
rect 11269 1050 11299 1450
rect 11791 1050 11821 1450
rect 11879 1050 11909 1450
rect 11967 1050 11997 1450
rect 12055 1050 12085 1450
rect 12143 1050 12173 1450
rect 12231 1050 12261 1450
rect 12753 1050 12783 1450
rect 12841 1050 12871 1450
rect 12929 1050 12959 1450
rect 13017 1050 13047 1450
rect 13105 1050 13135 1450
rect 13193 1050 13223 1450
rect 13715 1050 13745 1450
rect 13803 1050 13833 1450
rect 13891 1050 13921 1450
rect 13979 1050 14009 1450
rect 14067 1050 14097 1450
rect 14155 1050 14185 1450
rect 14677 1050 14707 1450
rect 14765 1050 14795 1450
rect 14853 1050 14883 1450
rect 14941 1050 14971 1450
rect 15029 1050 15059 1450
rect 15117 1050 15147 1450
rect 15639 1050 15669 1450
rect 15727 1050 15757 1450
rect 15815 1050 15845 1450
rect 15903 1050 15933 1450
rect 15991 1050 16021 1450
rect 16079 1050 16109 1450
rect 16601 1050 16631 1450
rect 16689 1050 16719 1450
rect 16777 1050 16807 1450
rect 16865 1050 16895 1450
rect 16953 1050 16983 1450
rect 17041 1050 17071 1450
rect 17503 1051 17533 1451
rect 17591 1051 17621 1451
rect 17679 1051 17709 1451
rect 17767 1051 17797 1451
rect 18167 1051 18197 1451
rect 18255 1051 18285 1451
rect 18343 1051 18373 1451
rect 18431 1051 18461 1451
rect 18835 1051 18865 1451
rect 18923 1051 18953 1451
rect 19011 1051 19041 1451
rect 19099 1051 19129 1451
<< ndiff >>
rect 91 363 147 379
rect 91 329 101 363
rect 135 329 147 363
rect 91 291 147 329
rect 177 363 447 379
rect 177 334 198 363
tri 177 318 193 334 ne
rect 193 329 198 334
rect 232 329 295 363
rect 329 329 392 363
rect 426 329 447 363
rect 193 318 447 329
rect 477 363 533 379
rect 477 329 489 363
rect 523 329 533 363
rect 91 257 101 291
rect 135 257 147 291
tri 253 288 283 318 ne
rect 283 291 342 318
rect 91 223 147 257
rect 91 189 101 223
rect 135 189 147 223
rect 91 157 147 189
tri 177 272 193 288 se
rect 193 272 237 288
tri 237 272 253 288 sw
rect 177 238 253 272
rect 177 204 198 238
rect 232 204 253 238
rect 177 203 253 204
tri 177 187 193 203 ne
rect 193 187 237 203
tri 237 187 253 203 nw
rect 283 257 295 291
rect 329 257 342 291
tri 342 288 372 318 nw
rect 283 223 342 257
rect 283 189 295 223
rect 329 189 342 223
tri 372 272 388 288 se
rect 388 272 431 288
tri 431 272 447 288 sw
rect 372 244 447 272
rect 372 210 393 244
rect 427 210 447 244
tri 372 194 388 210 ne
rect 388 194 431 210
tri 431 194 447 210 nw
tri 147 157 177 187 sw
tri 253 157 283 187 se
rect 283 164 342 189
tri 342 164 372 194 sw
tri 447 164 477 194 se
rect 477 164 533 329
rect 283 157 533 164
rect 91 153 533 157
rect 91 119 101 153
rect 135 119 295 153
rect 329 119 392 153
rect 426 119 489 153
rect 523 119 533 153
rect 91 103 533 119
rect 593 363 649 379
rect 593 329 603 363
rect 637 329 649 363
rect 593 291 649 329
rect 679 342 841 379
tri 679 326 695 342 ne
rect 695 326 841 342
tri 755 296 785 326 ne
rect 593 257 603 291
rect 637 257 649 291
rect 593 223 649 257
rect 593 189 603 223
rect 637 189 649 223
tri 679 280 695 296 se
rect 695 280 739 296
tri 739 280 755 296 sw
rect 679 247 755 280
rect 679 213 700 247
rect 734 213 755 247
rect 679 211 755 213
tri 679 195 695 211 ne
rect 695 195 739 211
tri 739 195 755 211 nw
rect 785 291 841 326
rect 785 257 797 291
rect 831 257 841 291
rect 785 223 841 257
rect 593 165 649 189
tri 649 165 679 195 sw
tri 755 165 785 195 se
rect 785 189 797 223
rect 831 189 841 223
rect 785 165 841 189
rect 593 153 841 165
rect 593 119 603 153
rect 637 119 700 153
rect 734 119 797 153
rect 831 119 841 153
rect 593 103 841 119
rect 1053 363 1109 379
rect 1053 329 1063 363
rect 1097 329 1109 363
rect 1053 291 1109 329
rect 1139 363 1409 379
rect 1139 334 1160 363
tri 1139 318 1155 334 ne
rect 1155 329 1160 334
rect 1194 329 1257 363
rect 1291 329 1354 363
rect 1388 329 1409 363
rect 1155 318 1409 329
rect 1439 363 1495 379
rect 1439 329 1451 363
rect 1485 329 1495 363
rect 1053 257 1063 291
rect 1097 257 1109 291
tri 1215 288 1245 318 ne
rect 1245 291 1304 318
rect 1053 223 1109 257
rect 1053 189 1063 223
rect 1097 189 1109 223
rect 1053 157 1109 189
tri 1139 272 1155 288 se
rect 1155 272 1199 288
tri 1199 272 1215 288 sw
rect 1139 238 1215 272
rect 1139 204 1160 238
rect 1194 204 1215 238
rect 1139 203 1215 204
tri 1139 187 1155 203 ne
rect 1155 187 1199 203
tri 1199 187 1215 203 nw
rect 1245 257 1257 291
rect 1291 257 1304 291
tri 1304 288 1334 318 nw
rect 1245 223 1304 257
rect 1245 189 1257 223
rect 1291 189 1304 223
tri 1334 272 1350 288 se
rect 1350 272 1393 288
tri 1393 272 1409 288 sw
rect 1334 244 1409 272
rect 1334 210 1355 244
rect 1389 210 1409 244
tri 1334 194 1350 210 ne
rect 1350 194 1393 210
tri 1393 194 1409 210 nw
tri 1109 157 1139 187 sw
tri 1215 157 1245 187 se
rect 1245 164 1304 189
tri 1304 164 1334 194 sw
tri 1409 164 1439 194 se
rect 1439 164 1495 329
rect 1245 157 1495 164
rect 1053 153 1495 157
rect 1053 119 1063 153
rect 1097 119 1257 153
rect 1291 119 1354 153
rect 1388 119 1451 153
rect 1485 119 1495 153
rect 1053 103 1495 119
rect 1555 363 1611 379
rect 1555 329 1565 363
rect 1599 329 1611 363
rect 1555 291 1611 329
rect 1641 342 1803 379
tri 1641 326 1657 342 ne
rect 1657 326 1803 342
tri 1717 296 1747 326 ne
rect 1555 257 1565 291
rect 1599 257 1611 291
rect 1555 223 1611 257
rect 1555 189 1565 223
rect 1599 189 1611 223
tri 1641 280 1657 296 se
rect 1657 280 1701 296
tri 1701 280 1717 296 sw
rect 1641 247 1717 280
rect 1641 213 1662 247
rect 1696 213 1717 247
rect 1641 211 1717 213
tri 1641 195 1657 211 ne
rect 1657 195 1701 211
tri 1701 195 1717 211 nw
rect 1747 291 1803 326
rect 1747 257 1759 291
rect 1793 257 1803 291
rect 1747 223 1803 257
rect 1555 165 1611 189
tri 1611 165 1641 195 sw
tri 1717 165 1747 195 se
rect 1747 189 1759 223
rect 1793 189 1803 223
rect 1747 165 1803 189
rect 1555 153 1803 165
rect 1555 119 1565 153
rect 1599 119 1662 153
rect 1696 119 1759 153
rect 1793 119 1803 153
rect 1555 103 1803 119
rect 2015 363 2071 379
rect 2015 329 2025 363
rect 2059 329 2071 363
rect 2015 291 2071 329
rect 2101 363 2371 379
rect 2101 334 2122 363
tri 2101 318 2117 334 ne
rect 2117 329 2122 334
rect 2156 329 2219 363
rect 2253 329 2316 363
rect 2350 329 2371 363
rect 2117 318 2371 329
rect 2401 363 2457 379
rect 2401 329 2413 363
rect 2447 329 2457 363
rect 2015 257 2025 291
rect 2059 257 2071 291
tri 2177 288 2207 318 ne
rect 2207 291 2266 318
rect 2015 223 2071 257
rect 2015 189 2025 223
rect 2059 189 2071 223
rect 2015 157 2071 189
tri 2101 272 2117 288 se
rect 2117 272 2161 288
tri 2161 272 2177 288 sw
rect 2101 238 2177 272
rect 2101 204 2122 238
rect 2156 204 2177 238
rect 2101 203 2177 204
tri 2101 187 2117 203 ne
rect 2117 187 2161 203
tri 2161 187 2177 203 nw
rect 2207 257 2219 291
rect 2253 257 2266 291
tri 2266 288 2296 318 nw
rect 2207 223 2266 257
rect 2207 189 2219 223
rect 2253 189 2266 223
tri 2296 272 2312 288 se
rect 2312 272 2355 288
tri 2355 272 2371 288 sw
rect 2296 244 2371 272
rect 2296 210 2317 244
rect 2351 210 2371 244
tri 2296 194 2312 210 ne
rect 2312 194 2355 210
tri 2355 194 2371 210 nw
tri 2071 157 2101 187 sw
tri 2177 157 2207 187 se
rect 2207 164 2266 189
tri 2266 164 2296 194 sw
tri 2371 164 2401 194 se
rect 2401 164 2457 329
rect 2207 157 2457 164
rect 2015 153 2457 157
rect 2015 119 2025 153
rect 2059 119 2219 153
rect 2253 119 2316 153
rect 2350 119 2413 153
rect 2447 119 2457 153
rect 2015 103 2457 119
rect 2517 363 2573 379
rect 2517 329 2527 363
rect 2561 329 2573 363
rect 2517 291 2573 329
rect 2603 342 2765 379
tri 2603 326 2619 342 ne
rect 2619 326 2765 342
tri 2679 296 2709 326 ne
rect 2517 257 2527 291
rect 2561 257 2573 291
rect 2517 223 2573 257
rect 2517 189 2527 223
rect 2561 189 2573 223
tri 2603 280 2619 296 se
rect 2619 280 2663 296
tri 2663 280 2679 296 sw
rect 2603 247 2679 280
rect 2603 213 2624 247
rect 2658 213 2679 247
rect 2603 211 2679 213
tri 2603 195 2619 211 ne
rect 2619 195 2663 211
tri 2663 195 2679 211 nw
rect 2709 291 2765 326
rect 2709 257 2721 291
rect 2755 257 2765 291
rect 2709 223 2765 257
rect 2517 165 2573 189
tri 2573 165 2603 195 sw
tri 2679 165 2709 195 se
rect 2709 189 2721 223
rect 2755 189 2765 223
rect 2709 165 2765 189
rect 2517 153 2765 165
rect 2517 119 2527 153
rect 2561 119 2624 153
rect 2658 119 2721 153
rect 2755 119 2765 153
rect 2517 103 2765 119
rect 2977 363 3033 379
rect 2977 329 2987 363
rect 3021 329 3033 363
rect 2977 291 3033 329
rect 3063 363 3333 379
rect 3063 334 3084 363
tri 3063 318 3079 334 ne
rect 3079 329 3084 334
rect 3118 329 3181 363
rect 3215 329 3278 363
rect 3312 329 3333 363
rect 3079 318 3333 329
rect 3363 363 3419 379
rect 3363 329 3375 363
rect 3409 329 3419 363
rect 2977 257 2987 291
rect 3021 257 3033 291
tri 3139 288 3169 318 ne
rect 3169 291 3228 318
rect 2977 223 3033 257
rect 2977 189 2987 223
rect 3021 189 3033 223
rect 2977 157 3033 189
tri 3063 272 3079 288 se
rect 3079 272 3123 288
tri 3123 272 3139 288 sw
rect 3063 238 3139 272
rect 3063 204 3084 238
rect 3118 204 3139 238
rect 3063 203 3139 204
tri 3063 187 3079 203 ne
rect 3079 187 3123 203
tri 3123 187 3139 203 nw
rect 3169 257 3181 291
rect 3215 257 3228 291
tri 3228 288 3258 318 nw
rect 3169 223 3228 257
rect 3169 189 3181 223
rect 3215 189 3228 223
tri 3258 272 3274 288 se
rect 3274 272 3317 288
tri 3317 272 3333 288 sw
rect 3258 244 3333 272
rect 3258 210 3279 244
rect 3313 210 3333 244
tri 3258 194 3274 210 ne
rect 3274 194 3317 210
tri 3317 194 3333 210 nw
tri 3033 157 3063 187 sw
tri 3139 157 3169 187 se
rect 3169 164 3228 189
tri 3228 164 3258 194 sw
tri 3333 164 3363 194 se
rect 3363 164 3419 329
rect 3169 157 3419 164
rect 2977 153 3419 157
rect 2977 119 2987 153
rect 3021 119 3181 153
rect 3215 119 3278 153
rect 3312 119 3375 153
rect 3409 119 3419 153
rect 2977 103 3419 119
rect 3479 363 3535 379
rect 3479 329 3489 363
rect 3523 329 3535 363
rect 3479 291 3535 329
rect 3565 342 3727 379
tri 3565 326 3581 342 ne
rect 3581 326 3727 342
tri 3641 296 3671 326 ne
rect 3479 257 3489 291
rect 3523 257 3535 291
rect 3479 223 3535 257
rect 3479 189 3489 223
rect 3523 189 3535 223
tri 3565 280 3581 296 se
rect 3581 280 3625 296
tri 3625 280 3641 296 sw
rect 3565 247 3641 280
rect 3565 213 3586 247
rect 3620 213 3641 247
rect 3565 211 3641 213
tri 3565 195 3581 211 ne
rect 3581 195 3625 211
tri 3625 195 3641 211 nw
rect 3671 291 3727 326
rect 3671 257 3683 291
rect 3717 257 3727 291
rect 3671 223 3727 257
rect 3479 165 3535 189
tri 3535 165 3565 195 sw
tri 3641 165 3671 195 se
rect 3671 189 3683 223
rect 3717 189 3727 223
rect 3671 165 3727 189
rect 3479 153 3727 165
rect 3479 119 3489 153
rect 3523 119 3586 153
rect 3620 119 3683 153
rect 3717 119 3727 153
rect 3479 103 3727 119
rect 3939 363 3995 379
rect 3939 329 3949 363
rect 3983 329 3995 363
rect 3939 291 3995 329
rect 4025 363 4295 379
rect 4025 334 4046 363
tri 4025 318 4041 334 ne
rect 4041 329 4046 334
rect 4080 329 4143 363
rect 4177 329 4240 363
rect 4274 329 4295 363
rect 4041 318 4295 329
rect 4325 363 4381 379
rect 4325 329 4337 363
rect 4371 329 4381 363
rect 3939 257 3949 291
rect 3983 257 3995 291
tri 4101 288 4131 318 ne
rect 4131 291 4190 318
rect 3939 223 3995 257
rect 3939 189 3949 223
rect 3983 189 3995 223
rect 3939 157 3995 189
tri 4025 272 4041 288 se
rect 4041 272 4085 288
tri 4085 272 4101 288 sw
rect 4025 238 4101 272
rect 4025 204 4046 238
rect 4080 204 4101 238
rect 4025 203 4101 204
tri 4025 187 4041 203 ne
rect 4041 187 4085 203
tri 4085 187 4101 203 nw
rect 4131 257 4143 291
rect 4177 257 4190 291
tri 4190 288 4220 318 nw
rect 4131 223 4190 257
rect 4131 189 4143 223
rect 4177 189 4190 223
tri 4220 272 4236 288 se
rect 4236 272 4279 288
tri 4279 272 4295 288 sw
rect 4220 244 4295 272
rect 4220 210 4241 244
rect 4275 210 4295 244
tri 4220 194 4236 210 ne
rect 4236 194 4279 210
tri 4279 194 4295 210 nw
tri 3995 157 4025 187 sw
tri 4101 157 4131 187 se
rect 4131 164 4190 189
tri 4190 164 4220 194 sw
tri 4295 164 4325 194 se
rect 4325 164 4381 329
rect 4131 157 4381 164
rect 3939 153 4381 157
rect 3939 119 3949 153
rect 3983 119 4143 153
rect 4177 119 4240 153
rect 4274 119 4337 153
rect 4371 119 4381 153
rect 3939 103 4381 119
rect 4441 363 4497 379
rect 4441 329 4451 363
rect 4485 329 4497 363
rect 4441 291 4497 329
rect 4527 342 4689 379
tri 4527 326 4543 342 ne
rect 4543 326 4689 342
tri 4603 296 4633 326 ne
rect 4441 257 4451 291
rect 4485 257 4497 291
rect 4441 223 4497 257
rect 4441 189 4451 223
rect 4485 189 4497 223
tri 4527 280 4543 296 se
rect 4543 280 4587 296
tri 4587 280 4603 296 sw
rect 4527 247 4603 280
rect 4527 213 4548 247
rect 4582 213 4603 247
rect 4527 211 4603 213
tri 4527 195 4543 211 ne
rect 4543 195 4587 211
tri 4587 195 4603 211 nw
rect 4633 291 4689 326
rect 4633 257 4645 291
rect 4679 257 4689 291
rect 4633 223 4689 257
rect 4441 165 4497 189
tri 4497 165 4527 195 sw
tri 4603 165 4633 195 se
rect 4633 189 4645 223
rect 4679 189 4689 223
rect 4633 165 4689 189
rect 4441 153 4689 165
rect 4441 119 4451 153
rect 4485 119 4548 153
rect 4582 119 4645 153
rect 4679 119 4689 153
rect 4441 103 4689 119
rect 4901 363 4957 379
rect 4901 329 4911 363
rect 4945 329 4957 363
rect 4901 291 4957 329
rect 4987 363 5257 379
rect 4987 334 5008 363
tri 4987 318 5003 334 ne
rect 5003 329 5008 334
rect 5042 329 5105 363
rect 5139 329 5202 363
rect 5236 329 5257 363
rect 5003 318 5257 329
rect 5287 363 5343 379
rect 5287 329 5299 363
rect 5333 329 5343 363
rect 4901 257 4911 291
rect 4945 257 4957 291
tri 5063 288 5093 318 ne
rect 5093 291 5152 318
rect 4901 223 4957 257
rect 4901 189 4911 223
rect 4945 189 4957 223
rect 4901 157 4957 189
tri 4987 272 5003 288 se
rect 5003 272 5047 288
tri 5047 272 5063 288 sw
rect 4987 238 5063 272
rect 4987 204 5008 238
rect 5042 204 5063 238
rect 4987 203 5063 204
tri 4987 187 5003 203 ne
rect 5003 187 5047 203
tri 5047 187 5063 203 nw
rect 5093 257 5105 291
rect 5139 257 5152 291
tri 5152 288 5182 318 nw
rect 5093 223 5152 257
rect 5093 189 5105 223
rect 5139 189 5152 223
tri 5182 272 5198 288 se
rect 5198 272 5241 288
tri 5241 272 5257 288 sw
rect 5182 244 5257 272
rect 5182 210 5203 244
rect 5237 210 5257 244
tri 5182 194 5198 210 ne
rect 5198 194 5241 210
tri 5241 194 5257 210 nw
tri 4957 157 4987 187 sw
tri 5063 157 5093 187 se
rect 5093 164 5152 189
tri 5152 164 5182 194 sw
tri 5257 164 5287 194 se
rect 5287 164 5343 329
rect 5093 157 5343 164
rect 4901 153 5343 157
rect 4901 119 4911 153
rect 4945 119 5105 153
rect 5139 119 5202 153
rect 5236 119 5299 153
rect 5333 119 5343 153
rect 4901 103 5343 119
rect 5403 363 5459 379
rect 5403 329 5413 363
rect 5447 329 5459 363
rect 5403 291 5459 329
rect 5489 342 5651 379
tri 5489 326 5505 342 ne
rect 5505 326 5651 342
tri 5565 296 5595 326 ne
rect 5403 257 5413 291
rect 5447 257 5459 291
rect 5403 223 5459 257
rect 5403 189 5413 223
rect 5447 189 5459 223
tri 5489 280 5505 296 se
rect 5505 280 5549 296
tri 5549 280 5565 296 sw
rect 5489 247 5565 280
rect 5489 213 5510 247
rect 5544 213 5565 247
rect 5489 211 5565 213
tri 5489 195 5505 211 ne
rect 5505 195 5549 211
tri 5549 195 5565 211 nw
rect 5595 291 5651 326
rect 5595 257 5607 291
rect 5641 257 5651 291
rect 5595 223 5651 257
rect 5403 165 5459 189
tri 5459 165 5489 195 sw
tri 5565 165 5595 195 se
rect 5595 189 5607 223
rect 5641 189 5651 223
rect 5595 165 5651 189
rect 5403 153 5651 165
rect 5403 119 5413 153
rect 5447 119 5510 153
rect 5544 119 5607 153
rect 5641 119 5651 153
rect 5403 103 5651 119
rect 5863 363 5919 379
rect 5863 329 5873 363
rect 5907 329 5919 363
rect 5863 291 5919 329
rect 5949 363 6219 379
rect 5949 334 5970 363
tri 5949 318 5965 334 ne
rect 5965 329 5970 334
rect 6004 329 6067 363
rect 6101 329 6164 363
rect 6198 329 6219 363
rect 5965 318 6219 329
rect 6249 363 6305 379
rect 6249 329 6261 363
rect 6295 329 6305 363
rect 5863 257 5873 291
rect 5907 257 5919 291
tri 6025 288 6055 318 ne
rect 6055 291 6114 318
rect 5863 223 5919 257
rect 5863 189 5873 223
rect 5907 189 5919 223
rect 5863 157 5919 189
tri 5949 272 5965 288 se
rect 5965 272 6009 288
tri 6009 272 6025 288 sw
rect 5949 238 6025 272
rect 5949 204 5970 238
rect 6004 204 6025 238
rect 5949 203 6025 204
tri 5949 187 5965 203 ne
rect 5965 187 6009 203
tri 6009 187 6025 203 nw
rect 6055 257 6067 291
rect 6101 257 6114 291
tri 6114 288 6144 318 nw
rect 6055 223 6114 257
rect 6055 189 6067 223
rect 6101 189 6114 223
tri 6144 272 6160 288 se
rect 6160 272 6203 288
tri 6203 272 6219 288 sw
rect 6144 244 6219 272
rect 6144 210 6165 244
rect 6199 210 6219 244
tri 6144 194 6160 210 ne
rect 6160 194 6203 210
tri 6203 194 6219 210 nw
tri 5919 157 5949 187 sw
tri 6025 157 6055 187 se
rect 6055 164 6114 189
tri 6114 164 6144 194 sw
tri 6219 164 6249 194 se
rect 6249 164 6305 329
rect 6055 157 6305 164
rect 5863 153 6305 157
rect 5863 119 5873 153
rect 5907 119 6067 153
rect 6101 119 6164 153
rect 6198 119 6261 153
rect 6295 119 6305 153
rect 5863 103 6305 119
rect 6365 363 6421 379
rect 6365 329 6375 363
rect 6409 329 6421 363
rect 6365 291 6421 329
rect 6451 342 6613 379
tri 6451 326 6467 342 ne
rect 6467 326 6613 342
tri 6527 296 6557 326 ne
rect 6365 257 6375 291
rect 6409 257 6421 291
rect 6365 223 6421 257
rect 6365 189 6375 223
rect 6409 189 6421 223
tri 6451 280 6467 296 se
rect 6467 280 6511 296
tri 6511 280 6527 296 sw
rect 6451 247 6527 280
rect 6451 213 6472 247
rect 6506 213 6527 247
rect 6451 211 6527 213
tri 6451 195 6467 211 ne
rect 6467 195 6511 211
tri 6511 195 6527 211 nw
rect 6557 291 6613 326
rect 6557 257 6569 291
rect 6603 257 6613 291
rect 6557 223 6613 257
rect 6365 165 6421 189
tri 6421 165 6451 195 sw
tri 6527 165 6557 195 se
rect 6557 189 6569 223
rect 6603 189 6613 223
rect 6557 165 6613 189
rect 6365 153 6613 165
rect 6365 119 6375 153
rect 6409 119 6472 153
rect 6506 119 6569 153
rect 6603 119 6613 153
rect 6365 103 6613 119
rect 6825 363 6881 379
rect 6825 329 6835 363
rect 6869 329 6881 363
rect 6825 291 6881 329
rect 6911 363 7181 379
rect 6911 334 6932 363
tri 6911 318 6927 334 ne
rect 6927 329 6932 334
rect 6966 329 7029 363
rect 7063 329 7126 363
rect 7160 329 7181 363
rect 6927 318 7181 329
rect 7211 363 7267 379
rect 7211 329 7223 363
rect 7257 329 7267 363
rect 6825 257 6835 291
rect 6869 257 6881 291
tri 6987 288 7017 318 ne
rect 7017 291 7076 318
rect 6825 223 6881 257
rect 6825 189 6835 223
rect 6869 189 6881 223
rect 6825 157 6881 189
tri 6911 272 6927 288 se
rect 6927 272 6971 288
tri 6971 272 6987 288 sw
rect 6911 238 6987 272
rect 6911 204 6932 238
rect 6966 204 6987 238
rect 6911 203 6987 204
tri 6911 187 6927 203 ne
rect 6927 187 6971 203
tri 6971 187 6987 203 nw
rect 7017 257 7029 291
rect 7063 257 7076 291
tri 7076 288 7106 318 nw
rect 7017 223 7076 257
rect 7017 189 7029 223
rect 7063 189 7076 223
tri 7106 272 7122 288 se
rect 7122 272 7165 288
tri 7165 272 7181 288 sw
rect 7106 244 7181 272
rect 7106 210 7127 244
rect 7161 210 7181 244
tri 7106 194 7122 210 ne
rect 7122 194 7165 210
tri 7165 194 7181 210 nw
tri 6881 157 6911 187 sw
tri 6987 157 7017 187 se
rect 7017 164 7076 189
tri 7076 164 7106 194 sw
tri 7181 164 7211 194 se
rect 7211 164 7267 329
rect 7017 157 7267 164
rect 6825 153 7267 157
rect 6825 119 6835 153
rect 6869 119 7029 153
rect 7063 119 7126 153
rect 7160 119 7223 153
rect 7257 119 7267 153
rect 6825 103 7267 119
rect 7327 363 7383 379
rect 7327 329 7337 363
rect 7371 329 7383 363
rect 7327 291 7383 329
rect 7413 342 7575 379
tri 7413 326 7429 342 ne
rect 7429 326 7575 342
tri 7489 296 7519 326 ne
rect 7327 257 7337 291
rect 7371 257 7383 291
rect 7327 223 7383 257
rect 7327 189 7337 223
rect 7371 189 7383 223
tri 7413 280 7429 296 se
rect 7429 280 7473 296
tri 7473 280 7489 296 sw
rect 7413 247 7489 280
rect 7413 213 7434 247
rect 7468 213 7489 247
rect 7413 211 7489 213
tri 7413 195 7429 211 ne
rect 7429 195 7473 211
tri 7473 195 7489 211 nw
rect 7519 291 7575 326
rect 7519 257 7531 291
rect 7565 257 7575 291
rect 7519 223 7575 257
rect 7327 165 7383 189
tri 7383 165 7413 195 sw
tri 7489 165 7519 195 se
rect 7519 189 7531 223
rect 7565 189 7575 223
rect 7519 165 7575 189
rect 7327 153 7575 165
rect 7327 119 7337 153
rect 7371 119 7434 153
rect 7468 119 7531 153
rect 7565 119 7575 153
rect 7327 103 7575 119
rect 7787 363 7843 379
rect 7787 329 7797 363
rect 7831 329 7843 363
rect 7787 291 7843 329
rect 7873 363 8143 379
rect 7873 334 7894 363
tri 7873 318 7889 334 ne
rect 7889 329 7894 334
rect 7928 329 7991 363
rect 8025 329 8088 363
rect 8122 329 8143 363
rect 7889 318 8143 329
rect 8173 363 8229 379
rect 8173 329 8185 363
rect 8219 329 8229 363
rect 7787 257 7797 291
rect 7831 257 7843 291
tri 7949 288 7979 318 ne
rect 7979 291 8038 318
rect 7787 223 7843 257
rect 7787 189 7797 223
rect 7831 189 7843 223
rect 7787 157 7843 189
tri 7873 272 7889 288 se
rect 7889 272 7933 288
tri 7933 272 7949 288 sw
rect 7873 238 7949 272
rect 7873 204 7894 238
rect 7928 204 7949 238
rect 7873 203 7949 204
tri 7873 187 7889 203 ne
rect 7889 187 7933 203
tri 7933 187 7949 203 nw
rect 7979 257 7991 291
rect 8025 257 8038 291
tri 8038 288 8068 318 nw
rect 7979 223 8038 257
rect 7979 189 7991 223
rect 8025 189 8038 223
tri 8068 272 8084 288 se
rect 8084 272 8127 288
tri 8127 272 8143 288 sw
rect 8068 244 8143 272
rect 8068 210 8089 244
rect 8123 210 8143 244
tri 8068 194 8084 210 ne
rect 8084 194 8127 210
tri 8127 194 8143 210 nw
tri 7843 157 7873 187 sw
tri 7949 157 7979 187 se
rect 7979 164 8038 189
tri 8038 164 8068 194 sw
tri 8143 164 8173 194 se
rect 8173 164 8229 329
rect 7979 157 8229 164
rect 7787 153 8229 157
rect 7787 119 7797 153
rect 7831 119 7991 153
rect 8025 119 8088 153
rect 8122 119 8185 153
rect 8219 119 8229 153
rect 7787 103 8229 119
rect 8289 363 8345 379
rect 8289 329 8299 363
rect 8333 329 8345 363
rect 8289 291 8345 329
rect 8375 342 8537 379
tri 8375 326 8391 342 ne
rect 8391 326 8537 342
tri 8451 296 8481 326 ne
rect 8289 257 8299 291
rect 8333 257 8345 291
rect 8289 223 8345 257
rect 8289 189 8299 223
rect 8333 189 8345 223
tri 8375 280 8391 296 se
rect 8391 280 8435 296
tri 8435 280 8451 296 sw
rect 8375 247 8451 280
rect 8375 213 8396 247
rect 8430 213 8451 247
rect 8375 211 8451 213
tri 8375 195 8391 211 ne
rect 8391 195 8435 211
tri 8435 195 8451 211 nw
rect 8481 291 8537 326
rect 8481 257 8493 291
rect 8527 257 8537 291
rect 8481 223 8537 257
rect 8289 165 8345 189
tri 8345 165 8375 195 sw
tri 8451 165 8481 195 se
rect 8481 189 8493 223
rect 8527 189 8537 223
rect 8481 165 8537 189
rect 8289 153 8537 165
rect 8289 119 8299 153
rect 8333 119 8396 153
rect 8430 119 8493 153
rect 8527 119 8537 153
rect 8289 103 8537 119
rect 8749 363 8805 379
rect 8749 329 8759 363
rect 8793 329 8805 363
rect 8749 291 8805 329
rect 8835 363 9105 379
rect 8835 334 8856 363
tri 8835 318 8851 334 ne
rect 8851 329 8856 334
rect 8890 329 8953 363
rect 8987 329 9050 363
rect 9084 329 9105 363
rect 8851 318 9105 329
rect 9135 363 9191 379
rect 9135 329 9147 363
rect 9181 329 9191 363
rect 8749 257 8759 291
rect 8793 257 8805 291
tri 8911 288 8941 318 ne
rect 8941 291 9000 318
rect 8749 223 8805 257
rect 8749 189 8759 223
rect 8793 189 8805 223
rect 8749 157 8805 189
tri 8835 272 8851 288 se
rect 8851 272 8895 288
tri 8895 272 8911 288 sw
rect 8835 238 8911 272
rect 8835 204 8856 238
rect 8890 204 8911 238
rect 8835 203 8911 204
tri 8835 187 8851 203 ne
rect 8851 187 8895 203
tri 8895 187 8911 203 nw
rect 8941 257 8953 291
rect 8987 257 9000 291
tri 9000 288 9030 318 nw
rect 8941 223 9000 257
rect 8941 189 8953 223
rect 8987 189 9000 223
tri 9030 272 9046 288 se
rect 9046 272 9089 288
tri 9089 272 9105 288 sw
rect 9030 244 9105 272
rect 9030 210 9051 244
rect 9085 210 9105 244
tri 9030 194 9046 210 ne
rect 9046 194 9089 210
tri 9089 194 9105 210 nw
tri 8805 157 8835 187 sw
tri 8911 157 8941 187 se
rect 8941 164 9000 189
tri 9000 164 9030 194 sw
tri 9105 164 9135 194 se
rect 9135 164 9191 329
rect 8941 157 9191 164
rect 8749 153 9191 157
rect 8749 119 8759 153
rect 8793 119 8953 153
rect 8987 119 9050 153
rect 9084 119 9147 153
rect 9181 119 9191 153
rect 8749 103 9191 119
rect 9251 363 9307 379
rect 9251 329 9261 363
rect 9295 329 9307 363
rect 9251 291 9307 329
rect 9337 342 9499 379
tri 9337 326 9353 342 ne
rect 9353 326 9499 342
tri 9413 296 9443 326 ne
rect 9251 257 9261 291
rect 9295 257 9307 291
rect 9251 223 9307 257
rect 9251 189 9261 223
rect 9295 189 9307 223
tri 9337 280 9353 296 se
rect 9353 280 9397 296
tri 9397 280 9413 296 sw
rect 9337 247 9413 280
rect 9337 213 9358 247
rect 9392 213 9413 247
rect 9337 211 9413 213
tri 9337 195 9353 211 ne
rect 9353 195 9397 211
tri 9397 195 9413 211 nw
rect 9443 291 9499 326
rect 9443 257 9455 291
rect 9489 257 9499 291
rect 9443 223 9499 257
rect 9251 165 9307 189
tri 9307 165 9337 195 sw
tri 9413 165 9443 195 se
rect 9443 189 9455 223
rect 9489 189 9499 223
rect 9443 165 9499 189
rect 9251 153 9499 165
rect 9251 119 9261 153
rect 9295 119 9358 153
rect 9392 119 9455 153
rect 9489 119 9499 153
rect 9251 103 9499 119
rect 9711 363 9767 379
rect 9711 329 9721 363
rect 9755 329 9767 363
rect 9711 291 9767 329
rect 9797 363 10067 379
rect 9797 334 9818 363
tri 9797 318 9813 334 ne
rect 9813 329 9818 334
rect 9852 329 9915 363
rect 9949 329 10012 363
rect 10046 329 10067 363
rect 9813 318 10067 329
rect 10097 363 10153 379
rect 10097 329 10109 363
rect 10143 329 10153 363
rect 9711 257 9721 291
rect 9755 257 9767 291
tri 9873 288 9903 318 ne
rect 9903 291 9962 318
rect 9711 223 9767 257
rect 9711 189 9721 223
rect 9755 189 9767 223
rect 9711 157 9767 189
tri 9797 272 9813 288 se
rect 9813 272 9857 288
tri 9857 272 9873 288 sw
rect 9797 238 9873 272
rect 9797 204 9818 238
rect 9852 204 9873 238
rect 9797 203 9873 204
tri 9797 187 9813 203 ne
rect 9813 187 9857 203
tri 9857 187 9873 203 nw
rect 9903 257 9915 291
rect 9949 257 9962 291
tri 9962 288 9992 318 nw
rect 9903 223 9962 257
rect 9903 189 9915 223
rect 9949 189 9962 223
tri 9992 272 10008 288 se
rect 10008 272 10051 288
tri 10051 272 10067 288 sw
rect 9992 244 10067 272
rect 9992 210 10013 244
rect 10047 210 10067 244
tri 9992 194 10008 210 ne
rect 10008 194 10051 210
tri 10051 194 10067 210 nw
tri 9767 157 9797 187 sw
tri 9873 157 9903 187 se
rect 9903 164 9962 189
tri 9962 164 9992 194 sw
tri 10067 164 10097 194 se
rect 10097 164 10153 329
rect 9903 157 10153 164
rect 9711 153 10153 157
rect 9711 119 9721 153
rect 9755 119 9915 153
rect 9949 119 10012 153
rect 10046 119 10109 153
rect 10143 119 10153 153
rect 9711 103 10153 119
rect 10213 363 10269 379
rect 10213 329 10223 363
rect 10257 329 10269 363
rect 10213 291 10269 329
rect 10299 342 10461 379
tri 10299 326 10315 342 ne
rect 10315 326 10461 342
tri 10375 296 10405 326 ne
rect 10213 257 10223 291
rect 10257 257 10269 291
rect 10213 223 10269 257
rect 10213 189 10223 223
rect 10257 189 10269 223
tri 10299 280 10315 296 se
rect 10315 280 10359 296
tri 10359 280 10375 296 sw
rect 10299 247 10375 280
rect 10299 213 10320 247
rect 10354 213 10375 247
rect 10299 211 10375 213
tri 10299 195 10315 211 ne
rect 10315 195 10359 211
tri 10359 195 10375 211 nw
rect 10405 291 10461 326
rect 10405 257 10417 291
rect 10451 257 10461 291
rect 10405 223 10461 257
rect 10213 165 10269 189
tri 10269 165 10299 195 sw
tri 10375 165 10405 195 se
rect 10405 189 10417 223
rect 10451 189 10461 223
rect 10405 165 10461 189
rect 10213 153 10461 165
rect 10213 119 10223 153
rect 10257 119 10320 153
rect 10354 119 10417 153
rect 10451 119 10461 153
rect 10213 103 10461 119
rect 10673 363 10729 379
rect 10673 329 10683 363
rect 10717 329 10729 363
rect 10673 291 10729 329
rect 10759 363 11029 379
rect 10759 334 10780 363
tri 10759 318 10775 334 ne
rect 10775 329 10780 334
rect 10814 329 10877 363
rect 10911 329 10974 363
rect 11008 329 11029 363
rect 10775 318 11029 329
rect 11059 363 11115 379
rect 11059 329 11071 363
rect 11105 329 11115 363
rect 10673 257 10683 291
rect 10717 257 10729 291
tri 10835 288 10865 318 ne
rect 10865 291 10924 318
rect 10673 223 10729 257
rect 10673 189 10683 223
rect 10717 189 10729 223
rect 10673 157 10729 189
tri 10759 272 10775 288 se
rect 10775 272 10819 288
tri 10819 272 10835 288 sw
rect 10759 238 10835 272
rect 10759 204 10780 238
rect 10814 204 10835 238
rect 10759 203 10835 204
tri 10759 187 10775 203 ne
rect 10775 187 10819 203
tri 10819 187 10835 203 nw
rect 10865 257 10877 291
rect 10911 257 10924 291
tri 10924 288 10954 318 nw
rect 10865 223 10924 257
rect 10865 189 10877 223
rect 10911 189 10924 223
tri 10954 272 10970 288 se
rect 10970 272 11013 288
tri 11013 272 11029 288 sw
rect 10954 244 11029 272
rect 10954 210 10975 244
rect 11009 210 11029 244
tri 10954 194 10970 210 ne
rect 10970 194 11013 210
tri 11013 194 11029 210 nw
tri 10729 157 10759 187 sw
tri 10835 157 10865 187 se
rect 10865 164 10924 189
tri 10924 164 10954 194 sw
tri 11029 164 11059 194 se
rect 11059 164 11115 329
rect 10865 157 11115 164
rect 10673 153 11115 157
rect 10673 119 10683 153
rect 10717 119 10877 153
rect 10911 119 10974 153
rect 11008 119 11071 153
rect 11105 119 11115 153
rect 10673 103 11115 119
rect 11175 363 11231 379
rect 11175 329 11185 363
rect 11219 329 11231 363
rect 11175 291 11231 329
rect 11261 342 11423 379
tri 11261 326 11277 342 ne
rect 11277 326 11423 342
tri 11337 296 11367 326 ne
rect 11175 257 11185 291
rect 11219 257 11231 291
rect 11175 223 11231 257
rect 11175 189 11185 223
rect 11219 189 11231 223
tri 11261 280 11277 296 se
rect 11277 280 11321 296
tri 11321 280 11337 296 sw
rect 11261 247 11337 280
rect 11261 213 11282 247
rect 11316 213 11337 247
rect 11261 211 11337 213
tri 11261 195 11277 211 ne
rect 11277 195 11321 211
tri 11321 195 11337 211 nw
rect 11367 291 11423 326
rect 11367 257 11379 291
rect 11413 257 11423 291
rect 11367 223 11423 257
rect 11175 165 11231 189
tri 11231 165 11261 195 sw
tri 11337 165 11367 195 se
rect 11367 189 11379 223
rect 11413 189 11423 223
rect 11367 165 11423 189
rect 11175 153 11423 165
rect 11175 119 11185 153
rect 11219 119 11282 153
rect 11316 119 11379 153
rect 11413 119 11423 153
rect 11175 103 11423 119
rect 11635 363 11691 379
rect 11635 329 11645 363
rect 11679 329 11691 363
rect 11635 291 11691 329
rect 11721 363 11991 379
rect 11721 334 11742 363
tri 11721 318 11737 334 ne
rect 11737 329 11742 334
rect 11776 329 11839 363
rect 11873 329 11936 363
rect 11970 329 11991 363
rect 11737 318 11991 329
rect 12021 363 12077 379
rect 12021 329 12033 363
rect 12067 329 12077 363
rect 11635 257 11645 291
rect 11679 257 11691 291
tri 11797 288 11827 318 ne
rect 11827 291 11886 318
rect 11635 223 11691 257
rect 11635 189 11645 223
rect 11679 189 11691 223
rect 11635 157 11691 189
tri 11721 272 11737 288 se
rect 11737 272 11781 288
tri 11781 272 11797 288 sw
rect 11721 238 11797 272
rect 11721 204 11742 238
rect 11776 204 11797 238
rect 11721 203 11797 204
tri 11721 187 11737 203 ne
rect 11737 187 11781 203
tri 11781 187 11797 203 nw
rect 11827 257 11839 291
rect 11873 257 11886 291
tri 11886 288 11916 318 nw
rect 11827 223 11886 257
rect 11827 189 11839 223
rect 11873 189 11886 223
tri 11916 272 11932 288 se
rect 11932 272 11975 288
tri 11975 272 11991 288 sw
rect 11916 244 11991 272
rect 11916 210 11937 244
rect 11971 210 11991 244
tri 11916 194 11932 210 ne
rect 11932 194 11975 210
tri 11975 194 11991 210 nw
tri 11691 157 11721 187 sw
tri 11797 157 11827 187 se
rect 11827 164 11886 189
tri 11886 164 11916 194 sw
tri 11991 164 12021 194 se
rect 12021 164 12077 329
rect 11827 157 12077 164
rect 11635 153 12077 157
rect 11635 119 11645 153
rect 11679 119 11839 153
rect 11873 119 11936 153
rect 11970 119 12033 153
rect 12067 119 12077 153
rect 11635 103 12077 119
rect 12137 363 12193 379
rect 12137 329 12147 363
rect 12181 329 12193 363
rect 12137 291 12193 329
rect 12223 342 12385 379
tri 12223 326 12239 342 ne
rect 12239 326 12385 342
tri 12299 296 12329 326 ne
rect 12137 257 12147 291
rect 12181 257 12193 291
rect 12137 223 12193 257
rect 12137 189 12147 223
rect 12181 189 12193 223
tri 12223 280 12239 296 se
rect 12239 280 12283 296
tri 12283 280 12299 296 sw
rect 12223 247 12299 280
rect 12223 213 12244 247
rect 12278 213 12299 247
rect 12223 211 12299 213
tri 12223 195 12239 211 ne
rect 12239 195 12283 211
tri 12283 195 12299 211 nw
rect 12329 291 12385 326
rect 12329 257 12341 291
rect 12375 257 12385 291
rect 12329 223 12385 257
rect 12137 165 12193 189
tri 12193 165 12223 195 sw
tri 12299 165 12329 195 se
rect 12329 189 12341 223
rect 12375 189 12385 223
rect 12329 165 12385 189
rect 12137 153 12385 165
rect 12137 119 12147 153
rect 12181 119 12244 153
rect 12278 119 12341 153
rect 12375 119 12385 153
rect 12137 103 12385 119
rect 12597 363 12653 379
rect 12597 329 12607 363
rect 12641 329 12653 363
rect 12597 291 12653 329
rect 12683 363 12953 379
rect 12683 334 12704 363
tri 12683 318 12699 334 ne
rect 12699 329 12704 334
rect 12738 329 12801 363
rect 12835 329 12898 363
rect 12932 329 12953 363
rect 12699 318 12953 329
rect 12983 363 13039 379
rect 12983 329 12995 363
rect 13029 329 13039 363
rect 12597 257 12607 291
rect 12641 257 12653 291
tri 12759 288 12789 318 ne
rect 12789 291 12848 318
rect 12597 223 12653 257
rect 12597 189 12607 223
rect 12641 189 12653 223
rect 12597 157 12653 189
tri 12683 272 12699 288 se
rect 12699 272 12743 288
tri 12743 272 12759 288 sw
rect 12683 238 12759 272
rect 12683 204 12704 238
rect 12738 204 12759 238
rect 12683 203 12759 204
tri 12683 187 12699 203 ne
rect 12699 187 12743 203
tri 12743 187 12759 203 nw
rect 12789 257 12801 291
rect 12835 257 12848 291
tri 12848 288 12878 318 nw
rect 12789 223 12848 257
rect 12789 189 12801 223
rect 12835 189 12848 223
tri 12878 272 12894 288 se
rect 12894 272 12937 288
tri 12937 272 12953 288 sw
rect 12878 244 12953 272
rect 12878 210 12899 244
rect 12933 210 12953 244
tri 12878 194 12894 210 ne
rect 12894 194 12937 210
tri 12937 194 12953 210 nw
tri 12653 157 12683 187 sw
tri 12759 157 12789 187 se
rect 12789 164 12848 189
tri 12848 164 12878 194 sw
tri 12953 164 12983 194 se
rect 12983 164 13039 329
rect 12789 157 13039 164
rect 12597 153 13039 157
rect 12597 119 12607 153
rect 12641 119 12801 153
rect 12835 119 12898 153
rect 12932 119 12995 153
rect 13029 119 13039 153
rect 12597 103 13039 119
rect 13099 363 13155 379
rect 13099 329 13109 363
rect 13143 329 13155 363
rect 13099 291 13155 329
rect 13185 342 13347 379
tri 13185 326 13201 342 ne
rect 13201 326 13347 342
tri 13261 296 13291 326 ne
rect 13099 257 13109 291
rect 13143 257 13155 291
rect 13099 223 13155 257
rect 13099 189 13109 223
rect 13143 189 13155 223
tri 13185 280 13201 296 se
rect 13201 280 13245 296
tri 13245 280 13261 296 sw
rect 13185 247 13261 280
rect 13185 213 13206 247
rect 13240 213 13261 247
rect 13185 211 13261 213
tri 13185 195 13201 211 ne
rect 13201 195 13245 211
tri 13245 195 13261 211 nw
rect 13291 291 13347 326
rect 13291 257 13303 291
rect 13337 257 13347 291
rect 13291 223 13347 257
rect 13099 165 13155 189
tri 13155 165 13185 195 sw
tri 13261 165 13291 195 se
rect 13291 189 13303 223
rect 13337 189 13347 223
rect 13291 165 13347 189
rect 13099 153 13347 165
rect 13099 119 13109 153
rect 13143 119 13206 153
rect 13240 119 13303 153
rect 13337 119 13347 153
rect 13099 103 13347 119
rect 13559 363 13615 379
rect 13559 329 13569 363
rect 13603 329 13615 363
rect 13559 291 13615 329
rect 13645 363 13915 379
rect 13645 334 13666 363
tri 13645 318 13661 334 ne
rect 13661 329 13666 334
rect 13700 329 13763 363
rect 13797 329 13860 363
rect 13894 329 13915 363
rect 13661 318 13915 329
rect 13945 363 14001 379
rect 13945 329 13957 363
rect 13991 329 14001 363
rect 13559 257 13569 291
rect 13603 257 13615 291
tri 13721 288 13751 318 ne
rect 13751 291 13810 318
rect 13559 223 13615 257
rect 13559 189 13569 223
rect 13603 189 13615 223
rect 13559 157 13615 189
tri 13645 272 13661 288 se
rect 13661 272 13705 288
tri 13705 272 13721 288 sw
rect 13645 238 13721 272
rect 13645 204 13666 238
rect 13700 204 13721 238
rect 13645 203 13721 204
tri 13645 187 13661 203 ne
rect 13661 187 13705 203
tri 13705 187 13721 203 nw
rect 13751 257 13763 291
rect 13797 257 13810 291
tri 13810 288 13840 318 nw
rect 13751 223 13810 257
rect 13751 189 13763 223
rect 13797 189 13810 223
tri 13840 272 13856 288 se
rect 13856 272 13899 288
tri 13899 272 13915 288 sw
rect 13840 244 13915 272
rect 13840 210 13861 244
rect 13895 210 13915 244
tri 13840 194 13856 210 ne
rect 13856 194 13899 210
tri 13899 194 13915 210 nw
tri 13615 157 13645 187 sw
tri 13721 157 13751 187 se
rect 13751 164 13810 189
tri 13810 164 13840 194 sw
tri 13915 164 13945 194 se
rect 13945 164 14001 329
rect 13751 157 14001 164
rect 13559 153 14001 157
rect 13559 119 13569 153
rect 13603 119 13763 153
rect 13797 119 13860 153
rect 13894 119 13957 153
rect 13991 119 14001 153
rect 13559 103 14001 119
rect 14061 363 14117 379
rect 14061 329 14071 363
rect 14105 329 14117 363
rect 14061 291 14117 329
rect 14147 342 14309 379
tri 14147 326 14163 342 ne
rect 14163 326 14309 342
tri 14223 296 14253 326 ne
rect 14061 257 14071 291
rect 14105 257 14117 291
rect 14061 223 14117 257
rect 14061 189 14071 223
rect 14105 189 14117 223
tri 14147 280 14163 296 se
rect 14163 280 14207 296
tri 14207 280 14223 296 sw
rect 14147 247 14223 280
rect 14147 213 14168 247
rect 14202 213 14223 247
rect 14147 211 14223 213
tri 14147 195 14163 211 ne
rect 14163 195 14207 211
tri 14207 195 14223 211 nw
rect 14253 291 14309 326
rect 14253 257 14265 291
rect 14299 257 14309 291
rect 14253 223 14309 257
rect 14061 165 14117 189
tri 14117 165 14147 195 sw
tri 14223 165 14253 195 se
rect 14253 189 14265 223
rect 14299 189 14309 223
rect 14253 165 14309 189
rect 14061 153 14309 165
rect 14061 119 14071 153
rect 14105 119 14168 153
rect 14202 119 14265 153
rect 14299 119 14309 153
rect 14061 103 14309 119
rect 14521 363 14577 379
rect 14521 329 14531 363
rect 14565 329 14577 363
rect 14521 291 14577 329
rect 14607 363 14877 379
rect 14607 334 14628 363
tri 14607 318 14623 334 ne
rect 14623 329 14628 334
rect 14662 329 14725 363
rect 14759 329 14822 363
rect 14856 329 14877 363
rect 14623 318 14877 329
rect 14907 363 14963 379
rect 14907 329 14919 363
rect 14953 329 14963 363
rect 14521 257 14531 291
rect 14565 257 14577 291
tri 14683 288 14713 318 ne
rect 14713 291 14772 318
rect 14521 223 14577 257
rect 14521 189 14531 223
rect 14565 189 14577 223
rect 14521 157 14577 189
tri 14607 272 14623 288 se
rect 14623 272 14667 288
tri 14667 272 14683 288 sw
rect 14607 238 14683 272
rect 14607 204 14628 238
rect 14662 204 14683 238
rect 14607 203 14683 204
tri 14607 187 14623 203 ne
rect 14623 187 14667 203
tri 14667 187 14683 203 nw
rect 14713 257 14725 291
rect 14759 257 14772 291
tri 14772 288 14802 318 nw
rect 14713 223 14772 257
rect 14713 189 14725 223
rect 14759 189 14772 223
tri 14802 272 14818 288 se
rect 14818 272 14861 288
tri 14861 272 14877 288 sw
rect 14802 244 14877 272
rect 14802 210 14823 244
rect 14857 210 14877 244
tri 14802 194 14818 210 ne
rect 14818 194 14861 210
tri 14861 194 14877 210 nw
tri 14577 157 14607 187 sw
tri 14683 157 14713 187 se
rect 14713 164 14772 189
tri 14772 164 14802 194 sw
tri 14877 164 14907 194 se
rect 14907 164 14963 329
rect 14713 157 14963 164
rect 14521 153 14963 157
rect 14521 119 14531 153
rect 14565 119 14725 153
rect 14759 119 14822 153
rect 14856 119 14919 153
rect 14953 119 14963 153
rect 14521 103 14963 119
rect 15023 363 15079 379
rect 15023 329 15033 363
rect 15067 329 15079 363
rect 15023 291 15079 329
rect 15109 342 15271 379
tri 15109 326 15125 342 ne
rect 15125 326 15271 342
tri 15185 296 15215 326 ne
rect 15023 257 15033 291
rect 15067 257 15079 291
rect 15023 223 15079 257
rect 15023 189 15033 223
rect 15067 189 15079 223
tri 15109 280 15125 296 se
rect 15125 280 15169 296
tri 15169 280 15185 296 sw
rect 15109 247 15185 280
rect 15109 213 15130 247
rect 15164 213 15185 247
rect 15109 211 15185 213
tri 15109 195 15125 211 ne
rect 15125 195 15169 211
tri 15169 195 15185 211 nw
rect 15215 291 15271 326
rect 15215 257 15227 291
rect 15261 257 15271 291
rect 15215 223 15271 257
rect 15023 165 15079 189
tri 15079 165 15109 195 sw
tri 15185 165 15215 195 se
rect 15215 189 15227 223
rect 15261 189 15271 223
rect 15215 165 15271 189
rect 15023 153 15271 165
rect 15023 119 15033 153
rect 15067 119 15130 153
rect 15164 119 15227 153
rect 15261 119 15271 153
rect 15023 103 15271 119
rect 15483 363 15539 379
rect 15483 329 15493 363
rect 15527 329 15539 363
rect 15483 291 15539 329
rect 15569 363 15839 379
rect 15569 334 15590 363
tri 15569 318 15585 334 ne
rect 15585 329 15590 334
rect 15624 329 15687 363
rect 15721 329 15784 363
rect 15818 329 15839 363
rect 15585 318 15839 329
rect 15869 363 15925 379
rect 15869 329 15881 363
rect 15915 329 15925 363
rect 15483 257 15493 291
rect 15527 257 15539 291
tri 15645 288 15675 318 ne
rect 15675 291 15734 318
rect 15483 223 15539 257
rect 15483 189 15493 223
rect 15527 189 15539 223
rect 15483 157 15539 189
tri 15569 272 15585 288 se
rect 15585 272 15629 288
tri 15629 272 15645 288 sw
rect 15569 238 15645 272
rect 15569 204 15590 238
rect 15624 204 15645 238
rect 15569 203 15645 204
tri 15569 187 15585 203 ne
rect 15585 187 15629 203
tri 15629 187 15645 203 nw
rect 15675 257 15687 291
rect 15721 257 15734 291
tri 15734 288 15764 318 nw
rect 15675 223 15734 257
rect 15675 189 15687 223
rect 15721 189 15734 223
tri 15764 272 15780 288 se
rect 15780 272 15823 288
tri 15823 272 15839 288 sw
rect 15764 244 15839 272
rect 15764 210 15785 244
rect 15819 210 15839 244
tri 15764 194 15780 210 ne
rect 15780 194 15823 210
tri 15823 194 15839 210 nw
tri 15539 157 15569 187 sw
tri 15645 157 15675 187 se
rect 15675 164 15734 189
tri 15734 164 15764 194 sw
tri 15839 164 15869 194 se
rect 15869 164 15925 329
rect 15675 157 15925 164
rect 15483 153 15925 157
rect 15483 119 15493 153
rect 15527 119 15687 153
rect 15721 119 15784 153
rect 15818 119 15881 153
rect 15915 119 15925 153
rect 15483 103 15925 119
rect 15985 363 16041 379
rect 15985 329 15995 363
rect 16029 329 16041 363
rect 15985 291 16041 329
rect 16071 342 16233 379
tri 16071 326 16087 342 ne
rect 16087 326 16233 342
tri 16147 296 16177 326 ne
rect 15985 257 15995 291
rect 16029 257 16041 291
rect 15985 223 16041 257
rect 15985 189 15995 223
rect 16029 189 16041 223
tri 16071 280 16087 296 se
rect 16087 280 16131 296
tri 16131 280 16147 296 sw
rect 16071 247 16147 280
rect 16071 213 16092 247
rect 16126 213 16147 247
rect 16071 211 16147 213
tri 16071 195 16087 211 ne
rect 16087 195 16131 211
tri 16131 195 16147 211 nw
rect 16177 291 16233 326
rect 16177 257 16189 291
rect 16223 257 16233 291
rect 16177 223 16233 257
rect 15985 165 16041 189
tri 16041 165 16071 195 sw
tri 16147 165 16177 195 se
rect 16177 189 16189 223
rect 16223 189 16233 223
rect 16177 165 16233 189
rect 15985 153 16233 165
rect 15985 119 15995 153
rect 16029 119 16092 153
rect 16126 119 16189 153
rect 16223 119 16233 153
rect 15985 103 16233 119
rect 16445 363 16501 379
rect 16445 329 16455 363
rect 16489 329 16501 363
rect 16445 291 16501 329
rect 16531 363 16801 379
rect 16531 334 16552 363
tri 16531 318 16547 334 ne
rect 16547 329 16552 334
rect 16586 329 16649 363
rect 16683 329 16746 363
rect 16780 329 16801 363
rect 16547 318 16801 329
rect 16831 363 16887 379
rect 16831 329 16843 363
rect 16877 329 16887 363
rect 16445 257 16455 291
rect 16489 257 16501 291
tri 16607 288 16637 318 ne
rect 16637 291 16696 318
rect 16445 223 16501 257
rect 16445 189 16455 223
rect 16489 189 16501 223
rect 16445 157 16501 189
tri 16531 272 16547 288 se
rect 16547 272 16591 288
tri 16591 272 16607 288 sw
rect 16531 238 16607 272
rect 16531 204 16552 238
rect 16586 204 16607 238
rect 16531 203 16607 204
tri 16531 187 16547 203 ne
rect 16547 187 16591 203
tri 16591 187 16607 203 nw
rect 16637 257 16649 291
rect 16683 257 16696 291
tri 16696 288 16726 318 nw
rect 16637 223 16696 257
rect 16637 189 16649 223
rect 16683 189 16696 223
tri 16726 272 16742 288 se
rect 16742 272 16785 288
tri 16785 272 16801 288 sw
rect 16726 244 16801 272
rect 16726 210 16747 244
rect 16781 210 16801 244
tri 16726 194 16742 210 ne
rect 16742 194 16785 210
tri 16785 194 16801 210 nw
tri 16501 157 16531 187 sw
tri 16607 157 16637 187 se
rect 16637 164 16696 189
tri 16696 164 16726 194 sw
tri 16801 164 16831 194 se
rect 16831 164 16887 329
rect 16637 157 16887 164
rect 16445 153 16887 157
rect 16445 119 16455 153
rect 16489 119 16649 153
rect 16683 119 16746 153
rect 16780 119 16843 153
rect 16877 119 16887 153
rect 16445 103 16887 119
rect 16947 363 17003 379
rect 16947 329 16957 363
rect 16991 329 17003 363
rect 16947 291 17003 329
rect 17033 342 17195 379
tri 17033 326 17049 342 ne
rect 17049 326 17195 342
tri 17109 296 17139 326 ne
rect 16947 257 16957 291
rect 16991 257 17003 291
rect 16947 223 17003 257
rect 16947 189 16957 223
rect 16991 189 17003 223
tri 17033 280 17049 296 se
rect 17049 280 17093 296
tri 17093 280 17109 296 sw
rect 17033 247 17109 280
rect 17033 213 17054 247
rect 17088 213 17109 247
rect 17033 211 17109 213
tri 17033 195 17049 211 ne
rect 17049 195 17093 211
tri 17093 195 17109 211 nw
rect 17139 291 17195 326
rect 17139 257 17151 291
rect 17185 257 17195 291
rect 17139 223 17195 257
rect 16947 165 17003 189
tri 17003 165 17033 195 sw
tri 17109 165 17139 195 se
rect 17139 189 17151 223
rect 17185 189 17195 223
rect 17139 165 17195 189
rect 16947 153 17195 165
rect 16947 119 16957 153
rect 16991 119 17054 153
rect 17088 119 17151 153
rect 17185 119 17195 153
rect 16947 103 17195 119
rect 17428 361 17484 377
rect 17428 327 17438 361
rect 17472 327 17484 361
rect 17428 289 17484 327
rect 17514 361 17678 377
rect 17514 332 17535 361
tri 17514 316 17530 332 ne
rect 17530 327 17535 332
rect 17569 327 17632 361
rect 17666 327 17678 361
rect 17530 316 17678 327
rect 17708 361 17868 377
rect 17708 340 17826 361
tri 17708 324 17724 340 ne
rect 17724 327 17826 340
rect 17860 327 17868 361
rect 17724 324 17868 327
rect 17428 255 17438 289
rect 17472 255 17484 289
tri 17590 286 17620 316 ne
rect 17620 289 17678 316
tri 17784 294 17814 324 ne
rect 17428 221 17484 255
rect 17428 187 17438 221
rect 17472 187 17484 221
rect 17428 155 17484 187
tri 17514 270 17530 286 se
rect 17530 270 17574 286
tri 17574 270 17590 286 sw
rect 17514 236 17590 270
rect 17514 202 17535 236
rect 17569 202 17590 236
rect 17514 201 17590 202
tri 17514 185 17530 201 ne
rect 17530 185 17574 201
tri 17574 185 17590 201 nw
rect 17620 255 17632 289
rect 17666 255 17678 289
rect 17620 221 17678 255
rect 17620 187 17632 221
rect 17666 187 17678 221
tri 17708 278 17724 294 se
rect 17724 278 17768 294
tri 17768 278 17784 294 sw
rect 17708 245 17784 278
rect 17708 211 17728 245
rect 17762 211 17784 245
rect 17708 209 17784 211
tri 17708 193 17724 209 ne
rect 17724 193 17768 209
tri 17768 193 17784 209 nw
rect 17814 289 17868 324
rect 17814 255 17826 289
rect 17860 255 17868 289
rect 17814 221 17868 255
tri 17484 155 17514 185 sw
tri 17590 155 17620 185 se
rect 17620 163 17678 187
tri 17678 163 17708 193 sw
tri 17784 163 17814 193 se
rect 17814 187 17826 221
rect 17860 187 17868 221
rect 17814 163 17868 187
rect 17620 155 17868 163
rect 17428 151 17868 155
rect 17428 117 17438 151
rect 17472 117 17632 151
rect 17666 117 17728 151
rect 17762 117 17826 151
rect 17860 117 17868 151
rect 17428 101 17868 117
rect 18094 361 18150 377
rect 18094 327 18104 361
rect 18138 327 18150 361
rect 18094 289 18150 327
rect 18180 361 18450 377
rect 18180 332 18201 361
tri 18180 316 18196 332 ne
rect 18196 327 18201 332
rect 18235 327 18298 361
rect 18332 340 18450 361
rect 18332 327 18434 340
rect 18196 324 18434 327
tri 18434 324 18450 340 nw
rect 18480 361 18536 377
rect 18480 327 18492 361
rect 18526 327 18536 361
rect 18196 316 18344 324
rect 18094 255 18104 289
rect 18138 255 18150 289
tri 18256 286 18286 316 ne
rect 18286 289 18344 316
tri 18344 294 18374 324 nw
rect 18094 221 18150 255
rect 18094 187 18104 221
rect 18138 187 18150 221
rect 18094 155 18150 187
tri 18180 270 18196 286 se
rect 18196 270 18240 286
tri 18240 270 18256 286 sw
rect 18180 236 18256 270
rect 18180 202 18201 236
rect 18235 202 18256 236
rect 18180 201 18256 202
tri 18180 185 18196 201 ne
rect 18196 185 18240 201
tri 18240 185 18256 201 nw
rect 18286 255 18298 289
rect 18332 255 18344 289
rect 18286 221 18344 255
rect 18286 187 18298 221
rect 18332 187 18344 221
tri 18374 278 18390 294 se
rect 18390 278 18434 294
tri 18434 278 18450 294 sw
rect 18374 245 18450 278
rect 18374 211 18395 245
rect 18429 211 18450 245
rect 18374 209 18450 211
tri 18374 193 18390 209 ne
rect 18390 193 18434 209
tri 18434 193 18450 209 nw
rect 18480 289 18536 327
rect 18480 255 18492 289
rect 18526 255 18536 289
rect 18480 221 18536 255
tri 18150 155 18180 185 sw
tri 18256 155 18286 185 se
rect 18286 163 18344 187
tri 18344 163 18374 193 sw
tri 18450 163 18480 193 se
rect 18480 187 18492 221
rect 18526 187 18536 221
rect 18480 163 18536 187
rect 18286 155 18536 163
rect 18094 151 18536 155
rect 18094 117 18104 151
rect 18138 117 18298 151
rect 18332 117 18395 151
rect 18429 117 18492 151
rect 18526 117 18536 151
rect 18094 101 18536 117
rect 18760 361 18816 377
rect 18760 327 18770 361
rect 18804 327 18816 361
rect 18760 289 18816 327
rect 18846 361 19010 377
rect 18846 332 18867 361
tri 18846 316 18862 332 ne
rect 18862 327 18867 332
rect 18901 327 18964 361
rect 18998 327 19010 361
rect 18862 316 19010 327
rect 19040 340 19202 377
tri 19040 324 19056 340 ne
rect 19056 324 19202 340
rect 18760 255 18770 289
rect 18804 255 18816 289
tri 18922 286 18952 316 ne
rect 18952 289 19010 316
tri 19116 294 19146 324 ne
rect 18760 221 18816 255
rect 18760 187 18770 221
rect 18804 187 18816 221
rect 18760 155 18816 187
tri 18846 270 18862 286 se
rect 18862 270 18906 286
tri 18906 270 18922 286 sw
rect 18846 236 18922 270
rect 18846 202 18867 236
rect 18901 202 18922 236
rect 18846 201 18922 202
tri 18846 185 18862 201 ne
rect 18862 185 18906 201
tri 18906 185 18922 201 nw
rect 18952 255 18964 289
rect 18998 255 19010 289
tri 19041 279 19056 294 se
rect 19056 279 19100 294
tri 19100 279 19115 294 sw
rect 19146 289 19202 324
rect 18952 221 19010 255
rect 18952 187 18964 221
rect 18998 187 19010 221
rect 19040 245 19116 279
rect 19040 211 19061 245
rect 19095 211 19116 245
rect 19040 209 19116 211
tri 19040 193 19056 209 ne
rect 19056 193 19100 209
tri 19100 193 19116 209 nw
rect 19146 255 19158 289
rect 19192 255 19202 289
rect 19146 221 19202 255
tri 18816 155 18846 185 sw
tri 18922 155 18952 185 se
rect 18952 163 19010 187
tri 19010 163 19040 193 sw
tri 19116 163 19146 193 se
rect 19146 187 19158 221
rect 19192 187 19202 221
rect 19146 163 19202 187
rect 18952 155 19202 163
rect 18760 151 19202 155
rect 18760 117 18770 151
rect 18804 117 18964 151
rect 18998 117 19061 151
rect 19095 117 19158 151
rect 19192 117 19202 151
rect 18760 101 19202 117
<< pdiff >>
rect 191 1412 247 1450
rect 191 1378 201 1412
rect 235 1378 247 1412
rect 191 1344 247 1378
rect 191 1310 201 1344
rect 235 1310 247 1344
rect 191 1276 247 1310
rect 191 1242 201 1276
rect 235 1242 247 1276
rect 191 1208 247 1242
rect 191 1174 201 1208
rect 235 1174 247 1208
rect 191 1139 247 1174
rect 191 1105 201 1139
rect 235 1105 247 1139
rect 191 1050 247 1105
rect 277 1412 335 1450
rect 277 1378 289 1412
rect 323 1378 335 1412
rect 277 1344 335 1378
rect 277 1310 289 1344
rect 323 1310 335 1344
rect 277 1276 335 1310
rect 277 1242 289 1276
rect 323 1242 335 1276
rect 277 1208 335 1242
rect 277 1174 289 1208
rect 323 1174 335 1208
rect 277 1139 335 1174
rect 277 1105 289 1139
rect 323 1105 335 1139
rect 277 1050 335 1105
rect 365 1412 423 1450
rect 365 1378 377 1412
rect 411 1378 423 1412
rect 365 1344 423 1378
rect 365 1310 377 1344
rect 411 1310 423 1344
rect 365 1276 423 1310
rect 365 1242 377 1276
rect 411 1242 423 1276
rect 365 1208 423 1242
rect 365 1174 377 1208
rect 411 1174 423 1208
rect 365 1050 423 1174
rect 453 1412 511 1450
rect 453 1378 465 1412
rect 499 1378 511 1412
rect 453 1344 511 1378
rect 453 1310 465 1344
rect 499 1310 511 1344
rect 453 1276 511 1310
rect 453 1242 465 1276
rect 499 1242 511 1276
rect 453 1208 511 1242
rect 453 1174 465 1208
rect 499 1174 511 1208
rect 453 1139 511 1174
rect 453 1105 465 1139
rect 499 1105 511 1139
rect 453 1050 511 1105
rect 541 1412 599 1450
rect 541 1378 553 1412
rect 587 1378 599 1412
rect 541 1344 599 1378
rect 541 1310 553 1344
rect 587 1310 599 1344
rect 541 1276 599 1310
rect 541 1242 553 1276
rect 587 1242 599 1276
rect 541 1208 599 1242
rect 541 1174 553 1208
rect 587 1174 599 1208
rect 541 1050 599 1174
rect 629 1412 687 1450
rect 629 1378 641 1412
rect 675 1378 687 1412
rect 629 1344 687 1378
rect 629 1310 641 1344
rect 675 1310 687 1344
rect 629 1276 687 1310
rect 629 1242 641 1276
rect 675 1242 687 1276
rect 629 1208 687 1242
rect 629 1174 641 1208
rect 675 1174 687 1208
rect 629 1139 687 1174
rect 629 1105 641 1139
rect 675 1105 687 1139
rect 629 1050 687 1105
rect 717 1412 771 1450
rect 717 1378 729 1412
rect 763 1378 771 1412
rect 717 1344 771 1378
rect 717 1310 729 1344
rect 763 1310 771 1344
rect 717 1276 771 1310
rect 717 1242 729 1276
rect 763 1242 771 1276
rect 717 1208 771 1242
rect 717 1174 729 1208
rect 763 1174 771 1208
rect 717 1050 771 1174
rect 1153 1412 1209 1450
rect 1153 1378 1163 1412
rect 1197 1378 1209 1412
rect 1153 1344 1209 1378
rect 1153 1310 1163 1344
rect 1197 1310 1209 1344
rect 1153 1276 1209 1310
rect 1153 1242 1163 1276
rect 1197 1242 1209 1276
rect 1153 1208 1209 1242
rect 1153 1174 1163 1208
rect 1197 1174 1209 1208
rect 1153 1139 1209 1174
rect 1153 1105 1163 1139
rect 1197 1105 1209 1139
rect 1153 1050 1209 1105
rect 1239 1412 1297 1450
rect 1239 1378 1251 1412
rect 1285 1378 1297 1412
rect 1239 1344 1297 1378
rect 1239 1310 1251 1344
rect 1285 1310 1297 1344
rect 1239 1276 1297 1310
rect 1239 1242 1251 1276
rect 1285 1242 1297 1276
rect 1239 1208 1297 1242
rect 1239 1174 1251 1208
rect 1285 1174 1297 1208
rect 1239 1139 1297 1174
rect 1239 1105 1251 1139
rect 1285 1105 1297 1139
rect 1239 1050 1297 1105
rect 1327 1412 1385 1450
rect 1327 1378 1339 1412
rect 1373 1378 1385 1412
rect 1327 1344 1385 1378
rect 1327 1310 1339 1344
rect 1373 1310 1385 1344
rect 1327 1276 1385 1310
rect 1327 1242 1339 1276
rect 1373 1242 1385 1276
rect 1327 1208 1385 1242
rect 1327 1174 1339 1208
rect 1373 1174 1385 1208
rect 1327 1050 1385 1174
rect 1415 1412 1473 1450
rect 1415 1378 1427 1412
rect 1461 1378 1473 1412
rect 1415 1344 1473 1378
rect 1415 1310 1427 1344
rect 1461 1310 1473 1344
rect 1415 1276 1473 1310
rect 1415 1242 1427 1276
rect 1461 1242 1473 1276
rect 1415 1208 1473 1242
rect 1415 1174 1427 1208
rect 1461 1174 1473 1208
rect 1415 1139 1473 1174
rect 1415 1105 1427 1139
rect 1461 1105 1473 1139
rect 1415 1050 1473 1105
rect 1503 1412 1561 1450
rect 1503 1378 1515 1412
rect 1549 1378 1561 1412
rect 1503 1344 1561 1378
rect 1503 1310 1515 1344
rect 1549 1310 1561 1344
rect 1503 1276 1561 1310
rect 1503 1242 1515 1276
rect 1549 1242 1561 1276
rect 1503 1208 1561 1242
rect 1503 1174 1515 1208
rect 1549 1174 1561 1208
rect 1503 1050 1561 1174
rect 1591 1412 1649 1450
rect 1591 1378 1603 1412
rect 1637 1378 1649 1412
rect 1591 1344 1649 1378
rect 1591 1310 1603 1344
rect 1637 1310 1649 1344
rect 1591 1276 1649 1310
rect 1591 1242 1603 1276
rect 1637 1242 1649 1276
rect 1591 1208 1649 1242
rect 1591 1174 1603 1208
rect 1637 1174 1649 1208
rect 1591 1139 1649 1174
rect 1591 1105 1603 1139
rect 1637 1105 1649 1139
rect 1591 1050 1649 1105
rect 1679 1412 1733 1450
rect 1679 1378 1691 1412
rect 1725 1378 1733 1412
rect 1679 1344 1733 1378
rect 1679 1310 1691 1344
rect 1725 1310 1733 1344
rect 1679 1276 1733 1310
rect 1679 1242 1691 1276
rect 1725 1242 1733 1276
rect 1679 1208 1733 1242
rect 1679 1174 1691 1208
rect 1725 1174 1733 1208
rect 1679 1050 1733 1174
rect 2115 1412 2171 1450
rect 2115 1378 2125 1412
rect 2159 1378 2171 1412
rect 2115 1344 2171 1378
rect 2115 1310 2125 1344
rect 2159 1310 2171 1344
rect 2115 1276 2171 1310
rect 2115 1242 2125 1276
rect 2159 1242 2171 1276
rect 2115 1208 2171 1242
rect 2115 1174 2125 1208
rect 2159 1174 2171 1208
rect 2115 1139 2171 1174
rect 2115 1105 2125 1139
rect 2159 1105 2171 1139
rect 2115 1050 2171 1105
rect 2201 1412 2259 1450
rect 2201 1378 2213 1412
rect 2247 1378 2259 1412
rect 2201 1344 2259 1378
rect 2201 1310 2213 1344
rect 2247 1310 2259 1344
rect 2201 1276 2259 1310
rect 2201 1242 2213 1276
rect 2247 1242 2259 1276
rect 2201 1208 2259 1242
rect 2201 1174 2213 1208
rect 2247 1174 2259 1208
rect 2201 1139 2259 1174
rect 2201 1105 2213 1139
rect 2247 1105 2259 1139
rect 2201 1050 2259 1105
rect 2289 1412 2347 1450
rect 2289 1378 2301 1412
rect 2335 1378 2347 1412
rect 2289 1344 2347 1378
rect 2289 1310 2301 1344
rect 2335 1310 2347 1344
rect 2289 1276 2347 1310
rect 2289 1242 2301 1276
rect 2335 1242 2347 1276
rect 2289 1208 2347 1242
rect 2289 1174 2301 1208
rect 2335 1174 2347 1208
rect 2289 1050 2347 1174
rect 2377 1412 2435 1450
rect 2377 1378 2389 1412
rect 2423 1378 2435 1412
rect 2377 1344 2435 1378
rect 2377 1310 2389 1344
rect 2423 1310 2435 1344
rect 2377 1276 2435 1310
rect 2377 1242 2389 1276
rect 2423 1242 2435 1276
rect 2377 1208 2435 1242
rect 2377 1174 2389 1208
rect 2423 1174 2435 1208
rect 2377 1139 2435 1174
rect 2377 1105 2389 1139
rect 2423 1105 2435 1139
rect 2377 1050 2435 1105
rect 2465 1412 2523 1450
rect 2465 1378 2477 1412
rect 2511 1378 2523 1412
rect 2465 1344 2523 1378
rect 2465 1310 2477 1344
rect 2511 1310 2523 1344
rect 2465 1276 2523 1310
rect 2465 1242 2477 1276
rect 2511 1242 2523 1276
rect 2465 1208 2523 1242
rect 2465 1174 2477 1208
rect 2511 1174 2523 1208
rect 2465 1050 2523 1174
rect 2553 1412 2611 1450
rect 2553 1378 2565 1412
rect 2599 1378 2611 1412
rect 2553 1344 2611 1378
rect 2553 1310 2565 1344
rect 2599 1310 2611 1344
rect 2553 1276 2611 1310
rect 2553 1242 2565 1276
rect 2599 1242 2611 1276
rect 2553 1208 2611 1242
rect 2553 1174 2565 1208
rect 2599 1174 2611 1208
rect 2553 1139 2611 1174
rect 2553 1105 2565 1139
rect 2599 1105 2611 1139
rect 2553 1050 2611 1105
rect 2641 1412 2695 1450
rect 2641 1378 2653 1412
rect 2687 1378 2695 1412
rect 2641 1344 2695 1378
rect 2641 1310 2653 1344
rect 2687 1310 2695 1344
rect 2641 1276 2695 1310
rect 2641 1242 2653 1276
rect 2687 1242 2695 1276
rect 2641 1208 2695 1242
rect 2641 1174 2653 1208
rect 2687 1174 2695 1208
rect 2641 1050 2695 1174
rect 3077 1412 3133 1450
rect 3077 1378 3087 1412
rect 3121 1378 3133 1412
rect 3077 1344 3133 1378
rect 3077 1310 3087 1344
rect 3121 1310 3133 1344
rect 3077 1276 3133 1310
rect 3077 1242 3087 1276
rect 3121 1242 3133 1276
rect 3077 1208 3133 1242
rect 3077 1174 3087 1208
rect 3121 1174 3133 1208
rect 3077 1139 3133 1174
rect 3077 1105 3087 1139
rect 3121 1105 3133 1139
rect 3077 1050 3133 1105
rect 3163 1412 3221 1450
rect 3163 1378 3175 1412
rect 3209 1378 3221 1412
rect 3163 1344 3221 1378
rect 3163 1310 3175 1344
rect 3209 1310 3221 1344
rect 3163 1276 3221 1310
rect 3163 1242 3175 1276
rect 3209 1242 3221 1276
rect 3163 1208 3221 1242
rect 3163 1174 3175 1208
rect 3209 1174 3221 1208
rect 3163 1139 3221 1174
rect 3163 1105 3175 1139
rect 3209 1105 3221 1139
rect 3163 1050 3221 1105
rect 3251 1412 3309 1450
rect 3251 1378 3263 1412
rect 3297 1378 3309 1412
rect 3251 1344 3309 1378
rect 3251 1310 3263 1344
rect 3297 1310 3309 1344
rect 3251 1276 3309 1310
rect 3251 1242 3263 1276
rect 3297 1242 3309 1276
rect 3251 1208 3309 1242
rect 3251 1174 3263 1208
rect 3297 1174 3309 1208
rect 3251 1050 3309 1174
rect 3339 1412 3397 1450
rect 3339 1378 3351 1412
rect 3385 1378 3397 1412
rect 3339 1344 3397 1378
rect 3339 1310 3351 1344
rect 3385 1310 3397 1344
rect 3339 1276 3397 1310
rect 3339 1242 3351 1276
rect 3385 1242 3397 1276
rect 3339 1208 3397 1242
rect 3339 1174 3351 1208
rect 3385 1174 3397 1208
rect 3339 1139 3397 1174
rect 3339 1105 3351 1139
rect 3385 1105 3397 1139
rect 3339 1050 3397 1105
rect 3427 1412 3485 1450
rect 3427 1378 3439 1412
rect 3473 1378 3485 1412
rect 3427 1344 3485 1378
rect 3427 1310 3439 1344
rect 3473 1310 3485 1344
rect 3427 1276 3485 1310
rect 3427 1242 3439 1276
rect 3473 1242 3485 1276
rect 3427 1208 3485 1242
rect 3427 1174 3439 1208
rect 3473 1174 3485 1208
rect 3427 1050 3485 1174
rect 3515 1412 3573 1450
rect 3515 1378 3527 1412
rect 3561 1378 3573 1412
rect 3515 1344 3573 1378
rect 3515 1310 3527 1344
rect 3561 1310 3573 1344
rect 3515 1276 3573 1310
rect 3515 1242 3527 1276
rect 3561 1242 3573 1276
rect 3515 1208 3573 1242
rect 3515 1174 3527 1208
rect 3561 1174 3573 1208
rect 3515 1139 3573 1174
rect 3515 1105 3527 1139
rect 3561 1105 3573 1139
rect 3515 1050 3573 1105
rect 3603 1412 3657 1450
rect 3603 1378 3615 1412
rect 3649 1378 3657 1412
rect 3603 1344 3657 1378
rect 3603 1310 3615 1344
rect 3649 1310 3657 1344
rect 3603 1276 3657 1310
rect 3603 1242 3615 1276
rect 3649 1242 3657 1276
rect 3603 1208 3657 1242
rect 3603 1174 3615 1208
rect 3649 1174 3657 1208
rect 3603 1050 3657 1174
rect 4039 1412 4095 1450
rect 4039 1378 4049 1412
rect 4083 1378 4095 1412
rect 4039 1344 4095 1378
rect 4039 1310 4049 1344
rect 4083 1310 4095 1344
rect 4039 1276 4095 1310
rect 4039 1242 4049 1276
rect 4083 1242 4095 1276
rect 4039 1208 4095 1242
rect 4039 1174 4049 1208
rect 4083 1174 4095 1208
rect 4039 1139 4095 1174
rect 4039 1105 4049 1139
rect 4083 1105 4095 1139
rect 4039 1050 4095 1105
rect 4125 1412 4183 1450
rect 4125 1378 4137 1412
rect 4171 1378 4183 1412
rect 4125 1344 4183 1378
rect 4125 1310 4137 1344
rect 4171 1310 4183 1344
rect 4125 1276 4183 1310
rect 4125 1242 4137 1276
rect 4171 1242 4183 1276
rect 4125 1208 4183 1242
rect 4125 1174 4137 1208
rect 4171 1174 4183 1208
rect 4125 1139 4183 1174
rect 4125 1105 4137 1139
rect 4171 1105 4183 1139
rect 4125 1050 4183 1105
rect 4213 1412 4271 1450
rect 4213 1378 4225 1412
rect 4259 1378 4271 1412
rect 4213 1344 4271 1378
rect 4213 1310 4225 1344
rect 4259 1310 4271 1344
rect 4213 1276 4271 1310
rect 4213 1242 4225 1276
rect 4259 1242 4271 1276
rect 4213 1208 4271 1242
rect 4213 1174 4225 1208
rect 4259 1174 4271 1208
rect 4213 1050 4271 1174
rect 4301 1412 4359 1450
rect 4301 1378 4313 1412
rect 4347 1378 4359 1412
rect 4301 1344 4359 1378
rect 4301 1310 4313 1344
rect 4347 1310 4359 1344
rect 4301 1276 4359 1310
rect 4301 1242 4313 1276
rect 4347 1242 4359 1276
rect 4301 1208 4359 1242
rect 4301 1174 4313 1208
rect 4347 1174 4359 1208
rect 4301 1139 4359 1174
rect 4301 1105 4313 1139
rect 4347 1105 4359 1139
rect 4301 1050 4359 1105
rect 4389 1412 4447 1450
rect 4389 1378 4401 1412
rect 4435 1378 4447 1412
rect 4389 1344 4447 1378
rect 4389 1310 4401 1344
rect 4435 1310 4447 1344
rect 4389 1276 4447 1310
rect 4389 1242 4401 1276
rect 4435 1242 4447 1276
rect 4389 1208 4447 1242
rect 4389 1174 4401 1208
rect 4435 1174 4447 1208
rect 4389 1050 4447 1174
rect 4477 1412 4535 1450
rect 4477 1378 4489 1412
rect 4523 1378 4535 1412
rect 4477 1344 4535 1378
rect 4477 1310 4489 1344
rect 4523 1310 4535 1344
rect 4477 1276 4535 1310
rect 4477 1242 4489 1276
rect 4523 1242 4535 1276
rect 4477 1208 4535 1242
rect 4477 1174 4489 1208
rect 4523 1174 4535 1208
rect 4477 1139 4535 1174
rect 4477 1105 4489 1139
rect 4523 1105 4535 1139
rect 4477 1050 4535 1105
rect 4565 1412 4619 1450
rect 4565 1378 4577 1412
rect 4611 1378 4619 1412
rect 4565 1344 4619 1378
rect 4565 1310 4577 1344
rect 4611 1310 4619 1344
rect 4565 1276 4619 1310
rect 4565 1242 4577 1276
rect 4611 1242 4619 1276
rect 4565 1208 4619 1242
rect 4565 1174 4577 1208
rect 4611 1174 4619 1208
rect 4565 1050 4619 1174
rect 5001 1412 5057 1450
rect 5001 1378 5011 1412
rect 5045 1378 5057 1412
rect 5001 1344 5057 1378
rect 5001 1310 5011 1344
rect 5045 1310 5057 1344
rect 5001 1276 5057 1310
rect 5001 1242 5011 1276
rect 5045 1242 5057 1276
rect 5001 1208 5057 1242
rect 5001 1174 5011 1208
rect 5045 1174 5057 1208
rect 5001 1139 5057 1174
rect 5001 1105 5011 1139
rect 5045 1105 5057 1139
rect 5001 1050 5057 1105
rect 5087 1412 5145 1450
rect 5087 1378 5099 1412
rect 5133 1378 5145 1412
rect 5087 1344 5145 1378
rect 5087 1310 5099 1344
rect 5133 1310 5145 1344
rect 5087 1276 5145 1310
rect 5087 1242 5099 1276
rect 5133 1242 5145 1276
rect 5087 1208 5145 1242
rect 5087 1174 5099 1208
rect 5133 1174 5145 1208
rect 5087 1139 5145 1174
rect 5087 1105 5099 1139
rect 5133 1105 5145 1139
rect 5087 1050 5145 1105
rect 5175 1412 5233 1450
rect 5175 1378 5187 1412
rect 5221 1378 5233 1412
rect 5175 1344 5233 1378
rect 5175 1310 5187 1344
rect 5221 1310 5233 1344
rect 5175 1276 5233 1310
rect 5175 1242 5187 1276
rect 5221 1242 5233 1276
rect 5175 1208 5233 1242
rect 5175 1174 5187 1208
rect 5221 1174 5233 1208
rect 5175 1050 5233 1174
rect 5263 1412 5321 1450
rect 5263 1378 5275 1412
rect 5309 1378 5321 1412
rect 5263 1344 5321 1378
rect 5263 1310 5275 1344
rect 5309 1310 5321 1344
rect 5263 1276 5321 1310
rect 5263 1242 5275 1276
rect 5309 1242 5321 1276
rect 5263 1208 5321 1242
rect 5263 1174 5275 1208
rect 5309 1174 5321 1208
rect 5263 1139 5321 1174
rect 5263 1105 5275 1139
rect 5309 1105 5321 1139
rect 5263 1050 5321 1105
rect 5351 1412 5409 1450
rect 5351 1378 5363 1412
rect 5397 1378 5409 1412
rect 5351 1344 5409 1378
rect 5351 1310 5363 1344
rect 5397 1310 5409 1344
rect 5351 1276 5409 1310
rect 5351 1242 5363 1276
rect 5397 1242 5409 1276
rect 5351 1208 5409 1242
rect 5351 1174 5363 1208
rect 5397 1174 5409 1208
rect 5351 1050 5409 1174
rect 5439 1412 5497 1450
rect 5439 1378 5451 1412
rect 5485 1378 5497 1412
rect 5439 1344 5497 1378
rect 5439 1310 5451 1344
rect 5485 1310 5497 1344
rect 5439 1276 5497 1310
rect 5439 1242 5451 1276
rect 5485 1242 5497 1276
rect 5439 1208 5497 1242
rect 5439 1174 5451 1208
rect 5485 1174 5497 1208
rect 5439 1139 5497 1174
rect 5439 1105 5451 1139
rect 5485 1105 5497 1139
rect 5439 1050 5497 1105
rect 5527 1412 5581 1450
rect 5527 1378 5539 1412
rect 5573 1378 5581 1412
rect 5527 1344 5581 1378
rect 5527 1310 5539 1344
rect 5573 1310 5581 1344
rect 5527 1276 5581 1310
rect 5527 1242 5539 1276
rect 5573 1242 5581 1276
rect 5527 1208 5581 1242
rect 5527 1174 5539 1208
rect 5573 1174 5581 1208
rect 5527 1050 5581 1174
rect 5963 1412 6019 1450
rect 5963 1378 5973 1412
rect 6007 1378 6019 1412
rect 5963 1344 6019 1378
rect 5963 1310 5973 1344
rect 6007 1310 6019 1344
rect 5963 1276 6019 1310
rect 5963 1242 5973 1276
rect 6007 1242 6019 1276
rect 5963 1208 6019 1242
rect 5963 1174 5973 1208
rect 6007 1174 6019 1208
rect 5963 1139 6019 1174
rect 5963 1105 5973 1139
rect 6007 1105 6019 1139
rect 5963 1050 6019 1105
rect 6049 1412 6107 1450
rect 6049 1378 6061 1412
rect 6095 1378 6107 1412
rect 6049 1344 6107 1378
rect 6049 1310 6061 1344
rect 6095 1310 6107 1344
rect 6049 1276 6107 1310
rect 6049 1242 6061 1276
rect 6095 1242 6107 1276
rect 6049 1208 6107 1242
rect 6049 1174 6061 1208
rect 6095 1174 6107 1208
rect 6049 1139 6107 1174
rect 6049 1105 6061 1139
rect 6095 1105 6107 1139
rect 6049 1050 6107 1105
rect 6137 1412 6195 1450
rect 6137 1378 6149 1412
rect 6183 1378 6195 1412
rect 6137 1344 6195 1378
rect 6137 1310 6149 1344
rect 6183 1310 6195 1344
rect 6137 1276 6195 1310
rect 6137 1242 6149 1276
rect 6183 1242 6195 1276
rect 6137 1208 6195 1242
rect 6137 1174 6149 1208
rect 6183 1174 6195 1208
rect 6137 1050 6195 1174
rect 6225 1412 6283 1450
rect 6225 1378 6237 1412
rect 6271 1378 6283 1412
rect 6225 1344 6283 1378
rect 6225 1310 6237 1344
rect 6271 1310 6283 1344
rect 6225 1276 6283 1310
rect 6225 1242 6237 1276
rect 6271 1242 6283 1276
rect 6225 1208 6283 1242
rect 6225 1174 6237 1208
rect 6271 1174 6283 1208
rect 6225 1139 6283 1174
rect 6225 1105 6237 1139
rect 6271 1105 6283 1139
rect 6225 1050 6283 1105
rect 6313 1412 6371 1450
rect 6313 1378 6325 1412
rect 6359 1378 6371 1412
rect 6313 1344 6371 1378
rect 6313 1310 6325 1344
rect 6359 1310 6371 1344
rect 6313 1276 6371 1310
rect 6313 1242 6325 1276
rect 6359 1242 6371 1276
rect 6313 1208 6371 1242
rect 6313 1174 6325 1208
rect 6359 1174 6371 1208
rect 6313 1050 6371 1174
rect 6401 1412 6459 1450
rect 6401 1378 6413 1412
rect 6447 1378 6459 1412
rect 6401 1344 6459 1378
rect 6401 1310 6413 1344
rect 6447 1310 6459 1344
rect 6401 1276 6459 1310
rect 6401 1242 6413 1276
rect 6447 1242 6459 1276
rect 6401 1208 6459 1242
rect 6401 1174 6413 1208
rect 6447 1174 6459 1208
rect 6401 1139 6459 1174
rect 6401 1105 6413 1139
rect 6447 1105 6459 1139
rect 6401 1050 6459 1105
rect 6489 1412 6543 1450
rect 6489 1378 6501 1412
rect 6535 1378 6543 1412
rect 6489 1344 6543 1378
rect 6489 1310 6501 1344
rect 6535 1310 6543 1344
rect 6489 1276 6543 1310
rect 6489 1242 6501 1276
rect 6535 1242 6543 1276
rect 6489 1208 6543 1242
rect 6489 1174 6501 1208
rect 6535 1174 6543 1208
rect 6489 1050 6543 1174
rect 6925 1412 6981 1450
rect 6925 1378 6935 1412
rect 6969 1378 6981 1412
rect 6925 1344 6981 1378
rect 6925 1310 6935 1344
rect 6969 1310 6981 1344
rect 6925 1276 6981 1310
rect 6925 1242 6935 1276
rect 6969 1242 6981 1276
rect 6925 1208 6981 1242
rect 6925 1174 6935 1208
rect 6969 1174 6981 1208
rect 6925 1139 6981 1174
rect 6925 1105 6935 1139
rect 6969 1105 6981 1139
rect 6925 1050 6981 1105
rect 7011 1412 7069 1450
rect 7011 1378 7023 1412
rect 7057 1378 7069 1412
rect 7011 1344 7069 1378
rect 7011 1310 7023 1344
rect 7057 1310 7069 1344
rect 7011 1276 7069 1310
rect 7011 1242 7023 1276
rect 7057 1242 7069 1276
rect 7011 1208 7069 1242
rect 7011 1174 7023 1208
rect 7057 1174 7069 1208
rect 7011 1139 7069 1174
rect 7011 1105 7023 1139
rect 7057 1105 7069 1139
rect 7011 1050 7069 1105
rect 7099 1412 7157 1450
rect 7099 1378 7111 1412
rect 7145 1378 7157 1412
rect 7099 1344 7157 1378
rect 7099 1310 7111 1344
rect 7145 1310 7157 1344
rect 7099 1276 7157 1310
rect 7099 1242 7111 1276
rect 7145 1242 7157 1276
rect 7099 1208 7157 1242
rect 7099 1174 7111 1208
rect 7145 1174 7157 1208
rect 7099 1050 7157 1174
rect 7187 1412 7245 1450
rect 7187 1378 7199 1412
rect 7233 1378 7245 1412
rect 7187 1344 7245 1378
rect 7187 1310 7199 1344
rect 7233 1310 7245 1344
rect 7187 1276 7245 1310
rect 7187 1242 7199 1276
rect 7233 1242 7245 1276
rect 7187 1208 7245 1242
rect 7187 1174 7199 1208
rect 7233 1174 7245 1208
rect 7187 1139 7245 1174
rect 7187 1105 7199 1139
rect 7233 1105 7245 1139
rect 7187 1050 7245 1105
rect 7275 1412 7333 1450
rect 7275 1378 7287 1412
rect 7321 1378 7333 1412
rect 7275 1344 7333 1378
rect 7275 1310 7287 1344
rect 7321 1310 7333 1344
rect 7275 1276 7333 1310
rect 7275 1242 7287 1276
rect 7321 1242 7333 1276
rect 7275 1208 7333 1242
rect 7275 1174 7287 1208
rect 7321 1174 7333 1208
rect 7275 1050 7333 1174
rect 7363 1412 7421 1450
rect 7363 1378 7375 1412
rect 7409 1378 7421 1412
rect 7363 1344 7421 1378
rect 7363 1310 7375 1344
rect 7409 1310 7421 1344
rect 7363 1276 7421 1310
rect 7363 1242 7375 1276
rect 7409 1242 7421 1276
rect 7363 1208 7421 1242
rect 7363 1174 7375 1208
rect 7409 1174 7421 1208
rect 7363 1139 7421 1174
rect 7363 1105 7375 1139
rect 7409 1105 7421 1139
rect 7363 1050 7421 1105
rect 7451 1412 7505 1450
rect 7451 1378 7463 1412
rect 7497 1378 7505 1412
rect 7451 1344 7505 1378
rect 7451 1310 7463 1344
rect 7497 1310 7505 1344
rect 7451 1276 7505 1310
rect 7451 1242 7463 1276
rect 7497 1242 7505 1276
rect 7451 1208 7505 1242
rect 7451 1174 7463 1208
rect 7497 1174 7505 1208
rect 7451 1050 7505 1174
rect 7887 1412 7943 1450
rect 7887 1378 7897 1412
rect 7931 1378 7943 1412
rect 7887 1344 7943 1378
rect 7887 1310 7897 1344
rect 7931 1310 7943 1344
rect 7887 1276 7943 1310
rect 7887 1242 7897 1276
rect 7931 1242 7943 1276
rect 7887 1208 7943 1242
rect 7887 1174 7897 1208
rect 7931 1174 7943 1208
rect 7887 1139 7943 1174
rect 7887 1105 7897 1139
rect 7931 1105 7943 1139
rect 7887 1050 7943 1105
rect 7973 1412 8031 1450
rect 7973 1378 7985 1412
rect 8019 1378 8031 1412
rect 7973 1344 8031 1378
rect 7973 1310 7985 1344
rect 8019 1310 8031 1344
rect 7973 1276 8031 1310
rect 7973 1242 7985 1276
rect 8019 1242 8031 1276
rect 7973 1208 8031 1242
rect 7973 1174 7985 1208
rect 8019 1174 8031 1208
rect 7973 1139 8031 1174
rect 7973 1105 7985 1139
rect 8019 1105 8031 1139
rect 7973 1050 8031 1105
rect 8061 1412 8119 1450
rect 8061 1378 8073 1412
rect 8107 1378 8119 1412
rect 8061 1344 8119 1378
rect 8061 1310 8073 1344
rect 8107 1310 8119 1344
rect 8061 1276 8119 1310
rect 8061 1242 8073 1276
rect 8107 1242 8119 1276
rect 8061 1208 8119 1242
rect 8061 1174 8073 1208
rect 8107 1174 8119 1208
rect 8061 1050 8119 1174
rect 8149 1412 8207 1450
rect 8149 1378 8161 1412
rect 8195 1378 8207 1412
rect 8149 1344 8207 1378
rect 8149 1310 8161 1344
rect 8195 1310 8207 1344
rect 8149 1276 8207 1310
rect 8149 1242 8161 1276
rect 8195 1242 8207 1276
rect 8149 1208 8207 1242
rect 8149 1174 8161 1208
rect 8195 1174 8207 1208
rect 8149 1139 8207 1174
rect 8149 1105 8161 1139
rect 8195 1105 8207 1139
rect 8149 1050 8207 1105
rect 8237 1412 8295 1450
rect 8237 1378 8249 1412
rect 8283 1378 8295 1412
rect 8237 1344 8295 1378
rect 8237 1310 8249 1344
rect 8283 1310 8295 1344
rect 8237 1276 8295 1310
rect 8237 1242 8249 1276
rect 8283 1242 8295 1276
rect 8237 1208 8295 1242
rect 8237 1174 8249 1208
rect 8283 1174 8295 1208
rect 8237 1050 8295 1174
rect 8325 1412 8383 1450
rect 8325 1378 8337 1412
rect 8371 1378 8383 1412
rect 8325 1344 8383 1378
rect 8325 1310 8337 1344
rect 8371 1310 8383 1344
rect 8325 1276 8383 1310
rect 8325 1242 8337 1276
rect 8371 1242 8383 1276
rect 8325 1208 8383 1242
rect 8325 1174 8337 1208
rect 8371 1174 8383 1208
rect 8325 1139 8383 1174
rect 8325 1105 8337 1139
rect 8371 1105 8383 1139
rect 8325 1050 8383 1105
rect 8413 1412 8467 1450
rect 8413 1378 8425 1412
rect 8459 1378 8467 1412
rect 8413 1344 8467 1378
rect 8413 1310 8425 1344
rect 8459 1310 8467 1344
rect 8413 1276 8467 1310
rect 8413 1242 8425 1276
rect 8459 1242 8467 1276
rect 8413 1208 8467 1242
rect 8413 1174 8425 1208
rect 8459 1174 8467 1208
rect 8413 1050 8467 1174
rect 8849 1412 8905 1450
rect 8849 1378 8859 1412
rect 8893 1378 8905 1412
rect 8849 1344 8905 1378
rect 8849 1310 8859 1344
rect 8893 1310 8905 1344
rect 8849 1276 8905 1310
rect 8849 1242 8859 1276
rect 8893 1242 8905 1276
rect 8849 1208 8905 1242
rect 8849 1174 8859 1208
rect 8893 1174 8905 1208
rect 8849 1139 8905 1174
rect 8849 1105 8859 1139
rect 8893 1105 8905 1139
rect 8849 1050 8905 1105
rect 8935 1412 8993 1450
rect 8935 1378 8947 1412
rect 8981 1378 8993 1412
rect 8935 1344 8993 1378
rect 8935 1310 8947 1344
rect 8981 1310 8993 1344
rect 8935 1276 8993 1310
rect 8935 1242 8947 1276
rect 8981 1242 8993 1276
rect 8935 1208 8993 1242
rect 8935 1174 8947 1208
rect 8981 1174 8993 1208
rect 8935 1139 8993 1174
rect 8935 1105 8947 1139
rect 8981 1105 8993 1139
rect 8935 1050 8993 1105
rect 9023 1412 9081 1450
rect 9023 1378 9035 1412
rect 9069 1378 9081 1412
rect 9023 1344 9081 1378
rect 9023 1310 9035 1344
rect 9069 1310 9081 1344
rect 9023 1276 9081 1310
rect 9023 1242 9035 1276
rect 9069 1242 9081 1276
rect 9023 1208 9081 1242
rect 9023 1174 9035 1208
rect 9069 1174 9081 1208
rect 9023 1050 9081 1174
rect 9111 1412 9169 1450
rect 9111 1378 9123 1412
rect 9157 1378 9169 1412
rect 9111 1344 9169 1378
rect 9111 1310 9123 1344
rect 9157 1310 9169 1344
rect 9111 1276 9169 1310
rect 9111 1242 9123 1276
rect 9157 1242 9169 1276
rect 9111 1208 9169 1242
rect 9111 1174 9123 1208
rect 9157 1174 9169 1208
rect 9111 1139 9169 1174
rect 9111 1105 9123 1139
rect 9157 1105 9169 1139
rect 9111 1050 9169 1105
rect 9199 1412 9257 1450
rect 9199 1378 9211 1412
rect 9245 1378 9257 1412
rect 9199 1344 9257 1378
rect 9199 1310 9211 1344
rect 9245 1310 9257 1344
rect 9199 1276 9257 1310
rect 9199 1242 9211 1276
rect 9245 1242 9257 1276
rect 9199 1208 9257 1242
rect 9199 1174 9211 1208
rect 9245 1174 9257 1208
rect 9199 1050 9257 1174
rect 9287 1412 9345 1450
rect 9287 1378 9299 1412
rect 9333 1378 9345 1412
rect 9287 1344 9345 1378
rect 9287 1310 9299 1344
rect 9333 1310 9345 1344
rect 9287 1276 9345 1310
rect 9287 1242 9299 1276
rect 9333 1242 9345 1276
rect 9287 1208 9345 1242
rect 9287 1174 9299 1208
rect 9333 1174 9345 1208
rect 9287 1139 9345 1174
rect 9287 1105 9299 1139
rect 9333 1105 9345 1139
rect 9287 1050 9345 1105
rect 9375 1412 9429 1450
rect 9375 1378 9387 1412
rect 9421 1378 9429 1412
rect 9375 1344 9429 1378
rect 9375 1310 9387 1344
rect 9421 1310 9429 1344
rect 9375 1276 9429 1310
rect 9375 1242 9387 1276
rect 9421 1242 9429 1276
rect 9375 1208 9429 1242
rect 9375 1174 9387 1208
rect 9421 1174 9429 1208
rect 9375 1050 9429 1174
rect 9811 1412 9867 1450
rect 9811 1378 9821 1412
rect 9855 1378 9867 1412
rect 9811 1344 9867 1378
rect 9811 1310 9821 1344
rect 9855 1310 9867 1344
rect 9811 1276 9867 1310
rect 9811 1242 9821 1276
rect 9855 1242 9867 1276
rect 9811 1208 9867 1242
rect 9811 1174 9821 1208
rect 9855 1174 9867 1208
rect 9811 1139 9867 1174
rect 9811 1105 9821 1139
rect 9855 1105 9867 1139
rect 9811 1050 9867 1105
rect 9897 1412 9955 1450
rect 9897 1378 9909 1412
rect 9943 1378 9955 1412
rect 9897 1344 9955 1378
rect 9897 1310 9909 1344
rect 9943 1310 9955 1344
rect 9897 1276 9955 1310
rect 9897 1242 9909 1276
rect 9943 1242 9955 1276
rect 9897 1208 9955 1242
rect 9897 1174 9909 1208
rect 9943 1174 9955 1208
rect 9897 1139 9955 1174
rect 9897 1105 9909 1139
rect 9943 1105 9955 1139
rect 9897 1050 9955 1105
rect 9985 1412 10043 1450
rect 9985 1378 9997 1412
rect 10031 1378 10043 1412
rect 9985 1344 10043 1378
rect 9985 1310 9997 1344
rect 10031 1310 10043 1344
rect 9985 1276 10043 1310
rect 9985 1242 9997 1276
rect 10031 1242 10043 1276
rect 9985 1208 10043 1242
rect 9985 1174 9997 1208
rect 10031 1174 10043 1208
rect 9985 1050 10043 1174
rect 10073 1412 10131 1450
rect 10073 1378 10085 1412
rect 10119 1378 10131 1412
rect 10073 1344 10131 1378
rect 10073 1310 10085 1344
rect 10119 1310 10131 1344
rect 10073 1276 10131 1310
rect 10073 1242 10085 1276
rect 10119 1242 10131 1276
rect 10073 1208 10131 1242
rect 10073 1174 10085 1208
rect 10119 1174 10131 1208
rect 10073 1139 10131 1174
rect 10073 1105 10085 1139
rect 10119 1105 10131 1139
rect 10073 1050 10131 1105
rect 10161 1412 10219 1450
rect 10161 1378 10173 1412
rect 10207 1378 10219 1412
rect 10161 1344 10219 1378
rect 10161 1310 10173 1344
rect 10207 1310 10219 1344
rect 10161 1276 10219 1310
rect 10161 1242 10173 1276
rect 10207 1242 10219 1276
rect 10161 1208 10219 1242
rect 10161 1174 10173 1208
rect 10207 1174 10219 1208
rect 10161 1050 10219 1174
rect 10249 1412 10307 1450
rect 10249 1378 10261 1412
rect 10295 1378 10307 1412
rect 10249 1344 10307 1378
rect 10249 1310 10261 1344
rect 10295 1310 10307 1344
rect 10249 1276 10307 1310
rect 10249 1242 10261 1276
rect 10295 1242 10307 1276
rect 10249 1208 10307 1242
rect 10249 1174 10261 1208
rect 10295 1174 10307 1208
rect 10249 1139 10307 1174
rect 10249 1105 10261 1139
rect 10295 1105 10307 1139
rect 10249 1050 10307 1105
rect 10337 1412 10391 1450
rect 10337 1378 10349 1412
rect 10383 1378 10391 1412
rect 10337 1344 10391 1378
rect 10337 1310 10349 1344
rect 10383 1310 10391 1344
rect 10337 1276 10391 1310
rect 10337 1242 10349 1276
rect 10383 1242 10391 1276
rect 10337 1208 10391 1242
rect 10337 1174 10349 1208
rect 10383 1174 10391 1208
rect 10337 1050 10391 1174
rect 10773 1412 10829 1450
rect 10773 1378 10783 1412
rect 10817 1378 10829 1412
rect 10773 1344 10829 1378
rect 10773 1310 10783 1344
rect 10817 1310 10829 1344
rect 10773 1276 10829 1310
rect 10773 1242 10783 1276
rect 10817 1242 10829 1276
rect 10773 1208 10829 1242
rect 10773 1174 10783 1208
rect 10817 1174 10829 1208
rect 10773 1139 10829 1174
rect 10773 1105 10783 1139
rect 10817 1105 10829 1139
rect 10773 1050 10829 1105
rect 10859 1412 10917 1450
rect 10859 1378 10871 1412
rect 10905 1378 10917 1412
rect 10859 1344 10917 1378
rect 10859 1310 10871 1344
rect 10905 1310 10917 1344
rect 10859 1276 10917 1310
rect 10859 1242 10871 1276
rect 10905 1242 10917 1276
rect 10859 1208 10917 1242
rect 10859 1174 10871 1208
rect 10905 1174 10917 1208
rect 10859 1139 10917 1174
rect 10859 1105 10871 1139
rect 10905 1105 10917 1139
rect 10859 1050 10917 1105
rect 10947 1412 11005 1450
rect 10947 1378 10959 1412
rect 10993 1378 11005 1412
rect 10947 1344 11005 1378
rect 10947 1310 10959 1344
rect 10993 1310 11005 1344
rect 10947 1276 11005 1310
rect 10947 1242 10959 1276
rect 10993 1242 11005 1276
rect 10947 1208 11005 1242
rect 10947 1174 10959 1208
rect 10993 1174 11005 1208
rect 10947 1050 11005 1174
rect 11035 1412 11093 1450
rect 11035 1378 11047 1412
rect 11081 1378 11093 1412
rect 11035 1344 11093 1378
rect 11035 1310 11047 1344
rect 11081 1310 11093 1344
rect 11035 1276 11093 1310
rect 11035 1242 11047 1276
rect 11081 1242 11093 1276
rect 11035 1208 11093 1242
rect 11035 1174 11047 1208
rect 11081 1174 11093 1208
rect 11035 1139 11093 1174
rect 11035 1105 11047 1139
rect 11081 1105 11093 1139
rect 11035 1050 11093 1105
rect 11123 1412 11181 1450
rect 11123 1378 11135 1412
rect 11169 1378 11181 1412
rect 11123 1344 11181 1378
rect 11123 1310 11135 1344
rect 11169 1310 11181 1344
rect 11123 1276 11181 1310
rect 11123 1242 11135 1276
rect 11169 1242 11181 1276
rect 11123 1208 11181 1242
rect 11123 1174 11135 1208
rect 11169 1174 11181 1208
rect 11123 1050 11181 1174
rect 11211 1412 11269 1450
rect 11211 1378 11223 1412
rect 11257 1378 11269 1412
rect 11211 1344 11269 1378
rect 11211 1310 11223 1344
rect 11257 1310 11269 1344
rect 11211 1276 11269 1310
rect 11211 1242 11223 1276
rect 11257 1242 11269 1276
rect 11211 1208 11269 1242
rect 11211 1174 11223 1208
rect 11257 1174 11269 1208
rect 11211 1139 11269 1174
rect 11211 1105 11223 1139
rect 11257 1105 11269 1139
rect 11211 1050 11269 1105
rect 11299 1412 11353 1450
rect 11299 1378 11311 1412
rect 11345 1378 11353 1412
rect 11299 1344 11353 1378
rect 11299 1310 11311 1344
rect 11345 1310 11353 1344
rect 11299 1276 11353 1310
rect 11299 1242 11311 1276
rect 11345 1242 11353 1276
rect 11299 1208 11353 1242
rect 11299 1174 11311 1208
rect 11345 1174 11353 1208
rect 11299 1050 11353 1174
rect 11735 1412 11791 1450
rect 11735 1378 11745 1412
rect 11779 1378 11791 1412
rect 11735 1344 11791 1378
rect 11735 1310 11745 1344
rect 11779 1310 11791 1344
rect 11735 1276 11791 1310
rect 11735 1242 11745 1276
rect 11779 1242 11791 1276
rect 11735 1208 11791 1242
rect 11735 1174 11745 1208
rect 11779 1174 11791 1208
rect 11735 1139 11791 1174
rect 11735 1105 11745 1139
rect 11779 1105 11791 1139
rect 11735 1050 11791 1105
rect 11821 1412 11879 1450
rect 11821 1378 11833 1412
rect 11867 1378 11879 1412
rect 11821 1344 11879 1378
rect 11821 1310 11833 1344
rect 11867 1310 11879 1344
rect 11821 1276 11879 1310
rect 11821 1242 11833 1276
rect 11867 1242 11879 1276
rect 11821 1208 11879 1242
rect 11821 1174 11833 1208
rect 11867 1174 11879 1208
rect 11821 1139 11879 1174
rect 11821 1105 11833 1139
rect 11867 1105 11879 1139
rect 11821 1050 11879 1105
rect 11909 1412 11967 1450
rect 11909 1378 11921 1412
rect 11955 1378 11967 1412
rect 11909 1344 11967 1378
rect 11909 1310 11921 1344
rect 11955 1310 11967 1344
rect 11909 1276 11967 1310
rect 11909 1242 11921 1276
rect 11955 1242 11967 1276
rect 11909 1208 11967 1242
rect 11909 1174 11921 1208
rect 11955 1174 11967 1208
rect 11909 1050 11967 1174
rect 11997 1412 12055 1450
rect 11997 1378 12009 1412
rect 12043 1378 12055 1412
rect 11997 1344 12055 1378
rect 11997 1310 12009 1344
rect 12043 1310 12055 1344
rect 11997 1276 12055 1310
rect 11997 1242 12009 1276
rect 12043 1242 12055 1276
rect 11997 1208 12055 1242
rect 11997 1174 12009 1208
rect 12043 1174 12055 1208
rect 11997 1139 12055 1174
rect 11997 1105 12009 1139
rect 12043 1105 12055 1139
rect 11997 1050 12055 1105
rect 12085 1412 12143 1450
rect 12085 1378 12097 1412
rect 12131 1378 12143 1412
rect 12085 1344 12143 1378
rect 12085 1310 12097 1344
rect 12131 1310 12143 1344
rect 12085 1276 12143 1310
rect 12085 1242 12097 1276
rect 12131 1242 12143 1276
rect 12085 1208 12143 1242
rect 12085 1174 12097 1208
rect 12131 1174 12143 1208
rect 12085 1050 12143 1174
rect 12173 1412 12231 1450
rect 12173 1378 12185 1412
rect 12219 1378 12231 1412
rect 12173 1344 12231 1378
rect 12173 1310 12185 1344
rect 12219 1310 12231 1344
rect 12173 1276 12231 1310
rect 12173 1242 12185 1276
rect 12219 1242 12231 1276
rect 12173 1208 12231 1242
rect 12173 1174 12185 1208
rect 12219 1174 12231 1208
rect 12173 1139 12231 1174
rect 12173 1105 12185 1139
rect 12219 1105 12231 1139
rect 12173 1050 12231 1105
rect 12261 1412 12315 1450
rect 12261 1378 12273 1412
rect 12307 1378 12315 1412
rect 12261 1344 12315 1378
rect 12261 1310 12273 1344
rect 12307 1310 12315 1344
rect 12261 1276 12315 1310
rect 12261 1242 12273 1276
rect 12307 1242 12315 1276
rect 12261 1208 12315 1242
rect 12261 1174 12273 1208
rect 12307 1174 12315 1208
rect 12261 1050 12315 1174
rect 12697 1412 12753 1450
rect 12697 1378 12707 1412
rect 12741 1378 12753 1412
rect 12697 1344 12753 1378
rect 12697 1310 12707 1344
rect 12741 1310 12753 1344
rect 12697 1276 12753 1310
rect 12697 1242 12707 1276
rect 12741 1242 12753 1276
rect 12697 1208 12753 1242
rect 12697 1174 12707 1208
rect 12741 1174 12753 1208
rect 12697 1139 12753 1174
rect 12697 1105 12707 1139
rect 12741 1105 12753 1139
rect 12697 1050 12753 1105
rect 12783 1412 12841 1450
rect 12783 1378 12795 1412
rect 12829 1378 12841 1412
rect 12783 1344 12841 1378
rect 12783 1310 12795 1344
rect 12829 1310 12841 1344
rect 12783 1276 12841 1310
rect 12783 1242 12795 1276
rect 12829 1242 12841 1276
rect 12783 1208 12841 1242
rect 12783 1174 12795 1208
rect 12829 1174 12841 1208
rect 12783 1139 12841 1174
rect 12783 1105 12795 1139
rect 12829 1105 12841 1139
rect 12783 1050 12841 1105
rect 12871 1412 12929 1450
rect 12871 1378 12883 1412
rect 12917 1378 12929 1412
rect 12871 1344 12929 1378
rect 12871 1310 12883 1344
rect 12917 1310 12929 1344
rect 12871 1276 12929 1310
rect 12871 1242 12883 1276
rect 12917 1242 12929 1276
rect 12871 1208 12929 1242
rect 12871 1174 12883 1208
rect 12917 1174 12929 1208
rect 12871 1050 12929 1174
rect 12959 1412 13017 1450
rect 12959 1378 12971 1412
rect 13005 1378 13017 1412
rect 12959 1344 13017 1378
rect 12959 1310 12971 1344
rect 13005 1310 13017 1344
rect 12959 1276 13017 1310
rect 12959 1242 12971 1276
rect 13005 1242 13017 1276
rect 12959 1208 13017 1242
rect 12959 1174 12971 1208
rect 13005 1174 13017 1208
rect 12959 1139 13017 1174
rect 12959 1105 12971 1139
rect 13005 1105 13017 1139
rect 12959 1050 13017 1105
rect 13047 1412 13105 1450
rect 13047 1378 13059 1412
rect 13093 1378 13105 1412
rect 13047 1344 13105 1378
rect 13047 1310 13059 1344
rect 13093 1310 13105 1344
rect 13047 1276 13105 1310
rect 13047 1242 13059 1276
rect 13093 1242 13105 1276
rect 13047 1208 13105 1242
rect 13047 1174 13059 1208
rect 13093 1174 13105 1208
rect 13047 1050 13105 1174
rect 13135 1412 13193 1450
rect 13135 1378 13147 1412
rect 13181 1378 13193 1412
rect 13135 1344 13193 1378
rect 13135 1310 13147 1344
rect 13181 1310 13193 1344
rect 13135 1276 13193 1310
rect 13135 1242 13147 1276
rect 13181 1242 13193 1276
rect 13135 1208 13193 1242
rect 13135 1174 13147 1208
rect 13181 1174 13193 1208
rect 13135 1139 13193 1174
rect 13135 1105 13147 1139
rect 13181 1105 13193 1139
rect 13135 1050 13193 1105
rect 13223 1412 13277 1450
rect 13223 1378 13235 1412
rect 13269 1378 13277 1412
rect 13223 1344 13277 1378
rect 13223 1310 13235 1344
rect 13269 1310 13277 1344
rect 13223 1276 13277 1310
rect 13223 1242 13235 1276
rect 13269 1242 13277 1276
rect 13223 1208 13277 1242
rect 13223 1174 13235 1208
rect 13269 1174 13277 1208
rect 13223 1050 13277 1174
rect 13659 1412 13715 1450
rect 13659 1378 13669 1412
rect 13703 1378 13715 1412
rect 13659 1344 13715 1378
rect 13659 1310 13669 1344
rect 13703 1310 13715 1344
rect 13659 1276 13715 1310
rect 13659 1242 13669 1276
rect 13703 1242 13715 1276
rect 13659 1208 13715 1242
rect 13659 1174 13669 1208
rect 13703 1174 13715 1208
rect 13659 1139 13715 1174
rect 13659 1105 13669 1139
rect 13703 1105 13715 1139
rect 13659 1050 13715 1105
rect 13745 1412 13803 1450
rect 13745 1378 13757 1412
rect 13791 1378 13803 1412
rect 13745 1344 13803 1378
rect 13745 1310 13757 1344
rect 13791 1310 13803 1344
rect 13745 1276 13803 1310
rect 13745 1242 13757 1276
rect 13791 1242 13803 1276
rect 13745 1208 13803 1242
rect 13745 1174 13757 1208
rect 13791 1174 13803 1208
rect 13745 1139 13803 1174
rect 13745 1105 13757 1139
rect 13791 1105 13803 1139
rect 13745 1050 13803 1105
rect 13833 1412 13891 1450
rect 13833 1378 13845 1412
rect 13879 1378 13891 1412
rect 13833 1344 13891 1378
rect 13833 1310 13845 1344
rect 13879 1310 13891 1344
rect 13833 1276 13891 1310
rect 13833 1242 13845 1276
rect 13879 1242 13891 1276
rect 13833 1208 13891 1242
rect 13833 1174 13845 1208
rect 13879 1174 13891 1208
rect 13833 1050 13891 1174
rect 13921 1412 13979 1450
rect 13921 1378 13933 1412
rect 13967 1378 13979 1412
rect 13921 1344 13979 1378
rect 13921 1310 13933 1344
rect 13967 1310 13979 1344
rect 13921 1276 13979 1310
rect 13921 1242 13933 1276
rect 13967 1242 13979 1276
rect 13921 1208 13979 1242
rect 13921 1174 13933 1208
rect 13967 1174 13979 1208
rect 13921 1139 13979 1174
rect 13921 1105 13933 1139
rect 13967 1105 13979 1139
rect 13921 1050 13979 1105
rect 14009 1412 14067 1450
rect 14009 1378 14021 1412
rect 14055 1378 14067 1412
rect 14009 1344 14067 1378
rect 14009 1310 14021 1344
rect 14055 1310 14067 1344
rect 14009 1276 14067 1310
rect 14009 1242 14021 1276
rect 14055 1242 14067 1276
rect 14009 1208 14067 1242
rect 14009 1174 14021 1208
rect 14055 1174 14067 1208
rect 14009 1050 14067 1174
rect 14097 1412 14155 1450
rect 14097 1378 14109 1412
rect 14143 1378 14155 1412
rect 14097 1344 14155 1378
rect 14097 1310 14109 1344
rect 14143 1310 14155 1344
rect 14097 1276 14155 1310
rect 14097 1242 14109 1276
rect 14143 1242 14155 1276
rect 14097 1208 14155 1242
rect 14097 1174 14109 1208
rect 14143 1174 14155 1208
rect 14097 1139 14155 1174
rect 14097 1105 14109 1139
rect 14143 1105 14155 1139
rect 14097 1050 14155 1105
rect 14185 1412 14239 1450
rect 14185 1378 14197 1412
rect 14231 1378 14239 1412
rect 14185 1344 14239 1378
rect 14185 1310 14197 1344
rect 14231 1310 14239 1344
rect 14185 1276 14239 1310
rect 14185 1242 14197 1276
rect 14231 1242 14239 1276
rect 14185 1208 14239 1242
rect 14185 1174 14197 1208
rect 14231 1174 14239 1208
rect 14185 1050 14239 1174
rect 14621 1412 14677 1450
rect 14621 1378 14631 1412
rect 14665 1378 14677 1412
rect 14621 1344 14677 1378
rect 14621 1310 14631 1344
rect 14665 1310 14677 1344
rect 14621 1276 14677 1310
rect 14621 1242 14631 1276
rect 14665 1242 14677 1276
rect 14621 1208 14677 1242
rect 14621 1174 14631 1208
rect 14665 1174 14677 1208
rect 14621 1139 14677 1174
rect 14621 1105 14631 1139
rect 14665 1105 14677 1139
rect 14621 1050 14677 1105
rect 14707 1412 14765 1450
rect 14707 1378 14719 1412
rect 14753 1378 14765 1412
rect 14707 1344 14765 1378
rect 14707 1310 14719 1344
rect 14753 1310 14765 1344
rect 14707 1276 14765 1310
rect 14707 1242 14719 1276
rect 14753 1242 14765 1276
rect 14707 1208 14765 1242
rect 14707 1174 14719 1208
rect 14753 1174 14765 1208
rect 14707 1139 14765 1174
rect 14707 1105 14719 1139
rect 14753 1105 14765 1139
rect 14707 1050 14765 1105
rect 14795 1412 14853 1450
rect 14795 1378 14807 1412
rect 14841 1378 14853 1412
rect 14795 1344 14853 1378
rect 14795 1310 14807 1344
rect 14841 1310 14853 1344
rect 14795 1276 14853 1310
rect 14795 1242 14807 1276
rect 14841 1242 14853 1276
rect 14795 1208 14853 1242
rect 14795 1174 14807 1208
rect 14841 1174 14853 1208
rect 14795 1050 14853 1174
rect 14883 1412 14941 1450
rect 14883 1378 14895 1412
rect 14929 1378 14941 1412
rect 14883 1344 14941 1378
rect 14883 1310 14895 1344
rect 14929 1310 14941 1344
rect 14883 1276 14941 1310
rect 14883 1242 14895 1276
rect 14929 1242 14941 1276
rect 14883 1208 14941 1242
rect 14883 1174 14895 1208
rect 14929 1174 14941 1208
rect 14883 1139 14941 1174
rect 14883 1105 14895 1139
rect 14929 1105 14941 1139
rect 14883 1050 14941 1105
rect 14971 1412 15029 1450
rect 14971 1378 14983 1412
rect 15017 1378 15029 1412
rect 14971 1344 15029 1378
rect 14971 1310 14983 1344
rect 15017 1310 15029 1344
rect 14971 1276 15029 1310
rect 14971 1242 14983 1276
rect 15017 1242 15029 1276
rect 14971 1208 15029 1242
rect 14971 1174 14983 1208
rect 15017 1174 15029 1208
rect 14971 1050 15029 1174
rect 15059 1412 15117 1450
rect 15059 1378 15071 1412
rect 15105 1378 15117 1412
rect 15059 1344 15117 1378
rect 15059 1310 15071 1344
rect 15105 1310 15117 1344
rect 15059 1276 15117 1310
rect 15059 1242 15071 1276
rect 15105 1242 15117 1276
rect 15059 1208 15117 1242
rect 15059 1174 15071 1208
rect 15105 1174 15117 1208
rect 15059 1139 15117 1174
rect 15059 1105 15071 1139
rect 15105 1105 15117 1139
rect 15059 1050 15117 1105
rect 15147 1412 15201 1450
rect 15147 1378 15159 1412
rect 15193 1378 15201 1412
rect 15147 1344 15201 1378
rect 15147 1310 15159 1344
rect 15193 1310 15201 1344
rect 15147 1276 15201 1310
rect 15147 1242 15159 1276
rect 15193 1242 15201 1276
rect 15147 1208 15201 1242
rect 15147 1174 15159 1208
rect 15193 1174 15201 1208
rect 15147 1050 15201 1174
rect 15583 1412 15639 1450
rect 15583 1378 15593 1412
rect 15627 1378 15639 1412
rect 15583 1344 15639 1378
rect 15583 1310 15593 1344
rect 15627 1310 15639 1344
rect 15583 1276 15639 1310
rect 15583 1242 15593 1276
rect 15627 1242 15639 1276
rect 15583 1208 15639 1242
rect 15583 1174 15593 1208
rect 15627 1174 15639 1208
rect 15583 1139 15639 1174
rect 15583 1105 15593 1139
rect 15627 1105 15639 1139
rect 15583 1050 15639 1105
rect 15669 1412 15727 1450
rect 15669 1378 15681 1412
rect 15715 1378 15727 1412
rect 15669 1344 15727 1378
rect 15669 1310 15681 1344
rect 15715 1310 15727 1344
rect 15669 1276 15727 1310
rect 15669 1242 15681 1276
rect 15715 1242 15727 1276
rect 15669 1208 15727 1242
rect 15669 1174 15681 1208
rect 15715 1174 15727 1208
rect 15669 1139 15727 1174
rect 15669 1105 15681 1139
rect 15715 1105 15727 1139
rect 15669 1050 15727 1105
rect 15757 1412 15815 1450
rect 15757 1378 15769 1412
rect 15803 1378 15815 1412
rect 15757 1344 15815 1378
rect 15757 1310 15769 1344
rect 15803 1310 15815 1344
rect 15757 1276 15815 1310
rect 15757 1242 15769 1276
rect 15803 1242 15815 1276
rect 15757 1208 15815 1242
rect 15757 1174 15769 1208
rect 15803 1174 15815 1208
rect 15757 1050 15815 1174
rect 15845 1412 15903 1450
rect 15845 1378 15857 1412
rect 15891 1378 15903 1412
rect 15845 1344 15903 1378
rect 15845 1310 15857 1344
rect 15891 1310 15903 1344
rect 15845 1276 15903 1310
rect 15845 1242 15857 1276
rect 15891 1242 15903 1276
rect 15845 1208 15903 1242
rect 15845 1174 15857 1208
rect 15891 1174 15903 1208
rect 15845 1139 15903 1174
rect 15845 1105 15857 1139
rect 15891 1105 15903 1139
rect 15845 1050 15903 1105
rect 15933 1412 15991 1450
rect 15933 1378 15945 1412
rect 15979 1378 15991 1412
rect 15933 1344 15991 1378
rect 15933 1310 15945 1344
rect 15979 1310 15991 1344
rect 15933 1276 15991 1310
rect 15933 1242 15945 1276
rect 15979 1242 15991 1276
rect 15933 1208 15991 1242
rect 15933 1174 15945 1208
rect 15979 1174 15991 1208
rect 15933 1050 15991 1174
rect 16021 1412 16079 1450
rect 16021 1378 16033 1412
rect 16067 1378 16079 1412
rect 16021 1344 16079 1378
rect 16021 1310 16033 1344
rect 16067 1310 16079 1344
rect 16021 1276 16079 1310
rect 16021 1242 16033 1276
rect 16067 1242 16079 1276
rect 16021 1208 16079 1242
rect 16021 1174 16033 1208
rect 16067 1174 16079 1208
rect 16021 1139 16079 1174
rect 16021 1105 16033 1139
rect 16067 1105 16079 1139
rect 16021 1050 16079 1105
rect 16109 1412 16163 1450
rect 16109 1378 16121 1412
rect 16155 1378 16163 1412
rect 16109 1344 16163 1378
rect 16109 1310 16121 1344
rect 16155 1310 16163 1344
rect 16109 1276 16163 1310
rect 16109 1242 16121 1276
rect 16155 1242 16163 1276
rect 16109 1208 16163 1242
rect 16109 1174 16121 1208
rect 16155 1174 16163 1208
rect 16109 1050 16163 1174
rect 16545 1412 16601 1450
rect 16545 1378 16555 1412
rect 16589 1378 16601 1412
rect 16545 1344 16601 1378
rect 16545 1310 16555 1344
rect 16589 1310 16601 1344
rect 16545 1276 16601 1310
rect 16545 1242 16555 1276
rect 16589 1242 16601 1276
rect 16545 1208 16601 1242
rect 16545 1174 16555 1208
rect 16589 1174 16601 1208
rect 16545 1139 16601 1174
rect 16545 1105 16555 1139
rect 16589 1105 16601 1139
rect 16545 1050 16601 1105
rect 16631 1412 16689 1450
rect 16631 1378 16643 1412
rect 16677 1378 16689 1412
rect 16631 1344 16689 1378
rect 16631 1310 16643 1344
rect 16677 1310 16689 1344
rect 16631 1276 16689 1310
rect 16631 1242 16643 1276
rect 16677 1242 16689 1276
rect 16631 1208 16689 1242
rect 16631 1174 16643 1208
rect 16677 1174 16689 1208
rect 16631 1139 16689 1174
rect 16631 1105 16643 1139
rect 16677 1105 16689 1139
rect 16631 1050 16689 1105
rect 16719 1412 16777 1450
rect 16719 1378 16731 1412
rect 16765 1378 16777 1412
rect 16719 1344 16777 1378
rect 16719 1310 16731 1344
rect 16765 1310 16777 1344
rect 16719 1276 16777 1310
rect 16719 1242 16731 1276
rect 16765 1242 16777 1276
rect 16719 1208 16777 1242
rect 16719 1174 16731 1208
rect 16765 1174 16777 1208
rect 16719 1050 16777 1174
rect 16807 1412 16865 1450
rect 16807 1378 16819 1412
rect 16853 1378 16865 1412
rect 16807 1344 16865 1378
rect 16807 1310 16819 1344
rect 16853 1310 16865 1344
rect 16807 1276 16865 1310
rect 16807 1242 16819 1276
rect 16853 1242 16865 1276
rect 16807 1208 16865 1242
rect 16807 1174 16819 1208
rect 16853 1174 16865 1208
rect 16807 1139 16865 1174
rect 16807 1105 16819 1139
rect 16853 1105 16865 1139
rect 16807 1050 16865 1105
rect 16895 1412 16953 1450
rect 16895 1378 16907 1412
rect 16941 1378 16953 1412
rect 16895 1344 16953 1378
rect 16895 1310 16907 1344
rect 16941 1310 16953 1344
rect 16895 1276 16953 1310
rect 16895 1242 16907 1276
rect 16941 1242 16953 1276
rect 16895 1208 16953 1242
rect 16895 1174 16907 1208
rect 16941 1174 16953 1208
rect 16895 1050 16953 1174
rect 16983 1412 17041 1450
rect 16983 1378 16995 1412
rect 17029 1378 17041 1412
rect 16983 1344 17041 1378
rect 16983 1310 16995 1344
rect 17029 1310 17041 1344
rect 16983 1276 17041 1310
rect 16983 1242 16995 1276
rect 17029 1242 17041 1276
rect 16983 1208 17041 1242
rect 16983 1174 16995 1208
rect 17029 1174 17041 1208
rect 16983 1139 17041 1174
rect 16983 1105 16995 1139
rect 17029 1105 17041 1139
rect 16983 1050 17041 1105
rect 17071 1412 17125 1450
rect 17071 1378 17083 1412
rect 17117 1378 17125 1412
rect 17071 1344 17125 1378
rect 17071 1310 17083 1344
rect 17117 1310 17125 1344
rect 17071 1276 17125 1310
rect 17071 1242 17083 1276
rect 17117 1242 17125 1276
rect 17071 1208 17125 1242
rect 17071 1174 17083 1208
rect 17117 1174 17125 1208
rect 17071 1050 17125 1174
rect 17447 1411 17503 1451
rect 17447 1377 17457 1411
rect 17491 1377 17503 1411
rect 17447 1343 17503 1377
rect 17447 1309 17457 1343
rect 17491 1309 17503 1343
rect 17447 1275 17503 1309
rect 17447 1241 17457 1275
rect 17491 1241 17503 1275
rect 17447 1207 17503 1241
rect 17447 1173 17457 1207
rect 17491 1173 17503 1207
rect 17447 1139 17503 1173
rect 17447 1105 17457 1139
rect 17491 1105 17503 1139
rect 17447 1051 17503 1105
rect 17533 1411 17591 1451
rect 17533 1377 17545 1411
rect 17579 1377 17591 1411
rect 17533 1343 17591 1377
rect 17533 1309 17545 1343
rect 17579 1309 17591 1343
rect 17533 1275 17591 1309
rect 17533 1241 17545 1275
rect 17579 1241 17591 1275
rect 17533 1207 17591 1241
rect 17533 1173 17545 1207
rect 17579 1173 17591 1207
rect 17533 1139 17591 1173
rect 17533 1105 17545 1139
rect 17579 1105 17591 1139
rect 17533 1051 17591 1105
rect 17621 1411 17679 1451
rect 17621 1377 17633 1411
rect 17667 1377 17679 1411
rect 17621 1343 17679 1377
rect 17621 1309 17633 1343
rect 17667 1309 17679 1343
rect 17621 1275 17679 1309
rect 17621 1241 17633 1275
rect 17667 1241 17679 1275
rect 17621 1207 17679 1241
rect 17621 1173 17633 1207
rect 17667 1173 17679 1207
rect 17621 1051 17679 1173
rect 17709 1411 17767 1451
rect 17709 1377 17721 1411
rect 17755 1377 17767 1411
rect 17709 1343 17767 1377
rect 17709 1309 17721 1343
rect 17755 1309 17767 1343
rect 17709 1275 17767 1309
rect 17709 1241 17721 1275
rect 17755 1241 17767 1275
rect 17709 1207 17767 1241
rect 17709 1173 17721 1207
rect 17755 1173 17767 1207
rect 17709 1051 17767 1173
rect 17797 1411 17851 1451
rect 17797 1377 17809 1411
rect 17843 1377 17851 1411
rect 17797 1343 17851 1377
rect 17797 1309 17809 1343
rect 17843 1309 17851 1343
rect 17797 1275 17851 1309
rect 17797 1241 17809 1275
rect 17843 1241 17851 1275
rect 17797 1207 17851 1241
rect 17797 1173 17809 1207
rect 17843 1173 17851 1207
rect 17797 1139 17851 1173
rect 17797 1105 17809 1139
rect 17843 1105 17851 1139
rect 17797 1051 17851 1105
rect 18113 1411 18167 1451
rect 18113 1377 18121 1411
rect 18155 1377 18167 1411
rect 18113 1343 18167 1377
rect 18113 1309 18121 1343
rect 18155 1309 18167 1343
rect 18113 1275 18167 1309
rect 18113 1241 18121 1275
rect 18155 1241 18167 1275
rect 18113 1207 18167 1241
rect 18113 1173 18121 1207
rect 18155 1173 18167 1207
rect 18113 1051 18167 1173
rect 18197 1343 18255 1451
rect 18197 1309 18209 1343
rect 18243 1309 18255 1343
rect 18197 1275 18255 1309
rect 18197 1241 18209 1275
rect 18243 1241 18255 1275
rect 18197 1207 18255 1241
rect 18197 1173 18209 1207
rect 18243 1173 18255 1207
rect 18197 1139 18255 1173
rect 18197 1105 18209 1139
rect 18243 1105 18255 1139
rect 18197 1051 18255 1105
rect 18285 1411 18343 1451
rect 18285 1377 18297 1411
rect 18331 1377 18343 1411
rect 18285 1343 18343 1377
rect 18285 1309 18297 1343
rect 18331 1309 18343 1343
rect 18285 1275 18343 1309
rect 18285 1241 18297 1275
rect 18331 1241 18343 1275
rect 18285 1207 18343 1241
rect 18285 1173 18297 1207
rect 18331 1173 18343 1207
rect 18285 1051 18343 1173
rect 18373 1343 18431 1451
rect 18373 1309 18385 1343
rect 18419 1309 18431 1343
rect 18373 1275 18431 1309
rect 18373 1241 18385 1275
rect 18419 1241 18431 1275
rect 18373 1207 18431 1241
rect 18373 1173 18385 1207
rect 18419 1173 18431 1207
rect 18373 1051 18431 1173
rect 18461 1411 18517 1451
rect 18461 1377 18473 1411
rect 18507 1377 18517 1411
rect 18461 1343 18517 1377
rect 18461 1309 18473 1343
rect 18507 1309 18517 1343
rect 18461 1275 18517 1309
rect 18461 1241 18473 1275
rect 18507 1241 18517 1275
rect 18461 1207 18517 1241
rect 18461 1173 18473 1207
rect 18507 1173 18517 1207
rect 18461 1051 18517 1173
rect 18779 1411 18835 1451
rect 18779 1377 18789 1411
rect 18823 1377 18835 1411
rect 18779 1343 18835 1377
rect 18779 1309 18789 1343
rect 18823 1309 18835 1343
rect 18779 1275 18835 1309
rect 18779 1241 18789 1275
rect 18823 1241 18835 1275
rect 18779 1207 18835 1241
rect 18779 1173 18789 1207
rect 18823 1173 18835 1207
rect 18779 1051 18835 1173
rect 18865 1343 18923 1451
rect 18865 1309 18877 1343
rect 18911 1309 18923 1343
rect 18865 1275 18923 1309
rect 18865 1241 18877 1275
rect 18911 1241 18923 1275
rect 18865 1207 18923 1241
rect 18865 1173 18877 1207
rect 18911 1173 18923 1207
rect 18865 1139 18923 1173
rect 18865 1105 18877 1139
rect 18911 1105 18923 1139
rect 18865 1051 18923 1105
rect 18953 1411 19011 1451
rect 18953 1377 18965 1411
rect 18999 1377 19011 1411
rect 18953 1343 19011 1377
rect 18953 1309 18965 1343
rect 18999 1309 19011 1343
rect 18953 1275 19011 1309
rect 18953 1241 18965 1275
rect 18999 1241 19011 1275
rect 18953 1207 19011 1241
rect 18953 1173 18965 1207
rect 18999 1173 19011 1207
rect 18953 1051 19011 1173
rect 19041 1343 19099 1451
rect 19041 1309 19053 1343
rect 19087 1309 19099 1343
rect 19041 1275 19099 1309
rect 19041 1241 19053 1275
rect 19087 1241 19099 1275
rect 19041 1207 19099 1241
rect 19041 1173 19053 1207
rect 19087 1173 19099 1207
rect 19041 1139 19099 1173
rect 19041 1105 19053 1139
rect 19087 1105 19099 1139
rect 19041 1051 19099 1105
rect 19129 1411 19183 1451
rect 19129 1377 19141 1411
rect 19175 1377 19183 1411
rect 19129 1343 19183 1377
rect 19129 1309 19141 1343
rect 19175 1309 19183 1343
rect 19129 1275 19183 1309
rect 19129 1241 19141 1275
rect 19175 1241 19183 1275
rect 19129 1207 19183 1241
rect 19129 1173 19141 1207
rect 19175 1173 19183 1207
rect 19129 1051 19183 1173
<< ndiffc >>
rect 101 329 135 363
rect 198 329 232 363
rect 295 329 329 363
rect 392 329 426 363
rect 489 329 523 363
rect 101 257 135 291
rect 101 189 135 223
rect 198 204 232 238
rect 295 257 329 291
rect 295 189 329 223
rect 393 210 427 244
rect 101 119 135 153
rect 295 119 329 153
rect 392 119 426 153
rect 489 119 523 153
rect 603 329 637 363
rect 603 257 637 291
rect 603 189 637 223
rect 700 213 734 247
rect 797 257 831 291
rect 797 189 831 223
rect 603 119 637 153
rect 700 119 734 153
rect 797 119 831 153
rect 1063 329 1097 363
rect 1160 329 1194 363
rect 1257 329 1291 363
rect 1354 329 1388 363
rect 1451 329 1485 363
rect 1063 257 1097 291
rect 1063 189 1097 223
rect 1160 204 1194 238
rect 1257 257 1291 291
rect 1257 189 1291 223
rect 1355 210 1389 244
rect 1063 119 1097 153
rect 1257 119 1291 153
rect 1354 119 1388 153
rect 1451 119 1485 153
rect 1565 329 1599 363
rect 1565 257 1599 291
rect 1565 189 1599 223
rect 1662 213 1696 247
rect 1759 257 1793 291
rect 1759 189 1793 223
rect 1565 119 1599 153
rect 1662 119 1696 153
rect 1759 119 1793 153
rect 2025 329 2059 363
rect 2122 329 2156 363
rect 2219 329 2253 363
rect 2316 329 2350 363
rect 2413 329 2447 363
rect 2025 257 2059 291
rect 2025 189 2059 223
rect 2122 204 2156 238
rect 2219 257 2253 291
rect 2219 189 2253 223
rect 2317 210 2351 244
rect 2025 119 2059 153
rect 2219 119 2253 153
rect 2316 119 2350 153
rect 2413 119 2447 153
rect 2527 329 2561 363
rect 2527 257 2561 291
rect 2527 189 2561 223
rect 2624 213 2658 247
rect 2721 257 2755 291
rect 2721 189 2755 223
rect 2527 119 2561 153
rect 2624 119 2658 153
rect 2721 119 2755 153
rect 2987 329 3021 363
rect 3084 329 3118 363
rect 3181 329 3215 363
rect 3278 329 3312 363
rect 3375 329 3409 363
rect 2987 257 3021 291
rect 2987 189 3021 223
rect 3084 204 3118 238
rect 3181 257 3215 291
rect 3181 189 3215 223
rect 3279 210 3313 244
rect 2987 119 3021 153
rect 3181 119 3215 153
rect 3278 119 3312 153
rect 3375 119 3409 153
rect 3489 329 3523 363
rect 3489 257 3523 291
rect 3489 189 3523 223
rect 3586 213 3620 247
rect 3683 257 3717 291
rect 3683 189 3717 223
rect 3489 119 3523 153
rect 3586 119 3620 153
rect 3683 119 3717 153
rect 3949 329 3983 363
rect 4046 329 4080 363
rect 4143 329 4177 363
rect 4240 329 4274 363
rect 4337 329 4371 363
rect 3949 257 3983 291
rect 3949 189 3983 223
rect 4046 204 4080 238
rect 4143 257 4177 291
rect 4143 189 4177 223
rect 4241 210 4275 244
rect 3949 119 3983 153
rect 4143 119 4177 153
rect 4240 119 4274 153
rect 4337 119 4371 153
rect 4451 329 4485 363
rect 4451 257 4485 291
rect 4451 189 4485 223
rect 4548 213 4582 247
rect 4645 257 4679 291
rect 4645 189 4679 223
rect 4451 119 4485 153
rect 4548 119 4582 153
rect 4645 119 4679 153
rect 4911 329 4945 363
rect 5008 329 5042 363
rect 5105 329 5139 363
rect 5202 329 5236 363
rect 5299 329 5333 363
rect 4911 257 4945 291
rect 4911 189 4945 223
rect 5008 204 5042 238
rect 5105 257 5139 291
rect 5105 189 5139 223
rect 5203 210 5237 244
rect 4911 119 4945 153
rect 5105 119 5139 153
rect 5202 119 5236 153
rect 5299 119 5333 153
rect 5413 329 5447 363
rect 5413 257 5447 291
rect 5413 189 5447 223
rect 5510 213 5544 247
rect 5607 257 5641 291
rect 5607 189 5641 223
rect 5413 119 5447 153
rect 5510 119 5544 153
rect 5607 119 5641 153
rect 5873 329 5907 363
rect 5970 329 6004 363
rect 6067 329 6101 363
rect 6164 329 6198 363
rect 6261 329 6295 363
rect 5873 257 5907 291
rect 5873 189 5907 223
rect 5970 204 6004 238
rect 6067 257 6101 291
rect 6067 189 6101 223
rect 6165 210 6199 244
rect 5873 119 5907 153
rect 6067 119 6101 153
rect 6164 119 6198 153
rect 6261 119 6295 153
rect 6375 329 6409 363
rect 6375 257 6409 291
rect 6375 189 6409 223
rect 6472 213 6506 247
rect 6569 257 6603 291
rect 6569 189 6603 223
rect 6375 119 6409 153
rect 6472 119 6506 153
rect 6569 119 6603 153
rect 6835 329 6869 363
rect 6932 329 6966 363
rect 7029 329 7063 363
rect 7126 329 7160 363
rect 7223 329 7257 363
rect 6835 257 6869 291
rect 6835 189 6869 223
rect 6932 204 6966 238
rect 7029 257 7063 291
rect 7029 189 7063 223
rect 7127 210 7161 244
rect 6835 119 6869 153
rect 7029 119 7063 153
rect 7126 119 7160 153
rect 7223 119 7257 153
rect 7337 329 7371 363
rect 7337 257 7371 291
rect 7337 189 7371 223
rect 7434 213 7468 247
rect 7531 257 7565 291
rect 7531 189 7565 223
rect 7337 119 7371 153
rect 7434 119 7468 153
rect 7531 119 7565 153
rect 7797 329 7831 363
rect 7894 329 7928 363
rect 7991 329 8025 363
rect 8088 329 8122 363
rect 8185 329 8219 363
rect 7797 257 7831 291
rect 7797 189 7831 223
rect 7894 204 7928 238
rect 7991 257 8025 291
rect 7991 189 8025 223
rect 8089 210 8123 244
rect 7797 119 7831 153
rect 7991 119 8025 153
rect 8088 119 8122 153
rect 8185 119 8219 153
rect 8299 329 8333 363
rect 8299 257 8333 291
rect 8299 189 8333 223
rect 8396 213 8430 247
rect 8493 257 8527 291
rect 8493 189 8527 223
rect 8299 119 8333 153
rect 8396 119 8430 153
rect 8493 119 8527 153
rect 8759 329 8793 363
rect 8856 329 8890 363
rect 8953 329 8987 363
rect 9050 329 9084 363
rect 9147 329 9181 363
rect 8759 257 8793 291
rect 8759 189 8793 223
rect 8856 204 8890 238
rect 8953 257 8987 291
rect 8953 189 8987 223
rect 9051 210 9085 244
rect 8759 119 8793 153
rect 8953 119 8987 153
rect 9050 119 9084 153
rect 9147 119 9181 153
rect 9261 329 9295 363
rect 9261 257 9295 291
rect 9261 189 9295 223
rect 9358 213 9392 247
rect 9455 257 9489 291
rect 9455 189 9489 223
rect 9261 119 9295 153
rect 9358 119 9392 153
rect 9455 119 9489 153
rect 9721 329 9755 363
rect 9818 329 9852 363
rect 9915 329 9949 363
rect 10012 329 10046 363
rect 10109 329 10143 363
rect 9721 257 9755 291
rect 9721 189 9755 223
rect 9818 204 9852 238
rect 9915 257 9949 291
rect 9915 189 9949 223
rect 10013 210 10047 244
rect 9721 119 9755 153
rect 9915 119 9949 153
rect 10012 119 10046 153
rect 10109 119 10143 153
rect 10223 329 10257 363
rect 10223 257 10257 291
rect 10223 189 10257 223
rect 10320 213 10354 247
rect 10417 257 10451 291
rect 10417 189 10451 223
rect 10223 119 10257 153
rect 10320 119 10354 153
rect 10417 119 10451 153
rect 10683 329 10717 363
rect 10780 329 10814 363
rect 10877 329 10911 363
rect 10974 329 11008 363
rect 11071 329 11105 363
rect 10683 257 10717 291
rect 10683 189 10717 223
rect 10780 204 10814 238
rect 10877 257 10911 291
rect 10877 189 10911 223
rect 10975 210 11009 244
rect 10683 119 10717 153
rect 10877 119 10911 153
rect 10974 119 11008 153
rect 11071 119 11105 153
rect 11185 329 11219 363
rect 11185 257 11219 291
rect 11185 189 11219 223
rect 11282 213 11316 247
rect 11379 257 11413 291
rect 11379 189 11413 223
rect 11185 119 11219 153
rect 11282 119 11316 153
rect 11379 119 11413 153
rect 11645 329 11679 363
rect 11742 329 11776 363
rect 11839 329 11873 363
rect 11936 329 11970 363
rect 12033 329 12067 363
rect 11645 257 11679 291
rect 11645 189 11679 223
rect 11742 204 11776 238
rect 11839 257 11873 291
rect 11839 189 11873 223
rect 11937 210 11971 244
rect 11645 119 11679 153
rect 11839 119 11873 153
rect 11936 119 11970 153
rect 12033 119 12067 153
rect 12147 329 12181 363
rect 12147 257 12181 291
rect 12147 189 12181 223
rect 12244 213 12278 247
rect 12341 257 12375 291
rect 12341 189 12375 223
rect 12147 119 12181 153
rect 12244 119 12278 153
rect 12341 119 12375 153
rect 12607 329 12641 363
rect 12704 329 12738 363
rect 12801 329 12835 363
rect 12898 329 12932 363
rect 12995 329 13029 363
rect 12607 257 12641 291
rect 12607 189 12641 223
rect 12704 204 12738 238
rect 12801 257 12835 291
rect 12801 189 12835 223
rect 12899 210 12933 244
rect 12607 119 12641 153
rect 12801 119 12835 153
rect 12898 119 12932 153
rect 12995 119 13029 153
rect 13109 329 13143 363
rect 13109 257 13143 291
rect 13109 189 13143 223
rect 13206 213 13240 247
rect 13303 257 13337 291
rect 13303 189 13337 223
rect 13109 119 13143 153
rect 13206 119 13240 153
rect 13303 119 13337 153
rect 13569 329 13603 363
rect 13666 329 13700 363
rect 13763 329 13797 363
rect 13860 329 13894 363
rect 13957 329 13991 363
rect 13569 257 13603 291
rect 13569 189 13603 223
rect 13666 204 13700 238
rect 13763 257 13797 291
rect 13763 189 13797 223
rect 13861 210 13895 244
rect 13569 119 13603 153
rect 13763 119 13797 153
rect 13860 119 13894 153
rect 13957 119 13991 153
rect 14071 329 14105 363
rect 14071 257 14105 291
rect 14071 189 14105 223
rect 14168 213 14202 247
rect 14265 257 14299 291
rect 14265 189 14299 223
rect 14071 119 14105 153
rect 14168 119 14202 153
rect 14265 119 14299 153
rect 14531 329 14565 363
rect 14628 329 14662 363
rect 14725 329 14759 363
rect 14822 329 14856 363
rect 14919 329 14953 363
rect 14531 257 14565 291
rect 14531 189 14565 223
rect 14628 204 14662 238
rect 14725 257 14759 291
rect 14725 189 14759 223
rect 14823 210 14857 244
rect 14531 119 14565 153
rect 14725 119 14759 153
rect 14822 119 14856 153
rect 14919 119 14953 153
rect 15033 329 15067 363
rect 15033 257 15067 291
rect 15033 189 15067 223
rect 15130 213 15164 247
rect 15227 257 15261 291
rect 15227 189 15261 223
rect 15033 119 15067 153
rect 15130 119 15164 153
rect 15227 119 15261 153
rect 15493 329 15527 363
rect 15590 329 15624 363
rect 15687 329 15721 363
rect 15784 329 15818 363
rect 15881 329 15915 363
rect 15493 257 15527 291
rect 15493 189 15527 223
rect 15590 204 15624 238
rect 15687 257 15721 291
rect 15687 189 15721 223
rect 15785 210 15819 244
rect 15493 119 15527 153
rect 15687 119 15721 153
rect 15784 119 15818 153
rect 15881 119 15915 153
rect 15995 329 16029 363
rect 15995 257 16029 291
rect 15995 189 16029 223
rect 16092 213 16126 247
rect 16189 257 16223 291
rect 16189 189 16223 223
rect 15995 119 16029 153
rect 16092 119 16126 153
rect 16189 119 16223 153
rect 16455 329 16489 363
rect 16552 329 16586 363
rect 16649 329 16683 363
rect 16746 329 16780 363
rect 16843 329 16877 363
rect 16455 257 16489 291
rect 16455 189 16489 223
rect 16552 204 16586 238
rect 16649 257 16683 291
rect 16649 189 16683 223
rect 16747 210 16781 244
rect 16455 119 16489 153
rect 16649 119 16683 153
rect 16746 119 16780 153
rect 16843 119 16877 153
rect 16957 329 16991 363
rect 16957 257 16991 291
rect 16957 189 16991 223
rect 17054 213 17088 247
rect 17151 257 17185 291
rect 17151 189 17185 223
rect 16957 119 16991 153
rect 17054 119 17088 153
rect 17151 119 17185 153
rect 17438 327 17472 361
rect 17535 327 17569 361
rect 17632 327 17666 361
rect 17826 327 17860 361
rect 17438 255 17472 289
rect 17438 187 17472 221
rect 17535 202 17569 236
rect 17632 255 17666 289
rect 17632 187 17666 221
rect 17728 211 17762 245
rect 17826 255 17860 289
rect 17826 187 17860 221
rect 17438 117 17472 151
rect 17632 117 17666 151
rect 17728 117 17762 151
rect 17826 117 17860 151
rect 18104 327 18138 361
rect 18201 327 18235 361
rect 18298 327 18332 361
rect 18492 327 18526 361
rect 18104 255 18138 289
rect 18104 187 18138 221
rect 18201 202 18235 236
rect 18298 255 18332 289
rect 18298 187 18332 221
rect 18395 211 18429 245
rect 18492 255 18526 289
rect 18492 187 18526 221
rect 18104 117 18138 151
rect 18298 117 18332 151
rect 18395 117 18429 151
rect 18492 117 18526 151
rect 18770 327 18804 361
rect 18867 327 18901 361
rect 18964 327 18998 361
rect 18770 255 18804 289
rect 18770 187 18804 221
rect 18867 202 18901 236
rect 18964 255 18998 289
rect 18964 187 18998 221
rect 19061 211 19095 245
rect 19158 255 19192 289
rect 19158 187 19192 221
rect 18770 117 18804 151
rect 18964 117 18998 151
rect 19061 117 19095 151
rect 19158 117 19192 151
<< pdiffc >>
rect 201 1378 235 1412
rect 201 1310 235 1344
rect 201 1242 235 1276
rect 201 1174 235 1208
rect 201 1105 235 1139
rect 289 1378 323 1412
rect 289 1310 323 1344
rect 289 1242 323 1276
rect 289 1174 323 1208
rect 289 1105 323 1139
rect 377 1378 411 1412
rect 377 1310 411 1344
rect 377 1242 411 1276
rect 377 1174 411 1208
rect 465 1378 499 1412
rect 465 1310 499 1344
rect 465 1242 499 1276
rect 465 1174 499 1208
rect 465 1105 499 1139
rect 553 1378 587 1412
rect 553 1310 587 1344
rect 553 1242 587 1276
rect 553 1174 587 1208
rect 641 1378 675 1412
rect 641 1310 675 1344
rect 641 1242 675 1276
rect 641 1174 675 1208
rect 641 1105 675 1139
rect 729 1378 763 1412
rect 729 1310 763 1344
rect 729 1242 763 1276
rect 729 1174 763 1208
rect 1163 1378 1197 1412
rect 1163 1310 1197 1344
rect 1163 1242 1197 1276
rect 1163 1174 1197 1208
rect 1163 1105 1197 1139
rect 1251 1378 1285 1412
rect 1251 1310 1285 1344
rect 1251 1242 1285 1276
rect 1251 1174 1285 1208
rect 1251 1105 1285 1139
rect 1339 1378 1373 1412
rect 1339 1310 1373 1344
rect 1339 1242 1373 1276
rect 1339 1174 1373 1208
rect 1427 1378 1461 1412
rect 1427 1310 1461 1344
rect 1427 1242 1461 1276
rect 1427 1174 1461 1208
rect 1427 1105 1461 1139
rect 1515 1378 1549 1412
rect 1515 1310 1549 1344
rect 1515 1242 1549 1276
rect 1515 1174 1549 1208
rect 1603 1378 1637 1412
rect 1603 1310 1637 1344
rect 1603 1242 1637 1276
rect 1603 1174 1637 1208
rect 1603 1105 1637 1139
rect 1691 1378 1725 1412
rect 1691 1310 1725 1344
rect 1691 1242 1725 1276
rect 1691 1174 1725 1208
rect 2125 1378 2159 1412
rect 2125 1310 2159 1344
rect 2125 1242 2159 1276
rect 2125 1174 2159 1208
rect 2125 1105 2159 1139
rect 2213 1378 2247 1412
rect 2213 1310 2247 1344
rect 2213 1242 2247 1276
rect 2213 1174 2247 1208
rect 2213 1105 2247 1139
rect 2301 1378 2335 1412
rect 2301 1310 2335 1344
rect 2301 1242 2335 1276
rect 2301 1174 2335 1208
rect 2389 1378 2423 1412
rect 2389 1310 2423 1344
rect 2389 1242 2423 1276
rect 2389 1174 2423 1208
rect 2389 1105 2423 1139
rect 2477 1378 2511 1412
rect 2477 1310 2511 1344
rect 2477 1242 2511 1276
rect 2477 1174 2511 1208
rect 2565 1378 2599 1412
rect 2565 1310 2599 1344
rect 2565 1242 2599 1276
rect 2565 1174 2599 1208
rect 2565 1105 2599 1139
rect 2653 1378 2687 1412
rect 2653 1310 2687 1344
rect 2653 1242 2687 1276
rect 2653 1174 2687 1208
rect 3087 1378 3121 1412
rect 3087 1310 3121 1344
rect 3087 1242 3121 1276
rect 3087 1174 3121 1208
rect 3087 1105 3121 1139
rect 3175 1378 3209 1412
rect 3175 1310 3209 1344
rect 3175 1242 3209 1276
rect 3175 1174 3209 1208
rect 3175 1105 3209 1139
rect 3263 1378 3297 1412
rect 3263 1310 3297 1344
rect 3263 1242 3297 1276
rect 3263 1174 3297 1208
rect 3351 1378 3385 1412
rect 3351 1310 3385 1344
rect 3351 1242 3385 1276
rect 3351 1174 3385 1208
rect 3351 1105 3385 1139
rect 3439 1378 3473 1412
rect 3439 1310 3473 1344
rect 3439 1242 3473 1276
rect 3439 1174 3473 1208
rect 3527 1378 3561 1412
rect 3527 1310 3561 1344
rect 3527 1242 3561 1276
rect 3527 1174 3561 1208
rect 3527 1105 3561 1139
rect 3615 1378 3649 1412
rect 3615 1310 3649 1344
rect 3615 1242 3649 1276
rect 3615 1174 3649 1208
rect 4049 1378 4083 1412
rect 4049 1310 4083 1344
rect 4049 1242 4083 1276
rect 4049 1174 4083 1208
rect 4049 1105 4083 1139
rect 4137 1378 4171 1412
rect 4137 1310 4171 1344
rect 4137 1242 4171 1276
rect 4137 1174 4171 1208
rect 4137 1105 4171 1139
rect 4225 1378 4259 1412
rect 4225 1310 4259 1344
rect 4225 1242 4259 1276
rect 4225 1174 4259 1208
rect 4313 1378 4347 1412
rect 4313 1310 4347 1344
rect 4313 1242 4347 1276
rect 4313 1174 4347 1208
rect 4313 1105 4347 1139
rect 4401 1378 4435 1412
rect 4401 1310 4435 1344
rect 4401 1242 4435 1276
rect 4401 1174 4435 1208
rect 4489 1378 4523 1412
rect 4489 1310 4523 1344
rect 4489 1242 4523 1276
rect 4489 1174 4523 1208
rect 4489 1105 4523 1139
rect 4577 1378 4611 1412
rect 4577 1310 4611 1344
rect 4577 1242 4611 1276
rect 4577 1174 4611 1208
rect 5011 1378 5045 1412
rect 5011 1310 5045 1344
rect 5011 1242 5045 1276
rect 5011 1174 5045 1208
rect 5011 1105 5045 1139
rect 5099 1378 5133 1412
rect 5099 1310 5133 1344
rect 5099 1242 5133 1276
rect 5099 1174 5133 1208
rect 5099 1105 5133 1139
rect 5187 1378 5221 1412
rect 5187 1310 5221 1344
rect 5187 1242 5221 1276
rect 5187 1174 5221 1208
rect 5275 1378 5309 1412
rect 5275 1310 5309 1344
rect 5275 1242 5309 1276
rect 5275 1174 5309 1208
rect 5275 1105 5309 1139
rect 5363 1378 5397 1412
rect 5363 1310 5397 1344
rect 5363 1242 5397 1276
rect 5363 1174 5397 1208
rect 5451 1378 5485 1412
rect 5451 1310 5485 1344
rect 5451 1242 5485 1276
rect 5451 1174 5485 1208
rect 5451 1105 5485 1139
rect 5539 1378 5573 1412
rect 5539 1310 5573 1344
rect 5539 1242 5573 1276
rect 5539 1174 5573 1208
rect 5973 1378 6007 1412
rect 5973 1310 6007 1344
rect 5973 1242 6007 1276
rect 5973 1174 6007 1208
rect 5973 1105 6007 1139
rect 6061 1378 6095 1412
rect 6061 1310 6095 1344
rect 6061 1242 6095 1276
rect 6061 1174 6095 1208
rect 6061 1105 6095 1139
rect 6149 1378 6183 1412
rect 6149 1310 6183 1344
rect 6149 1242 6183 1276
rect 6149 1174 6183 1208
rect 6237 1378 6271 1412
rect 6237 1310 6271 1344
rect 6237 1242 6271 1276
rect 6237 1174 6271 1208
rect 6237 1105 6271 1139
rect 6325 1378 6359 1412
rect 6325 1310 6359 1344
rect 6325 1242 6359 1276
rect 6325 1174 6359 1208
rect 6413 1378 6447 1412
rect 6413 1310 6447 1344
rect 6413 1242 6447 1276
rect 6413 1174 6447 1208
rect 6413 1105 6447 1139
rect 6501 1378 6535 1412
rect 6501 1310 6535 1344
rect 6501 1242 6535 1276
rect 6501 1174 6535 1208
rect 6935 1378 6969 1412
rect 6935 1310 6969 1344
rect 6935 1242 6969 1276
rect 6935 1174 6969 1208
rect 6935 1105 6969 1139
rect 7023 1378 7057 1412
rect 7023 1310 7057 1344
rect 7023 1242 7057 1276
rect 7023 1174 7057 1208
rect 7023 1105 7057 1139
rect 7111 1378 7145 1412
rect 7111 1310 7145 1344
rect 7111 1242 7145 1276
rect 7111 1174 7145 1208
rect 7199 1378 7233 1412
rect 7199 1310 7233 1344
rect 7199 1242 7233 1276
rect 7199 1174 7233 1208
rect 7199 1105 7233 1139
rect 7287 1378 7321 1412
rect 7287 1310 7321 1344
rect 7287 1242 7321 1276
rect 7287 1174 7321 1208
rect 7375 1378 7409 1412
rect 7375 1310 7409 1344
rect 7375 1242 7409 1276
rect 7375 1174 7409 1208
rect 7375 1105 7409 1139
rect 7463 1378 7497 1412
rect 7463 1310 7497 1344
rect 7463 1242 7497 1276
rect 7463 1174 7497 1208
rect 7897 1378 7931 1412
rect 7897 1310 7931 1344
rect 7897 1242 7931 1276
rect 7897 1174 7931 1208
rect 7897 1105 7931 1139
rect 7985 1378 8019 1412
rect 7985 1310 8019 1344
rect 7985 1242 8019 1276
rect 7985 1174 8019 1208
rect 7985 1105 8019 1139
rect 8073 1378 8107 1412
rect 8073 1310 8107 1344
rect 8073 1242 8107 1276
rect 8073 1174 8107 1208
rect 8161 1378 8195 1412
rect 8161 1310 8195 1344
rect 8161 1242 8195 1276
rect 8161 1174 8195 1208
rect 8161 1105 8195 1139
rect 8249 1378 8283 1412
rect 8249 1310 8283 1344
rect 8249 1242 8283 1276
rect 8249 1174 8283 1208
rect 8337 1378 8371 1412
rect 8337 1310 8371 1344
rect 8337 1242 8371 1276
rect 8337 1174 8371 1208
rect 8337 1105 8371 1139
rect 8425 1378 8459 1412
rect 8425 1310 8459 1344
rect 8425 1242 8459 1276
rect 8425 1174 8459 1208
rect 8859 1378 8893 1412
rect 8859 1310 8893 1344
rect 8859 1242 8893 1276
rect 8859 1174 8893 1208
rect 8859 1105 8893 1139
rect 8947 1378 8981 1412
rect 8947 1310 8981 1344
rect 8947 1242 8981 1276
rect 8947 1174 8981 1208
rect 8947 1105 8981 1139
rect 9035 1378 9069 1412
rect 9035 1310 9069 1344
rect 9035 1242 9069 1276
rect 9035 1174 9069 1208
rect 9123 1378 9157 1412
rect 9123 1310 9157 1344
rect 9123 1242 9157 1276
rect 9123 1174 9157 1208
rect 9123 1105 9157 1139
rect 9211 1378 9245 1412
rect 9211 1310 9245 1344
rect 9211 1242 9245 1276
rect 9211 1174 9245 1208
rect 9299 1378 9333 1412
rect 9299 1310 9333 1344
rect 9299 1242 9333 1276
rect 9299 1174 9333 1208
rect 9299 1105 9333 1139
rect 9387 1378 9421 1412
rect 9387 1310 9421 1344
rect 9387 1242 9421 1276
rect 9387 1174 9421 1208
rect 9821 1378 9855 1412
rect 9821 1310 9855 1344
rect 9821 1242 9855 1276
rect 9821 1174 9855 1208
rect 9821 1105 9855 1139
rect 9909 1378 9943 1412
rect 9909 1310 9943 1344
rect 9909 1242 9943 1276
rect 9909 1174 9943 1208
rect 9909 1105 9943 1139
rect 9997 1378 10031 1412
rect 9997 1310 10031 1344
rect 9997 1242 10031 1276
rect 9997 1174 10031 1208
rect 10085 1378 10119 1412
rect 10085 1310 10119 1344
rect 10085 1242 10119 1276
rect 10085 1174 10119 1208
rect 10085 1105 10119 1139
rect 10173 1378 10207 1412
rect 10173 1310 10207 1344
rect 10173 1242 10207 1276
rect 10173 1174 10207 1208
rect 10261 1378 10295 1412
rect 10261 1310 10295 1344
rect 10261 1242 10295 1276
rect 10261 1174 10295 1208
rect 10261 1105 10295 1139
rect 10349 1378 10383 1412
rect 10349 1310 10383 1344
rect 10349 1242 10383 1276
rect 10349 1174 10383 1208
rect 10783 1378 10817 1412
rect 10783 1310 10817 1344
rect 10783 1242 10817 1276
rect 10783 1174 10817 1208
rect 10783 1105 10817 1139
rect 10871 1378 10905 1412
rect 10871 1310 10905 1344
rect 10871 1242 10905 1276
rect 10871 1174 10905 1208
rect 10871 1105 10905 1139
rect 10959 1378 10993 1412
rect 10959 1310 10993 1344
rect 10959 1242 10993 1276
rect 10959 1174 10993 1208
rect 11047 1378 11081 1412
rect 11047 1310 11081 1344
rect 11047 1242 11081 1276
rect 11047 1174 11081 1208
rect 11047 1105 11081 1139
rect 11135 1378 11169 1412
rect 11135 1310 11169 1344
rect 11135 1242 11169 1276
rect 11135 1174 11169 1208
rect 11223 1378 11257 1412
rect 11223 1310 11257 1344
rect 11223 1242 11257 1276
rect 11223 1174 11257 1208
rect 11223 1105 11257 1139
rect 11311 1378 11345 1412
rect 11311 1310 11345 1344
rect 11311 1242 11345 1276
rect 11311 1174 11345 1208
rect 11745 1378 11779 1412
rect 11745 1310 11779 1344
rect 11745 1242 11779 1276
rect 11745 1174 11779 1208
rect 11745 1105 11779 1139
rect 11833 1378 11867 1412
rect 11833 1310 11867 1344
rect 11833 1242 11867 1276
rect 11833 1174 11867 1208
rect 11833 1105 11867 1139
rect 11921 1378 11955 1412
rect 11921 1310 11955 1344
rect 11921 1242 11955 1276
rect 11921 1174 11955 1208
rect 12009 1378 12043 1412
rect 12009 1310 12043 1344
rect 12009 1242 12043 1276
rect 12009 1174 12043 1208
rect 12009 1105 12043 1139
rect 12097 1378 12131 1412
rect 12097 1310 12131 1344
rect 12097 1242 12131 1276
rect 12097 1174 12131 1208
rect 12185 1378 12219 1412
rect 12185 1310 12219 1344
rect 12185 1242 12219 1276
rect 12185 1174 12219 1208
rect 12185 1105 12219 1139
rect 12273 1378 12307 1412
rect 12273 1310 12307 1344
rect 12273 1242 12307 1276
rect 12273 1174 12307 1208
rect 12707 1378 12741 1412
rect 12707 1310 12741 1344
rect 12707 1242 12741 1276
rect 12707 1174 12741 1208
rect 12707 1105 12741 1139
rect 12795 1378 12829 1412
rect 12795 1310 12829 1344
rect 12795 1242 12829 1276
rect 12795 1174 12829 1208
rect 12795 1105 12829 1139
rect 12883 1378 12917 1412
rect 12883 1310 12917 1344
rect 12883 1242 12917 1276
rect 12883 1174 12917 1208
rect 12971 1378 13005 1412
rect 12971 1310 13005 1344
rect 12971 1242 13005 1276
rect 12971 1174 13005 1208
rect 12971 1105 13005 1139
rect 13059 1378 13093 1412
rect 13059 1310 13093 1344
rect 13059 1242 13093 1276
rect 13059 1174 13093 1208
rect 13147 1378 13181 1412
rect 13147 1310 13181 1344
rect 13147 1242 13181 1276
rect 13147 1174 13181 1208
rect 13147 1105 13181 1139
rect 13235 1378 13269 1412
rect 13235 1310 13269 1344
rect 13235 1242 13269 1276
rect 13235 1174 13269 1208
rect 13669 1378 13703 1412
rect 13669 1310 13703 1344
rect 13669 1242 13703 1276
rect 13669 1174 13703 1208
rect 13669 1105 13703 1139
rect 13757 1378 13791 1412
rect 13757 1310 13791 1344
rect 13757 1242 13791 1276
rect 13757 1174 13791 1208
rect 13757 1105 13791 1139
rect 13845 1378 13879 1412
rect 13845 1310 13879 1344
rect 13845 1242 13879 1276
rect 13845 1174 13879 1208
rect 13933 1378 13967 1412
rect 13933 1310 13967 1344
rect 13933 1242 13967 1276
rect 13933 1174 13967 1208
rect 13933 1105 13967 1139
rect 14021 1378 14055 1412
rect 14021 1310 14055 1344
rect 14021 1242 14055 1276
rect 14021 1174 14055 1208
rect 14109 1378 14143 1412
rect 14109 1310 14143 1344
rect 14109 1242 14143 1276
rect 14109 1174 14143 1208
rect 14109 1105 14143 1139
rect 14197 1378 14231 1412
rect 14197 1310 14231 1344
rect 14197 1242 14231 1276
rect 14197 1174 14231 1208
rect 14631 1378 14665 1412
rect 14631 1310 14665 1344
rect 14631 1242 14665 1276
rect 14631 1174 14665 1208
rect 14631 1105 14665 1139
rect 14719 1378 14753 1412
rect 14719 1310 14753 1344
rect 14719 1242 14753 1276
rect 14719 1174 14753 1208
rect 14719 1105 14753 1139
rect 14807 1378 14841 1412
rect 14807 1310 14841 1344
rect 14807 1242 14841 1276
rect 14807 1174 14841 1208
rect 14895 1378 14929 1412
rect 14895 1310 14929 1344
rect 14895 1242 14929 1276
rect 14895 1174 14929 1208
rect 14895 1105 14929 1139
rect 14983 1378 15017 1412
rect 14983 1310 15017 1344
rect 14983 1242 15017 1276
rect 14983 1174 15017 1208
rect 15071 1378 15105 1412
rect 15071 1310 15105 1344
rect 15071 1242 15105 1276
rect 15071 1174 15105 1208
rect 15071 1105 15105 1139
rect 15159 1378 15193 1412
rect 15159 1310 15193 1344
rect 15159 1242 15193 1276
rect 15159 1174 15193 1208
rect 15593 1378 15627 1412
rect 15593 1310 15627 1344
rect 15593 1242 15627 1276
rect 15593 1174 15627 1208
rect 15593 1105 15627 1139
rect 15681 1378 15715 1412
rect 15681 1310 15715 1344
rect 15681 1242 15715 1276
rect 15681 1174 15715 1208
rect 15681 1105 15715 1139
rect 15769 1378 15803 1412
rect 15769 1310 15803 1344
rect 15769 1242 15803 1276
rect 15769 1174 15803 1208
rect 15857 1378 15891 1412
rect 15857 1310 15891 1344
rect 15857 1242 15891 1276
rect 15857 1174 15891 1208
rect 15857 1105 15891 1139
rect 15945 1378 15979 1412
rect 15945 1310 15979 1344
rect 15945 1242 15979 1276
rect 15945 1174 15979 1208
rect 16033 1378 16067 1412
rect 16033 1310 16067 1344
rect 16033 1242 16067 1276
rect 16033 1174 16067 1208
rect 16033 1105 16067 1139
rect 16121 1378 16155 1412
rect 16121 1310 16155 1344
rect 16121 1242 16155 1276
rect 16121 1174 16155 1208
rect 16555 1378 16589 1412
rect 16555 1310 16589 1344
rect 16555 1242 16589 1276
rect 16555 1174 16589 1208
rect 16555 1105 16589 1139
rect 16643 1378 16677 1412
rect 16643 1310 16677 1344
rect 16643 1242 16677 1276
rect 16643 1174 16677 1208
rect 16643 1105 16677 1139
rect 16731 1378 16765 1412
rect 16731 1310 16765 1344
rect 16731 1242 16765 1276
rect 16731 1174 16765 1208
rect 16819 1378 16853 1412
rect 16819 1310 16853 1344
rect 16819 1242 16853 1276
rect 16819 1174 16853 1208
rect 16819 1105 16853 1139
rect 16907 1378 16941 1412
rect 16907 1310 16941 1344
rect 16907 1242 16941 1276
rect 16907 1174 16941 1208
rect 16995 1378 17029 1412
rect 16995 1310 17029 1344
rect 16995 1242 17029 1276
rect 16995 1174 17029 1208
rect 16995 1105 17029 1139
rect 17083 1378 17117 1412
rect 17083 1310 17117 1344
rect 17083 1242 17117 1276
rect 17083 1174 17117 1208
rect 17457 1377 17491 1411
rect 17457 1309 17491 1343
rect 17457 1241 17491 1275
rect 17457 1173 17491 1207
rect 17457 1105 17491 1139
rect 17545 1377 17579 1411
rect 17545 1309 17579 1343
rect 17545 1241 17579 1275
rect 17545 1173 17579 1207
rect 17545 1105 17579 1139
rect 17633 1377 17667 1411
rect 17633 1309 17667 1343
rect 17633 1241 17667 1275
rect 17633 1173 17667 1207
rect 17721 1377 17755 1411
rect 17721 1309 17755 1343
rect 17721 1241 17755 1275
rect 17721 1173 17755 1207
rect 17809 1377 17843 1411
rect 17809 1309 17843 1343
rect 17809 1241 17843 1275
rect 17809 1173 17843 1207
rect 17809 1105 17843 1139
rect 18121 1377 18155 1411
rect 18121 1309 18155 1343
rect 18121 1241 18155 1275
rect 18121 1173 18155 1207
rect 18209 1309 18243 1343
rect 18209 1241 18243 1275
rect 18209 1173 18243 1207
rect 18209 1105 18243 1139
rect 18297 1377 18331 1411
rect 18297 1309 18331 1343
rect 18297 1241 18331 1275
rect 18297 1173 18331 1207
rect 18385 1309 18419 1343
rect 18385 1241 18419 1275
rect 18385 1173 18419 1207
rect 18473 1377 18507 1411
rect 18473 1309 18507 1343
rect 18473 1241 18507 1275
rect 18473 1173 18507 1207
rect 18789 1377 18823 1411
rect 18789 1309 18823 1343
rect 18789 1241 18823 1275
rect 18789 1173 18823 1207
rect 18877 1309 18911 1343
rect 18877 1241 18911 1275
rect 18877 1173 18911 1207
rect 18877 1105 18911 1139
rect 18965 1377 18999 1411
rect 18965 1309 18999 1343
rect 18965 1241 18999 1275
rect 18965 1173 18999 1207
rect 19053 1309 19087 1343
rect 19053 1241 19087 1275
rect 19053 1173 19087 1207
rect 19053 1105 19087 1139
rect 19141 1377 19175 1411
rect 19141 1309 19175 1343
rect 19141 1241 19175 1275
rect 19141 1173 19175 1207
<< psubdiff >>
rect -31 546 19345 572
rect -31 512 -17 546
rect 17 512 945 546
rect 979 512 1907 546
rect 1941 512 2869 546
rect 2903 512 3831 546
rect 3865 512 4793 546
rect 4827 512 5755 546
rect 5789 512 6717 546
rect 6751 512 7679 546
rect 7713 512 8641 546
rect 8675 512 9603 546
rect 9637 512 10565 546
rect 10599 512 11527 546
rect 11561 512 12489 546
rect 12523 512 13451 546
rect 13485 512 14413 546
rect 14447 512 15375 546
rect 15409 512 16337 546
rect 16371 512 17299 546
rect 17333 512 17965 546
rect 17999 512 18631 546
rect 18665 512 19297 546
rect 19331 512 19345 546
rect -31 510 19345 512
rect -31 474 31 510
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect -31 368 -17 402
rect 17 368 31 402
rect 931 474 993 510
rect 931 440 945 474
rect 979 440 993 474
rect 931 402 993 440
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect 931 368 945 402
rect 979 368 993 402
rect 1893 474 1955 510
rect 1893 440 1907 474
rect 1941 440 1955 474
rect 1893 402 1955 440
rect 931 330 993 368
rect 931 296 945 330
rect 979 296 993 330
rect 931 258 993 296
rect 931 224 945 258
rect 979 224 993 258
rect 931 186 993 224
rect 931 152 945 186
rect 979 152 993 186
rect 931 114 993 152
rect -31 47 31 80
rect 931 80 945 114
rect 979 80 993 114
rect 1893 368 1907 402
rect 1941 368 1955 402
rect 2855 474 2917 510
rect 2855 440 2869 474
rect 2903 440 2917 474
rect 2855 402 2917 440
rect 1893 330 1955 368
rect 1893 296 1907 330
rect 1941 296 1955 330
rect 1893 258 1955 296
rect 1893 224 1907 258
rect 1941 224 1955 258
rect 1893 186 1955 224
rect 1893 152 1907 186
rect 1941 152 1955 186
rect 1893 114 1955 152
rect 931 47 993 80
rect 1893 80 1907 114
rect 1941 80 1955 114
rect 2855 368 2869 402
rect 2903 368 2917 402
rect 3817 474 3879 510
rect 3817 440 3831 474
rect 3865 440 3879 474
rect 3817 402 3879 440
rect 2855 330 2917 368
rect 2855 296 2869 330
rect 2903 296 2917 330
rect 2855 258 2917 296
rect 2855 224 2869 258
rect 2903 224 2917 258
rect 2855 186 2917 224
rect 2855 152 2869 186
rect 2903 152 2917 186
rect 2855 114 2917 152
rect 1893 47 1955 80
rect 2855 80 2869 114
rect 2903 80 2917 114
rect 3817 368 3831 402
rect 3865 368 3879 402
rect 4779 474 4841 510
rect 4779 440 4793 474
rect 4827 440 4841 474
rect 4779 402 4841 440
rect 3817 330 3879 368
rect 3817 296 3831 330
rect 3865 296 3879 330
rect 3817 258 3879 296
rect 3817 224 3831 258
rect 3865 224 3879 258
rect 3817 186 3879 224
rect 3817 152 3831 186
rect 3865 152 3879 186
rect 3817 114 3879 152
rect 2855 47 2917 80
rect 3817 80 3831 114
rect 3865 80 3879 114
rect 4779 368 4793 402
rect 4827 368 4841 402
rect 5741 474 5803 510
rect 5741 440 5755 474
rect 5789 440 5803 474
rect 5741 402 5803 440
rect 4779 330 4841 368
rect 4779 296 4793 330
rect 4827 296 4841 330
rect 4779 258 4841 296
rect 4779 224 4793 258
rect 4827 224 4841 258
rect 4779 186 4841 224
rect 4779 152 4793 186
rect 4827 152 4841 186
rect 4779 114 4841 152
rect 3817 47 3879 80
rect 4779 80 4793 114
rect 4827 80 4841 114
rect 5741 368 5755 402
rect 5789 368 5803 402
rect 6703 474 6765 510
rect 6703 440 6717 474
rect 6751 440 6765 474
rect 6703 402 6765 440
rect 5741 330 5803 368
rect 5741 296 5755 330
rect 5789 296 5803 330
rect 5741 258 5803 296
rect 5741 224 5755 258
rect 5789 224 5803 258
rect 5741 186 5803 224
rect 5741 152 5755 186
rect 5789 152 5803 186
rect 5741 114 5803 152
rect 4779 47 4841 80
rect 5741 80 5755 114
rect 5789 80 5803 114
rect 6703 368 6717 402
rect 6751 368 6765 402
rect 7665 474 7727 510
rect 7665 440 7679 474
rect 7713 440 7727 474
rect 7665 402 7727 440
rect 6703 330 6765 368
rect 6703 296 6717 330
rect 6751 296 6765 330
rect 6703 258 6765 296
rect 6703 224 6717 258
rect 6751 224 6765 258
rect 6703 186 6765 224
rect 6703 152 6717 186
rect 6751 152 6765 186
rect 6703 114 6765 152
rect 5741 47 5803 80
rect 6703 80 6717 114
rect 6751 80 6765 114
rect 7665 368 7679 402
rect 7713 368 7727 402
rect 8627 474 8689 510
rect 8627 440 8641 474
rect 8675 440 8689 474
rect 8627 402 8689 440
rect 7665 330 7727 368
rect 7665 296 7679 330
rect 7713 296 7727 330
rect 7665 258 7727 296
rect 7665 224 7679 258
rect 7713 224 7727 258
rect 7665 186 7727 224
rect 7665 152 7679 186
rect 7713 152 7727 186
rect 7665 114 7727 152
rect 6703 47 6765 80
rect 7665 80 7679 114
rect 7713 80 7727 114
rect 8627 368 8641 402
rect 8675 368 8689 402
rect 9589 474 9651 510
rect 9589 440 9603 474
rect 9637 440 9651 474
rect 9589 402 9651 440
rect 8627 330 8689 368
rect 8627 296 8641 330
rect 8675 296 8689 330
rect 8627 258 8689 296
rect 8627 224 8641 258
rect 8675 224 8689 258
rect 8627 186 8689 224
rect 8627 152 8641 186
rect 8675 152 8689 186
rect 8627 114 8689 152
rect 7665 47 7727 80
rect 8627 80 8641 114
rect 8675 80 8689 114
rect 9589 368 9603 402
rect 9637 368 9651 402
rect 10551 474 10613 510
rect 10551 440 10565 474
rect 10599 440 10613 474
rect 10551 402 10613 440
rect 9589 330 9651 368
rect 9589 296 9603 330
rect 9637 296 9651 330
rect 9589 258 9651 296
rect 9589 224 9603 258
rect 9637 224 9651 258
rect 9589 186 9651 224
rect 9589 152 9603 186
rect 9637 152 9651 186
rect 9589 114 9651 152
rect 8627 47 8689 80
rect 9589 80 9603 114
rect 9637 80 9651 114
rect 10551 368 10565 402
rect 10599 368 10613 402
rect 11513 474 11575 510
rect 11513 440 11527 474
rect 11561 440 11575 474
rect 11513 402 11575 440
rect 10551 330 10613 368
rect 10551 296 10565 330
rect 10599 296 10613 330
rect 10551 258 10613 296
rect 10551 224 10565 258
rect 10599 224 10613 258
rect 10551 186 10613 224
rect 10551 152 10565 186
rect 10599 152 10613 186
rect 10551 114 10613 152
rect 9589 47 9651 80
rect 10551 80 10565 114
rect 10599 80 10613 114
rect 11513 368 11527 402
rect 11561 368 11575 402
rect 12475 474 12537 510
rect 12475 440 12489 474
rect 12523 440 12537 474
rect 12475 402 12537 440
rect 11513 330 11575 368
rect 11513 296 11527 330
rect 11561 296 11575 330
rect 11513 258 11575 296
rect 11513 224 11527 258
rect 11561 224 11575 258
rect 11513 186 11575 224
rect 11513 152 11527 186
rect 11561 152 11575 186
rect 11513 114 11575 152
rect 10551 47 10613 80
rect 11513 80 11527 114
rect 11561 80 11575 114
rect 12475 368 12489 402
rect 12523 368 12537 402
rect 13437 474 13499 510
rect 13437 440 13451 474
rect 13485 440 13499 474
rect 13437 402 13499 440
rect 12475 330 12537 368
rect 12475 296 12489 330
rect 12523 296 12537 330
rect 12475 258 12537 296
rect 12475 224 12489 258
rect 12523 224 12537 258
rect 12475 186 12537 224
rect 12475 152 12489 186
rect 12523 152 12537 186
rect 12475 114 12537 152
rect 11513 47 11575 80
rect 12475 80 12489 114
rect 12523 80 12537 114
rect 13437 368 13451 402
rect 13485 368 13499 402
rect 14399 474 14461 510
rect 14399 440 14413 474
rect 14447 440 14461 474
rect 14399 402 14461 440
rect 13437 330 13499 368
rect 13437 296 13451 330
rect 13485 296 13499 330
rect 13437 258 13499 296
rect 13437 224 13451 258
rect 13485 224 13499 258
rect 13437 186 13499 224
rect 13437 152 13451 186
rect 13485 152 13499 186
rect 13437 114 13499 152
rect 12475 47 12537 80
rect 13437 80 13451 114
rect 13485 80 13499 114
rect 14399 368 14413 402
rect 14447 368 14461 402
rect 15361 474 15423 510
rect 15361 440 15375 474
rect 15409 440 15423 474
rect 15361 402 15423 440
rect 14399 330 14461 368
rect 14399 296 14413 330
rect 14447 296 14461 330
rect 14399 258 14461 296
rect 14399 224 14413 258
rect 14447 224 14461 258
rect 14399 186 14461 224
rect 14399 152 14413 186
rect 14447 152 14461 186
rect 14399 114 14461 152
rect 13437 47 13499 80
rect 14399 80 14413 114
rect 14447 80 14461 114
rect 15361 368 15375 402
rect 15409 368 15423 402
rect 16323 474 16385 510
rect 16323 440 16337 474
rect 16371 440 16385 474
rect 16323 402 16385 440
rect 15361 330 15423 368
rect 15361 296 15375 330
rect 15409 296 15423 330
rect 15361 258 15423 296
rect 15361 224 15375 258
rect 15409 224 15423 258
rect 15361 186 15423 224
rect 15361 152 15375 186
rect 15409 152 15423 186
rect 15361 114 15423 152
rect 14399 47 14461 80
rect 15361 80 15375 114
rect 15409 80 15423 114
rect 16323 368 16337 402
rect 16371 368 16385 402
rect 17285 474 17347 510
rect 17285 440 17299 474
rect 17333 440 17347 474
rect 17285 402 17347 440
rect 17951 474 18013 510
rect 17951 440 17965 474
rect 17999 440 18013 474
rect 16323 330 16385 368
rect 16323 296 16337 330
rect 16371 296 16385 330
rect 16323 258 16385 296
rect 16323 224 16337 258
rect 16371 224 16385 258
rect 16323 186 16385 224
rect 16323 152 16337 186
rect 16371 152 16385 186
rect 16323 114 16385 152
rect 15361 47 15423 80
rect 16323 80 16337 114
rect 16371 80 16385 114
rect 17285 368 17299 402
rect 17333 368 17347 402
rect 17951 402 18013 440
rect 17285 330 17347 368
rect 17285 296 17299 330
rect 17333 296 17347 330
rect 17285 258 17347 296
rect 17285 224 17299 258
rect 17333 224 17347 258
rect 17285 186 17347 224
rect 17285 152 17299 186
rect 17333 152 17347 186
rect 17285 114 17347 152
rect 16323 47 16385 80
rect 17285 80 17299 114
rect 17333 80 17347 114
rect 17951 368 17965 402
rect 17999 368 18013 402
rect 18617 474 18679 510
rect 18617 440 18631 474
rect 18665 440 18679 474
rect 18617 402 18679 440
rect 19283 474 19345 510
rect 19283 440 19297 474
rect 19331 440 19345 474
rect 17951 330 18013 368
rect 17951 296 17965 330
rect 17999 296 18013 330
rect 17951 258 18013 296
rect 17951 224 17965 258
rect 17999 224 18013 258
rect 17951 186 18013 224
rect 17951 152 17965 186
rect 17999 152 18013 186
rect 17951 114 18013 152
rect 17285 47 17347 80
rect 17951 80 17965 114
rect 17999 80 18013 114
rect 18617 368 18631 402
rect 18665 368 18679 402
rect 19283 402 19345 440
rect 18617 330 18679 368
rect 18617 296 18631 330
rect 18665 296 18679 330
rect 18617 258 18679 296
rect 18617 224 18631 258
rect 18665 224 18679 258
rect 18617 186 18679 224
rect 18617 152 18631 186
rect 18665 152 18679 186
rect 18617 114 18679 152
rect 17951 47 18013 80
rect 18617 80 18631 114
rect 18665 80 18679 114
rect 19283 368 19297 402
rect 19331 368 19345 402
rect 19283 330 19345 368
rect 19283 296 19297 330
rect 19331 296 19345 330
rect 19283 258 19345 296
rect 19283 224 19297 258
rect 19331 224 19345 258
rect 19283 186 19345 224
rect 19283 152 19297 186
rect 19331 152 19345 186
rect 19283 114 19345 152
rect 18617 47 18679 80
rect 19283 80 19297 114
rect 19331 80 19345 114
rect 19283 47 19345 80
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 343 47
rect 377 13 415 47
rect 449 13 513 47
rect 547 13 585 47
rect 619 13 657 47
rect 691 13 729 47
rect 763 13 801 47
rect 835 13 873 47
rect 907 13 1017 47
rect 1051 13 1089 47
rect 1123 13 1161 47
rect 1195 13 1233 47
rect 1267 13 1305 47
rect 1339 13 1377 47
rect 1411 13 1475 47
rect 1509 13 1547 47
rect 1581 13 1619 47
rect 1653 13 1691 47
rect 1725 13 1763 47
rect 1797 13 1835 47
rect 1869 13 1979 47
rect 2013 13 2051 47
rect 2085 13 2123 47
rect 2157 13 2195 47
rect 2229 13 2267 47
rect 2301 13 2339 47
rect 2373 13 2437 47
rect 2471 13 2509 47
rect 2543 13 2581 47
rect 2615 13 2653 47
rect 2687 13 2725 47
rect 2759 13 2797 47
rect 2831 13 2941 47
rect 2975 13 3013 47
rect 3047 13 3085 47
rect 3119 13 3157 47
rect 3191 13 3229 47
rect 3263 13 3301 47
rect 3335 13 3399 47
rect 3433 13 3471 47
rect 3505 13 3543 47
rect 3577 13 3615 47
rect 3649 13 3687 47
rect 3721 13 3759 47
rect 3793 13 3903 47
rect 3937 13 3975 47
rect 4009 13 4047 47
rect 4081 13 4119 47
rect 4153 13 4191 47
rect 4225 13 4263 47
rect 4297 13 4361 47
rect 4395 13 4433 47
rect 4467 13 4505 47
rect 4539 13 4577 47
rect 4611 13 4649 47
rect 4683 13 4721 47
rect 4755 13 4865 47
rect 4899 13 4937 47
rect 4971 13 5009 47
rect 5043 13 5081 47
rect 5115 13 5153 47
rect 5187 13 5225 47
rect 5259 13 5323 47
rect 5357 13 5395 47
rect 5429 13 5467 47
rect 5501 13 5539 47
rect 5573 13 5611 47
rect 5645 13 5683 47
rect 5717 13 5827 47
rect 5861 13 5899 47
rect 5933 13 5971 47
rect 6005 13 6043 47
rect 6077 13 6115 47
rect 6149 13 6187 47
rect 6221 13 6285 47
rect 6319 13 6357 47
rect 6391 13 6429 47
rect 6463 13 6501 47
rect 6535 13 6573 47
rect 6607 13 6645 47
rect 6679 13 6789 47
rect 6823 13 6861 47
rect 6895 13 6933 47
rect 6967 13 7005 47
rect 7039 13 7077 47
rect 7111 13 7149 47
rect 7183 13 7247 47
rect 7281 13 7319 47
rect 7353 13 7391 47
rect 7425 13 7463 47
rect 7497 13 7535 47
rect 7569 13 7607 47
rect 7641 13 7751 47
rect 7785 13 7823 47
rect 7857 13 7895 47
rect 7929 13 7967 47
rect 8001 13 8039 47
rect 8073 13 8111 47
rect 8145 13 8209 47
rect 8243 13 8281 47
rect 8315 13 8353 47
rect 8387 13 8425 47
rect 8459 13 8497 47
rect 8531 13 8569 47
rect 8603 13 8713 47
rect 8747 13 8785 47
rect 8819 13 8857 47
rect 8891 13 8929 47
rect 8963 13 9001 47
rect 9035 13 9073 47
rect 9107 13 9171 47
rect 9205 13 9243 47
rect 9277 13 9315 47
rect 9349 13 9387 47
rect 9421 13 9459 47
rect 9493 13 9531 47
rect 9565 13 9675 47
rect 9709 13 9747 47
rect 9781 13 9819 47
rect 9853 13 9891 47
rect 9925 13 9963 47
rect 9997 13 10035 47
rect 10069 13 10133 47
rect 10167 13 10205 47
rect 10239 13 10277 47
rect 10311 13 10349 47
rect 10383 13 10421 47
rect 10455 13 10493 47
rect 10527 13 10637 47
rect 10671 13 10709 47
rect 10743 13 10781 47
rect 10815 13 10853 47
rect 10887 13 10925 47
rect 10959 13 10997 47
rect 11031 13 11095 47
rect 11129 13 11167 47
rect 11201 13 11239 47
rect 11273 13 11311 47
rect 11345 13 11383 47
rect 11417 13 11455 47
rect 11489 13 11599 47
rect 11633 13 11671 47
rect 11705 13 11743 47
rect 11777 13 11815 47
rect 11849 13 11887 47
rect 11921 13 11959 47
rect 11993 13 12057 47
rect 12091 13 12129 47
rect 12163 13 12201 47
rect 12235 13 12273 47
rect 12307 13 12345 47
rect 12379 13 12417 47
rect 12451 13 12561 47
rect 12595 13 12633 47
rect 12667 13 12705 47
rect 12739 13 12777 47
rect 12811 13 12849 47
rect 12883 13 12921 47
rect 12955 13 13019 47
rect 13053 13 13091 47
rect 13125 13 13163 47
rect 13197 13 13235 47
rect 13269 13 13307 47
rect 13341 13 13379 47
rect 13413 13 13523 47
rect 13557 13 13595 47
rect 13629 13 13667 47
rect 13701 13 13739 47
rect 13773 13 13811 47
rect 13845 13 13883 47
rect 13917 13 13981 47
rect 14015 13 14053 47
rect 14087 13 14125 47
rect 14159 13 14197 47
rect 14231 13 14269 47
rect 14303 13 14341 47
rect 14375 13 14485 47
rect 14519 13 14557 47
rect 14591 13 14629 47
rect 14663 13 14701 47
rect 14735 13 14773 47
rect 14807 13 14845 47
rect 14879 13 14943 47
rect 14977 13 15015 47
rect 15049 13 15087 47
rect 15121 13 15159 47
rect 15193 13 15231 47
rect 15265 13 15303 47
rect 15337 13 15447 47
rect 15481 13 15519 47
rect 15553 13 15591 47
rect 15625 13 15663 47
rect 15697 13 15735 47
rect 15769 13 15807 47
rect 15841 13 15905 47
rect 15939 13 15977 47
rect 16011 13 16049 47
rect 16083 13 16121 47
rect 16155 13 16193 47
rect 16227 13 16265 47
rect 16299 13 16409 47
rect 16443 13 16481 47
rect 16515 13 16553 47
rect 16587 13 16625 47
rect 16659 13 16697 47
rect 16731 13 16769 47
rect 16803 13 16867 47
rect 16901 13 16939 47
rect 16973 13 17011 47
rect 17045 13 17083 47
rect 17117 13 17155 47
rect 17189 13 17227 47
rect 17261 13 17371 47
rect 17405 13 17443 47
rect 17477 13 17515 47
rect 17549 13 17587 47
rect 17621 13 17677 47
rect 17711 13 17749 47
rect 17783 13 17821 47
rect 17855 13 17893 47
rect 17927 13 18037 47
rect 18071 13 18109 47
rect 18143 13 18181 47
rect 18215 13 18253 47
rect 18287 13 18343 47
rect 18377 13 18415 47
rect 18449 13 18487 47
rect 18521 13 18559 47
rect 18593 13 18703 47
rect 18737 13 18775 47
rect 18809 13 18847 47
rect 18881 13 18919 47
rect 18953 13 19009 47
rect 19043 13 19081 47
rect 19115 13 19153 47
rect 19187 13 19225 47
rect 19259 13 19345 47
rect -31 11 31 13
rect 931 11 993 13
rect 1893 11 1955 13
rect 2855 11 2917 13
rect 3817 11 3879 13
rect 4779 11 4841 13
rect 5741 11 5803 13
rect 6703 11 6765 13
rect 7665 11 7727 13
rect 8627 11 8689 13
rect 9589 11 9651 13
rect 10551 11 10613 13
rect 11513 11 11575 13
rect 12475 11 12537 13
rect 13437 11 13499 13
rect 14399 11 14461 13
rect 15361 11 15423 13
rect 16323 11 16385 13
rect 17285 11 17347 13
rect 17951 11 18013 13
rect 18617 11 18679 13
rect 19283 11 19345 13
<< nsubdiff >>
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 343 1539
rect 377 1505 415 1539
rect 449 1505 513 1539
rect 547 1505 585 1539
rect 619 1505 657 1539
rect 691 1505 729 1539
rect 763 1505 801 1539
rect 835 1505 873 1539
rect 907 1505 1017 1539
rect 1051 1505 1089 1539
rect 1123 1505 1161 1539
rect 1195 1505 1233 1539
rect 1267 1505 1305 1539
rect 1339 1505 1377 1539
rect 1411 1505 1475 1539
rect 1509 1505 1547 1539
rect 1581 1505 1619 1539
rect 1653 1505 1691 1539
rect 1725 1505 1763 1539
rect 1797 1505 1835 1539
rect 1869 1505 1979 1539
rect 2013 1505 2051 1539
rect 2085 1505 2123 1539
rect 2157 1505 2195 1539
rect 2229 1505 2267 1539
rect 2301 1505 2339 1539
rect 2373 1505 2437 1539
rect 2471 1505 2509 1539
rect 2543 1505 2581 1539
rect 2615 1505 2653 1539
rect 2687 1505 2725 1539
rect 2759 1505 2797 1539
rect 2831 1505 2941 1539
rect 2975 1505 3013 1539
rect 3047 1505 3085 1539
rect 3119 1505 3157 1539
rect 3191 1505 3229 1539
rect 3263 1505 3301 1539
rect 3335 1505 3399 1539
rect 3433 1505 3471 1539
rect 3505 1505 3543 1539
rect 3577 1505 3615 1539
rect 3649 1505 3687 1539
rect 3721 1505 3759 1539
rect 3793 1505 3903 1539
rect 3937 1505 3975 1539
rect 4009 1505 4047 1539
rect 4081 1505 4119 1539
rect 4153 1505 4191 1539
rect 4225 1505 4263 1539
rect 4297 1505 4361 1539
rect 4395 1505 4433 1539
rect 4467 1505 4505 1539
rect 4539 1505 4577 1539
rect 4611 1505 4649 1539
rect 4683 1505 4721 1539
rect 4755 1505 4865 1539
rect 4899 1505 4937 1539
rect 4971 1505 5009 1539
rect 5043 1505 5081 1539
rect 5115 1505 5153 1539
rect 5187 1505 5225 1539
rect 5259 1505 5323 1539
rect 5357 1505 5395 1539
rect 5429 1505 5467 1539
rect 5501 1505 5539 1539
rect 5573 1505 5611 1539
rect 5645 1505 5683 1539
rect 5717 1505 5827 1539
rect 5861 1505 5899 1539
rect 5933 1505 5971 1539
rect 6005 1505 6043 1539
rect 6077 1505 6115 1539
rect 6149 1505 6187 1539
rect 6221 1505 6285 1539
rect 6319 1505 6357 1539
rect 6391 1505 6429 1539
rect 6463 1505 6501 1539
rect 6535 1505 6573 1539
rect 6607 1505 6645 1539
rect 6679 1505 6789 1539
rect 6823 1505 6861 1539
rect 6895 1505 6933 1539
rect 6967 1505 7005 1539
rect 7039 1505 7077 1539
rect 7111 1505 7149 1539
rect 7183 1505 7247 1539
rect 7281 1505 7319 1539
rect 7353 1505 7391 1539
rect 7425 1505 7463 1539
rect 7497 1505 7535 1539
rect 7569 1505 7607 1539
rect 7641 1505 7751 1539
rect 7785 1505 7823 1539
rect 7857 1505 7895 1539
rect 7929 1505 7967 1539
rect 8001 1505 8039 1539
rect 8073 1505 8111 1539
rect 8145 1505 8209 1539
rect 8243 1505 8281 1539
rect 8315 1505 8353 1539
rect 8387 1505 8425 1539
rect 8459 1505 8497 1539
rect 8531 1505 8569 1539
rect 8603 1505 8713 1539
rect 8747 1505 8785 1539
rect 8819 1505 8857 1539
rect 8891 1505 8929 1539
rect 8963 1505 9001 1539
rect 9035 1505 9073 1539
rect 9107 1505 9171 1539
rect 9205 1505 9243 1539
rect 9277 1505 9315 1539
rect 9349 1505 9387 1539
rect 9421 1505 9459 1539
rect 9493 1505 9531 1539
rect 9565 1505 9675 1539
rect 9709 1505 9747 1539
rect 9781 1505 9819 1539
rect 9853 1505 9891 1539
rect 9925 1505 9963 1539
rect 9997 1505 10035 1539
rect 10069 1505 10133 1539
rect 10167 1505 10205 1539
rect 10239 1505 10277 1539
rect 10311 1505 10349 1539
rect 10383 1505 10421 1539
rect 10455 1505 10493 1539
rect 10527 1505 10637 1539
rect 10671 1505 10709 1539
rect 10743 1505 10781 1539
rect 10815 1505 10853 1539
rect 10887 1505 10925 1539
rect 10959 1505 10997 1539
rect 11031 1505 11095 1539
rect 11129 1505 11167 1539
rect 11201 1505 11239 1539
rect 11273 1505 11311 1539
rect 11345 1505 11383 1539
rect 11417 1505 11455 1539
rect 11489 1505 11599 1539
rect 11633 1505 11671 1539
rect 11705 1505 11743 1539
rect 11777 1505 11815 1539
rect 11849 1505 11887 1539
rect 11921 1505 11959 1539
rect 11993 1505 12057 1539
rect 12091 1505 12129 1539
rect 12163 1505 12201 1539
rect 12235 1505 12273 1539
rect 12307 1505 12345 1539
rect 12379 1505 12417 1539
rect 12451 1505 12561 1539
rect 12595 1505 12633 1539
rect 12667 1505 12705 1539
rect 12739 1505 12777 1539
rect 12811 1505 12849 1539
rect 12883 1505 12921 1539
rect 12955 1505 13019 1539
rect 13053 1505 13091 1539
rect 13125 1505 13163 1539
rect 13197 1505 13235 1539
rect 13269 1505 13307 1539
rect 13341 1505 13379 1539
rect 13413 1505 13523 1539
rect 13557 1505 13595 1539
rect 13629 1505 13667 1539
rect 13701 1505 13739 1539
rect 13773 1505 13811 1539
rect 13845 1505 13883 1539
rect 13917 1505 13981 1539
rect 14015 1505 14053 1539
rect 14087 1505 14125 1539
rect 14159 1505 14197 1539
rect 14231 1505 14269 1539
rect 14303 1505 14341 1539
rect 14375 1505 14485 1539
rect 14519 1505 14557 1539
rect 14591 1505 14629 1539
rect 14663 1505 14701 1539
rect 14735 1505 14773 1539
rect 14807 1505 14845 1539
rect 14879 1505 14943 1539
rect 14977 1505 15015 1539
rect 15049 1505 15087 1539
rect 15121 1505 15159 1539
rect 15193 1505 15231 1539
rect 15265 1505 15303 1539
rect 15337 1505 15447 1539
rect 15481 1505 15519 1539
rect 15553 1505 15591 1539
rect 15625 1505 15663 1539
rect 15697 1505 15735 1539
rect 15769 1505 15807 1539
rect 15841 1505 15905 1539
rect 15939 1505 15977 1539
rect 16011 1505 16049 1539
rect 16083 1505 16121 1539
rect 16155 1505 16193 1539
rect 16227 1505 16265 1539
rect 16299 1505 16409 1539
rect 16443 1505 16481 1539
rect 16515 1505 16553 1539
rect 16587 1505 16625 1539
rect 16659 1505 16697 1539
rect 16731 1505 16769 1539
rect 16803 1505 16867 1539
rect 16901 1505 16939 1539
rect 16973 1505 17011 1539
rect 17045 1505 17083 1539
rect 17117 1505 17155 1539
rect 17189 1505 17227 1539
rect 17261 1505 17371 1539
rect 17405 1505 17443 1539
rect 17477 1505 17515 1539
rect 17549 1505 17587 1539
rect 17621 1505 17677 1539
rect 17711 1505 17749 1539
rect 17783 1505 17821 1539
rect 17855 1505 17893 1539
rect 17927 1505 18037 1539
rect 18071 1505 18109 1539
rect 18143 1505 18181 1539
rect 18215 1505 18253 1539
rect 18287 1505 18343 1539
rect 18377 1505 18415 1539
rect 18449 1505 18487 1539
rect 18521 1505 18559 1539
rect 18593 1505 18703 1539
rect 18737 1505 18775 1539
rect 18809 1505 18847 1539
rect 18881 1505 18919 1539
rect 18953 1505 19009 1539
rect 19043 1505 19081 1539
rect 19115 1505 19153 1539
rect 19187 1505 19225 1539
rect 19259 1505 19345 1539
rect -31 1470 31 1505
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect 931 1470 993 1505
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect -31 1038 31 1076
rect 931 1436 945 1470
rect 979 1436 993 1470
rect 1893 1470 1955 1505
rect 931 1398 993 1436
rect 931 1364 945 1398
rect 979 1364 993 1398
rect 931 1326 993 1364
rect 931 1292 945 1326
rect 979 1292 993 1326
rect 931 1254 993 1292
rect 931 1220 945 1254
rect 979 1220 993 1254
rect 931 1182 993 1220
rect 931 1148 945 1182
rect 979 1148 993 1182
rect 931 1110 993 1148
rect 931 1076 945 1110
rect 979 1076 993 1110
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect 931 1038 993 1076
rect 1893 1436 1907 1470
rect 1941 1436 1955 1470
rect 2855 1470 2917 1505
rect 1893 1398 1955 1436
rect 1893 1364 1907 1398
rect 1941 1364 1955 1398
rect 1893 1326 1955 1364
rect 1893 1292 1907 1326
rect 1941 1292 1955 1326
rect 1893 1254 1955 1292
rect 1893 1220 1907 1254
rect 1941 1220 1955 1254
rect 1893 1182 1955 1220
rect 1893 1148 1907 1182
rect 1941 1148 1955 1182
rect 1893 1110 1955 1148
rect 1893 1076 1907 1110
rect 1941 1076 1955 1110
rect 931 1004 945 1038
rect 979 1004 993 1038
rect 931 966 993 1004
rect -31 930 31 932
rect 931 932 945 966
rect 979 932 993 966
rect 1893 1038 1955 1076
rect 2855 1436 2869 1470
rect 2903 1436 2917 1470
rect 3817 1470 3879 1505
rect 2855 1398 2917 1436
rect 2855 1364 2869 1398
rect 2903 1364 2917 1398
rect 2855 1326 2917 1364
rect 2855 1292 2869 1326
rect 2903 1292 2917 1326
rect 2855 1254 2917 1292
rect 2855 1220 2869 1254
rect 2903 1220 2917 1254
rect 2855 1182 2917 1220
rect 2855 1148 2869 1182
rect 2903 1148 2917 1182
rect 2855 1110 2917 1148
rect 2855 1076 2869 1110
rect 2903 1076 2917 1110
rect 1893 1004 1907 1038
rect 1941 1004 1955 1038
rect 1893 966 1955 1004
rect 931 930 993 932
rect 1893 932 1907 966
rect 1941 932 1955 966
rect 2855 1038 2917 1076
rect 3817 1436 3831 1470
rect 3865 1436 3879 1470
rect 4779 1470 4841 1505
rect 3817 1398 3879 1436
rect 3817 1364 3831 1398
rect 3865 1364 3879 1398
rect 3817 1326 3879 1364
rect 3817 1292 3831 1326
rect 3865 1292 3879 1326
rect 3817 1254 3879 1292
rect 3817 1220 3831 1254
rect 3865 1220 3879 1254
rect 3817 1182 3879 1220
rect 3817 1148 3831 1182
rect 3865 1148 3879 1182
rect 3817 1110 3879 1148
rect 3817 1076 3831 1110
rect 3865 1076 3879 1110
rect 2855 1004 2869 1038
rect 2903 1004 2917 1038
rect 2855 966 2917 1004
rect 1893 930 1955 932
rect 2855 932 2869 966
rect 2903 932 2917 966
rect 3817 1038 3879 1076
rect 4779 1436 4793 1470
rect 4827 1436 4841 1470
rect 5741 1470 5803 1505
rect 4779 1398 4841 1436
rect 4779 1364 4793 1398
rect 4827 1364 4841 1398
rect 4779 1326 4841 1364
rect 4779 1292 4793 1326
rect 4827 1292 4841 1326
rect 4779 1254 4841 1292
rect 4779 1220 4793 1254
rect 4827 1220 4841 1254
rect 4779 1182 4841 1220
rect 4779 1148 4793 1182
rect 4827 1148 4841 1182
rect 4779 1110 4841 1148
rect 4779 1076 4793 1110
rect 4827 1076 4841 1110
rect 3817 1004 3831 1038
rect 3865 1004 3879 1038
rect 3817 966 3879 1004
rect 2855 930 2917 932
rect 3817 932 3831 966
rect 3865 932 3879 966
rect 4779 1038 4841 1076
rect 5741 1436 5755 1470
rect 5789 1436 5803 1470
rect 6703 1470 6765 1505
rect 5741 1398 5803 1436
rect 5741 1364 5755 1398
rect 5789 1364 5803 1398
rect 5741 1326 5803 1364
rect 5741 1292 5755 1326
rect 5789 1292 5803 1326
rect 5741 1254 5803 1292
rect 5741 1220 5755 1254
rect 5789 1220 5803 1254
rect 5741 1182 5803 1220
rect 5741 1148 5755 1182
rect 5789 1148 5803 1182
rect 5741 1110 5803 1148
rect 5741 1076 5755 1110
rect 5789 1076 5803 1110
rect 4779 1004 4793 1038
rect 4827 1004 4841 1038
rect 4779 966 4841 1004
rect 3817 930 3879 932
rect 4779 932 4793 966
rect 4827 932 4841 966
rect 5741 1038 5803 1076
rect 6703 1436 6717 1470
rect 6751 1436 6765 1470
rect 7665 1470 7727 1505
rect 6703 1398 6765 1436
rect 6703 1364 6717 1398
rect 6751 1364 6765 1398
rect 6703 1326 6765 1364
rect 6703 1292 6717 1326
rect 6751 1292 6765 1326
rect 6703 1254 6765 1292
rect 6703 1220 6717 1254
rect 6751 1220 6765 1254
rect 6703 1182 6765 1220
rect 6703 1148 6717 1182
rect 6751 1148 6765 1182
rect 6703 1110 6765 1148
rect 6703 1076 6717 1110
rect 6751 1076 6765 1110
rect 5741 1004 5755 1038
rect 5789 1004 5803 1038
rect 5741 966 5803 1004
rect 4779 930 4841 932
rect 5741 932 5755 966
rect 5789 932 5803 966
rect 6703 1038 6765 1076
rect 7665 1436 7679 1470
rect 7713 1436 7727 1470
rect 8627 1470 8689 1505
rect 7665 1398 7727 1436
rect 7665 1364 7679 1398
rect 7713 1364 7727 1398
rect 7665 1326 7727 1364
rect 7665 1292 7679 1326
rect 7713 1292 7727 1326
rect 7665 1254 7727 1292
rect 7665 1220 7679 1254
rect 7713 1220 7727 1254
rect 7665 1182 7727 1220
rect 7665 1148 7679 1182
rect 7713 1148 7727 1182
rect 7665 1110 7727 1148
rect 7665 1076 7679 1110
rect 7713 1076 7727 1110
rect 6703 1004 6717 1038
rect 6751 1004 6765 1038
rect 6703 966 6765 1004
rect 5741 930 5803 932
rect 6703 932 6717 966
rect 6751 932 6765 966
rect 7665 1038 7727 1076
rect 8627 1436 8641 1470
rect 8675 1436 8689 1470
rect 9589 1470 9651 1505
rect 8627 1398 8689 1436
rect 8627 1364 8641 1398
rect 8675 1364 8689 1398
rect 8627 1326 8689 1364
rect 8627 1292 8641 1326
rect 8675 1292 8689 1326
rect 8627 1254 8689 1292
rect 8627 1220 8641 1254
rect 8675 1220 8689 1254
rect 8627 1182 8689 1220
rect 8627 1148 8641 1182
rect 8675 1148 8689 1182
rect 8627 1110 8689 1148
rect 8627 1076 8641 1110
rect 8675 1076 8689 1110
rect 7665 1004 7679 1038
rect 7713 1004 7727 1038
rect 7665 966 7727 1004
rect 6703 930 6765 932
rect 7665 932 7679 966
rect 7713 932 7727 966
rect 8627 1038 8689 1076
rect 9589 1436 9603 1470
rect 9637 1436 9651 1470
rect 10551 1470 10613 1505
rect 9589 1398 9651 1436
rect 9589 1364 9603 1398
rect 9637 1364 9651 1398
rect 9589 1326 9651 1364
rect 9589 1292 9603 1326
rect 9637 1292 9651 1326
rect 9589 1254 9651 1292
rect 9589 1220 9603 1254
rect 9637 1220 9651 1254
rect 9589 1182 9651 1220
rect 9589 1148 9603 1182
rect 9637 1148 9651 1182
rect 9589 1110 9651 1148
rect 9589 1076 9603 1110
rect 9637 1076 9651 1110
rect 8627 1004 8641 1038
rect 8675 1004 8689 1038
rect 8627 966 8689 1004
rect 7665 930 7727 932
rect 8627 932 8641 966
rect 8675 932 8689 966
rect 9589 1038 9651 1076
rect 10551 1436 10565 1470
rect 10599 1436 10613 1470
rect 11513 1470 11575 1505
rect 10551 1398 10613 1436
rect 10551 1364 10565 1398
rect 10599 1364 10613 1398
rect 10551 1326 10613 1364
rect 10551 1292 10565 1326
rect 10599 1292 10613 1326
rect 10551 1254 10613 1292
rect 10551 1220 10565 1254
rect 10599 1220 10613 1254
rect 10551 1182 10613 1220
rect 10551 1148 10565 1182
rect 10599 1148 10613 1182
rect 10551 1110 10613 1148
rect 10551 1076 10565 1110
rect 10599 1076 10613 1110
rect 9589 1004 9603 1038
rect 9637 1004 9651 1038
rect 9589 966 9651 1004
rect 8627 930 8689 932
rect 9589 932 9603 966
rect 9637 932 9651 966
rect 10551 1038 10613 1076
rect 11513 1436 11527 1470
rect 11561 1436 11575 1470
rect 12475 1470 12537 1505
rect 11513 1398 11575 1436
rect 11513 1364 11527 1398
rect 11561 1364 11575 1398
rect 11513 1326 11575 1364
rect 11513 1292 11527 1326
rect 11561 1292 11575 1326
rect 11513 1254 11575 1292
rect 11513 1220 11527 1254
rect 11561 1220 11575 1254
rect 11513 1182 11575 1220
rect 11513 1148 11527 1182
rect 11561 1148 11575 1182
rect 11513 1110 11575 1148
rect 11513 1076 11527 1110
rect 11561 1076 11575 1110
rect 10551 1004 10565 1038
rect 10599 1004 10613 1038
rect 10551 966 10613 1004
rect 9589 930 9651 932
rect 10551 932 10565 966
rect 10599 932 10613 966
rect 11513 1038 11575 1076
rect 12475 1436 12489 1470
rect 12523 1436 12537 1470
rect 13437 1470 13499 1505
rect 12475 1398 12537 1436
rect 12475 1364 12489 1398
rect 12523 1364 12537 1398
rect 12475 1326 12537 1364
rect 12475 1292 12489 1326
rect 12523 1292 12537 1326
rect 12475 1254 12537 1292
rect 12475 1220 12489 1254
rect 12523 1220 12537 1254
rect 12475 1182 12537 1220
rect 12475 1148 12489 1182
rect 12523 1148 12537 1182
rect 12475 1110 12537 1148
rect 12475 1076 12489 1110
rect 12523 1076 12537 1110
rect 11513 1004 11527 1038
rect 11561 1004 11575 1038
rect 11513 966 11575 1004
rect 10551 930 10613 932
rect 11513 932 11527 966
rect 11561 932 11575 966
rect 12475 1038 12537 1076
rect 13437 1436 13451 1470
rect 13485 1436 13499 1470
rect 14399 1470 14461 1505
rect 13437 1398 13499 1436
rect 13437 1364 13451 1398
rect 13485 1364 13499 1398
rect 13437 1326 13499 1364
rect 13437 1292 13451 1326
rect 13485 1292 13499 1326
rect 13437 1254 13499 1292
rect 13437 1220 13451 1254
rect 13485 1220 13499 1254
rect 13437 1182 13499 1220
rect 13437 1148 13451 1182
rect 13485 1148 13499 1182
rect 13437 1110 13499 1148
rect 13437 1076 13451 1110
rect 13485 1076 13499 1110
rect 12475 1004 12489 1038
rect 12523 1004 12537 1038
rect 12475 966 12537 1004
rect 11513 930 11575 932
rect 12475 932 12489 966
rect 12523 932 12537 966
rect 13437 1038 13499 1076
rect 14399 1436 14413 1470
rect 14447 1436 14461 1470
rect 15361 1470 15423 1505
rect 14399 1398 14461 1436
rect 14399 1364 14413 1398
rect 14447 1364 14461 1398
rect 14399 1326 14461 1364
rect 14399 1292 14413 1326
rect 14447 1292 14461 1326
rect 14399 1254 14461 1292
rect 14399 1220 14413 1254
rect 14447 1220 14461 1254
rect 14399 1182 14461 1220
rect 14399 1148 14413 1182
rect 14447 1148 14461 1182
rect 14399 1110 14461 1148
rect 14399 1076 14413 1110
rect 14447 1076 14461 1110
rect 13437 1004 13451 1038
rect 13485 1004 13499 1038
rect 13437 966 13499 1004
rect 12475 930 12537 932
rect 13437 932 13451 966
rect 13485 932 13499 966
rect 14399 1038 14461 1076
rect 15361 1436 15375 1470
rect 15409 1436 15423 1470
rect 16323 1470 16385 1505
rect 15361 1398 15423 1436
rect 15361 1364 15375 1398
rect 15409 1364 15423 1398
rect 15361 1326 15423 1364
rect 15361 1292 15375 1326
rect 15409 1292 15423 1326
rect 15361 1254 15423 1292
rect 15361 1220 15375 1254
rect 15409 1220 15423 1254
rect 15361 1182 15423 1220
rect 15361 1148 15375 1182
rect 15409 1148 15423 1182
rect 15361 1110 15423 1148
rect 15361 1076 15375 1110
rect 15409 1076 15423 1110
rect 14399 1004 14413 1038
rect 14447 1004 14461 1038
rect 14399 966 14461 1004
rect 13437 930 13499 932
rect 14399 932 14413 966
rect 14447 932 14461 966
rect 15361 1038 15423 1076
rect 16323 1436 16337 1470
rect 16371 1436 16385 1470
rect 17285 1470 17347 1505
rect 16323 1398 16385 1436
rect 16323 1364 16337 1398
rect 16371 1364 16385 1398
rect 16323 1326 16385 1364
rect 16323 1292 16337 1326
rect 16371 1292 16385 1326
rect 16323 1254 16385 1292
rect 16323 1220 16337 1254
rect 16371 1220 16385 1254
rect 16323 1182 16385 1220
rect 16323 1148 16337 1182
rect 16371 1148 16385 1182
rect 16323 1110 16385 1148
rect 16323 1076 16337 1110
rect 16371 1076 16385 1110
rect 15361 1004 15375 1038
rect 15409 1004 15423 1038
rect 15361 966 15423 1004
rect 14399 930 14461 932
rect 15361 932 15375 966
rect 15409 932 15423 966
rect 16323 1038 16385 1076
rect 17285 1436 17299 1470
rect 17333 1436 17347 1470
rect 17951 1470 18013 1505
rect 17285 1398 17347 1436
rect 17285 1364 17299 1398
rect 17333 1364 17347 1398
rect 17285 1326 17347 1364
rect 17285 1292 17299 1326
rect 17333 1292 17347 1326
rect 17285 1254 17347 1292
rect 17285 1220 17299 1254
rect 17333 1220 17347 1254
rect 17285 1182 17347 1220
rect 17285 1148 17299 1182
rect 17333 1148 17347 1182
rect 17285 1110 17347 1148
rect 17285 1076 17299 1110
rect 17333 1076 17347 1110
rect 16323 1004 16337 1038
rect 16371 1004 16385 1038
rect 16323 966 16385 1004
rect 15361 930 15423 932
rect 16323 932 16337 966
rect 16371 932 16385 966
rect 17285 1038 17347 1076
rect 17951 1436 17965 1470
rect 17999 1436 18013 1470
rect 18617 1470 18679 1505
rect 17951 1398 18013 1436
rect 17951 1364 17965 1398
rect 17999 1364 18013 1398
rect 17951 1326 18013 1364
rect 17951 1292 17965 1326
rect 17999 1292 18013 1326
rect 17951 1254 18013 1292
rect 17951 1220 17965 1254
rect 17999 1220 18013 1254
rect 17951 1182 18013 1220
rect 17951 1148 17965 1182
rect 17999 1148 18013 1182
rect 17951 1110 18013 1148
rect 17951 1076 17965 1110
rect 17999 1076 18013 1110
rect 17285 1004 17299 1038
rect 17333 1004 17347 1038
rect 17285 966 17347 1004
rect 16323 930 16385 932
rect 17285 932 17299 966
rect 17333 932 17347 966
rect 17951 1038 18013 1076
rect 18617 1436 18631 1470
rect 18665 1436 18679 1470
rect 19283 1470 19345 1505
rect 18617 1398 18679 1436
rect 18617 1364 18631 1398
rect 18665 1364 18679 1398
rect 18617 1326 18679 1364
rect 18617 1292 18631 1326
rect 18665 1292 18679 1326
rect 18617 1254 18679 1292
rect 18617 1220 18631 1254
rect 18665 1220 18679 1254
rect 18617 1182 18679 1220
rect 18617 1148 18631 1182
rect 18665 1148 18679 1182
rect 18617 1110 18679 1148
rect 18617 1076 18631 1110
rect 18665 1076 18679 1110
rect 17951 1004 17965 1038
rect 17999 1004 18013 1038
rect 17951 966 18013 1004
rect 17285 930 17347 932
rect 17951 932 17965 966
rect 17999 932 18013 966
rect 18617 1038 18679 1076
rect 19283 1436 19297 1470
rect 19331 1436 19345 1470
rect 19283 1398 19345 1436
rect 19283 1364 19297 1398
rect 19331 1364 19345 1398
rect 19283 1326 19345 1364
rect 19283 1292 19297 1326
rect 19331 1292 19345 1326
rect 19283 1254 19345 1292
rect 19283 1220 19297 1254
rect 19331 1220 19345 1254
rect 19283 1182 19345 1220
rect 19283 1148 19297 1182
rect 19331 1148 19345 1182
rect 19283 1110 19345 1148
rect 19283 1076 19297 1110
rect 19331 1076 19345 1110
rect 18617 1004 18631 1038
rect 18665 1004 18679 1038
rect 18617 966 18679 1004
rect 17951 930 18013 932
rect 18617 932 18631 966
rect 18665 932 18679 966
rect 19283 1038 19345 1076
rect 19283 1004 19297 1038
rect 19331 1004 19345 1038
rect 19283 966 19345 1004
rect 18617 930 18679 932
rect 19283 932 19297 966
rect 19331 932 19345 966
rect 19283 930 19345 932
rect -31 868 19345 930
<< psubdiffcont >>
rect -17 512 17 546
rect 945 512 979 546
rect 1907 512 1941 546
rect 2869 512 2903 546
rect 3831 512 3865 546
rect 4793 512 4827 546
rect 5755 512 5789 546
rect 6717 512 6751 546
rect 7679 512 7713 546
rect 8641 512 8675 546
rect 9603 512 9637 546
rect 10565 512 10599 546
rect 11527 512 11561 546
rect 12489 512 12523 546
rect 13451 512 13485 546
rect 14413 512 14447 546
rect 15375 512 15409 546
rect 16337 512 16371 546
rect 17299 512 17333 546
rect 17965 512 17999 546
rect 18631 512 18665 546
rect 19297 512 19331 546
rect -17 440 17 474
rect -17 368 17 402
rect 945 440 979 474
rect -17 296 17 330
rect -17 224 17 258
rect -17 152 17 186
rect -17 80 17 114
rect 945 368 979 402
rect 1907 440 1941 474
rect 945 296 979 330
rect 945 224 979 258
rect 945 152 979 186
rect 945 80 979 114
rect 1907 368 1941 402
rect 2869 440 2903 474
rect 1907 296 1941 330
rect 1907 224 1941 258
rect 1907 152 1941 186
rect 1907 80 1941 114
rect 2869 368 2903 402
rect 3831 440 3865 474
rect 2869 296 2903 330
rect 2869 224 2903 258
rect 2869 152 2903 186
rect 2869 80 2903 114
rect 3831 368 3865 402
rect 4793 440 4827 474
rect 3831 296 3865 330
rect 3831 224 3865 258
rect 3831 152 3865 186
rect 3831 80 3865 114
rect 4793 368 4827 402
rect 5755 440 5789 474
rect 4793 296 4827 330
rect 4793 224 4827 258
rect 4793 152 4827 186
rect 4793 80 4827 114
rect 5755 368 5789 402
rect 6717 440 6751 474
rect 5755 296 5789 330
rect 5755 224 5789 258
rect 5755 152 5789 186
rect 5755 80 5789 114
rect 6717 368 6751 402
rect 7679 440 7713 474
rect 6717 296 6751 330
rect 6717 224 6751 258
rect 6717 152 6751 186
rect 6717 80 6751 114
rect 7679 368 7713 402
rect 8641 440 8675 474
rect 7679 296 7713 330
rect 7679 224 7713 258
rect 7679 152 7713 186
rect 7679 80 7713 114
rect 8641 368 8675 402
rect 9603 440 9637 474
rect 8641 296 8675 330
rect 8641 224 8675 258
rect 8641 152 8675 186
rect 8641 80 8675 114
rect 9603 368 9637 402
rect 10565 440 10599 474
rect 9603 296 9637 330
rect 9603 224 9637 258
rect 9603 152 9637 186
rect 9603 80 9637 114
rect 10565 368 10599 402
rect 11527 440 11561 474
rect 10565 296 10599 330
rect 10565 224 10599 258
rect 10565 152 10599 186
rect 10565 80 10599 114
rect 11527 368 11561 402
rect 12489 440 12523 474
rect 11527 296 11561 330
rect 11527 224 11561 258
rect 11527 152 11561 186
rect 11527 80 11561 114
rect 12489 368 12523 402
rect 13451 440 13485 474
rect 12489 296 12523 330
rect 12489 224 12523 258
rect 12489 152 12523 186
rect 12489 80 12523 114
rect 13451 368 13485 402
rect 14413 440 14447 474
rect 13451 296 13485 330
rect 13451 224 13485 258
rect 13451 152 13485 186
rect 13451 80 13485 114
rect 14413 368 14447 402
rect 15375 440 15409 474
rect 14413 296 14447 330
rect 14413 224 14447 258
rect 14413 152 14447 186
rect 14413 80 14447 114
rect 15375 368 15409 402
rect 16337 440 16371 474
rect 15375 296 15409 330
rect 15375 224 15409 258
rect 15375 152 15409 186
rect 15375 80 15409 114
rect 16337 368 16371 402
rect 17299 440 17333 474
rect 17965 440 17999 474
rect 16337 296 16371 330
rect 16337 224 16371 258
rect 16337 152 16371 186
rect 16337 80 16371 114
rect 17299 368 17333 402
rect 17299 296 17333 330
rect 17299 224 17333 258
rect 17299 152 17333 186
rect 17299 80 17333 114
rect 17965 368 17999 402
rect 18631 440 18665 474
rect 19297 440 19331 474
rect 17965 296 17999 330
rect 17965 224 17999 258
rect 17965 152 17999 186
rect 17965 80 17999 114
rect 18631 368 18665 402
rect 18631 296 18665 330
rect 18631 224 18665 258
rect 18631 152 18665 186
rect 18631 80 18665 114
rect 19297 368 19331 402
rect 19297 296 19331 330
rect 19297 224 19331 258
rect 19297 152 19331 186
rect 19297 80 19331 114
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 343 13 377 47
rect 415 13 449 47
rect 513 13 547 47
rect 585 13 619 47
rect 657 13 691 47
rect 729 13 763 47
rect 801 13 835 47
rect 873 13 907 47
rect 1017 13 1051 47
rect 1089 13 1123 47
rect 1161 13 1195 47
rect 1233 13 1267 47
rect 1305 13 1339 47
rect 1377 13 1411 47
rect 1475 13 1509 47
rect 1547 13 1581 47
rect 1619 13 1653 47
rect 1691 13 1725 47
rect 1763 13 1797 47
rect 1835 13 1869 47
rect 1979 13 2013 47
rect 2051 13 2085 47
rect 2123 13 2157 47
rect 2195 13 2229 47
rect 2267 13 2301 47
rect 2339 13 2373 47
rect 2437 13 2471 47
rect 2509 13 2543 47
rect 2581 13 2615 47
rect 2653 13 2687 47
rect 2725 13 2759 47
rect 2797 13 2831 47
rect 2941 13 2975 47
rect 3013 13 3047 47
rect 3085 13 3119 47
rect 3157 13 3191 47
rect 3229 13 3263 47
rect 3301 13 3335 47
rect 3399 13 3433 47
rect 3471 13 3505 47
rect 3543 13 3577 47
rect 3615 13 3649 47
rect 3687 13 3721 47
rect 3759 13 3793 47
rect 3903 13 3937 47
rect 3975 13 4009 47
rect 4047 13 4081 47
rect 4119 13 4153 47
rect 4191 13 4225 47
rect 4263 13 4297 47
rect 4361 13 4395 47
rect 4433 13 4467 47
rect 4505 13 4539 47
rect 4577 13 4611 47
rect 4649 13 4683 47
rect 4721 13 4755 47
rect 4865 13 4899 47
rect 4937 13 4971 47
rect 5009 13 5043 47
rect 5081 13 5115 47
rect 5153 13 5187 47
rect 5225 13 5259 47
rect 5323 13 5357 47
rect 5395 13 5429 47
rect 5467 13 5501 47
rect 5539 13 5573 47
rect 5611 13 5645 47
rect 5683 13 5717 47
rect 5827 13 5861 47
rect 5899 13 5933 47
rect 5971 13 6005 47
rect 6043 13 6077 47
rect 6115 13 6149 47
rect 6187 13 6221 47
rect 6285 13 6319 47
rect 6357 13 6391 47
rect 6429 13 6463 47
rect 6501 13 6535 47
rect 6573 13 6607 47
rect 6645 13 6679 47
rect 6789 13 6823 47
rect 6861 13 6895 47
rect 6933 13 6967 47
rect 7005 13 7039 47
rect 7077 13 7111 47
rect 7149 13 7183 47
rect 7247 13 7281 47
rect 7319 13 7353 47
rect 7391 13 7425 47
rect 7463 13 7497 47
rect 7535 13 7569 47
rect 7607 13 7641 47
rect 7751 13 7785 47
rect 7823 13 7857 47
rect 7895 13 7929 47
rect 7967 13 8001 47
rect 8039 13 8073 47
rect 8111 13 8145 47
rect 8209 13 8243 47
rect 8281 13 8315 47
rect 8353 13 8387 47
rect 8425 13 8459 47
rect 8497 13 8531 47
rect 8569 13 8603 47
rect 8713 13 8747 47
rect 8785 13 8819 47
rect 8857 13 8891 47
rect 8929 13 8963 47
rect 9001 13 9035 47
rect 9073 13 9107 47
rect 9171 13 9205 47
rect 9243 13 9277 47
rect 9315 13 9349 47
rect 9387 13 9421 47
rect 9459 13 9493 47
rect 9531 13 9565 47
rect 9675 13 9709 47
rect 9747 13 9781 47
rect 9819 13 9853 47
rect 9891 13 9925 47
rect 9963 13 9997 47
rect 10035 13 10069 47
rect 10133 13 10167 47
rect 10205 13 10239 47
rect 10277 13 10311 47
rect 10349 13 10383 47
rect 10421 13 10455 47
rect 10493 13 10527 47
rect 10637 13 10671 47
rect 10709 13 10743 47
rect 10781 13 10815 47
rect 10853 13 10887 47
rect 10925 13 10959 47
rect 10997 13 11031 47
rect 11095 13 11129 47
rect 11167 13 11201 47
rect 11239 13 11273 47
rect 11311 13 11345 47
rect 11383 13 11417 47
rect 11455 13 11489 47
rect 11599 13 11633 47
rect 11671 13 11705 47
rect 11743 13 11777 47
rect 11815 13 11849 47
rect 11887 13 11921 47
rect 11959 13 11993 47
rect 12057 13 12091 47
rect 12129 13 12163 47
rect 12201 13 12235 47
rect 12273 13 12307 47
rect 12345 13 12379 47
rect 12417 13 12451 47
rect 12561 13 12595 47
rect 12633 13 12667 47
rect 12705 13 12739 47
rect 12777 13 12811 47
rect 12849 13 12883 47
rect 12921 13 12955 47
rect 13019 13 13053 47
rect 13091 13 13125 47
rect 13163 13 13197 47
rect 13235 13 13269 47
rect 13307 13 13341 47
rect 13379 13 13413 47
rect 13523 13 13557 47
rect 13595 13 13629 47
rect 13667 13 13701 47
rect 13739 13 13773 47
rect 13811 13 13845 47
rect 13883 13 13917 47
rect 13981 13 14015 47
rect 14053 13 14087 47
rect 14125 13 14159 47
rect 14197 13 14231 47
rect 14269 13 14303 47
rect 14341 13 14375 47
rect 14485 13 14519 47
rect 14557 13 14591 47
rect 14629 13 14663 47
rect 14701 13 14735 47
rect 14773 13 14807 47
rect 14845 13 14879 47
rect 14943 13 14977 47
rect 15015 13 15049 47
rect 15087 13 15121 47
rect 15159 13 15193 47
rect 15231 13 15265 47
rect 15303 13 15337 47
rect 15447 13 15481 47
rect 15519 13 15553 47
rect 15591 13 15625 47
rect 15663 13 15697 47
rect 15735 13 15769 47
rect 15807 13 15841 47
rect 15905 13 15939 47
rect 15977 13 16011 47
rect 16049 13 16083 47
rect 16121 13 16155 47
rect 16193 13 16227 47
rect 16265 13 16299 47
rect 16409 13 16443 47
rect 16481 13 16515 47
rect 16553 13 16587 47
rect 16625 13 16659 47
rect 16697 13 16731 47
rect 16769 13 16803 47
rect 16867 13 16901 47
rect 16939 13 16973 47
rect 17011 13 17045 47
rect 17083 13 17117 47
rect 17155 13 17189 47
rect 17227 13 17261 47
rect 17371 13 17405 47
rect 17443 13 17477 47
rect 17515 13 17549 47
rect 17587 13 17621 47
rect 17677 13 17711 47
rect 17749 13 17783 47
rect 17821 13 17855 47
rect 17893 13 17927 47
rect 18037 13 18071 47
rect 18109 13 18143 47
rect 18181 13 18215 47
rect 18253 13 18287 47
rect 18343 13 18377 47
rect 18415 13 18449 47
rect 18487 13 18521 47
rect 18559 13 18593 47
rect 18703 13 18737 47
rect 18775 13 18809 47
rect 18847 13 18881 47
rect 18919 13 18953 47
rect 19009 13 19043 47
rect 19081 13 19115 47
rect 19153 13 19187 47
rect 19225 13 19259 47
<< nsubdiffcont >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 343 1505 377 1539
rect 415 1505 449 1539
rect 513 1505 547 1539
rect 585 1505 619 1539
rect 657 1505 691 1539
rect 729 1505 763 1539
rect 801 1505 835 1539
rect 873 1505 907 1539
rect 1017 1505 1051 1539
rect 1089 1505 1123 1539
rect 1161 1505 1195 1539
rect 1233 1505 1267 1539
rect 1305 1505 1339 1539
rect 1377 1505 1411 1539
rect 1475 1505 1509 1539
rect 1547 1505 1581 1539
rect 1619 1505 1653 1539
rect 1691 1505 1725 1539
rect 1763 1505 1797 1539
rect 1835 1505 1869 1539
rect 1979 1505 2013 1539
rect 2051 1505 2085 1539
rect 2123 1505 2157 1539
rect 2195 1505 2229 1539
rect 2267 1505 2301 1539
rect 2339 1505 2373 1539
rect 2437 1505 2471 1539
rect 2509 1505 2543 1539
rect 2581 1505 2615 1539
rect 2653 1505 2687 1539
rect 2725 1505 2759 1539
rect 2797 1505 2831 1539
rect 2941 1505 2975 1539
rect 3013 1505 3047 1539
rect 3085 1505 3119 1539
rect 3157 1505 3191 1539
rect 3229 1505 3263 1539
rect 3301 1505 3335 1539
rect 3399 1505 3433 1539
rect 3471 1505 3505 1539
rect 3543 1505 3577 1539
rect 3615 1505 3649 1539
rect 3687 1505 3721 1539
rect 3759 1505 3793 1539
rect 3903 1505 3937 1539
rect 3975 1505 4009 1539
rect 4047 1505 4081 1539
rect 4119 1505 4153 1539
rect 4191 1505 4225 1539
rect 4263 1505 4297 1539
rect 4361 1505 4395 1539
rect 4433 1505 4467 1539
rect 4505 1505 4539 1539
rect 4577 1505 4611 1539
rect 4649 1505 4683 1539
rect 4721 1505 4755 1539
rect 4865 1505 4899 1539
rect 4937 1505 4971 1539
rect 5009 1505 5043 1539
rect 5081 1505 5115 1539
rect 5153 1505 5187 1539
rect 5225 1505 5259 1539
rect 5323 1505 5357 1539
rect 5395 1505 5429 1539
rect 5467 1505 5501 1539
rect 5539 1505 5573 1539
rect 5611 1505 5645 1539
rect 5683 1505 5717 1539
rect 5827 1505 5861 1539
rect 5899 1505 5933 1539
rect 5971 1505 6005 1539
rect 6043 1505 6077 1539
rect 6115 1505 6149 1539
rect 6187 1505 6221 1539
rect 6285 1505 6319 1539
rect 6357 1505 6391 1539
rect 6429 1505 6463 1539
rect 6501 1505 6535 1539
rect 6573 1505 6607 1539
rect 6645 1505 6679 1539
rect 6789 1505 6823 1539
rect 6861 1505 6895 1539
rect 6933 1505 6967 1539
rect 7005 1505 7039 1539
rect 7077 1505 7111 1539
rect 7149 1505 7183 1539
rect 7247 1505 7281 1539
rect 7319 1505 7353 1539
rect 7391 1505 7425 1539
rect 7463 1505 7497 1539
rect 7535 1505 7569 1539
rect 7607 1505 7641 1539
rect 7751 1505 7785 1539
rect 7823 1505 7857 1539
rect 7895 1505 7929 1539
rect 7967 1505 8001 1539
rect 8039 1505 8073 1539
rect 8111 1505 8145 1539
rect 8209 1505 8243 1539
rect 8281 1505 8315 1539
rect 8353 1505 8387 1539
rect 8425 1505 8459 1539
rect 8497 1505 8531 1539
rect 8569 1505 8603 1539
rect 8713 1505 8747 1539
rect 8785 1505 8819 1539
rect 8857 1505 8891 1539
rect 8929 1505 8963 1539
rect 9001 1505 9035 1539
rect 9073 1505 9107 1539
rect 9171 1505 9205 1539
rect 9243 1505 9277 1539
rect 9315 1505 9349 1539
rect 9387 1505 9421 1539
rect 9459 1505 9493 1539
rect 9531 1505 9565 1539
rect 9675 1505 9709 1539
rect 9747 1505 9781 1539
rect 9819 1505 9853 1539
rect 9891 1505 9925 1539
rect 9963 1505 9997 1539
rect 10035 1505 10069 1539
rect 10133 1505 10167 1539
rect 10205 1505 10239 1539
rect 10277 1505 10311 1539
rect 10349 1505 10383 1539
rect 10421 1505 10455 1539
rect 10493 1505 10527 1539
rect 10637 1505 10671 1539
rect 10709 1505 10743 1539
rect 10781 1505 10815 1539
rect 10853 1505 10887 1539
rect 10925 1505 10959 1539
rect 10997 1505 11031 1539
rect 11095 1505 11129 1539
rect 11167 1505 11201 1539
rect 11239 1505 11273 1539
rect 11311 1505 11345 1539
rect 11383 1505 11417 1539
rect 11455 1505 11489 1539
rect 11599 1505 11633 1539
rect 11671 1505 11705 1539
rect 11743 1505 11777 1539
rect 11815 1505 11849 1539
rect 11887 1505 11921 1539
rect 11959 1505 11993 1539
rect 12057 1505 12091 1539
rect 12129 1505 12163 1539
rect 12201 1505 12235 1539
rect 12273 1505 12307 1539
rect 12345 1505 12379 1539
rect 12417 1505 12451 1539
rect 12561 1505 12595 1539
rect 12633 1505 12667 1539
rect 12705 1505 12739 1539
rect 12777 1505 12811 1539
rect 12849 1505 12883 1539
rect 12921 1505 12955 1539
rect 13019 1505 13053 1539
rect 13091 1505 13125 1539
rect 13163 1505 13197 1539
rect 13235 1505 13269 1539
rect 13307 1505 13341 1539
rect 13379 1505 13413 1539
rect 13523 1505 13557 1539
rect 13595 1505 13629 1539
rect 13667 1505 13701 1539
rect 13739 1505 13773 1539
rect 13811 1505 13845 1539
rect 13883 1505 13917 1539
rect 13981 1505 14015 1539
rect 14053 1505 14087 1539
rect 14125 1505 14159 1539
rect 14197 1505 14231 1539
rect 14269 1505 14303 1539
rect 14341 1505 14375 1539
rect 14485 1505 14519 1539
rect 14557 1505 14591 1539
rect 14629 1505 14663 1539
rect 14701 1505 14735 1539
rect 14773 1505 14807 1539
rect 14845 1505 14879 1539
rect 14943 1505 14977 1539
rect 15015 1505 15049 1539
rect 15087 1505 15121 1539
rect 15159 1505 15193 1539
rect 15231 1505 15265 1539
rect 15303 1505 15337 1539
rect 15447 1505 15481 1539
rect 15519 1505 15553 1539
rect 15591 1505 15625 1539
rect 15663 1505 15697 1539
rect 15735 1505 15769 1539
rect 15807 1505 15841 1539
rect 15905 1505 15939 1539
rect 15977 1505 16011 1539
rect 16049 1505 16083 1539
rect 16121 1505 16155 1539
rect 16193 1505 16227 1539
rect 16265 1505 16299 1539
rect 16409 1505 16443 1539
rect 16481 1505 16515 1539
rect 16553 1505 16587 1539
rect 16625 1505 16659 1539
rect 16697 1505 16731 1539
rect 16769 1505 16803 1539
rect 16867 1505 16901 1539
rect 16939 1505 16973 1539
rect 17011 1505 17045 1539
rect 17083 1505 17117 1539
rect 17155 1505 17189 1539
rect 17227 1505 17261 1539
rect 17371 1505 17405 1539
rect 17443 1505 17477 1539
rect 17515 1505 17549 1539
rect 17587 1505 17621 1539
rect 17677 1505 17711 1539
rect 17749 1505 17783 1539
rect 17821 1505 17855 1539
rect 17893 1505 17927 1539
rect 18037 1505 18071 1539
rect 18109 1505 18143 1539
rect 18181 1505 18215 1539
rect 18253 1505 18287 1539
rect 18343 1505 18377 1539
rect 18415 1505 18449 1539
rect 18487 1505 18521 1539
rect 18559 1505 18593 1539
rect 18703 1505 18737 1539
rect 18775 1505 18809 1539
rect 18847 1505 18881 1539
rect 18919 1505 18953 1539
rect 19009 1505 19043 1539
rect 19081 1505 19115 1539
rect 19153 1505 19187 1539
rect 19225 1505 19259 1539
rect -17 1436 17 1470
rect -17 1364 17 1398
rect -17 1292 17 1326
rect -17 1220 17 1254
rect -17 1148 17 1182
rect -17 1076 17 1110
rect 945 1436 979 1470
rect 945 1364 979 1398
rect 945 1292 979 1326
rect 945 1220 979 1254
rect 945 1148 979 1182
rect 945 1076 979 1110
rect -17 1004 17 1038
rect -17 932 17 966
rect 1907 1436 1941 1470
rect 1907 1364 1941 1398
rect 1907 1292 1941 1326
rect 1907 1220 1941 1254
rect 1907 1148 1941 1182
rect 1907 1076 1941 1110
rect 945 1004 979 1038
rect 945 932 979 966
rect 2869 1436 2903 1470
rect 2869 1364 2903 1398
rect 2869 1292 2903 1326
rect 2869 1220 2903 1254
rect 2869 1148 2903 1182
rect 2869 1076 2903 1110
rect 1907 1004 1941 1038
rect 1907 932 1941 966
rect 3831 1436 3865 1470
rect 3831 1364 3865 1398
rect 3831 1292 3865 1326
rect 3831 1220 3865 1254
rect 3831 1148 3865 1182
rect 3831 1076 3865 1110
rect 2869 1004 2903 1038
rect 2869 932 2903 966
rect 4793 1436 4827 1470
rect 4793 1364 4827 1398
rect 4793 1292 4827 1326
rect 4793 1220 4827 1254
rect 4793 1148 4827 1182
rect 4793 1076 4827 1110
rect 3831 1004 3865 1038
rect 3831 932 3865 966
rect 5755 1436 5789 1470
rect 5755 1364 5789 1398
rect 5755 1292 5789 1326
rect 5755 1220 5789 1254
rect 5755 1148 5789 1182
rect 5755 1076 5789 1110
rect 4793 1004 4827 1038
rect 4793 932 4827 966
rect 6717 1436 6751 1470
rect 6717 1364 6751 1398
rect 6717 1292 6751 1326
rect 6717 1220 6751 1254
rect 6717 1148 6751 1182
rect 6717 1076 6751 1110
rect 5755 1004 5789 1038
rect 5755 932 5789 966
rect 7679 1436 7713 1470
rect 7679 1364 7713 1398
rect 7679 1292 7713 1326
rect 7679 1220 7713 1254
rect 7679 1148 7713 1182
rect 7679 1076 7713 1110
rect 6717 1004 6751 1038
rect 6717 932 6751 966
rect 8641 1436 8675 1470
rect 8641 1364 8675 1398
rect 8641 1292 8675 1326
rect 8641 1220 8675 1254
rect 8641 1148 8675 1182
rect 8641 1076 8675 1110
rect 7679 1004 7713 1038
rect 7679 932 7713 966
rect 9603 1436 9637 1470
rect 9603 1364 9637 1398
rect 9603 1292 9637 1326
rect 9603 1220 9637 1254
rect 9603 1148 9637 1182
rect 9603 1076 9637 1110
rect 8641 1004 8675 1038
rect 8641 932 8675 966
rect 10565 1436 10599 1470
rect 10565 1364 10599 1398
rect 10565 1292 10599 1326
rect 10565 1220 10599 1254
rect 10565 1148 10599 1182
rect 10565 1076 10599 1110
rect 9603 1004 9637 1038
rect 9603 932 9637 966
rect 11527 1436 11561 1470
rect 11527 1364 11561 1398
rect 11527 1292 11561 1326
rect 11527 1220 11561 1254
rect 11527 1148 11561 1182
rect 11527 1076 11561 1110
rect 10565 1004 10599 1038
rect 10565 932 10599 966
rect 12489 1436 12523 1470
rect 12489 1364 12523 1398
rect 12489 1292 12523 1326
rect 12489 1220 12523 1254
rect 12489 1148 12523 1182
rect 12489 1076 12523 1110
rect 11527 1004 11561 1038
rect 11527 932 11561 966
rect 13451 1436 13485 1470
rect 13451 1364 13485 1398
rect 13451 1292 13485 1326
rect 13451 1220 13485 1254
rect 13451 1148 13485 1182
rect 13451 1076 13485 1110
rect 12489 1004 12523 1038
rect 12489 932 12523 966
rect 14413 1436 14447 1470
rect 14413 1364 14447 1398
rect 14413 1292 14447 1326
rect 14413 1220 14447 1254
rect 14413 1148 14447 1182
rect 14413 1076 14447 1110
rect 13451 1004 13485 1038
rect 13451 932 13485 966
rect 15375 1436 15409 1470
rect 15375 1364 15409 1398
rect 15375 1292 15409 1326
rect 15375 1220 15409 1254
rect 15375 1148 15409 1182
rect 15375 1076 15409 1110
rect 14413 1004 14447 1038
rect 14413 932 14447 966
rect 16337 1436 16371 1470
rect 16337 1364 16371 1398
rect 16337 1292 16371 1326
rect 16337 1220 16371 1254
rect 16337 1148 16371 1182
rect 16337 1076 16371 1110
rect 15375 1004 15409 1038
rect 15375 932 15409 966
rect 17299 1436 17333 1470
rect 17299 1364 17333 1398
rect 17299 1292 17333 1326
rect 17299 1220 17333 1254
rect 17299 1148 17333 1182
rect 17299 1076 17333 1110
rect 16337 1004 16371 1038
rect 16337 932 16371 966
rect 17965 1436 17999 1470
rect 17965 1364 17999 1398
rect 17965 1292 17999 1326
rect 17965 1220 17999 1254
rect 17965 1148 17999 1182
rect 17965 1076 17999 1110
rect 17299 1004 17333 1038
rect 17299 932 17333 966
rect 18631 1436 18665 1470
rect 18631 1364 18665 1398
rect 18631 1292 18665 1326
rect 18631 1220 18665 1254
rect 18631 1148 18665 1182
rect 18631 1076 18665 1110
rect 17965 1004 17999 1038
rect 17965 932 17999 966
rect 19297 1436 19331 1470
rect 19297 1364 19331 1398
rect 19297 1292 19331 1326
rect 19297 1220 19331 1254
rect 19297 1148 19331 1182
rect 19297 1076 19331 1110
rect 18631 1004 18665 1038
rect 18631 932 18665 966
rect 19297 1004 19331 1038
rect 19297 932 19331 966
<< poly >>
rect 247 1450 277 1476
rect 335 1450 365 1476
rect 423 1450 453 1476
rect 511 1450 541 1476
rect 599 1450 629 1476
rect 687 1450 717 1476
rect 1209 1450 1239 1476
rect 1297 1450 1327 1476
rect 1385 1450 1415 1476
rect 1473 1450 1503 1476
rect 1561 1450 1591 1476
rect 1649 1450 1679 1476
rect 247 1019 277 1050
rect 335 1019 365 1050
rect 423 1019 453 1050
rect 511 1019 541 1050
rect 195 1003 365 1019
rect 195 969 205 1003
rect 239 989 365 1003
rect 417 1003 541 1019
rect 239 969 249 989
rect 195 953 249 969
rect 417 969 427 1003
rect 461 989 541 1003
rect 599 1019 629 1050
rect 687 1019 717 1050
rect 599 1003 717 1019
rect 599 989 649 1003
rect 461 969 471 989
rect 417 953 471 969
rect 639 969 649 989
rect 683 989 717 1003
rect 2171 1450 2201 1476
rect 2259 1450 2289 1476
rect 2347 1450 2377 1476
rect 2435 1450 2465 1476
rect 2523 1450 2553 1476
rect 2611 1450 2641 1476
rect 1209 1019 1239 1050
rect 1297 1019 1327 1050
rect 1385 1019 1415 1050
rect 1473 1019 1503 1050
rect 683 969 693 989
rect 639 953 693 969
rect 1157 1003 1327 1019
rect 1157 969 1167 1003
rect 1201 989 1327 1003
rect 1379 1003 1503 1019
rect 1201 969 1211 989
rect 1157 953 1211 969
rect 1379 969 1389 1003
rect 1423 989 1503 1003
rect 1561 1019 1591 1050
rect 1649 1019 1679 1050
rect 1561 1003 1679 1019
rect 1561 989 1611 1003
rect 1423 969 1433 989
rect 1379 953 1433 969
rect 1601 969 1611 989
rect 1645 989 1679 1003
rect 3133 1450 3163 1476
rect 3221 1450 3251 1476
rect 3309 1450 3339 1476
rect 3397 1450 3427 1476
rect 3485 1450 3515 1476
rect 3573 1450 3603 1476
rect 2171 1019 2201 1050
rect 2259 1019 2289 1050
rect 2347 1019 2377 1050
rect 2435 1019 2465 1050
rect 1645 969 1655 989
rect 1601 953 1655 969
rect 2119 1003 2289 1019
rect 2119 969 2129 1003
rect 2163 989 2289 1003
rect 2341 1003 2465 1019
rect 2163 969 2173 989
rect 2119 953 2173 969
rect 2341 969 2351 1003
rect 2385 989 2465 1003
rect 2523 1019 2553 1050
rect 2611 1019 2641 1050
rect 2523 1003 2641 1019
rect 2523 989 2573 1003
rect 2385 969 2395 989
rect 2341 953 2395 969
rect 2563 969 2573 989
rect 2607 989 2641 1003
rect 4095 1450 4125 1476
rect 4183 1450 4213 1476
rect 4271 1450 4301 1476
rect 4359 1450 4389 1476
rect 4447 1450 4477 1476
rect 4535 1450 4565 1476
rect 3133 1019 3163 1050
rect 3221 1019 3251 1050
rect 3309 1019 3339 1050
rect 3397 1019 3427 1050
rect 2607 969 2617 989
rect 2563 953 2617 969
rect 3081 1003 3251 1019
rect 3081 969 3091 1003
rect 3125 989 3251 1003
rect 3303 1003 3427 1019
rect 3125 969 3135 989
rect 3081 953 3135 969
rect 3303 969 3313 1003
rect 3347 989 3427 1003
rect 3485 1019 3515 1050
rect 3573 1019 3603 1050
rect 3485 1003 3603 1019
rect 3485 989 3535 1003
rect 3347 969 3357 989
rect 3303 953 3357 969
rect 3525 969 3535 989
rect 3569 989 3603 1003
rect 5057 1450 5087 1476
rect 5145 1450 5175 1476
rect 5233 1450 5263 1476
rect 5321 1450 5351 1476
rect 5409 1450 5439 1476
rect 5497 1450 5527 1476
rect 4095 1019 4125 1050
rect 4183 1019 4213 1050
rect 4271 1019 4301 1050
rect 4359 1019 4389 1050
rect 3569 969 3579 989
rect 3525 953 3579 969
rect 4043 1003 4213 1019
rect 4043 969 4053 1003
rect 4087 989 4213 1003
rect 4265 1003 4389 1019
rect 4087 969 4097 989
rect 4043 953 4097 969
rect 4265 969 4275 1003
rect 4309 989 4389 1003
rect 4447 1019 4477 1050
rect 4535 1019 4565 1050
rect 4447 1003 4565 1019
rect 4447 989 4497 1003
rect 4309 969 4319 989
rect 4265 953 4319 969
rect 4487 969 4497 989
rect 4531 989 4565 1003
rect 6019 1450 6049 1476
rect 6107 1450 6137 1476
rect 6195 1450 6225 1476
rect 6283 1450 6313 1476
rect 6371 1450 6401 1476
rect 6459 1450 6489 1476
rect 5057 1019 5087 1050
rect 5145 1019 5175 1050
rect 5233 1019 5263 1050
rect 5321 1019 5351 1050
rect 4531 969 4541 989
rect 4487 953 4541 969
rect 5005 1003 5175 1019
rect 5005 969 5015 1003
rect 5049 989 5175 1003
rect 5227 1003 5351 1019
rect 5049 969 5059 989
rect 5005 953 5059 969
rect 5227 969 5237 1003
rect 5271 989 5351 1003
rect 5409 1019 5439 1050
rect 5497 1019 5527 1050
rect 5409 1003 5527 1019
rect 5409 989 5459 1003
rect 5271 969 5281 989
rect 5227 953 5281 969
rect 5449 969 5459 989
rect 5493 989 5527 1003
rect 6981 1450 7011 1476
rect 7069 1450 7099 1476
rect 7157 1450 7187 1476
rect 7245 1450 7275 1476
rect 7333 1450 7363 1476
rect 7421 1450 7451 1476
rect 6019 1019 6049 1050
rect 6107 1019 6137 1050
rect 6195 1019 6225 1050
rect 6283 1019 6313 1050
rect 5493 969 5503 989
rect 5449 953 5503 969
rect 5967 1003 6137 1019
rect 5967 969 5977 1003
rect 6011 989 6137 1003
rect 6189 1003 6313 1019
rect 6011 969 6021 989
rect 5967 953 6021 969
rect 6189 969 6199 1003
rect 6233 989 6313 1003
rect 6371 1019 6401 1050
rect 6459 1019 6489 1050
rect 6371 1003 6489 1019
rect 6371 989 6421 1003
rect 6233 969 6243 989
rect 6189 953 6243 969
rect 6411 969 6421 989
rect 6455 989 6489 1003
rect 7943 1450 7973 1476
rect 8031 1450 8061 1476
rect 8119 1450 8149 1476
rect 8207 1450 8237 1476
rect 8295 1450 8325 1476
rect 8383 1450 8413 1476
rect 6981 1019 7011 1050
rect 7069 1019 7099 1050
rect 7157 1019 7187 1050
rect 7245 1019 7275 1050
rect 6455 969 6465 989
rect 6411 953 6465 969
rect 6929 1003 7099 1019
rect 6929 969 6939 1003
rect 6973 989 7099 1003
rect 7151 1003 7275 1019
rect 6973 969 6983 989
rect 6929 953 6983 969
rect 7151 969 7161 1003
rect 7195 989 7275 1003
rect 7333 1019 7363 1050
rect 7421 1019 7451 1050
rect 7333 1003 7451 1019
rect 7333 989 7383 1003
rect 7195 969 7205 989
rect 7151 953 7205 969
rect 7373 969 7383 989
rect 7417 989 7451 1003
rect 8905 1450 8935 1476
rect 8993 1450 9023 1476
rect 9081 1450 9111 1476
rect 9169 1450 9199 1476
rect 9257 1450 9287 1476
rect 9345 1450 9375 1476
rect 7943 1019 7973 1050
rect 8031 1019 8061 1050
rect 8119 1019 8149 1050
rect 8207 1019 8237 1050
rect 7417 969 7427 989
rect 7373 953 7427 969
rect 7891 1003 8061 1019
rect 7891 969 7901 1003
rect 7935 989 8061 1003
rect 8113 1003 8237 1019
rect 7935 969 7945 989
rect 7891 953 7945 969
rect 8113 969 8123 1003
rect 8157 989 8237 1003
rect 8295 1019 8325 1050
rect 8383 1019 8413 1050
rect 8295 1003 8413 1019
rect 8295 989 8345 1003
rect 8157 969 8167 989
rect 8113 953 8167 969
rect 8335 969 8345 989
rect 8379 989 8413 1003
rect 9867 1450 9897 1476
rect 9955 1450 9985 1476
rect 10043 1450 10073 1476
rect 10131 1450 10161 1476
rect 10219 1450 10249 1476
rect 10307 1450 10337 1476
rect 8905 1019 8935 1050
rect 8993 1019 9023 1050
rect 9081 1019 9111 1050
rect 9169 1019 9199 1050
rect 8379 969 8389 989
rect 8335 953 8389 969
rect 8853 1003 9023 1019
rect 8853 969 8863 1003
rect 8897 989 9023 1003
rect 9075 1003 9199 1019
rect 8897 969 8907 989
rect 8853 953 8907 969
rect 9075 969 9085 1003
rect 9119 989 9199 1003
rect 9257 1019 9287 1050
rect 9345 1019 9375 1050
rect 9257 1003 9375 1019
rect 9257 989 9307 1003
rect 9119 969 9129 989
rect 9075 953 9129 969
rect 9297 969 9307 989
rect 9341 989 9375 1003
rect 10829 1450 10859 1476
rect 10917 1450 10947 1476
rect 11005 1450 11035 1476
rect 11093 1450 11123 1476
rect 11181 1450 11211 1476
rect 11269 1450 11299 1476
rect 9867 1019 9897 1050
rect 9955 1019 9985 1050
rect 10043 1019 10073 1050
rect 10131 1019 10161 1050
rect 9341 969 9351 989
rect 9297 953 9351 969
rect 9815 1003 9985 1019
rect 9815 969 9825 1003
rect 9859 989 9985 1003
rect 10037 1003 10161 1019
rect 9859 969 9869 989
rect 9815 953 9869 969
rect 10037 969 10047 1003
rect 10081 989 10161 1003
rect 10219 1019 10249 1050
rect 10307 1019 10337 1050
rect 10219 1003 10337 1019
rect 10219 989 10269 1003
rect 10081 969 10091 989
rect 10037 953 10091 969
rect 10259 969 10269 989
rect 10303 989 10337 1003
rect 11791 1450 11821 1476
rect 11879 1450 11909 1476
rect 11967 1450 11997 1476
rect 12055 1450 12085 1476
rect 12143 1450 12173 1476
rect 12231 1450 12261 1476
rect 10829 1019 10859 1050
rect 10917 1019 10947 1050
rect 11005 1019 11035 1050
rect 11093 1019 11123 1050
rect 10303 969 10313 989
rect 10259 953 10313 969
rect 10777 1003 10947 1019
rect 10777 969 10787 1003
rect 10821 989 10947 1003
rect 10999 1003 11123 1019
rect 10821 969 10831 989
rect 10777 953 10831 969
rect 10999 969 11009 1003
rect 11043 989 11123 1003
rect 11181 1019 11211 1050
rect 11269 1019 11299 1050
rect 11181 1003 11299 1019
rect 11181 989 11231 1003
rect 11043 969 11053 989
rect 10999 953 11053 969
rect 11221 969 11231 989
rect 11265 989 11299 1003
rect 12753 1450 12783 1476
rect 12841 1450 12871 1476
rect 12929 1450 12959 1476
rect 13017 1450 13047 1476
rect 13105 1450 13135 1476
rect 13193 1450 13223 1476
rect 11791 1019 11821 1050
rect 11879 1019 11909 1050
rect 11967 1019 11997 1050
rect 12055 1019 12085 1050
rect 11265 969 11275 989
rect 11221 953 11275 969
rect 11739 1003 11909 1019
rect 11739 969 11749 1003
rect 11783 989 11909 1003
rect 11961 1003 12085 1019
rect 11783 969 11793 989
rect 11739 953 11793 969
rect 11961 969 11971 1003
rect 12005 989 12085 1003
rect 12143 1019 12173 1050
rect 12231 1019 12261 1050
rect 12143 1003 12261 1019
rect 12143 989 12193 1003
rect 12005 969 12015 989
rect 11961 953 12015 969
rect 12183 969 12193 989
rect 12227 989 12261 1003
rect 13715 1450 13745 1476
rect 13803 1450 13833 1476
rect 13891 1450 13921 1476
rect 13979 1450 14009 1476
rect 14067 1450 14097 1476
rect 14155 1450 14185 1476
rect 12753 1019 12783 1050
rect 12841 1019 12871 1050
rect 12929 1019 12959 1050
rect 13017 1019 13047 1050
rect 12227 969 12237 989
rect 12183 953 12237 969
rect 12701 1003 12871 1019
rect 12701 969 12711 1003
rect 12745 989 12871 1003
rect 12923 1003 13047 1019
rect 12745 969 12755 989
rect 12701 953 12755 969
rect 12923 969 12933 1003
rect 12967 989 13047 1003
rect 13105 1019 13135 1050
rect 13193 1019 13223 1050
rect 13105 1003 13223 1019
rect 13105 989 13155 1003
rect 12967 969 12977 989
rect 12923 953 12977 969
rect 13145 969 13155 989
rect 13189 989 13223 1003
rect 14677 1450 14707 1476
rect 14765 1450 14795 1476
rect 14853 1450 14883 1476
rect 14941 1450 14971 1476
rect 15029 1450 15059 1476
rect 15117 1450 15147 1476
rect 13715 1019 13745 1050
rect 13803 1019 13833 1050
rect 13891 1019 13921 1050
rect 13979 1019 14009 1050
rect 13189 969 13199 989
rect 13145 953 13199 969
rect 13663 1003 13833 1019
rect 13663 969 13673 1003
rect 13707 989 13833 1003
rect 13885 1003 14009 1019
rect 13707 969 13717 989
rect 13663 953 13717 969
rect 13885 969 13895 1003
rect 13929 989 14009 1003
rect 14067 1019 14097 1050
rect 14155 1019 14185 1050
rect 14067 1003 14185 1019
rect 14067 989 14117 1003
rect 13929 969 13939 989
rect 13885 953 13939 969
rect 14107 969 14117 989
rect 14151 989 14185 1003
rect 15639 1450 15669 1476
rect 15727 1450 15757 1476
rect 15815 1450 15845 1476
rect 15903 1450 15933 1476
rect 15991 1450 16021 1476
rect 16079 1450 16109 1476
rect 14677 1019 14707 1050
rect 14765 1019 14795 1050
rect 14853 1019 14883 1050
rect 14941 1019 14971 1050
rect 14151 969 14161 989
rect 14107 953 14161 969
rect 14625 1003 14795 1019
rect 14625 969 14635 1003
rect 14669 989 14795 1003
rect 14847 1003 14971 1019
rect 14669 969 14679 989
rect 14625 953 14679 969
rect 14847 969 14857 1003
rect 14891 989 14971 1003
rect 15029 1019 15059 1050
rect 15117 1019 15147 1050
rect 15029 1003 15147 1019
rect 15029 989 15079 1003
rect 14891 969 14901 989
rect 14847 953 14901 969
rect 15069 969 15079 989
rect 15113 989 15147 1003
rect 16601 1450 16631 1476
rect 16689 1450 16719 1476
rect 16777 1450 16807 1476
rect 16865 1450 16895 1476
rect 16953 1450 16983 1476
rect 17041 1450 17071 1476
rect 15639 1019 15669 1050
rect 15727 1019 15757 1050
rect 15815 1019 15845 1050
rect 15903 1019 15933 1050
rect 15113 969 15123 989
rect 15069 953 15123 969
rect 15587 1003 15757 1019
rect 15587 969 15597 1003
rect 15631 989 15757 1003
rect 15809 1003 15933 1019
rect 15631 969 15641 989
rect 15587 953 15641 969
rect 15809 969 15819 1003
rect 15853 989 15933 1003
rect 15991 1019 16021 1050
rect 16079 1019 16109 1050
rect 15991 1003 16109 1019
rect 15991 989 16041 1003
rect 15853 969 15863 989
rect 15809 953 15863 969
rect 16031 969 16041 989
rect 16075 989 16109 1003
rect 17503 1451 17533 1477
rect 17591 1451 17621 1477
rect 17679 1451 17709 1477
rect 17767 1451 17797 1477
rect 16601 1019 16631 1050
rect 16689 1019 16719 1050
rect 16777 1019 16807 1050
rect 16865 1019 16895 1050
rect 16075 969 16085 989
rect 16031 953 16085 969
rect 16549 1003 16719 1019
rect 16549 969 16559 1003
rect 16593 989 16719 1003
rect 16771 1003 16895 1019
rect 16593 969 16603 989
rect 16549 953 16603 969
rect 16771 969 16781 1003
rect 16815 989 16895 1003
rect 16953 1019 16983 1050
rect 17041 1019 17071 1050
rect 16953 1003 17071 1019
rect 16953 989 17003 1003
rect 16815 969 16825 989
rect 16771 953 16825 969
rect 16993 969 17003 989
rect 17037 989 17071 1003
rect 18167 1451 18197 1477
rect 18255 1451 18285 1477
rect 18343 1451 18373 1477
rect 18431 1451 18461 1477
rect 17503 1020 17533 1051
rect 17591 1020 17621 1051
rect 17679 1020 17709 1051
rect 17767 1020 17797 1051
rect 17037 969 17047 989
rect 16993 953 17047 969
rect 17437 1004 17621 1020
rect 17437 970 17447 1004
rect 17481 990 17621 1004
rect 17667 1004 17797 1020
rect 17481 970 17491 990
rect 17437 954 17491 970
rect 17667 970 17677 1004
rect 17711 990 17797 1004
rect 18835 1451 18865 1477
rect 18923 1451 18953 1477
rect 19011 1451 19041 1477
rect 19099 1451 19129 1477
rect 17711 970 17721 990
rect 17667 954 17721 970
rect 18167 1020 18197 1051
rect 18255 1020 18285 1051
rect 18167 1004 18285 1020
rect 18167 990 18187 1004
rect 18177 970 18187 990
rect 18221 990 18285 1004
rect 18343 1020 18373 1051
rect 18431 1020 18461 1051
rect 18343 1004 18527 1020
rect 18343 990 18483 1004
rect 18221 970 18231 990
rect 18177 954 18231 970
rect 18473 970 18483 990
rect 18517 970 18527 1004
rect 18473 954 18527 970
rect 18835 1020 18865 1051
rect 18923 1020 18953 1051
rect 19011 1020 19041 1051
rect 19099 1020 19129 1051
rect 18769 1004 18953 1020
rect 18769 970 18779 1004
rect 18813 990 18953 1004
rect 18995 1004 19129 1020
rect 18813 970 18823 990
rect 18769 954 18823 970
rect 18995 970 19005 1004
rect 19039 990 19129 1004
rect 19039 970 19049 990
rect 18995 954 19049 970
rect 195 461 249 477
rect 195 441 205 461
rect 147 427 205 441
rect 239 427 249 461
rect 147 411 249 427
rect 417 461 471 477
rect 417 427 427 461
rect 461 441 471 461
rect 639 461 693 477
rect 461 427 477 441
rect 417 411 477 427
rect 639 427 649 461
rect 683 427 693 461
rect 639 411 693 427
rect 1157 461 1211 477
rect 1157 441 1167 461
rect 147 379 177 411
rect 447 379 477 411
rect 649 379 679 411
rect 1109 427 1167 441
rect 1201 427 1211 461
rect 1109 411 1211 427
rect 1379 461 1433 477
rect 1379 427 1389 461
rect 1423 441 1433 461
rect 1601 461 1655 477
rect 1423 427 1439 441
rect 1379 411 1439 427
rect 1601 427 1611 461
rect 1645 427 1655 461
rect 1601 411 1655 427
rect 2119 461 2173 477
rect 2119 441 2129 461
rect 1109 379 1139 411
rect 1409 379 1439 411
rect 1611 379 1641 411
rect 2071 427 2129 441
rect 2163 427 2173 461
rect 2071 411 2173 427
rect 2341 461 2395 477
rect 2341 427 2351 461
rect 2385 441 2395 461
rect 2563 461 2617 477
rect 2385 427 2401 441
rect 2341 411 2401 427
rect 2563 427 2573 461
rect 2607 427 2617 461
rect 2563 411 2617 427
rect 3081 461 3135 477
rect 3081 441 3091 461
rect 2071 379 2101 411
rect 2371 379 2401 411
rect 2573 379 2603 411
rect 3033 427 3091 441
rect 3125 427 3135 461
rect 3033 411 3135 427
rect 3303 461 3357 477
rect 3303 427 3313 461
rect 3347 441 3357 461
rect 3525 461 3579 477
rect 3347 427 3363 441
rect 3303 411 3363 427
rect 3525 427 3535 461
rect 3569 427 3579 461
rect 3525 411 3579 427
rect 4043 461 4097 477
rect 4043 441 4053 461
rect 3033 379 3063 411
rect 3333 379 3363 411
rect 3535 379 3565 411
rect 3995 427 4053 441
rect 4087 427 4097 461
rect 3995 411 4097 427
rect 4265 461 4319 477
rect 4265 427 4275 461
rect 4309 441 4319 461
rect 4487 461 4541 477
rect 4309 427 4325 441
rect 4265 411 4325 427
rect 4487 427 4497 461
rect 4531 427 4541 461
rect 4487 411 4541 427
rect 5005 461 5059 477
rect 5005 441 5015 461
rect 3995 379 4025 411
rect 4295 379 4325 411
rect 4497 379 4527 411
rect 4957 427 5015 441
rect 5049 427 5059 461
rect 4957 411 5059 427
rect 5227 461 5281 477
rect 5227 427 5237 461
rect 5271 441 5281 461
rect 5449 461 5503 477
rect 5271 427 5287 441
rect 5227 411 5287 427
rect 5449 427 5459 461
rect 5493 427 5503 461
rect 5449 411 5503 427
rect 5967 461 6021 477
rect 5967 441 5977 461
rect 4957 379 4987 411
rect 5257 379 5287 411
rect 5459 379 5489 411
rect 5919 427 5977 441
rect 6011 427 6021 461
rect 5919 411 6021 427
rect 6189 461 6243 477
rect 6189 427 6199 461
rect 6233 441 6243 461
rect 6411 461 6465 477
rect 6233 427 6249 441
rect 6189 411 6249 427
rect 6411 427 6421 461
rect 6455 427 6465 461
rect 6411 411 6465 427
rect 6929 461 6983 477
rect 6929 441 6939 461
rect 5919 379 5949 411
rect 6219 379 6249 411
rect 6421 379 6451 411
rect 6881 427 6939 441
rect 6973 427 6983 461
rect 6881 411 6983 427
rect 7151 461 7205 477
rect 7151 427 7161 461
rect 7195 441 7205 461
rect 7373 461 7427 477
rect 7195 427 7211 441
rect 7151 411 7211 427
rect 7373 427 7383 461
rect 7417 427 7427 461
rect 7373 411 7427 427
rect 7891 461 7945 477
rect 7891 441 7901 461
rect 6881 379 6911 411
rect 7181 379 7211 411
rect 7383 379 7413 411
rect 7843 427 7901 441
rect 7935 427 7945 461
rect 7843 411 7945 427
rect 8113 461 8167 477
rect 8113 427 8123 461
rect 8157 441 8167 461
rect 8335 461 8389 477
rect 8157 427 8173 441
rect 8113 411 8173 427
rect 8335 427 8345 461
rect 8379 427 8389 461
rect 8335 411 8389 427
rect 8853 461 8907 477
rect 8853 441 8863 461
rect 7843 379 7873 411
rect 8143 379 8173 411
rect 8345 379 8375 411
rect 8805 427 8863 441
rect 8897 427 8907 461
rect 8805 411 8907 427
rect 9075 461 9129 477
rect 9075 427 9085 461
rect 9119 441 9129 461
rect 9297 461 9351 477
rect 9119 427 9135 441
rect 9075 411 9135 427
rect 9297 427 9307 461
rect 9341 427 9351 461
rect 9297 411 9351 427
rect 9815 461 9869 477
rect 9815 441 9825 461
rect 8805 379 8835 411
rect 9105 379 9135 411
rect 9307 379 9337 411
rect 9767 427 9825 441
rect 9859 427 9869 461
rect 9767 411 9869 427
rect 10037 461 10091 477
rect 10037 427 10047 461
rect 10081 441 10091 461
rect 10259 461 10313 477
rect 10081 427 10097 441
rect 10037 411 10097 427
rect 10259 427 10269 461
rect 10303 427 10313 461
rect 10259 411 10313 427
rect 10777 461 10831 477
rect 10777 441 10787 461
rect 9767 379 9797 411
rect 10067 379 10097 411
rect 10269 379 10299 411
rect 10729 427 10787 441
rect 10821 427 10831 461
rect 10729 411 10831 427
rect 10999 461 11053 477
rect 10999 427 11009 461
rect 11043 441 11053 461
rect 11221 461 11275 477
rect 11043 427 11059 441
rect 10999 411 11059 427
rect 11221 427 11231 461
rect 11265 427 11275 461
rect 11221 411 11275 427
rect 11739 461 11793 477
rect 11739 441 11749 461
rect 10729 379 10759 411
rect 11029 379 11059 411
rect 11231 379 11261 411
rect 11691 427 11749 441
rect 11783 427 11793 461
rect 11691 411 11793 427
rect 11961 461 12015 477
rect 11961 427 11971 461
rect 12005 441 12015 461
rect 12183 461 12237 477
rect 12005 427 12021 441
rect 11961 411 12021 427
rect 12183 427 12193 461
rect 12227 427 12237 461
rect 12183 411 12237 427
rect 12701 461 12755 477
rect 12701 441 12711 461
rect 11691 379 11721 411
rect 11991 379 12021 411
rect 12193 379 12223 411
rect 12653 427 12711 441
rect 12745 427 12755 461
rect 12653 411 12755 427
rect 12923 461 12977 477
rect 12923 427 12933 461
rect 12967 441 12977 461
rect 13145 461 13199 477
rect 12967 427 12983 441
rect 12923 411 12983 427
rect 13145 427 13155 461
rect 13189 427 13199 461
rect 13145 411 13199 427
rect 13663 461 13717 477
rect 13663 441 13673 461
rect 12653 379 12683 411
rect 12953 379 12983 411
rect 13155 379 13185 411
rect 13615 427 13673 441
rect 13707 427 13717 461
rect 13615 411 13717 427
rect 13885 461 13939 477
rect 13885 427 13895 461
rect 13929 441 13939 461
rect 14107 461 14161 477
rect 13929 427 13945 441
rect 13885 411 13945 427
rect 14107 427 14117 461
rect 14151 427 14161 461
rect 14107 411 14161 427
rect 14625 461 14679 477
rect 14625 441 14635 461
rect 13615 379 13645 411
rect 13915 379 13945 411
rect 14117 379 14147 411
rect 14577 427 14635 441
rect 14669 427 14679 461
rect 14577 411 14679 427
rect 14847 461 14901 477
rect 14847 427 14857 461
rect 14891 441 14901 461
rect 15069 461 15123 477
rect 14891 427 14907 441
rect 14847 411 14907 427
rect 15069 427 15079 461
rect 15113 427 15123 461
rect 15069 411 15123 427
rect 15587 461 15641 477
rect 15587 441 15597 461
rect 14577 379 14607 411
rect 14877 379 14907 411
rect 15079 379 15109 411
rect 15539 427 15597 441
rect 15631 427 15641 461
rect 15539 411 15641 427
rect 15809 461 15863 477
rect 15809 427 15819 461
rect 15853 441 15863 461
rect 16031 461 16085 477
rect 15853 427 15869 441
rect 15809 411 15869 427
rect 16031 427 16041 461
rect 16075 427 16085 461
rect 16031 411 16085 427
rect 16549 461 16603 477
rect 16549 441 16559 461
rect 15539 379 15569 411
rect 15839 379 15869 411
rect 16041 379 16071 411
rect 16501 427 16559 441
rect 16593 427 16603 461
rect 16501 411 16603 427
rect 16771 461 16825 477
rect 16771 427 16781 461
rect 16815 441 16825 461
rect 16993 461 17047 477
rect 16815 427 16831 441
rect 16771 411 16831 427
rect 16993 427 17003 461
rect 17037 427 17047 461
rect 16993 411 17047 427
rect 16501 379 16531 411
rect 16801 379 16831 411
rect 17003 379 17033 411
rect 17437 461 17491 477
rect 17437 427 17447 461
rect 17481 441 17491 461
rect 17659 461 17713 477
rect 17481 427 17514 441
rect 17437 411 17514 427
rect 17659 427 17669 461
rect 17703 427 17713 461
rect 17659 411 17713 427
rect 18177 461 18231 477
rect 18177 441 18187 461
rect 17484 377 17514 411
rect 17678 377 17708 411
rect 18150 427 18187 441
rect 18221 427 18231 461
rect 18473 461 18527 477
rect 18473 441 18483 461
rect 18150 411 18231 427
rect 18450 427 18483 441
rect 18517 427 18527 461
rect 18450 411 18527 427
rect 18150 377 18180 411
rect 18450 377 18480 411
rect 18769 461 18823 477
rect 18769 427 18779 461
rect 18813 441 18823 461
rect 18991 461 19045 477
rect 18813 427 18846 441
rect 18769 411 18846 427
rect 18991 427 19001 461
rect 19035 427 19045 461
rect 18991 411 19045 427
rect 18816 377 18846 411
rect 19010 377 19040 411
<< polycont >>
rect 205 969 239 1003
rect 427 969 461 1003
rect 649 969 683 1003
rect 1167 969 1201 1003
rect 1389 969 1423 1003
rect 1611 969 1645 1003
rect 2129 969 2163 1003
rect 2351 969 2385 1003
rect 2573 969 2607 1003
rect 3091 969 3125 1003
rect 3313 969 3347 1003
rect 3535 969 3569 1003
rect 4053 969 4087 1003
rect 4275 969 4309 1003
rect 4497 969 4531 1003
rect 5015 969 5049 1003
rect 5237 969 5271 1003
rect 5459 969 5493 1003
rect 5977 969 6011 1003
rect 6199 969 6233 1003
rect 6421 969 6455 1003
rect 6939 969 6973 1003
rect 7161 969 7195 1003
rect 7383 969 7417 1003
rect 7901 969 7935 1003
rect 8123 969 8157 1003
rect 8345 969 8379 1003
rect 8863 969 8897 1003
rect 9085 969 9119 1003
rect 9307 969 9341 1003
rect 9825 969 9859 1003
rect 10047 969 10081 1003
rect 10269 969 10303 1003
rect 10787 969 10821 1003
rect 11009 969 11043 1003
rect 11231 969 11265 1003
rect 11749 969 11783 1003
rect 11971 969 12005 1003
rect 12193 969 12227 1003
rect 12711 969 12745 1003
rect 12933 969 12967 1003
rect 13155 969 13189 1003
rect 13673 969 13707 1003
rect 13895 969 13929 1003
rect 14117 969 14151 1003
rect 14635 969 14669 1003
rect 14857 969 14891 1003
rect 15079 969 15113 1003
rect 15597 969 15631 1003
rect 15819 969 15853 1003
rect 16041 969 16075 1003
rect 16559 969 16593 1003
rect 16781 969 16815 1003
rect 17003 969 17037 1003
rect 17447 970 17481 1004
rect 17677 970 17711 1004
rect 18187 970 18221 1004
rect 18483 970 18517 1004
rect 18779 970 18813 1004
rect 19005 970 19039 1004
rect 205 427 239 461
rect 427 427 461 461
rect 649 427 683 461
rect 1167 427 1201 461
rect 1389 427 1423 461
rect 1611 427 1645 461
rect 2129 427 2163 461
rect 2351 427 2385 461
rect 2573 427 2607 461
rect 3091 427 3125 461
rect 3313 427 3347 461
rect 3535 427 3569 461
rect 4053 427 4087 461
rect 4275 427 4309 461
rect 4497 427 4531 461
rect 5015 427 5049 461
rect 5237 427 5271 461
rect 5459 427 5493 461
rect 5977 427 6011 461
rect 6199 427 6233 461
rect 6421 427 6455 461
rect 6939 427 6973 461
rect 7161 427 7195 461
rect 7383 427 7417 461
rect 7901 427 7935 461
rect 8123 427 8157 461
rect 8345 427 8379 461
rect 8863 427 8897 461
rect 9085 427 9119 461
rect 9307 427 9341 461
rect 9825 427 9859 461
rect 10047 427 10081 461
rect 10269 427 10303 461
rect 10787 427 10821 461
rect 11009 427 11043 461
rect 11231 427 11265 461
rect 11749 427 11783 461
rect 11971 427 12005 461
rect 12193 427 12227 461
rect 12711 427 12745 461
rect 12933 427 12967 461
rect 13155 427 13189 461
rect 13673 427 13707 461
rect 13895 427 13929 461
rect 14117 427 14151 461
rect 14635 427 14669 461
rect 14857 427 14891 461
rect 15079 427 15113 461
rect 15597 427 15631 461
rect 15819 427 15853 461
rect 16041 427 16075 461
rect 16559 427 16593 461
rect 16781 427 16815 461
rect 17003 427 17037 461
rect 17447 427 17481 461
rect 17669 427 17703 461
rect 18187 427 18221 461
rect 18483 427 18517 461
rect 18779 427 18813 461
rect 19001 427 19035 461
<< locali >>
rect -31 1539 19345 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 343 1539
rect 377 1505 415 1539
rect 449 1505 513 1539
rect 547 1505 585 1539
rect 619 1505 657 1539
rect 691 1505 729 1539
rect 763 1505 801 1539
rect 835 1505 873 1539
rect 907 1505 1017 1539
rect 1051 1505 1089 1539
rect 1123 1505 1161 1539
rect 1195 1505 1233 1539
rect 1267 1505 1305 1539
rect 1339 1505 1377 1539
rect 1411 1505 1475 1539
rect 1509 1505 1547 1539
rect 1581 1505 1619 1539
rect 1653 1505 1691 1539
rect 1725 1505 1763 1539
rect 1797 1505 1835 1539
rect 1869 1505 1979 1539
rect 2013 1505 2051 1539
rect 2085 1505 2123 1539
rect 2157 1505 2195 1539
rect 2229 1505 2267 1539
rect 2301 1505 2339 1539
rect 2373 1505 2437 1539
rect 2471 1505 2509 1539
rect 2543 1505 2581 1539
rect 2615 1505 2653 1539
rect 2687 1505 2725 1539
rect 2759 1505 2797 1539
rect 2831 1505 2941 1539
rect 2975 1505 3013 1539
rect 3047 1505 3085 1539
rect 3119 1505 3157 1539
rect 3191 1505 3229 1539
rect 3263 1505 3301 1539
rect 3335 1505 3399 1539
rect 3433 1505 3471 1539
rect 3505 1505 3543 1539
rect 3577 1505 3615 1539
rect 3649 1505 3687 1539
rect 3721 1505 3759 1539
rect 3793 1505 3903 1539
rect 3937 1505 3975 1539
rect 4009 1505 4047 1539
rect 4081 1505 4119 1539
rect 4153 1505 4191 1539
rect 4225 1505 4263 1539
rect 4297 1505 4361 1539
rect 4395 1505 4433 1539
rect 4467 1505 4505 1539
rect 4539 1505 4577 1539
rect 4611 1505 4649 1539
rect 4683 1505 4721 1539
rect 4755 1505 4865 1539
rect 4899 1505 4937 1539
rect 4971 1505 5009 1539
rect 5043 1505 5081 1539
rect 5115 1505 5153 1539
rect 5187 1505 5225 1539
rect 5259 1505 5323 1539
rect 5357 1505 5395 1539
rect 5429 1505 5467 1539
rect 5501 1505 5539 1539
rect 5573 1505 5611 1539
rect 5645 1505 5683 1539
rect 5717 1505 5827 1539
rect 5861 1505 5899 1539
rect 5933 1505 5971 1539
rect 6005 1505 6043 1539
rect 6077 1505 6115 1539
rect 6149 1505 6187 1539
rect 6221 1505 6285 1539
rect 6319 1505 6357 1539
rect 6391 1505 6429 1539
rect 6463 1505 6501 1539
rect 6535 1505 6573 1539
rect 6607 1505 6645 1539
rect 6679 1505 6789 1539
rect 6823 1505 6861 1539
rect 6895 1505 6933 1539
rect 6967 1505 7005 1539
rect 7039 1505 7077 1539
rect 7111 1505 7149 1539
rect 7183 1505 7247 1539
rect 7281 1505 7319 1539
rect 7353 1505 7391 1539
rect 7425 1505 7463 1539
rect 7497 1505 7535 1539
rect 7569 1505 7607 1539
rect 7641 1505 7751 1539
rect 7785 1505 7823 1539
rect 7857 1505 7895 1539
rect 7929 1505 7967 1539
rect 8001 1505 8039 1539
rect 8073 1505 8111 1539
rect 8145 1505 8209 1539
rect 8243 1505 8281 1539
rect 8315 1505 8353 1539
rect 8387 1505 8425 1539
rect 8459 1505 8497 1539
rect 8531 1505 8569 1539
rect 8603 1505 8713 1539
rect 8747 1505 8785 1539
rect 8819 1505 8857 1539
rect 8891 1505 8929 1539
rect 8963 1505 9001 1539
rect 9035 1505 9073 1539
rect 9107 1505 9171 1539
rect 9205 1505 9243 1539
rect 9277 1505 9315 1539
rect 9349 1505 9387 1539
rect 9421 1505 9459 1539
rect 9493 1505 9531 1539
rect 9565 1505 9675 1539
rect 9709 1505 9747 1539
rect 9781 1505 9819 1539
rect 9853 1505 9891 1539
rect 9925 1505 9963 1539
rect 9997 1505 10035 1539
rect 10069 1505 10133 1539
rect 10167 1505 10205 1539
rect 10239 1505 10277 1539
rect 10311 1505 10349 1539
rect 10383 1505 10421 1539
rect 10455 1505 10493 1539
rect 10527 1505 10637 1539
rect 10671 1505 10709 1539
rect 10743 1505 10781 1539
rect 10815 1505 10853 1539
rect 10887 1505 10925 1539
rect 10959 1505 10997 1539
rect 11031 1505 11095 1539
rect 11129 1505 11167 1539
rect 11201 1505 11239 1539
rect 11273 1505 11311 1539
rect 11345 1505 11383 1539
rect 11417 1505 11455 1539
rect 11489 1505 11599 1539
rect 11633 1505 11671 1539
rect 11705 1505 11743 1539
rect 11777 1505 11815 1539
rect 11849 1505 11887 1539
rect 11921 1505 11959 1539
rect 11993 1505 12057 1539
rect 12091 1505 12129 1539
rect 12163 1505 12201 1539
rect 12235 1505 12273 1539
rect 12307 1505 12345 1539
rect 12379 1505 12417 1539
rect 12451 1505 12561 1539
rect 12595 1505 12633 1539
rect 12667 1505 12705 1539
rect 12739 1505 12777 1539
rect 12811 1505 12849 1539
rect 12883 1505 12921 1539
rect 12955 1505 13019 1539
rect 13053 1505 13091 1539
rect 13125 1505 13163 1539
rect 13197 1505 13235 1539
rect 13269 1505 13307 1539
rect 13341 1505 13379 1539
rect 13413 1505 13523 1539
rect 13557 1505 13595 1539
rect 13629 1505 13667 1539
rect 13701 1505 13739 1539
rect 13773 1505 13811 1539
rect 13845 1505 13883 1539
rect 13917 1505 13981 1539
rect 14015 1505 14053 1539
rect 14087 1505 14125 1539
rect 14159 1505 14197 1539
rect 14231 1505 14269 1539
rect 14303 1505 14341 1539
rect 14375 1505 14485 1539
rect 14519 1505 14557 1539
rect 14591 1505 14629 1539
rect 14663 1505 14701 1539
rect 14735 1505 14773 1539
rect 14807 1505 14845 1539
rect 14879 1505 14943 1539
rect 14977 1505 15015 1539
rect 15049 1505 15087 1539
rect 15121 1505 15159 1539
rect 15193 1505 15231 1539
rect 15265 1505 15303 1539
rect 15337 1505 15447 1539
rect 15481 1505 15519 1539
rect 15553 1505 15591 1539
rect 15625 1505 15663 1539
rect 15697 1505 15735 1539
rect 15769 1505 15807 1539
rect 15841 1505 15905 1539
rect 15939 1505 15977 1539
rect 16011 1505 16049 1539
rect 16083 1505 16121 1539
rect 16155 1505 16193 1539
rect 16227 1505 16265 1539
rect 16299 1505 16409 1539
rect 16443 1505 16481 1539
rect 16515 1505 16553 1539
rect 16587 1505 16625 1539
rect 16659 1505 16697 1539
rect 16731 1505 16769 1539
rect 16803 1505 16867 1539
rect 16901 1505 16939 1539
rect 16973 1505 17011 1539
rect 17045 1505 17083 1539
rect 17117 1505 17155 1539
rect 17189 1505 17227 1539
rect 17261 1505 17371 1539
rect 17405 1505 17443 1539
rect 17477 1505 17515 1539
rect 17549 1505 17587 1539
rect 17621 1505 17677 1539
rect 17711 1505 17749 1539
rect 17783 1505 17821 1539
rect 17855 1505 17893 1539
rect 17927 1505 18037 1539
rect 18071 1505 18109 1539
rect 18143 1505 18181 1539
rect 18215 1505 18253 1539
rect 18287 1505 18343 1539
rect 18377 1505 18415 1539
rect 18449 1505 18487 1539
rect 18521 1505 18559 1539
rect 18593 1505 18703 1539
rect 18737 1505 18775 1539
rect 18809 1505 18847 1539
rect 18881 1505 18919 1539
rect 18953 1505 19009 1539
rect 19043 1505 19081 1539
rect 19115 1505 19153 1539
rect 19187 1505 19225 1539
rect 19259 1505 19345 1539
rect -31 1492 19345 1505
rect -31 1470 31 1492
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect 201 1412 235 1492
rect 201 1344 235 1378
rect 201 1276 235 1310
rect 201 1208 235 1242
rect 201 1139 235 1174
rect 201 1089 235 1105
rect 289 1412 323 1450
rect 289 1344 323 1378
rect 289 1276 323 1310
rect 289 1208 323 1242
rect 289 1139 323 1174
rect 377 1412 411 1492
rect 377 1344 411 1378
rect 377 1276 411 1310
rect 377 1208 411 1242
rect 377 1157 411 1174
rect 465 1412 499 1450
rect 465 1344 499 1378
rect 465 1276 499 1310
rect 465 1208 499 1242
rect 289 1094 323 1105
rect 465 1139 499 1174
rect 553 1412 587 1492
rect 553 1344 587 1378
rect 553 1276 587 1310
rect 553 1208 587 1242
rect 553 1157 587 1174
rect 641 1412 675 1450
rect 641 1344 675 1378
rect 641 1276 675 1310
rect 641 1208 675 1242
rect 465 1094 499 1105
rect 641 1139 675 1174
rect 729 1412 763 1492
rect 729 1344 763 1378
rect 729 1276 763 1310
rect 729 1208 763 1242
rect 729 1157 763 1174
rect 931 1470 993 1492
rect 931 1436 945 1470
rect 979 1436 993 1470
rect 931 1398 993 1436
rect 931 1364 945 1398
rect 979 1364 993 1398
rect 931 1326 993 1364
rect 931 1292 945 1326
rect 979 1292 993 1326
rect 931 1254 993 1292
rect 931 1220 945 1254
rect 979 1220 993 1254
rect 931 1182 993 1220
rect 641 1094 675 1105
rect 931 1148 945 1182
rect 979 1148 993 1182
rect 931 1110 993 1148
rect -31 1038 31 1076
rect 289 1060 831 1094
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect -31 868 31 932
rect 205 1003 239 1019
rect 205 905 239 969
rect -31 546 31 572
rect -31 512 -17 546
rect 17 512 31 546
rect -31 474 31 512
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect 205 461 239 871
rect 205 411 239 427
rect 427 1003 461 1019
rect 427 535 461 969
rect 427 461 461 501
rect 427 411 461 427
rect 649 1003 683 1019
rect 649 757 683 969
rect 649 461 683 723
rect 649 411 683 427
rect 797 610 831 1060
rect 931 1076 945 1110
rect 979 1076 993 1110
rect 1163 1412 1197 1492
rect 1163 1344 1197 1378
rect 1163 1276 1197 1310
rect 1163 1208 1197 1242
rect 1163 1139 1197 1174
rect 1163 1089 1197 1105
rect 1251 1412 1285 1450
rect 1251 1344 1285 1378
rect 1251 1276 1285 1310
rect 1251 1208 1285 1242
rect 1251 1139 1285 1174
rect 1339 1412 1373 1492
rect 1339 1344 1373 1378
rect 1339 1276 1373 1310
rect 1339 1208 1373 1242
rect 1339 1157 1373 1174
rect 1427 1412 1461 1450
rect 1427 1344 1461 1378
rect 1427 1276 1461 1310
rect 1427 1208 1461 1242
rect 1251 1094 1285 1105
rect 1427 1139 1461 1174
rect 1515 1412 1549 1492
rect 1515 1344 1549 1378
rect 1515 1276 1549 1310
rect 1515 1208 1549 1242
rect 1515 1157 1549 1174
rect 1603 1412 1637 1450
rect 1603 1344 1637 1378
rect 1603 1276 1637 1310
rect 1603 1208 1637 1242
rect 1427 1094 1461 1105
rect 1603 1139 1637 1174
rect 1691 1412 1725 1492
rect 1691 1344 1725 1378
rect 1691 1276 1725 1310
rect 1691 1208 1725 1242
rect 1691 1157 1725 1174
rect 1893 1470 1955 1492
rect 1893 1436 1907 1470
rect 1941 1436 1955 1470
rect 1893 1398 1955 1436
rect 1893 1364 1907 1398
rect 1941 1364 1955 1398
rect 1893 1326 1955 1364
rect 1893 1292 1907 1326
rect 1941 1292 1955 1326
rect 1893 1254 1955 1292
rect 1893 1220 1907 1254
rect 1941 1220 1955 1254
rect 1893 1182 1955 1220
rect 1603 1094 1637 1105
rect 1893 1148 1907 1182
rect 1941 1148 1955 1182
rect 1893 1110 1955 1148
rect 931 1038 993 1076
rect 1251 1060 1793 1094
rect 931 1004 945 1038
rect 979 1004 993 1038
rect 931 966 993 1004
rect 931 932 945 966
rect 979 932 993 966
rect 931 868 993 932
rect 1167 1003 1201 1019
rect 1389 1003 1423 1019
rect -31 368 -17 402
rect 17 368 31 402
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect 101 363 135 379
rect 295 363 329 379
rect 489 363 523 379
rect 135 329 198 363
rect 232 329 295 363
rect 329 329 392 363
rect 426 329 489 363
rect 101 291 135 329
rect 101 223 135 257
rect 295 291 329 329
rect 489 313 523 329
rect 603 363 637 379
rect 797 378 831 576
rect 1167 610 1201 969
rect 1388 979 1389 995
rect 1422 945 1423 969
rect 1388 929 1423 945
rect 603 291 637 329
rect 101 153 135 189
rect 101 103 135 119
rect 198 238 232 254
rect -31 62 31 80
rect 198 62 232 204
rect 295 223 329 257
rect 393 244 427 260
rect 603 244 637 257
rect 427 223 637 244
rect 427 210 603 223
rect 393 194 427 210
rect 295 153 329 189
rect 700 344 831 378
rect 931 546 993 572
rect 931 512 945 546
rect 979 512 993 546
rect 931 474 993 512
rect 931 440 945 474
rect 979 440 993 474
rect 931 402 993 440
rect 1167 461 1201 576
rect 1167 411 1201 427
rect 1389 461 1423 929
rect 1611 1003 1645 1019
rect 1611 847 1645 969
rect 1610 831 1645 847
rect 1644 797 1645 831
rect 1610 781 1645 797
rect 1389 411 1423 427
rect 1611 461 1645 781
rect 1611 411 1645 427
rect 1759 757 1793 1060
rect 1893 1076 1907 1110
rect 1941 1076 1955 1110
rect 2125 1412 2159 1492
rect 2125 1344 2159 1378
rect 2125 1276 2159 1310
rect 2125 1208 2159 1242
rect 2125 1139 2159 1174
rect 2125 1089 2159 1105
rect 2213 1412 2247 1450
rect 2213 1344 2247 1378
rect 2213 1276 2247 1310
rect 2213 1208 2247 1242
rect 2213 1139 2247 1174
rect 2301 1412 2335 1492
rect 2301 1344 2335 1378
rect 2301 1276 2335 1310
rect 2301 1208 2335 1242
rect 2301 1157 2335 1174
rect 2389 1412 2423 1450
rect 2389 1344 2423 1378
rect 2389 1276 2423 1310
rect 2389 1208 2423 1242
rect 2213 1094 2247 1105
rect 2389 1139 2423 1174
rect 2477 1412 2511 1492
rect 2477 1344 2511 1378
rect 2477 1276 2511 1310
rect 2477 1208 2511 1242
rect 2477 1157 2511 1174
rect 2565 1412 2599 1450
rect 2565 1344 2599 1378
rect 2565 1276 2599 1310
rect 2565 1208 2599 1242
rect 2389 1094 2423 1105
rect 2565 1139 2599 1174
rect 2653 1412 2687 1492
rect 2653 1344 2687 1378
rect 2653 1276 2687 1310
rect 2653 1208 2687 1242
rect 2653 1157 2687 1174
rect 2855 1470 2917 1492
rect 2855 1436 2869 1470
rect 2903 1436 2917 1470
rect 2855 1398 2917 1436
rect 2855 1364 2869 1398
rect 2903 1364 2917 1398
rect 2855 1326 2917 1364
rect 2855 1292 2869 1326
rect 2903 1292 2917 1326
rect 2855 1254 2917 1292
rect 2855 1220 2869 1254
rect 2903 1220 2917 1254
rect 2855 1182 2917 1220
rect 2565 1094 2599 1105
rect 2855 1148 2869 1182
rect 2903 1148 2917 1182
rect 2855 1110 2917 1148
rect 1893 1038 1955 1076
rect 2213 1060 2755 1094
rect 1893 1004 1907 1038
rect 1941 1004 1955 1038
rect 1893 966 1955 1004
rect 1893 932 1907 966
rect 1941 932 1955 966
rect 1893 868 1955 932
rect 2129 1003 2163 1019
rect 931 368 945 402
rect 979 368 993 402
rect 700 247 734 344
rect 931 330 993 368
rect 700 197 734 213
rect 797 291 831 307
rect 797 223 831 257
rect 489 153 523 169
rect 329 119 392 153
rect 426 119 489 153
rect 295 103 329 119
rect 489 103 523 119
rect 603 153 637 189
rect 797 153 831 189
rect 637 119 700 153
rect 734 119 797 153
rect 603 103 637 119
rect 797 103 831 119
rect 931 296 945 330
rect 979 296 993 330
rect 931 258 993 296
rect 931 224 945 258
rect 979 224 993 258
rect 931 186 993 224
rect 931 152 945 186
rect 979 152 993 186
rect 931 114 993 152
rect 931 80 945 114
rect 979 80 993 114
rect 1063 363 1097 379
rect 1257 363 1291 379
rect 1451 363 1485 379
rect 1097 329 1160 363
rect 1194 329 1257 363
rect 1291 329 1354 363
rect 1388 329 1451 363
rect 1063 291 1097 329
rect 1063 223 1097 257
rect 1257 291 1291 329
rect 1451 313 1485 329
rect 1565 363 1599 379
rect 1759 378 1793 723
rect 2129 610 2163 969
rect 1565 291 1599 329
rect 1063 153 1097 189
rect 1063 103 1097 119
rect 1160 238 1194 254
rect 931 62 993 80
rect 1160 62 1194 204
rect 1257 223 1291 257
rect 1355 244 1389 260
rect 1565 244 1599 257
rect 1389 223 1599 244
rect 1389 210 1565 223
rect 1355 194 1389 210
rect 1257 153 1291 189
rect 1662 344 1793 378
rect 1893 546 1955 572
rect 1893 512 1907 546
rect 1941 512 1955 546
rect 1893 474 1955 512
rect 1893 440 1907 474
rect 1941 440 1955 474
rect 1893 402 1955 440
rect 2129 461 2163 576
rect 2129 411 2163 427
rect 2351 1003 2385 1019
rect 2351 462 2385 969
rect 2351 411 2385 427
rect 2573 1003 2607 1019
rect 2573 831 2607 969
rect 2573 461 2607 797
rect 2573 411 2607 427
rect 2721 609 2755 1060
rect 2855 1076 2869 1110
rect 2903 1076 2917 1110
rect 3087 1412 3121 1492
rect 3087 1344 3121 1378
rect 3087 1276 3121 1310
rect 3087 1208 3121 1242
rect 3087 1139 3121 1174
rect 3087 1089 3121 1105
rect 3175 1412 3209 1450
rect 3175 1344 3209 1378
rect 3175 1276 3209 1310
rect 3175 1208 3209 1242
rect 3175 1139 3209 1174
rect 3263 1412 3297 1492
rect 3263 1344 3297 1378
rect 3263 1276 3297 1310
rect 3263 1208 3297 1242
rect 3263 1157 3297 1174
rect 3351 1412 3385 1450
rect 3351 1344 3385 1378
rect 3351 1276 3385 1310
rect 3351 1208 3385 1242
rect 3175 1094 3209 1105
rect 3351 1139 3385 1174
rect 3439 1412 3473 1492
rect 3439 1344 3473 1378
rect 3439 1276 3473 1310
rect 3439 1208 3473 1242
rect 3439 1157 3473 1174
rect 3527 1412 3561 1450
rect 3527 1344 3561 1378
rect 3527 1276 3561 1310
rect 3527 1208 3561 1242
rect 3351 1094 3385 1105
rect 3527 1139 3561 1174
rect 3615 1412 3649 1492
rect 3615 1344 3649 1378
rect 3615 1276 3649 1310
rect 3615 1208 3649 1242
rect 3615 1157 3649 1174
rect 3817 1470 3879 1492
rect 3817 1436 3831 1470
rect 3865 1436 3879 1470
rect 3817 1398 3879 1436
rect 3817 1364 3831 1398
rect 3865 1364 3879 1398
rect 3817 1326 3879 1364
rect 3817 1292 3831 1326
rect 3865 1292 3879 1326
rect 3817 1254 3879 1292
rect 3817 1220 3831 1254
rect 3865 1220 3879 1254
rect 3817 1182 3879 1220
rect 3527 1094 3561 1105
rect 3817 1148 3831 1182
rect 3865 1148 3879 1182
rect 3817 1110 3879 1148
rect 2855 1038 2917 1076
rect 3175 1060 3717 1094
rect 2855 1004 2869 1038
rect 2903 1004 2917 1038
rect 2855 966 2917 1004
rect 2855 932 2869 966
rect 2903 932 2917 966
rect 2855 868 2917 932
rect 3091 1003 3125 1019
rect 1893 368 1907 402
rect 1941 368 1955 402
rect 1662 247 1696 344
rect 1893 330 1955 368
rect 1662 197 1696 213
rect 1759 291 1793 307
rect 1759 223 1793 257
rect 1451 153 1485 169
rect 1291 119 1354 153
rect 1388 119 1451 153
rect 1257 103 1291 119
rect 1451 103 1485 119
rect 1565 153 1599 189
rect 1759 153 1793 189
rect 1599 119 1662 153
rect 1696 119 1759 153
rect 1565 103 1599 119
rect 1759 103 1793 119
rect 1893 296 1907 330
rect 1941 296 1955 330
rect 1893 258 1955 296
rect 1893 224 1907 258
rect 1941 224 1955 258
rect 1893 186 1955 224
rect 1893 152 1907 186
rect 1941 152 1955 186
rect 1893 114 1955 152
rect 1893 80 1907 114
rect 1941 80 1955 114
rect 2025 363 2059 379
rect 2219 363 2253 379
rect 2413 363 2447 379
rect 2059 329 2122 363
rect 2156 329 2219 363
rect 2253 329 2316 363
rect 2350 329 2413 363
rect 2025 291 2059 329
rect 2025 223 2059 257
rect 2219 291 2253 329
rect 2413 313 2447 329
rect 2527 363 2561 379
rect 2721 378 2755 575
rect 3091 609 3125 969
rect 2527 291 2561 329
rect 2025 153 2059 189
rect 2025 103 2059 119
rect 2122 238 2156 254
rect 1893 62 1955 80
rect 2122 62 2156 204
rect 2219 223 2253 257
rect 2317 244 2351 260
rect 2527 244 2561 257
rect 2351 223 2561 244
rect 2351 210 2527 223
rect 2317 194 2351 210
rect 2219 153 2253 189
rect 2624 344 2755 378
rect 2855 546 2917 572
rect 2855 512 2869 546
rect 2903 512 2917 546
rect 2855 474 2917 512
rect 2855 440 2869 474
rect 2903 440 2917 474
rect 2855 402 2917 440
rect 3091 461 3125 575
rect 3091 411 3125 427
rect 3313 1003 3347 1019
rect 3313 461 3347 945
rect 3313 411 3347 427
rect 3535 1003 3569 1019
rect 3535 535 3569 969
rect 3535 461 3569 501
rect 3535 411 3569 427
rect 3683 831 3717 1060
rect 3817 1076 3831 1110
rect 3865 1076 3879 1110
rect 4049 1412 4083 1492
rect 4049 1344 4083 1378
rect 4049 1276 4083 1310
rect 4049 1208 4083 1242
rect 4049 1139 4083 1174
rect 4049 1089 4083 1105
rect 4137 1412 4171 1450
rect 4137 1344 4171 1378
rect 4137 1276 4171 1310
rect 4137 1208 4171 1242
rect 4137 1139 4171 1174
rect 4225 1412 4259 1492
rect 4225 1344 4259 1378
rect 4225 1276 4259 1310
rect 4225 1208 4259 1242
rect 4225 1157 4259 1174
rect 4313 1412 4347 1450
rect 4313 1344 4347 1378
rect 4313 1276 4347 1310
rect 4313 1208 4347 1242
rect 4137 1094 4171 1105
rect 4313 1139 4347 1174
rect 4401 1412 4435 1492
rect 4401 1344 4435 1378
rect 4401 1276 4435 1310
rect 4401 1208 4435 1242
rect 4401 1157 4435 1174
rect 4489 1412 4523 1450
rect 4489 1344 4523 1378
rect 4489 1276 4523 1310
rect 4489 1208 4523 1242
rect 4313 1094 4347 1105
rect 4489 1139 4523 1174
rect 4577 1412 4611 1492
rect 4577 1344 4611 1378
rect 4577 1276 4611 1310
rect 4577 1208 4611 1242
rect 4577 1157 4611 1174
rect 4779 1470 4841 1492
rect 4779 1436 4793 1470
rect 4827 1436 4841 1470
rect 4779 1398 4841 1436
rect 4779 1364 4793 1398
rect 4827 1364 4841 1398
rect 4779 1326 4841 1364
rect 4779 1292 4793 1326
rect 4827 1292 4841 1326
rect 4779 1254 4841 1292
rect 4779 1220 4793 1254
rect 4827 1220 4841 1254
rect 4779 1182 4841 1220
rect 4489 1094 4523 1105
rect 4779 1148 4793 1182
rect 4827 1148 4841 1182
rect 4779 1110 4841 1148
rect 3817 1038 3879 1076
rect 4137 1060 4679 1094
rect 3817 1004 3831 1038
rect 3865 1004 3879 1038
rect 3817 966 3879 1004
rect 3817 932 3831 966
rect 3865 932 3879 966
rect 3817 868 3879 932
rect 4053 1003 4087 1019
rect 2855 368 2869 402
rect 2903 368 2917 402
rect 2624 247 2658 344
rect 2855 330 2917 368
rect 2624 197 2658 213
rect 2721 291 2755 307
rect 2721 223 2755 257
rect 2413 153 2447 169
rect 2253 119 2316 153
rect 2350 119 2413 153
rect 2219 103 2253 119
rect 2413 103 2447 119
rect 2527 153 2561 189
rect 2721 153 2755 189
rect 2561 119 2624 153
rect 2658 119 2721 153
rect 2527 103 2561 119
rect 2721 103 2755 119
rect 2855 296 2869 330
rect 2903 296 2917 330
rect 2855 258 2917 296
rect 2855 224 2869 258
rect 2903 224 2917 258
rect 2855 186 2917 224
rect 2855 152 2869 186
rect 2903 152 2917 186
rect 2855 114 2917 152
rect 2855 80 2869 114
rect 2903 80 2917 114
rect 2987 363 3021 379
rect 3181 363 3215 379
rect 3375 363 3409 379
rect 3021 329 3084 363
rect 3118 329 3181 363
rect 3215 329 3278 363
rect 3312 329 3375 363
rect 2987 291 3021 329
rect 2987 223 3021 257
rect 3181 291 3215 329
rect 3375 313 3409 329
rect 3489 363 3523 379
rect 3683 378 3717 797
rect 4053 757 4087 969
rect 3489 291 3523 329
rect 2987 153 3021 189
rect 2987 103 3021 119
rect 3084 238 3118 254
rect 2855 62 2917 80
rect 3084 62 3118 204
rect 3181 223 3215 257
rect 3279 244 3313 260
rect 3489 244 3523 257
rect 3313 223 3523 244
rect 3313 210 3489 223
rect 3279 194 3313 210
rect 3181 153 3215 189
rect 3586 344 3717 378
rect 3817 546 3879 572
rect 3817 512 3831 546
rect 3865 512 3879 546
rect 3817 474 3879 512
rect 3817 440 3831 474
rect 3865 440 3879 474
rect 3817 402 3879 440
rect 4053 461 4087 723
rect 4053 411 4087 427
rect 4275 1003 4309 1019
rect 4275 535 4309 969
rect 4275 461 4309 501
rect 4275 411 4309 427
rect 4497 1003 4531 1019
rect 4497 683 4531 969
rect 4497 461 4531 649
rect 4497 411 4531 427
rect 4645 757 4679 1060
rect 4779 1076 4793 1110
rect 4827 1076 4841 1110
rect 5011 1412 5045 1492
rect 5011 1344 5045 1378
rect 5011 1276 5045 1310
rect 5011 1208 5045 1242
rect 5011 1139 5045 1174
rect 5011 1089 5045 1105
rect 5099 1412 5133 1450
rect 5099 1344 5133 1378
rect 5099 1276 5133 1310
rect 5099 1208 5133 1242
rect 5099 1139 5133 1174
rect 5187 1412 5221 1492
rect 5187 1344 5221 1378
rect 5187 1276 5221 1310
rect 5187 1208 5221 1242
rect 5187 1157 5221 1174
rect 5275 1412 5309 1450
rect 5275 1344 5309 1378
rect 5275 1276 5309 1310
rect 5275 1208 5309 1242
rect 5099 1094 5133 1105
rect 5275 1139 5309 1174
rect 5363 1412 5397 1492
rect 5363 1344 5397 1378
rect 5363 1276 5397 1310
rect 5363 1208 5397 1242
rect 5363 1157 5397 1174
rect 5451 1412 5485 1450
rect 5451 1344 5485 1378
rect 5451 1276 5485 1310
rect 5451 1208 5485 1242
rect 5275 1094 5309 1105
rect 5451 1139 5485 1174
rect 5539 1412 5573 1492
rect 5539 1344 5573 1378
rect 5539 1276 5573 1310
rect 5539 1208 5573 1242
rect 5539 1157 5573 1174
rect 5741 1470 5803 1492
rect 5741 1436 5755 1470
rect 5789 1436 5803 1470
rect 5741 1398 5803 1436
rect 5741 1364 5755 1398
rect 5789 1364 5803 1398
rect 5741 1326 5803 1364
rect 5741 1292 5755 1326
rect 5789 1292 5803 1326
rect 5741 1254 5803 1292
rect 5741 1220 5755 1254
rect 5789 1220 5803 1254
rect 5741 1182 5803 1220
rect 5451 1094 5485 1105
rect 5741 1148 5755 1182
rect 5789 1148 5803 1182
rect 5741 1110 5803 1148
rect 4779 1038 4841 1076
rect 5099 1060 5641 1094
rect 4779 1004 4793 1038
rect 4827 1004 4841 1038
rect 4779 966 4841 1004
rect 4779 932 4793 966
rect 4827 932 4841 966
rect 4779 868 4841 932
rect 5015 1003 5049 1019
rect 3817 368 3831 402
rect 3865 368 3879 402
rect 3586 247 3620 344
rect 3817 330 3879 368
rect 3586 197 3620 213
rect 3683 291 3717 307
rect 3683 223 3717 257
rect 3375 153 3409 169
rect 3215 119 3278 153
rect 3312 119 3375 153
rect 3181 103 3215 119
rect 3375 103 3409 119
rect 3489 153 3523 189
rect 3683 153 3717 189
rect 3523 119 3586 153
rect 3620 119 3683 153
rect 3489 103 3523 119
rect 3683 103 3717 119
rect 3817 296 3831 330
rect 3865 296 3879 330
rect 3817 258 3879 296
rect 3817 224 3831 258
rect 3865 224 3879 258
rect 3817 186 3879 224
rect 3817 152 3831 186
rect 3865 152 3879 186
rect 3817 114 3879 152
rect 3817 80 3831 114
rect 3865 80 3879 114
rect 3949 363 3983 379
rect 4143 363 4177 379
rect 4337 363 4371 379
rect 3983 329 4046 363
rect 4080 329 4143 363
rect 4177 329 4240 363
rect 4274 329 4337 363
rect 3949 291 3983 329
rect 3949 223 3983 257
rect 4143 291 4177 329
rect 4337 313 4371 329
rect 4451 363 4485 379
rect 4645 378 4679 723
rect 5015 757 5049 969
rect 4451 291 4485 329
rect 3949 153 3983 189
rect 3949 103 3983 119
rect 4046 238 4080 254
rect 3817 62 3879 80
rect 4046 62 4080 204
rect 4143 223 4177 257
rect 4241 244 4275 260
rect 4451 244 4485 257
rect 4275 223 4485 244
rect 4275 210 4451 223
rect 4241 194 4275 210
rect 4143 153 4177 189
rect 4548 344 4679 378
rect 4779 546 4841 572
rect 4779 512 4793 546
rect 4827 512 4841 546
rect 4779 474 4841 512
rect 4779 440 4793 474
rect 4827 440 4841 474
rect 4779 402 4841 440
rect 5015 461 5049 723
rect 5015 411 5049 427
rect 5237 1003 5271 1019
rect 5237 461 5271 969
rect 5237 411 5271 427
rect 5459 1003 5493 1019
rect 5459 831 5493 969
rect 5459 461 5493 797
rect 5459 411 5493 427
rect 5607 683 5641 1060
rect 5741 1076 5755 1110
rect 5789 1076 5803 1110
rect 5973 1412 6007 1492
rect 5973 1344 6007 1378
rect 5973 1276 6007 1310
rect 5973 1208 6007 1242
rect 5973 1139 6007 1174
rect 5973 1089 6007 1105
rect 6061 1412 6095 1450
rect 6061 1344 6095 1378
rect 6061 1276 6095 1310
rect 6061 1208 6095 1242
rect 6061 1139 6095 1174
rect 6149 1412 6183 1492
rect 6149 1344 6183 1378
rect 6149 1276 6183 1310
rect 6149 1208 6183 1242
rect 6149 1157 6183 1174
rect 6237 1412 6271 1450
rect 6237 1344 6271 1378
rect 6237 1276 6271 1310
rect 6237 1208 6271 1242
rect 6061 1094 6095 1105
rect 6237 1139 6271 1174
rect 6325 1412 6359 1492
rect 6325 1344 6359 1378
rect 6325 1276 6359 1310
rect 6325 1208 6359 1242
rect 6325 1157 6359 1174
rect 6413 1412 6447 1450
rect 6413 1344 6447 1378
rect 6413 1276 6447 1310
rect 6413 1208 6447 1242
rect 6237 1094 6271 1105
rect 6413 1139 6447 1174
rect 6501 1412 6535 1492
rect 6501 1344 6535 1378
rect 6501 1276 6535 1310
rect 6501 1208 6535 1242
rect 6501 1157 6535 1174
rect 6703 1470 6765 1492
rect 6703 1436 6717 1470
rect 6751 1436 6765 1470
rect 6703 1398 6765 1436
rect 6703 1364 6717 1398
rect 6751 1364 6765 1398
rect 6703 1326 6765 1364
rect 6703 1292 6717 1326
rect 6751 1292 6765 1326
rect 6703 1254 6765 1292
rect 6703 1220 6717 1254
rect 6751 1220 6765 1254
rect 6703 1182 6765 1220
rect 6413 1094 6447 1105
rect 6703 1148 6717 1182
rect 6751 1148 6765 1182
rect 6703 1110 6765 1148
rect 5741 1038 5803 1076
rect 6061 1060 6603 1094
rect 5741 1004 5755 1038
rect 5789 1004 5803 1038
rect 5741 966 5803 1004
rect 5741 932 5755 966
rect 5789 932 5803 966
rect 5741 868 5803 932
rect 5977 1003 6011 1019
rect 5977 905 6011 969
rect 4779 368 4793 402
rect 4827 368 4841 402
rect 4548 247 4582 344
rect 4779 330 4841 368
rect 4548 197 4582 213
rect 4645 291 4679 307
rect 4645 223 4679 257
rect 4337 153 4371 169
rect 4177 119 4240 153
rect 4274 119 4337 153
rect 4143 103 4177 119
rect 4337 103 4371 119
rect 4451 153 4485 189
rect 4645 153 4679 189
rect 4485 119 4548 153
rect 4582 119 4645 153
rect 4451 103 4485 119
rect 4645 103 4679 119
rect 4779 296 4793 330
rect 4827 296 4841 330
rect 4779 258 4841 296
rect 4779 224 4793 258
rect 4827 224 4841 258
rect 4779 186 4841 224
rect 4779 152 4793 186
rect 4827 152 4841 186
rect 4779 114 4841 152
rect 4779 80 4793 114
rect 4827 80 4841 114
rect 4911 363 4945 379
rect 5105 363 5139 379
rect 5299 363 5333 379
rect 4945 329 5008 363
rect 5042 329 5105 363
rect 5139 329 5202 363
rect 5236 329 5299 363
rect 4911 291 4945 329
rect 4911 223 4945 257
rect 5105 291 5139 329
rect 5299 313 5333 329
rect 5413 363 5447 379
rect 5607 378 5641 649
rect 5413 291 5447 329
rect 4911 153 4945 189
rect 4911 103 4945 119
rect 5008 238 5042 254
rect 4779 62 4841 80
rect 5008 62 5042 204
rect 5105 223 5139 257
rect 5203 244 5237 260
rect 5413 244 5447 257
rect 5237 223 5447 244
rect 5237 210 5413 223
rect 5203 194 5237 210
rect 5105 153 5139 189
rect 5510 344 5641 378
rect 5741 546 5803 572
rect 5741 512 5755 546
rect 5789 512 5803 546
rect 5741 474 5803 512
rect 5741 440 5755 474
rect 5789 440 5803 474
rect 5741 402 5803 440
rect 5977 461 6011 871
rect 5977 411 6011 427
rect 6199 1003 6233 1019
rect 6199 535 6233 969
rect 6199 461 6233 501
rect 6199 411 6233 427
rect 6421 1003 6455 1019
rect 6421 757 6455 969
rect 6421 461 6455 723
rect 6421 411 6455 427
rect 6569 610 6603 1060
rect 6703 1076 6717 1110
rect 6751 1076 6765 1110
rect 6935 1412 6969 1492
rect 6935 1344 6969 1378
rect 6935 1276 6969 1310
rect 6935 1208 6969 1242
rect 6935 1139 6969 1174
rect 6935 1089 6969 1105
rect 7023 1412 7057 1450
rect 7023 1344 7057 1378
rect 7023 1276 7057 1310
rect 7023 1208 7057 1242
rect 7023 1139 7057 1174
rect 7111 1412 7145 1492
rect 7111 1344 7145 1378
rect 7111 1276 7145 1310
rect 7111 1208 7145 1242
rect 7111 1157 7145 1174
rect 7199 1412 7233 1450
rect 7199 1344 7233 1378
rect 7199 1276 7233 1310
rect 7199 1208 7233 1242
rect 7023 1094 7057 1105
rect 7199 1139 7233 1174
rect 7287 1412 7321 1492
rect 7287 1344 7321 1378
rect 7287 1276 7321 1310
rect 7287 1208 7321 1242
rect 7287 1157 7321 1174
rect 7375 1412 7409 1450
rect 7375 1344 7409 1378
rect 7375 1276 7409 1310
rect 7375 1208 7409 1242
rect 7199 1094 7233 1105
rect 7375 1139 7409 1174
rect 7463 1412 7497 1492
rect 7463 1344 7497 1378
rect 7463 1276 7497 1310
rect 7463 1208 7497 1242
rect 7463 1157 7497 1174
rect 7665 1470 7727 1492
rect 7665 1436 7679 1470
rect 7713 1436 7727 1470
rect 7665 1398 7727 1436
rect 7665 1364 7679 1398
rect 7713 1364 7727 1398
rect 7665 1326 7727 1364
rect 7665 1292 7679 1326
rect 7713 1292 7727 1326
rect 7665 1254 7727 1292
rect 7665 1220 7679 1254
rect 7713 1220 7727 1254
rect 7665 1182 7727 1220
rect 7375 1094 7409 1105
rect 7665 1148 7679 1182
rect 7713 1148 7727 1182
rect 7665 1110 7727 1148
rect 6703 1038 6765 1076
rect 7023 1060 7565 1094
rect 6703 1004 6717 1038
rect 6751 1004 6765 1038
rect 6703 966 6765 1004
rect 6703 932 6717 966
rect 6751 932 6765 966
rect 6703 868 6765 932
rect 6939 1003 6973 1019
rect 7161 1003 7195 1019
rect 5741 368 5755 402
rect 5789 368 5803 402
rect 5510 247 5544 344
rect 5741 330 5803 368
rect 5510 197 5544 213
rect 5607 291 5641 307
rect 5607 223 5641 257
rect 5299 153 5333 169
rect 5139 119 5202 153
rect 5236 119 5299 153
rect 5105 103 5139 119
rect 5299 103 5333 119
rect 5413 153 5447 189
rect 5607 153 5641 189
rect 5447 119 5510 153
rect 5544 119 5607 153
rect 5413 103 5447 119
rect 5607 103 5641 119
rect 5741 296 5755 330
rect 5789 296 5803 330
rect 5741 258 5803 296
rect 5741 224 5755 258
rect 5789 224 5803 258
rect 5741 186 5803 224
rect 5741 152 5755 186
rect 5789 152 5803 186
rect 5741 114 5803 152
rect 5741 80 5755 114
rect 5789 80 5803 114
rect 5873 363 5907 379
rect 6067 363 6101 379
rect 6261 363 6295 379
rect 5907 329 5970 363
rect 6004 329 6067 363
rect 6101 329 6164 363
rect 6198 329 6261 363
rect 5873 291 5907 329
rect 5873 223 5907 257
rect 6067 291 6101 329
rect 6261 313 6295 329
rect 6375 363 6409 379
rect 6569 378 6603 576
rect 6939 610 6973 969
rect 7160 979 7161 995
rect 7194 945 7195 969
rect 7160 929 7195 945
rect 6375 291 6409 329
rect 5873 153 5907 189
rect 5873 103 5907 119
rect 5970 238 6004 254
rect 5741 62 5803 80
rect 5970 62 6004 204
rect 6067 223 6101 257
rect 6165 244 6199 260
rect 6375 244 6409 257
rect 6199 223 6409 244
rect 6199 210 6375 223
rect 6165 194 6199 210
rect 6067 153 6101 189
rect 6472 344 6603 378
rect 6703 546 6765 572
rect 6703 512 6717 546
rect 6751 512 6765 546
rect 6703 474 6765 512
rect 6703 440 6717 474
rect 6751 440 6765 474
rect 6703 402 6765 440
rect 6939 461 6973 576
rect 6939 411 6973 427
rect 7161 461 7195 929
rect 7383 1003 7417 1019
rect 7383 847 7417 969
rect 7382 831 7417 847
rect 7416 797 7417 831
rect 7382 781 7417 797
rect 7161 411 7195 427
rect 7383 461 7417 781
rect 7383 411 7417 427
rect 7531 757 7565 1060
rect 7665 1076 7679 1110
rect 7713 1076 7727 1110
rect 7897 1412 7931 1492
rect 7897 1344 7931 1378
rect 7897 1276 7931 1310
rect 7897 1208 7931 1242
rect 7897 1139 7931 1174
rect 7897 1089 7931 1105
rect 7985 1412 8019 1450
rect 7985 1344 8019 1378
rect 7985 1276 8019 1310
rect 7985 1208 8019 1242
rect 7985 1139 8019 1174
rect 8073 1412 8107 1492
rect 8073 1344 8107 1378
rect 8073 1276 8107 1310
rect 8073 1208 8107 1242
rect 8073 1157 8107 1174
rect 8161 1412 8195 1450
rect 8161 1344 8195 1378
rect 8161 1276 8195 1310
rect 8161 1208 8195 1242
rect 7985 1094 8019 1105
rect 8161 1139 8195 1174
rect 8249 1412 8283 1492
rect 8249 1344 8283 1378
rect 8249 1276 8283 1310
rect 8249 1208 8283 1242
rect 8249 1157 8283 1174
rect 8337 1412 8371 1450
rect 8337 1344 8371 1378
rect 8337 1276 8371 1310
rect 8337 1208 8371 1242
rect 8161 1094 8195 1105
rect 8337 1139 8371 1174
rect 8425 1412 8459 1492
rect 8425 1344 8459 1378
rect 8425 1276 8459 1310
rect 8425 1208 8459 1242
rect 8425 1157 8459 1174
rect 8627 1470 8689 1492
rect 8627 1436 8641 1470
rect 8675 1436 8689 1470
rect 8627 1398 8689 1436
rect 8627 1364 8641 1398
rect 8675 1364 8689 1398
rect 8627 1326 8689 1364
rect 8627 1292 8641 1326
rect 8675 1292 8689 1326
rect 8627 1254 8689 1292
rect 8627 1220 8641 1254
rect 8675 1220 8689 1254
rect 8627 1182 8689 1220
rect 8337 1094 8371 1105
rect 8627 1148 8641 1182
rect 8675 1148 8689 1182
rect 8627 1110 8689 1148
rect 7665 1038 7727 1076
rect 7985 1060 8527 1094
rect 7665 1004 7679 1038
rect 7713 1004 7727 1038
rect 7665 966 7727 1004
rect 7665 932 7679 966
rect 7713 932 7727 966
rect 7665 868 7727 932
rect 7901 1003 7935 1019
rect 6703 368 6717 402
rect 6751 368 6765 402
rect 6472 247 6506 344
rect 6703 330 6765 368
rect 6472 197 6506 213
rect 6569 291 6603 307
rect 6569 223 6603 257
rect 6261 153 6295 169
rect 6101 119 6164 153
rect 6198 119 6261 153
rect 6067 103 6101 119
rect 6261 103 6295 119
rect 6375 153 6409 189
rect 6569 153 6603 189
rect 6409 119 6472 153
rect 6506 119 6569 153
rect 6375 103 6409 119
rect 6569 103 6603 119
rect 6703 296 6717 330
rect 6751 296 6765 330
rect 6703 258 6765 296
rect 6703 224 6717 258
rect 6751 224 6765 258
rect 6703 186 6765 224
rect 6703 152 6717 186
rect 6751 152 6765 186
rect 6703 114 6765 152
rect 6703 80 6717 114
rect 6751 80 6765 114
rect 6835 363 6869 379
rect 7029 363 7063 379
rect 7223 363 7257 379
rect 6869 329 6932 363
rect 6966 329 7029 363
rect 7063 329 7126 363
rect 7160 329 7223 363
rect 6835 291 6869 329
rect 6835 223 6869 257
rect 7029 291 7063 329
rect 7223 313 7257 329
rect 7337 363 7371 379
rect 7531 378 7565 723
rect 7901 610 7935 969
rect 7337 291 7371 329
rect 6835 153 6869 189
rect 6835 103 6869 119
rect 6932 238 6966 254
rect 6703 62 6765 80
rect 6932 62 6966 204
rect 7029 223 7063 257
rect 7127 244 7161 260
rect 7337 244 7371 257
rect 7161 223 7371 244
rect 7161 210 7337 223
rect 7127 194 7161 210
rect 7029 153 7063 189
rect 7434 344 7565 378
rect 7665 546 7727 572
rect 7665 512 7679 546
rect 7713 512 7727 546
rect 7665 474 7727 512
rect 7665 440 7679 474
rect 7713 440 7727 474
rect 7665 402 7727 440
rect 7901 461 7935 576
rect 7901 411 7935 427
rect 8123 1003 8157 1019
rect 8123 462 8157 969
rect 8123 411 8157 427
rect 8345 1003 8379 1019
rect 8345 831 8379 969
rect 8345 461 8379 797
rect 8345 411 8379 427
rect 8493 609 8527 1060
rect 8627 1076 8641 1110
rect 8675 1076 8689 1110
rect 8859 1412 8893 1492
rect 8859 1344 8893 1378
rect 8859 1276 8893 1310
rect 8859 1208 8893 1242
rect 8859 1139 8893 1174
rect 8859 1089 8893 1105
rect 8947 1412 8981 1450
rect 8947 1344 8981 1378
rect 8947 1276 8981 1310
rect 8947 1208 8981 1242
rect 8947 1139 8981 1174
rect 9035 1412 9069 1492
rect 9035 1344 9069 1378
rect 9035 1276 9069 1310
rect 9035 1208 9069 1242
rect 9035 1157 9069 1174
rect 9123 1412 9157 1450
rect 9123 1344 9157 1378
rect 9123 1276 9157 1310
rect 9123 1208 9157 1242
rect 8947 1094 8981 1105
rect 9123 1139 9157 1174
rect 9211 1412 9245 1492
rect 9211 1344 9245 1378
rect 9211 1276 9245 1310
rect 9211 1208 9245 1242
rect 9211 1157 9245 1174
rect 9299 1412 9333 1450
rect 9299 1344 9333 1378
rect 9299 1276 9333 1310
rect 9299 1208 9333 1242
rect 9123 1094 9157 1105
rect 9299 1139 9333 1174
rect 9387 1412 9421 1492
rect 9387 1344 9421 1378
rect 9387 1276 9421 1310
rect 9387 1208 9421 1242
rect 9387 1157 9421 1174
rect 9589 1470 9651 1492
rect 9589 1436 9603 1470
rect 9637 1436 9651 1470
rect 9589 1398 9651 1436
rect 9589 1364 9603 1398
rect 9637 1364 9651 1398
rect 9589 1326 9651 1364
rect 9589 1292 9603 1326
rect 9637 1292 9651 1326
rect 9589 1254 9651 1292
rect 9589 1220 9603 1254
rect 9637 1220 9651 1254
rect 9589 1182 9651 1220
rect 9299 1094 9333 1105
rect 9589 1148 9603 1182
rect 9637 1148 9651 1182
rect 9589 1110 9651 1148
rect 8627 1038 8689 1076
rect 8947 1060 9489 1094
rect 8627 1004 8641 1038
rect 8675 1004 8689 1038
rect 8627 966 8689 1004
rect 8627 932 8641 966
rect 8675 932 8689 966
rect 8627 868 8689 932
rect 8863 1003 8897 1019
rect 7665 368 7679 402
rect 7713 368 7727 402
rect 7434 247 7468 344
rect 7665 330 7727 368
rect 7434 197 7468 213
rect 7531 291 7565 307
rect 7531 223 7565 257
rect 7223 153 7257 169
rect 7063 119 7126 153
rect 7160 119 7223 153
rect 7029 103 7063 119
rect 7223 103 7257 119
rect 7337 153 7371 189
rect 7531 153 7565 189
rect 7371 119 7434 153
rect 7468 119 7531 153
rect 7337 103 7371 119
rect 7531 103 7565 119
rect 7665 296 7679 330
rect 7713 296 7727 330
rect 7665 258 7727 296
rect 7665 224 7679 258
rect 7713 224 7727 258
rect 7665 186 7727 224
rect 7665 152 7679 186
rect 7713 152 7727 186
rect 7665 114 7727 152
rect 7665 80 7679 114
rect 7713 80 7727 114
rect 7797 363 7831 379
rect 7991 363 8025 379
rect 8185 363 8219 379
rect 7831 329 7894 363
rect 7928 329 7991 363
rect 8025 329 8088 363
rect 8122 329 8185 363
rect 7797 291 7831 329
rect 7797 223 7831 257
rect 7991 291 8025 329
rect 8185 313 8219 329
rect 8299 363 8333 379
rect 8493 378 8527 575
rect 8863 609 8897 969
rect 8299 291 8333 329
rect 7797 153 7831 189
rect 7797 103 7831 119
rect 7894 238 7928 254
rect 7665 62 7727 80
rect 7894 62 7928 204
rect 7991 223 8025 257
rect 8089 244 8123 260
rect 8299 244 8333 257
rect 8123 223 8333 244
rect 8123 210 8299 223
rect 8089 194 8123 210
rect 7991 153 8025 189
rect 8396 344 8527 378
rect 8627 546 8689 572
rect 8627 512 8641 546
rect 8675 512 8689 546
rect 8627 474 8689 512
rect 8627 440 8641 474
rect 8675 440 8689 474
rect 8627 402 8689 440
rect 8863 461 8897 575
rect 8863 411 8897 427
rect 9085 1003 9119 1019
rect 9085 461 9119 945
rect 9085 411 9119 427
rect 9307 1003 9341 1019
rect 9307 535 9341 969
rect 9307 461 9341 501
rect 9307 411 9341 427
rect 9455 831 9489 1060
rect 9589 1076 9603 1110
rect 9637 1076 9651 1110
rect 9821 1412 9855 1492
rect 9821 1344 9855 1378
rect 9821 1276 9855 1310
rect 9821 1208 9855 1242
rect 9821 1139 9855 1174
rect 9821 1089 9855 1105
rect 9909 1412 9943 1450
rect 9909 1344 9943 1378
rect 9909 1276 9943 1310
rect 9909 1208 9943 1242
rect 9909 1139 9943 1174
rect 9997 1412 10031 1492
rect 9997 1344 10031 1378
rect 9997 1276 10031 1310
rect 9997 1208 10031 1242
rect 9997 1157 10031 1174
rect 10085 1412 10119 1450
rect 10085 1344 10119 1378
rect 10085 1276 10119 1310
rect 10085 1208 10119 1242
rect 9909 1094 9943 1105
rect 10085 1139 10119 1174
rect 10173 1412 10207 1492
rect 10173 1344 10207 1378
rect 10173 1276 10207 1310
rect 10173 1208 10207 1242
rect 10173 1157 10207 1174
rect 10261 1412 10295 1450
rect 10261 1344 10295 1378
rect 10261 1276 10295 1310
rect 10261 1208 10295 1242
rect 10085 1094 10119 1105
rect 10261 1139 10295 1174
rect 10349 1412 10383 1492
rect 10349 1344 10383 1378
rect 10349 1276 10383 1310
rect 10349 1208 10383 1242
rect 10349 1157 10383 1174
rect 10551 1470 10613 1492
rect 10551 1436 10565 1470
rect 10599 1436 10613 1470
rect 10551 1398 10613 1436
rect 10551 1364 10565 1398
rect 10599 1364 10613 1398
rect 10551 1326 10613 1364
rect 10551 1292 10565 1326
rect 10599 1292 10613 1326
rect 10551 1254 10613 1292
rect 10551 1220 10565 1254
rect 10599 1220 10613 1254
rect 10551 1182 10613 1220
rect 10261 1094 10295 1105
rect 10551 1148 10565 1182
rect 10599 1148 10613 1182
rect 10551 1110 10613 1148
rect 9589 1038 9651 1076
rect 9909 1060 10451 1094
rect 9589 1004 9603 1038
rect 9637 1004 9651 1038
rect 9589 966 9651 1004
rect 9589 932 9603 966
rect 9637 932 9651 966
rect 9589 868 9651 932
rect 9825 1003 9859 1019
rect 8627 368 8641 402
rect 8675 368 8689 402
rect 8396 247 8430 344
rect 8627 330 8689 368
rect 8396 197 8430 213
rect 8493 291 8527 307
rect 8493 223 8527 257
rect 8185 153 8219 169
rect 8025 119 8088 153
rect 8122 119 8185 153
rect 7991 103 8025 119
rect 8185 103 8219 119
rect 8299 153 8333 189
rect 8493 153 8527 189
rect 8333 119 8396 153
rect 8430 119 8493 153
rect 8299 103 8333 119
rect 8493 103 8527 119
rect 8627 296 8641 330
rect 8675 296 8689 330
rect 8627 258 8689 296
rect 8627 224 8641 258
rect 8675 224 8689 258
rect 8627 186 8689 224
rect 8627 152 8641 186
rect 8675 152 8689 186
rect 8627 114 8689 152
rect 8627 80 8641 114
rect 8675 80 8689 114
rect 8759 363 8793 379
rect 8953 363 8987 379
rect 9147 363 9181 379
rect 8793 329 8856 363
rect 8890 329 8953 363
rect 8987 329 9050 363
rect 9084 329 9147 363
rect 8759 291 8793 329
rect 8759 223 8793 257
rect 8953 291 8987 329
rect 9147 313 9181 329
rect 9261 363 9295 379
rect 9455 378 9489 797
rect 9825 757 9859 969
rect 9261 291 9295 329
rect 8759 153 8793 189
rect 8759 103 8793 119
rect 8856 238 8890 254
rect 8627 62 8689 80
rect 8856 62 8890 204
rect 8953 223 8987 257
rect 9051 244 9085 260
rect 9261 244 9295 257
rect 9085 223 9295 244
rect 9085 210 9261 223
rect 9051 194 9085 210
rect 8953 153 8987 189
rect 9358 344 9489 378
rect 9589 546 9651 572
rect 9589 512 9603 546
rect 9637 512 9651 546
rect 9589 474 9651 512
rect 9589 440 9603 474
rect 9637 440 9651 474
rect 9589 402 9651 440
rect 9825 461 9859 723
rect 9825 411 9859 427
rect 10047 1003 10081 1019
rect 10047 535 10081 969
rect 10047 461 10081 501
rect 10047 411 10081 427
rect 10269 1003 10303 1019
rect 10269 609 10303 969
rect 10269 461 10303 575
rect 10269 411 10303 427
rect 10417 757 10451 1060
rect 10551 1076 10565 1110
rect 10599 1076 10613 1110
rect 10783 1412 10817 1492
rect 10783 1344 10817 1378
rect 10783 1276 10817 1310
rect 10783 1208 10817 1242
rect 10783 1139 10817 1174
rect 10783 1089 10817 1105
rect 10871 1412 10905 1450
rect 10871 1344 10905 1378
rect 10871 1276 10905 1310
rect 10871 1208 10905 1242
rect 10871 1139 10905 1174
rect 10959 1412 10993 1492
rect 10959 1344 10993 1378
rect 10959 1276 10993 1310
rect 10959 1208 10993 1242
rect 10959 1157 10993 1174
rect 11047 1412 11081 1450
rect 11047 1344 11081 1378
rect 11047 1276 11081 1310
rect 11047 1208 11081 1242
rect 10871 1094 10905 1105
rect 11047 1139 11081 1174
rect 11135 1412 11169 1492
rect 11135 1344 11169 1378
rect 11135 1276 11169 1310
rect 11135 1208 11169 1242
rect 11135 1157 11169 1174
rect 11223 1412 11257 1450
rect 11223 1344 11257 1378
rect 11223 1276 11257 1310
rect 11223 1208 11257 1242
rect 11047 1094 11081 1105
rect 11223 1139 11257 1174
rect 11311 1412 11345 1492
rect 11311 1344 11345 1378
rect 11311 1276 11345 1310
rect 11311 1208 11345 1242
rect 11311 1157 11345 1174
rect 11513 1470 11575 1492
rect 11513 1436 11527 1470
rect 11561 1436 11575 1470
rect 11513 1398 11575 1436
rect 11513 1364 11527 1398
rect 11561 1364 11575 1398
rect 11513 1326 11575 1364
rect 11513 1292 11527 1326
rect 11561 1292 11575 1326
rect 11513 1254 11575 1292
rect 11513 1220 11527 1254
rect 11561 1220 11575 1254
rect 11513 1182 11575 1220
rect 11223 1094 11257 1105
rect 11513 1148 11527 1182
rect 11561 1148 11575 1182
rect 11513 1110 11575 1148
rect 10551 1038 10613 1076
rect 10871 1060 11413 1094
rect 10551 1004 10565 1038
rect 10599 1004 10613 1038
rect 10551 966 10613 1004
rect 10551 932 10565 966
rect 10599 932 10613 966
rect 10551 868 10613 932
rect 10787 1003 10821 1019
rect 9589 368 9603 402
rect 9637 368 9651 402
rect 9358 247 9392 344
rect 9589 330 9651 368
rect 9358 197 9392 213
rect 9455 291 9489 307
rect 9455 223 9489 257
rect 9147 153 9181 169
rect 8987 119 9050 153
rect 9084 119 9147 153
rect 8953 103 8987 119
rect 9147 103 9181 119
rect 9261 153 9295 189
rect 9455 153 9489 189
rect 9295 119 9358 153
rect 9392 119 9455 153
rect 9261 103 9295 119
rect 9455 103 9489 119
rect 9589 296 9603 330
rect 9637 296 9651 330
rect 9589 258 9651 296
rect 9589 224 9603 258
rect 9637 224 9651 258
rect 9589 186 9651 224
rect 9589 152 9603 186
rect 9637 152 9651 186
rect 9589 114 9651 152
rect 9589 80 9603 114
rect 9637 80 9651 114
rect 9721 363 9755 379
rect 9915 363 9949 379
rect 10109 363 10143 379
rect 9755 329 9818 363
rect 9852 329 9915 363
rect 9949 329 10012 363
rect 10046 329 10109 363
rect 9721 291 9755 329
rect 9721 223 9755 257
rect 9915 291 9949 329
rect 10109 313 10143 329
rect 10223 363 10257 379
rect 10417 378 10451 723
rect 10787 757 10821 969
rect 10223 291 10257 329
rect 9721 153 9755 189
rect 9721 103 9755 119
rect 9818 238 9852 254
rect 9589 62 9651 80
rect 9818 62 9852 204
rect 9915 223 9949 257
rect 10013 244 10047 260
rect 10223 244 10257 257
rect 10047 223 10257 244
rect 10047 210 10223 223
rect 10013 194 10047 210
rect 9915 153 9949 189
rect 10320 344 10451 378
rect 10551 546 10613 572
rect 10551 512 10565 546
rect 10599 512 10613 546
rect 10551 474 10613 512
rect 10551 440 10565 474
rect 10599 440 10613 474
rect 10551 402 10613 440
rect 10787 461 10821 723
rect 10787 411 10821 427
rect 11009 1003 11043 1019
rect 11009 461 11043 969
rect 11009 411 11043 427
rect 11231 1003 11265 1019
rect 11231 831 11265 969
rect 11231 461 11265 797
rect 11231 411 11265 427
rect 11379 831 11413 1060
rect 11513 1076 11527 1110
rect 11561 1076 11575 1110
rect 11745 1412 11779 1492
rect 11745 1344 11779 1378
rect 11745 1276 11779 1310
rect 11745 1208 11779 1242
rect 11745 1139 11779 1174
rect 11745 1089 11779 1105
rect 11833 1412 11867 1450
rect 11833 1344 11867 1378
rect 11833 1276 11867 1310
rect 11833 1208 11867 1242
rect 11833 1139 11867 1174
rect 11921 1412 11955 1492
rect 11921 1344 11955 1378
rect 11921 1276 11955 1310
rect 11921 1208 11955 1242
rect 11921 1157 11955 1174
rect 12009 1412 12043 1450
rect 12009 1344 12043 1378
rect 12009 1276 12043 1310
rect 12009 1208 12043 1242
rect 11833 1094 11867 1105
rect 12009 1139 12043 1174
rect 12097 1412 12131 1492
rect 12097 1344 12131 1378
rect 12097 1276 12131 1310
rect 12097 1208 12131 1242
rect 12097 1157 12131 1174
rect 12185 1412 12219 1450
rect 12185 1344 12219 1378
rect 12185 1276 12219 1310
rect 12185 1208 12219 1242
rect 12009 1094 12043 1105
rect 12185 1139 12219 1174
rect 12273 1412 12307 1492
rect 12273 1344 12307 1378
rect 12273 1276 12307 1310
rect 12273 1208 12307 1242
rect 12273 1157 12307 1174
rect 12475 1470 12537 1492
rect 12475 1436 12489 1470
rect 12523 1436 12537 1470
rect 12475 1398 12537 1436
rect 12475 1364 12489 1398
rect 12523 1364 12537 1398
rect 12475 1326 12537 1364
rect 12475 1292 12489 1326
rect 12523 1292 12537 1326
rect 12475 1254 12537 1292
rect 12475 1220 12489 1254
rect 12523 1220 12537 1254
rect 12475 1182 12537 1220
rect 12185 1094 12219 1105
rect 12475 1148 12489 1182
rect 12523 1148 12537 1182
rect 12475 1110 12537 1148
rect 11513 1038 11575 1076
rect 11833 1060 12375 1094
rect 11513 1004 11527 1038
rect 11561 1004 11575 1038
rect 11513 966 11575 1004
rect 11513 932 11527 966
rect 11561 932 11575 966
rect 11513 868 11575 932
rect 11749 1003 11783 1019
rect 11749 905 11783 969
rect 11379 609 11413 797
rect 10551 368 10565 402
rect 10599 368 10613 402
rect 10320 247 10354 344
rect 10551 330 10613 368
rect 10320 197 10354 213
rect 10417 291 10451 307
rect 10417 223 10451 257
rect 10109 153 10143 169
rect 9949 119 10012 153
rect 10046 119 10109 153
rect 9915 103 9949 119
rect 10109 103 10143 119
rect 10223 153 10257 189
rect 10417 153 10451 189
rect 10257 119 10320 153
rect 10354 119 10417 153
rect 10223 103 10257 119
rect 10417 103 10451 119
rect 10551 296 10565 330
rect 10599 296 10613 330
rect 10551 258 10613 296
rect 10551 224 10565 258
rect 10599 224 10613 258
rect 10551 186 10613 224
rect 10551 152 10565 186
rect 10599 152 10613 186
rect 10551 114 10613 152
rect 10551 80 10565 114
rect 10599 80 10613 114
rect 10683 363 10717 379
rect 10877 363 10911 379
rect 11071 363 11105 379
rect 10717 329 10780 363
rect 10814 329 10877 363
rect 10911 329 10974 363
rect 11008 329 11071 363
rect 10683 291 10717 329
rect 10683 223 10717 257
rect 10877 291 10911 329
rect 11071 313 11105 329
rect 11185 363 11219 379
rect 11379 378 11413 575
rect 11185 291 11219 329
rect 10683 153 10717 189
rect 10683 103 10717 119
rect 10780 238 10814 254
rect 10551 62 10613 80
rect 10780 62 10814 204
rect 10877 223 10911 257
rect 10975 244 11009 260
rect 11185 244 11219 257
rect 11009 223 11219 244
rect 11009 210 11185 223
rect 10975 194 11009 210
rect 10877 153 10911 189
rect 11282 344 11413 378
rect 11513 546 11575 572
rect 11513 512 11527 546
rect 11561 512 11575 546
rect 11513 474 11575 512
rect 11513 440 11527 474
rect 11561 440 11575 474
rect 11513 402 11575 440
rect 11749 461 11783 871
rect 11749 411 11783 427
rect 11971 1003 12005 1019
rect 11971 535 12005 969
rect 11971 461 12005 501
rect 11971 411 12005 427
rect 12193 1003 12227 1019
rect 12193 757 12227 969
rect 12193 461 12227 723
rect 12193 411 12227 427
rect 12341 610 12375 1060
rect 12475 1076 12489 1110
rect 12523 1076 12537 1110
rect 12707 1412 12741 1492
rect 12707 1344 12741 1378
rect 12707 1276 12741 1310
rect 12707 1208 12741 1242
rect 12707 1139 12741 1174
rect 12707 1089 12741 1105
rect 12795 1412 12829 1450
rect 12795 1344 12829 1378
rect 12795 1276 12829 1310
rect 12795 1208 12829 1242
rect 12795 1139 12829 1174
rect 12883 1412 12917 1492
rect 12883 1344 12917 1378
rect 12883 1276 12917 1310
rect 12883 1208 12917 1242
rect 12883 1157 12917 1174
rect 12971 1412 13005 1450
rect 12971 1344 13005 1378
rect 12971 1276 13005 1310
rect 12971 1208 13005 1242
rect 12795 1094 12829 1105
rect 12971 1139 13005 1174
rect 13059 1412 13093 1492
rect 13059 1344 13093 1378
rect 13059 1276 13093 1310
rect 13059 1208 13093 1242
rect 13059 1157 13093 1174
rect 13147 1412 13181 1450
rect 13147 1344 13181 1378
rect 13147 1276 13181 1310
rect 13147 1208 13181 1242
rect 12971 1094 13005 1105
rect 13147 1139 13181 1174
rect 13235 1412 13269 1492
rect 13235 1344 13269 1378
rect 13235 1276 13269 1310
rect 13235 1208 13269 1242
rect 13235 1157 13269 1174
rect 13437 1470 13499 1492
rect 13437 1436 13451 1470
rect 13485 1436 13499 1470
rect 13437 1398 13499 1436
rect 13437 1364 13451 1398
rect 13485 1364 13499 1398
rect 13437 1326 13499 1364
rect 13437 1292 13451 1326
rect 13485 1292 13499 1326
rect 13437 1254 13499 1292
rect 13437 1220 13451 1254
rect 13485 1220 13499 1254
rect 13437 1182 13499 1220
rect 13147 1094 13181 1105
rect 13437 1148 13451 1182
rect 13485 1148 13499 1182
rect 13437 1110 13499 1148
rect 12475 1038 12537 1076
rect 12795 1060 13337 1094
rect 12475 1004 12489 1038
rect 12523 1004 12537 1038
rect 12475 966 12537 1004
rect 12475 932 12489 966
rect 12523 932 12537 966
rect 12475 868 12537 932
rect 12711 1003 12745 1019
rect 12933 1003 12967 1019
rect 11513 368 11527 402
rect 11561 368 11575 402
rect 11282 247 11316 344
rect 11513 330 11575 368
rect 11282 197 11316 213
rect 11379 291 11413 307
rect 11379 223 11413 257
rect 11071 153 11105 169
rect 10911 119 10974 153
rect 11008 119 11071 153
rect 10877 103 10911 119
rect 11071 103 11105 119
rect 11185 153 11219 189
rect 11379 153 11413 189
rect 11219 119 11282 153
rect 11316 119 11379 153
rect 11185 103 11219 119
rect 11379 103 11413 119
rect 11513 296 11527 330
rect 11561 296 11575 330
rect 11513 258 11575 296
rect 11513 224 11527 258
rect 11561 224 11575 258
rect 11513 186 11575 224
rect 11513 152 11527 186
rect 11561 152 11575 186
rect 11513 114 11575 152
rect 11513 80 11527 114
rect 11561 80 11575 114
rect 11645 363 11679 379
rect 11839 363 11873 379
rect 12033 363 12067 379
rect 11679 329 11742 363
rect 11776 329 11839 363
rect 11873 329 11936 363
rect 11970 329 12033 363
rect 11645 291 11679 329
rect 11645 223 11679 257
rect 11839 291 11873 329
rect 12033 313 12067 329
rect 12147 363 12181 379
rect 12341 378 12375 576
rect 12711 610 12745 969
rect 12932 979 12933 995
rect 12966 945 12967 969
rect 12932 929 12967 945
rect 12147 291 12181 329
rect 11645 153 11679 189
rect 11645 103 11679 119
rect 11742 238 11776 254
rect 11513 62 11575 80
rect 11742 62 11776 204
rect 11839 223 11873 257
rect 11937 244 11971 260
rect 12147 244 12181 257
rect 11971 223 12181 244
rect 11971 210 12147 223
rect 11937 194 11971 210
rect 11839 153 11873 189
rect 12244 344 12375 378
rect 12475 546 12537 572
rect 12475 512 12489 546
rect 12523 512 12537 546
rect 12475 474 12537 512
rect 12475 440 12489 474
rect 12523 440 12537 474
rect 12475 402 12537 440
rect 12711 461 12745 576
rect 12711 411 12745 427
rect 12933 461 12967 929
rect 13155 1003 13189 1019
rect 13155 847 13189 969
rect 13154 831 13189 847
rect 13188 797 13189 831
rect 13154 781 13189 797
rect 12933 411 12967 427
rect 13155 461 13189 781
rect 13155 411 13189 427
rect 13303 757 13337 1060
rect 13437 1076 13451 1110
rect 13485 1076 13499 1110
rect 13669 1412 13703 1492
rect 13669 1344 13703 1378
rect 13669 1276 13703 1310
rect 13669 1208 13703 1242
rect 13669 1139 13703 1174
rect 13669 1089 13703 1105
rect 13757 1412 13791 1450
rect 13757 1344 13791 1378
rect 13757 1276 13791 1310
rect 13757 1208 13791 1242
rect 13757 1139 13791 1174
rect 13845 1412 13879 1492
rect 13845 1344 13879 1378
rect 13845 1276 13879 1310
rect 13845 1208 13879 1242
rect 13845 1157 13879 1174
rect 13933 1412 13967 1450
rect 13933 1344 13967 1378
rect 13933 1276 13967 1310
rect 13933 1208 13967 1242
rect 13757 1094 13791 1105
rect 13933 1139 13967 1174
rect 14021 1412 14055 1492
rect 14021 1344 14055 1378
rect 14021 1276 14055 1310
rect 14021 1208 14055 1242
rect 14021 1157 14055 1174
rect 14109 1412 14143 1450
rect 14109 1344 14143 1378
rect 14109 1276 14143 1310
rect 14109 1208 14143 1242
rect 13933 1094 13967 1105
rect 14109 1139 14143 1174
rect 14197 1412 14231 1492
rect 14197 1344 14231 1378
rect 14197 1276 14231 1310
rect 14197 1208 14231 1242
rect 14197 1157 14231 1174
rect 14399 1470 14461 1492
rect 14399 1436 14413 1470
rect 14447 1436 14461 1470
rect 14399 1398 14461 1436
rect 14399 1364 14413 1398
rect 14447 1364 14461 1398
rect 14399 1326 14461 1364
rect 14399 1292 14413 1326
rect 14447 1292 14461 1326
rect 14399 1254 14461 1292
rect 14399 1220 14413 1254
rect 14447 1220 14461 1254
rect 14399 1182 14461 1220
rect 14109 1094 14143 1105
rect 14399 1148 14413 1182
rect 14447 1148 14461 1182
rect 14399 1110 14461 1148
rect 13437 1038 13499 1076
rect 13757 1060 14299 1094
rect 13437 1004 13451 1038
rect 13485 1004 13499 1038
rect 13437 966 13499 1004
rect 13437 932 13451 966
rect 13485 932 13499 966
rect 13437 868 13499 932
rect 13673 1003 13707 1019
rect 12475 368 12489 402
rect 12523 368 12537 402
rect 12244 247 12278 344
rect 12475 330 12537 368
rect 12244 197 12278 213
rect 12341 291 12375 307
rect 12341 223 12375 257
rect 12033 153 12067 169
rect 11873 119 11936 153
rect 11970 119 12033 153
rect 11839 103 11873 119
rect 12033 103 12067 119
rect 12147 153 12181 189
rect 12341 153 12375 189
rect 12181 119 12244 153
rect 12278 119 12341 153
rect 12147 103 12181 119
rect 12341 103 12375 119
rect 12475 296 12489 330
rect 12523 296 12537 330
rect 12475 258 12537 296
rect 12475 224 12489 258
rect 12523 224 12537 258
rect 12475 186 12537 224
rect 12475 152 12489 186
rect 12523 152 12537 186
rect 12475 114 12537 152
rect 12475 80 12489 114
rect 12523 80 12537 114
rect 12607 363 12641 379
rect 12801 363 12835 379
rect 12995 363 13029 379
rect 12641 329 12704 363
rect 12738 329 12801 363
rect 12835 329 12898 363
rect 12932 329 12995 363
rect 12607 291 12641 329
rect 12607 223 12641 257
rect 12801 291 12835 329
rect 12995 313 13029 329
rect 13109 363 13143 379
rect 13303 378 13337 723
rect 13673 610 13707 969
rect 13109 291 13143 329
rect 12607 153 12641 189
rect 12607 103 12641 119
rect 12704 238 12738 254
rect 12475 62 12537 80
rect 12704 62 12738 204
rect 12801 223 12835 257
rect 12899 244 12933 260
rect 13109 244 13143 257
rect 12933 223 13143 244
rect 12933 210 13109 223
rect 12899 194 12933 210
rect 12801 153 12835 189
rect 13206 344 13337 378
rect 13437 546 13499 572
rect 13437 512 13451 546
rect 13485 512 13499 546
rect 13437 474 13499 512
rect 13437 440 13451 474
rect 13485 440 13499 474
rect 13437 402 13499 440
rect 13673 461 13707 576
rect 13673 411 13707 427
rect 13895 1003 13929 1019
rect 13895 462 13929 969
rect 13895 411 13929 427
rect 14117 1003 14151 1019
rect 14117 831 14151 969
rect 14117 461 14151 797
rect 14117 411 14151 427
rect 14265 609 14299 1060
rect 14399 1076 14413 1110
rect 14447 1076 14461 1110
rect 14631 1412 14665 1492
rect 14631 1344 14665 1378
rect 14631 1276 14665 1310
rect 14631 1208 14665 1242
rect 14631 1139 14665 1174
rect 14631 1089 14665 1105
rect 14719 1412 14753 1450
rect 14719 1344 14753 1378
rect 14719 1276 14753 1310
rect 14719 1208 14753 1242
rect 14719 1139 14753 1174
rect 14807 1412 14841 1492
rect 14807 1344 14841 1378
rect 14807 1276 14841 1310
rect 14807 1208 14841 1242
rect 14807 1157 14841 1174
rect 14895 1412 14929 1450
rect 14895 1344 14929 1378
rect 14895 1276 14929 1310
rect 14895 1208 14929 1242
rect 14719 1094 14753 1105
rect 14895 1139 14929 1174
rect 14983 1412 15017 1492
rect 14983 1344 15017 1378
rect 14983 1276 15017 1310
rect 14983 1208 15017 1242
rect 14983 1157 15017 1174
rect 15071 1412 15105 1450
rect 15071 1344 15105 1378
rect 15071 1276 15105 1310
rect 15071 1208 15105 1242
rect 14895 1094 14929 1105
rect 15071 1139 15105 1174
rect 15159 1412 15193 1492
rect 15159 1344 15193 1378
rect 15159 1276 15193 1310
rect 15159 1208 15193 1242
rect 15159 1157 15193 1174
rect 15361 1470 15423 1492
rect 15361 1436 15375 1470
rect 15409 1436 15423 1470
rect 15361 1398 15423 1436
rect 15361 1364 15375 1398
rect 15409 1364 15423 1398
rect 15361 1326 15423 1364
rect 15361 1292 15375 1326
rect 15409 1292 15423 1326
rect 15361 1254 15423 1292
rect 15361 1220 15375 1254
rect 15409 1220 15423 1254
rect 15361 1182 15423 1220
rect 15071 1094 15105 1105
rect 15361 1148 15375 1182
rect 15409 1148 15423 1182
rect 15361 1110 15423 1148
rect 14399 1038 14461 1076
rect 14719 1060 15261 1094
rect 14399 1004 14413 1038
rect 14447 1004 14461 1038
rect 14399 966 14461 1004
rect 14399 932 14413 966
rect 14447 932 14461 966
rect 14399 868 14461 932
rect 14635 1003 14669 1019
rect 13437 368 13451 402
rect 13485 368 13499 402
rect 13206 247 13240 344
rect 13437 330 13499 368
rect 13206 197 13240 213
rect 13303 291 13337 307
rect 13303 223 13337 257
rect 12995 153 13029 169
rect 12835 119 12898 153
rect 12932 119 12995 153
rect 12801 103 12835 119
rect 12995 103 13029 119
rect 13109 153 13143 189
rect 13303 153 13337 189
rect 13143 119 13206 153
rect 13240 119 13303 153
rect 13109 103 13143 119
rect 13303 103 13337 119
rect 13437 296 13451 330
rect 13485 296 13499 330
rect 13437 258 13499 296
rect 13437 224 13451 258
rect 13485 224 13499 258
rect 13437 186 13499 224
rect 13437 152 13451 186
rect 13485 152 13499 186
rect 13437 114 13499 152
rect 13437 80 13451 114
rect 13485 80 13499 114
rect 13569 363 13603 379
rect 13763 363 13797 379
rect 13957 363 13991 379
rect 13603 329 13666 363
rect 13700 329 13763 363
rect 13797 329 13860 363
rect 13894 329 13957 363
rect 13569 291 13603 329
rect 13569 223 13603 257
rect 13763 291 13797 329
rect 13957 313 13991 329
rect 14071 363 14105 379
rect 14265 378 14299 575
rect 14635 609 14669 969
rect 14071 291 14105 329
rect 13569 153 13603 189
rect 13569 103 13603 119
rect 13666 238 13700 254
rect 13437 62 13499 80
rect 13666 62 13700 204
rect 13763 223 13797 257
rect 13861 244 13895 260
rect 14071 244 14105 257
rect 13895 223 14105 244
rect 13895 210 14071 223
rect 13861 194 13895 210
rect 13763 153 13797 189
rect 14168 344 14299 378
rect 14399 546 14461 572
rect 14399 512 14413 546
rect 14447 512 14461 546
rect 14399 474 14461 512
rect 14399 440 14413 474
rect 14447 440 14461 474
rect 14399 402 14461 440
rect 14635 461 14669 575
rect 14635 411 14669 427
rect 14857 1003 14891 1019
rect 14857 461 14891 945
rect 14857 411 14891 427
rect 15079 1003 15113 1019
rect 15079 535 15113 969
rect 15079 461 15113 501
rect 15079 411 15113 427
rect 15227 831 15261 1060
rect 15361 1076 15375 1110
rect 15409 1076 15423 1110
rect 15593 1412 15627 1492
rect 15593 1344 15627 1378
rect 15593 1276 15627 1310
rect 15593 1208 15627 1242
rect 15593 1139 15627 1174
rect 15593 1089 15627 1105
rect 15681 1412 15715 1450
rect 15681 1344 15715 1378
rect 15681 1276 15715 1310
rect 15681 1208 15715 1242
rect 15681 1139 15715 1174
rect 15769 1412 15803 1492
rect 15769 1344 15803 1378
rect 15769 1276 15803 1310
rect 15769 1208 15803 1242
rect 15769 1157 15803 1174
rect 15857 1412 15891 1450
rect 15857 1344 15891 1378
rect 15857 1276 15891 1310
rect 15857 1208 15891 1242
rect 15681 1094 15715 1105
rect 15857 1139 15891 1174
rect 15945 1412 15979 1492
rect 15945 1344 15979 1378
rect 15945 1276 15979 1310
rect 15945 1208 15979 1242
rect 15945 1157 15979 1174
rect 16033 1412 16067 1450
rect 16033 1344 16067 1378
rect 16033 1276 16067 1310
rect 16033 1208 16067 1242
rect 15857 1094 15891 1105
rect 16033 1139 16067 1174
rect 16121 1412 16155 1492
rect 16121 1344 16155 1378
rect 16121 1276 16155 1310
rect 16121 1208 16155 1242
rect 16121 1157 16155 1174
rect 16323 1470 16385 1492
rect 16323 1436 16337 1470
rect 16371 1436 16385 1470
rect 16323 1398 16385 1436
rect 16323 1364 16337 1398
rect 16371 1364 16385 1398
rect 16323 1326 16385 1364
rect 16323 1292 16337 1326
rect 16371 1292 16385 1326
rect 16323 1254 16385 1292
rect 16323 1220 16337 1254
rect 16371 1220 16385 1254
rect 16323 1182 16385 1220
rect 16033 1094 16067 1105
rect 16323 1148 16337 1182
rect 16371 1148 16385 1182
rect 16323 1110 16385 1148
rect 15361 1038 15423 1076
rect 15681 1060 16223 1094
rect 15361 1004 15375 1038
rect 15409 1004 15423 1038
rect 15361 966 15423 1004
rect 15361 932 15375 966
rect 15409 932 15423 966
rect 15361 868 15423 932
rect 15597 1003 15631 1019
rect 14399 368 14413 402
rect 14447 368 14461 402
rect 14168 247 14202 344
rect 14399 330 14461 368
rect 14168 197 14202 213
rect 14265 291 14299 307
rect 14265 223 14299 257
rect 13957 153 13991 169
rect 13797 119 13860 153
rect 13894 119 13957 153
rect 13763 103 13797 119
rect 13957 103 13991 119
rect 14071 153 14105 189
rect 14265 153 14299 189
rect 14105 119 14168 153
rect 14202 119 14265 153
rect 14071 103 14105 119
rect 14265 103 14299 119
rect 14399 296 14413 330
rect 14447 296 14461 330
rect 14399 258 14461 296
rect 14399 224 14413 258
rect 14447 224 14461 258
rect 14399 186 14461 224
rect 14399 152 14413 186
rect 14447 152 14461 186
rect 14399 114 14461 152
rect 14399 80 14413 114
rect 14447 80 14461 114
rect 14531 363 14565 379
rect 14725 363 14759 379
rect 14919 363 14953 379
rect 14565 329 14628 363
rect 14662 329 14725 363
rect 14759 329 14822 363
rect 14856 329 14919 363
rect 14531 291 14565 329
rect 14531 223 14565 257
rect 14725 291 14759 329
rect 14919 313 14953 329
rect 15033 363 15067 379
rect 15227 378 15261 797
rect 15597 757 15631 969
rect 15033 291 15067 329
rect 14531 153 14565 189
rect 14531 103 14565 119
rect 14628 238 14662 254
rect 14399 62 14461 80
rect 14628 62 14662 204
rect 14725 223 14759 257
rect 14823 244 14857 260
rect 15033 244 15067 257
rect 14857 223 15067 244
rect 14857 210 15033 223
rect 14823 194 14857 210
rect 14725 153 14759 189
rect 15130 344 15261 378
rect 15361 546 15423 572
rect 15361 512 15375 546
rect 15409 512 15423 546
rect 15361 474 15423 512
rect 15361 440 15375 474
rect 15409 440 15423 474
rect 15361 402 15423 440
rect 15597 461 15631 723
rect 15597 411 15631 427
rect 15819 1003 15853 1019
rect 15819 535 15853 969
rect 15819 461 15853 501
rect 15819 411 15853 427
rect 16041 1003 16075 1019
rect 16041 609 16075 969
rect 16041 461 16075 575
rect 16041 411 16075 427
rect 16189 757 16223 1060
rect 16323 1076 16337 1110
rect 16371 1076 16385 1110
rect 16555 1412 16589 1492
rect 16555 1344 16589 1378
rect 16555 1276 16589 1310
rect 16555 1208 16589 1242
rect 16555 1139 16589 1174
rect 16555 1089 16589 1105
rect 16643 1412 16677 1450
rect 16643 1344 16677 1378
rect 16643 1276 16677 1310
rect 16643 1208 16677 1242
rect 16643 1139 16677 1174
rect 16731 1412 16765 1492
rect 16731 1344 16765 1378
rect 16731 1276 16765 1310
rect 16731 1208 16765 1242
rect 16731 1157 16765 1174
rect 16819 1412 16853 1450
rect 16819 1344 16853 1378
rect 16819 1276 16853 1310
rect 16819 1208 16853 1242
rect 16643 1094 16677 1105
rect 16819 1139 16853 1174
rect 16907 1412 16941 1492
rect 16907 1344 16941 1378
rect 16907 1276 16941 1310
rect 16907 1208 16941 1242
rect 16907 1157 16941 1174
rect 16995 1412 17029 1450
rect 16995 1344 17029 1378
rect 16995 1276 17029 1310
rect 16995 1208 17029 1242
rect 16819 1094 16853 1105
rect 16995 1139 17029 1174
rect 17083 1412 17117 1492
rect 17083 1344 17117 1378
rect 17083 1276 17117 1310
rect 17083 1208 17117 1242
rect 17083 1157 17117 1174
rect 17285 1470 17347 1492
rect 17285 1436 17299 1470
rect 17333 1436 17347 1470
rect 17285 1398 17347 1436
rect 17285 1364 17299 1398
rect 17333 1364 17347 1398
rect 17285 1326 17347 1364
rect 17285 1292 17299 1326
rect 17333 1292 17347 1326
rect 17285 1254 17347 1292
rect 17285 1220 17299 1254
rect 17333 1220 17347 1254
rect 17285 1182 17347 1220
rect 16995 1094 17029 1105
rect 17285 1148 17299 1182
rect 17333 1148 17347 1182
rect 17285 1110 17347 1148
rect 16323 1038 16385 1076
rect 16643 1060 17185 1094
rect 16323 1004 16337 1038
rect 16371 1004 16385 1038
rect 16323 966 16385 1004
rect 16323 932 16337 966
rect 16371 932 16385 966
rect 16323 868 16385 932
rect 16559 1003 16593 1019
rect 15361 368 15375 402
rect 15409 368 15423 402
rect 15130 247 15164 344
rect 15361 330 15423 368
rect 15130 197 15164 213
rect 15227 291 15261 307
rect 15227 223 15261 257
rect 14919 153 14953 169
rect 14759 119 14822 153
rect 14856 119 14919 153
rect 14725 103 14759 119
rect 14919 103 14953 119
rect 15033 153 15067 189
rect 15227 153 15261 189
rect 15067 119 15130 153
rect 15164 119 15227 153
rect 15033 103 15067 119
rect 15227 103 15261 119
rect 15361 296 15375 330
rect 15409 296 15423 330
rect 15361 258 15423 296
rect 15361 224 15375 258
rect 15409 224 15423 258
rect 15361 186 15423 224
rect 15361 152 15375 186
rect 15409 152 15423 186
rect 15361 114 15423 152
rect 15361 80 15375 114
rect 15409 80 15423 114
rect 15493 363 15527 379
rect 15687 363 15721 379
rect 15881 363 15915 379
rect 15527 329 15590 363
rect 15624 329 15687 363
rect 15721 329 15784 363
rect 15818 329 15881 363
rect 15493 291 15527 329
rect 15493 223 15527 257
rect 15687 291 15721 329
rect 15881 313 15915 329
rect 15995 363 16029 379
rect 16189 378 16223 723
rect 16559 757 16593 969
rect 15995 291 16029 329
rect 15493 153 15527 189
rect 15493 103 15527 119
rect 15590 238 15624 254
rect 15361 62 15423 80
rect 15590 62 15624 204
rect 15687 223 15721 257
rect 15785 244 15819 260
rect 15995 244 16029 257
rect 15819 223 16029 244
rect 15819 210 15995 223
rect 15785 194 15819 210
rect 15687 153 15721 189
rect 16092 344 16223 378
rect 16323 546 16385 572
rect 16323 512 16337 546
rect 16371 512 16385 546
rect 16323 474 16385 512
rect 16323 440 16337 474
rect 16371 440 16385 474
rect 16323 402 16385 440
rect 16559 461 16593 723
rect 16559 411 16593 427
rect 16781 1003 16815 1019
rect 16781 461 16815 969
rect 16781 411 16815 427
rect 17003 1003 17037 1019
rect 17003 831 17037 969
rect 17003 461 17037 797
rect 17003 411 17037 427
rect 17151 831 17185 1060
rect 17285 1076 17299 1110
rect 17333 1076 17347 1110
rect 17285 1038 17347 1076
rect 17457 1411 17491 1492
rect 17457 1343 17491 1377
rect 17457 1275 17491 1309
rect 17457 1207 17491 1241
rect 17457 1139 17491 1173
rect 17457 1071 17491 1105
rect 17545 1411 17581 1445
rect 17633 1411 17667 1492
rect 17545 1343 17579 1377
rect 17545 1275 17579 1309
rect 17545 1207 17579 1241
rect 17545 1139 17579 1173
rect 17633 1343 17667 1377
rect 17633 1275 17667 1309
rect 17633 1207 17667 1241
rect 17633 1157 17667 1173
rect 17721 1411 17755 1445
rect 17721 1343 17755 1377
rect 17721 1275 17755 1309
rect 17721 1207 17755 1241
rect 17721 1105 17755 1173
rect 17545 1071 17721 1105
rect 17809 1411 17843 1492
rect 17809 1343 17843 1377
rect 17809 1275 17843 1309
rect 17809 1207 17843 1241
rect 17809 1139 17843 1173
rect 17809 1071 17843 1105
rect 17951 1470 18013 1492
rect 17951 1436 17965 1470
rect 17999 1436 18013 1470
rect 18617 1470 18679 1492
rect 17951 1398 18013 1436
rect 17951 1364 17965 1398
rect 17999 1364 18013 1398
rect 17951 1326 18013 1364
rect 17951 1292 17965 1326
rect 17999 1292 18013 1326
rect 17951 1254 18013 1292
rect 17951 1220 17965 1254
rect 17999 1220 18013 1254
rect 17951 1182 18013 1220
rect 17951 1148 17965 1182
rect 17999 1148 18013 1182
rect 17951 1110 18013 1148
rect 17951 1076 17965 1110
rect 17999 1076 18013 1110
rect 17721 1055 17755 1071
rect 17285 1004 17299 1038
rect 17333 1004 17347 1038
rect 17951 1038 18013 1076
rect 18121 1411 18507 1445
rect 18121 1343 18155 1377
rect 18121 1275 18155 1309
rect 18121 1207 18155 1241
rect 18121 1105 18155 1173
rect 18209 1343 18243 1359
rect 18209 1275 18243 1309
rect 18209 1207 18243 1241
rect 18209 1139 18243 1173
rect 18297 1343 18331 1377
rect 18297 1275 18331 1309
rect 18297 1207 18331 1241
rect 18297 1157 18331 1173
rect 18385 1343 18419 1359
rect 18385 1275 18419 1309
rect 18385 1207 18419 1241
rect 18385 1105 18419 1173
rect 18473 1343 18507 1377
rect 18473 1275 18507 1309
rect 18473 1207 18507 1241
rect 18473 1121 18507 1173
rect 18617 1436 18631 1470
rect 18665 1436 18679 1470
rect 19283 1470 19345 1492
rect 18617 1398 18679 1436
rect 18617 1364 18631 1398
rect 18665 1364 18679 1398
rect 18617 1326 18679 1364
rect 18617 1292 18631 1326
rect 18665 1292 18679 1326
rect 18617 1254 18679 1292
rect 18617 1220 18631 1254
rect 18665 1220 18679 1254
rect 18617 1182 18679 1220
rect 18617 1148 18631 1182
rect 18665 1148 18679 1182
rect 18209 1071 18385 1105
rect 18121 1055 18155 1071
rect 18385 1055 18419 1071
rect 18617 1110 18679 1148
rect 18617 1076 18631 1110
rect 18665 1076 18679 1110
rect 17285 966 17347 1004
rect 17285 932 17299 966
rect 17333 932 17347 966
rect 17285 868 17347 932
rect 17447 1004 17481 1020
rect 17677 1004 17711 1020
rect 17151 609 17185 797
rect 16323 368 16337 402
rect 16371 368 16385 402
rect 16092 247 16126 344
rect 16323 330 16385 368
rect 16092 197 16126 213
rect 16189 291 16223 307
rect 16189 223 16223 257
rect 15881 153 15915 169
rect 15721 119 15784 153
rect 15818 119 15881 153
rect 15687 103 15721 119
rect 15881 103 15915 119
rect 15995 153 16029 189
rect 16189 153 16223 189
rect 16029 119 16092 153
rect 16126 119 16189 153
rect 15995 103 16029 119
rect 16189 103 16223 119
rect 16323 296 16337 330
rect 16371 296 16385 330
rect 16323 258 16385 296
rect 16323 224 16337 258
rect 16371 224 16385 258
rect 16323 186 16385 224
rect 16323 152 16337 186
rect 16371 152 16385 186
rect 16323 114 16385 152
rect 16323 80 16337 114
rect 16371 80 16385 114
rect 16455 363 16489 379
rect 16649 363 16683 379
rect 16843 363 16877 379
rect 16489 329 16552 363
rect 16586 329 16649 363
rect 16683 329 16746 363
rect 16780 329 16843 363
rect 16455 291 16489 329
rect 16455 223 16489 257
rect 16649 291 16683 329
rect 16843 313 16877 329
rect 16957 363 16991 379
rect 17151 378 17185 575
rect 17447 831 17481 945
rect 16957 291 16991 329
rect 16455 153 16489 189
rect 16455 103 16489 119
rect 16552 238 16586 254
rect 16323 62 16385 80
rect 16552 62 16586 204
rect 16649 223 16683 257
rect 16747 244 16781 260
rect 16957 244 16991 257
rect 16781 223 16991 244
rect 16781 210 16957 223
rect 16747 194 16781 210
rect 16649 153 16683 189
rect 17054 344 17185 378
rect 17285 546 17347 572
rect 17285 512 17299 546
rect 17333 512 17347 546
rect 17285 474 17347 512
rect 17285 440 17299 474
rect 17333 440 17347 474
rect 17285 402 17347 440
rect 17447 461 17481 797
rect 17447 411 17481 427
rect 17669 970 17677 988
rect 17669 954 17711 970
rect 17951 1004 17965 1038
rect 17999 1004 18013 1038
rect 18617 1038 18679 1076
rect 18789 1411 19175 1445
rect 18789 1343 18823 1377
rect 18789 1275 18823 1309
rect 18789 1207 18823 1241
rect 18789 1105 18823 1173
rect 18877 1343 18911 1359
rect 18877 1275 18911 1309
rect 18877 1207 18911 1241
rect 18877 1139 18911 1173
rect 18965 1343 18999 1377
rect 18965 1275 18999 1309
rect 18965 1207 18999 1241
rect 18965 1157 18999 1173
rect 19053 1343 19087 1359
rect 19053 1275 19087 1309
rect 19053 1207 19087 1241
rect 19053 1139 19087 1173
rect 19141 1343 19175 1377
rect 19141 1275 19175 1309
rect 19141 1207 19175 1241
rect 19141 1157 19175 1173
rect 19283 1436 19297 1470
rect 19331 1436 19345 1470
rect 19283 1398 19345 1436
rect 19283 1364 19297 1398
rect 19331 1364 19345 1398
rect 19283 1326 19345 1364
rect 19283 1292 19297 1326
rect 19331 1292 19345 1326
rect 19283 1254 19345 1292
rect 19283 1220 19297 1254
rect 19331 1220 19345 1254
rect 19283 1182 19345 1220
rect 19283 1148 19297 1182
rect 19331 1148 19345 1182
rect 19283 1110 19345 1148
rect 18877 1071 19183 1105
rect 18789 1055 18823 1071
rect 17951 966 18013 1004
rect 17669 905 17703 954
rect 17669 461 17703 871
rect 17951 932 17965 966
rect 17999 932 18013 966
rect 17951 868 18013 932
rect 18187 1004 18221 1020
rect 17669 411 17703 427
rect 17951 546 18013 572
rect 17951 512 17965 546
rect 17999 512 18013 546
rect 17951 474 18013 512
rect 17951 440 17965 474
rect 17999 440 18013 474
rect 17285 368 17299 402
rect 17333 368 17347 402
rect 17951 402 18013 440
rect 18187 461 18221 945
rect 18187 411 18221 427
rect 18483 1004 18517 1020
rect 18483 683 18517 970
rect 18617 1004 18631 1038
rect 18665 1004 18679 1038
rect 18617 966 18679 1004
rect 18617 932 18631 966
rect 18665 932 18679 966
rect 18617 868 18679 932
rect 18779 1004 18813 1020
rect 18483 461 18517 649
rect 18483 411 18517 427
rect 18617 546 18679 572
rect 18617 512 18631 546
rect 18665 512 18679 546
rect 18617 474 18679 512
rect 18617 440 18631 474
rect 18665 440 18679 474
rect 17054 247 17088 344
rect 17285 330 17347 368
rect 17054 197 17088 213
rect 17151 291 17185 307
rect 17151 223 17185 257
rect 16843 153 16877 169
rect 16683 119 16746 153
rect 16780 119 16843 153
rect 16649 103 16683 119
rect 16843 103 16877 119
rect 16957 153 16991 189
rect 17151 153 17185 189
rect 16991 119 17054 153
rect 17088 119 17151 153
rect 16957 103 16991 119
rect 17151 103 17185 119
rect 17285 296 17299 330
rect 17333 296 17347 330
rect 17285 258 17347 296
rect 17285 224 17299 258
rect 17333 224 17347 258
rect 17285 186 17347 224
rect 17285 152 17299 186
rect 17333 152 17347 186
rect 17285 114 17347 152
rect 17285 80 17299 114
rect 17333 80 17347 114
rect 17438 361 17472 377
rect 17632 361 17666 377
rect 17472 327 17535 361
rect 17569 327 17632 361
rect 17438 289 17472 327
rect 17438 221 17472 255
rect 17632 289 17666 327
rect 17826 361 17860 377
rect 17729 281 17763 297
rect 17438 151 17472 187
rect 17438 101 17472 117
rect 17535 236 17569 252
rect 17285 62 17347 80
rect 17535 62 17569 202
rect 17632 221 17666 255
rect 17728 247 17729 262
rect 17728 245 17763 247
rect 17762 231 17763 245
rect 17826 289 17860 327
rect 17728 195 17762 211
rect 17826 221 17860 255
rect 17632 151 17666 187
rect 17826 151 17860 187
rect 17666 117 17728 151
rect 17762 117 17826 151
rect 17632 101 17666 117
rect 17826 101 17860 117
rect 17951 368 17965 402
rect 17999 368 18013 402
rect 18617 402 18679 440
rect 18779 461 18813 970
rect 18779 411 18813 427
rect 19001 1004 19039 1020
rect 19001 970 19005 1004
rect 19001 954 19039 970
rect 19001 905 19035 954
rect 19001 461 19035 871
rect 19001 411 19035 427
rect 19149 831 19183 1071
rect 19283 1076 19297 1110
rect 19331 1076 19345 1110
rect 19283 1038 19345 1076
rect 19283 1004 19297 1038
rect 19331 1004 19345 1038
rect 19283 966 19345 1004
rect 19283 932 19297 966
rect 19331 932 19345 966
rect 19283 868 19345 932
rect 17951 330 18013 368
rect 17951 296 17965 330
rect 17999 296 18013 330
rect 17951 258 18013 296
rect 17951 224 17965 258
rect 17999 224 18013 258
rect 17951 186 18013 224
rect 17951 152 17965 186
rect 17999 152 18013 186
rect 17951 114 18013 152
rect 17951 80 17965 114
rect 17999 80 18013 114
rect 18104 361 18138 377
rect 18298 361 18332 377
rect 18138 327 18201 361
rect 18235 327 18298 361
rect 18104 289 18138 327
rect 18104 221 18138 255
rect 18298 289 18332 327
rect 18492 361 18526 377
rect 18104 151 18138 187
rect 18104 101 18138 117
rect 18201 236 18235 252
rect 17951 62 18013 80
rect 18201 62 18235 202
rect 18298 221 18332 255
rect 18395 281 18429 297
rect 18395 245 18429 247
rect 18395 195 18429 211
rect 18492 289 18526 327
rect 18492 221 18526 255
rect 18298 151 18332 187
rect 18492 151 18526 187
rect 18332 117 18395 151
rect 18429 117 18492 151
rect 18298 101 18332 117
rect 18492 101 18526 117
rect 18617 368 18631 402
rect 18665 368 18679 402
rect 18617 330 18679 368
rect 18617 296 18631 330
rect 18665 296 18679 330
rect 18617 258 18679 296
rect 18617 224 18631 258
rect 18665 224 18679 258
rect 18617 186 18679 224
rect 18617 152 18631 186
rect 18665 152 18679 186
rect 18617 114 18679 152
rect 18617 80 18631 114
rect 18665 80 18679 114
rect 18770 361 18804 377
rect 18964 361 18998 377
rect 19149 374 19183 797
rect 18804 327 18867 361
rect 18901 327 18964 361
rect 18770 289 18804 327
rect 18770 221 18804 255
rect 18964 289 18998 327
rect 18770 151 18804 187
rect 18770 101 18804 117
rect 18867 236 18901 252
rect 18617 62 18679 80
rect 18867 62 18901 202
rect 18964 221 18998 255
rect 19061 340 19183 374
rect 19283 546 19345 572
rect 19283 512 19297 546
rect 19331 512 19345 546
rect 19283 474 19345 512
rect 19283 440 19297 474
rect 19331 440 19345 474
rect 19283 402 19345 440
rect 19283 368 19297 402
rect 19331 368 19345 402
rect 19061 281 19095 340
rect 19283 330 19345 368
rect 19061 245 19095 247
rect 19061 195 19095 211
rect 19158 289 19192 306
rect 19158 221 19192 255
rect 18964 151 18998 187
rect 19158 151 19192 187
rect 18998 117 19061 151
rect 19095 117 19158 151
rect 18964 101 18998 117
rect 19158 101 19192 117
rect 19283 296 19297 330
rect 19331 296 19345 330
rect 19283 258 19345 296
rect 19283 224 19297 258
rect 19331 224 19345 258
rect 19283 186 19345 224
rect 19283 152 19297 186
rect 19331 152 19345 186
rect 19283 114 19345 152
rect 19283 80 19297 114
rect 19331 80 19345 114
rect 19283 62 19345 80
rect -31 47 18395 62
rect 18429 47 19345 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 343 47
rect 377 13 415 47
rect 449 13 513 47
rect 547 13 585 47
rect 619 13 657 47
rect 691 13 729 47
rect 763 13 801 47
rect 835 13 873 47
rect 907 13 1017 47
rect 1051 13 1089 47
rect 1123 13 1161 47
rect 1195 13 1233 47
rect 1267 13 1305 47
rect 1339 13 1377 47
rect 1411 13 1475 47
rect 1509 13 1547 47
rect 1581 13 1619 47
rect 1653 13 1691 47
rect 1725 13 1763 47
rect 1797 13 1835 47
rect 1869 13 1979 47
rect 2013 13 2051 47
rect 2085 13 2123 47
rect 2157 13 2195 47
rect 2229 13 2267 47
rect 2301 13 2339 47
rect 2373 13 2437 47
rect 2471 13 2509 47
rect 2543 13 2581 47
rect 2615 13 2653 47
rect 2687 13 2725 47
rect 2759 13 2797 47
rect 2831 13 2941 47
rect 2975 13 3013 47
rect 3047 13 3085 47
rect 3119 13 3157 47
rect 3191 13 3229 47
rect 3263 13 3301 47
rect 3335 13 3399 47
rect 3433 13 3471 47
rect 3505 13 3543 47
rect 3577 13 3615 47
rect 3649 13 3687 47
rect 3721 13 3759 47
rect 3793 13 3903 47
rect 3937 13 3975 47
rect 4009 13 4047 47
rect 4081 13 4119 47
rect 4153 13 4191 47
rect 4225 13 4263 47
rect 4297 13 4361 47
rect 4395 13 4433 47
rect 4467 13 4505 47
rect 4539 13 4577 47
rect 4611 13 4649 47
rect 4683 13 4721 47
rect 4755 13 4865 47
rect 4899 13 4937 47
rect 4971 13 5009 47
rect 5043 13 5081 47
rect 5115 13 5153 47
rect 5187 13 5225 47
rect 5259 13 5323 47
rect 5357 13 5395 47
rect 5429 13 5467 47
rect 5501 13 5539 47
rect 5573 13 5611 47
rect 5645 13 5683 47
rect 5717 13 5827 47
rect 5861 13 5899 47
rect 5933 13 5971 47
rect 6005 13 6043 47
rect 6077 13 6115 47
rect 6149 13 6187 47
rect 6221 13 6285 47
rect 6319 13 6357 47
rect 6391 13 6429 47
rect 6463 13 6501 47
rect 6535 13 6573 47
rect 6607 13 6645 47
rect 6679 13 6789 47
rect 6823 13 6861 47
rect 6895 13 6933 47
rect 6967 13 7005 47
rect 7039 13 7077 47
rect 7111 13 7149 47
rect 7183 13 7247 47
rect 7281 13 7319 47
rect 7353 13 7391 47
rect 7425 13 7463 47
rect 7497 13 7535 47
rect 7569 13 7607 47
rect 7641 13 7751 47
rect 7785 13 7823 47
rect 7857 13 7895 47
rect 7929 13 7967 47
rect 8001 13 8039 47
rect 8073 13 8111 47
rect 8145 13 8209 47
rect 8243 13 8281 47
rect 8315 13 8353 47
rect 8387 13 8425 47
rect 8459 13 8497 47
rect 8531 13 8569 47
rect 8603 13 8713 47
rect 8747 13 8785 47
rect 8819 13 8857 47
rect 8891 13 8929 47
rect 8963 13 9001 47
rect 9035 13 9073 47
rect 9107 13 9171 47
rect 9205 13 9243 47
rect 9277 13 9315 47
rect 9349 13 9387 47
rect 9421 13 9459 47
rect 9493 13 9531 47
rect 9565 13 9675 47
rect 9709 13 9747 47
rect 9781 13 9819 47
rect 9853 13 9891 47
rect 9925 13 9963 47
rect 9997 13 10035 47
rect 10069 13 10133 47
rect 10167 13 10205 47
rect 10239 13 10277 47
rect 10311 13 10349 47
rect 10383 13 10421 47
rect 10455 13 10493 47
rect 10527 13 10637 47
rect 10671 13 10709 47
rect 10743 13 10781 47
rect 10815 13 10853 47
rect 10887 13 10925 47
rect 10959 13 10997 47
rect 11031 13 11095 47
rect 11129 13 11167 47
rect 11201 13 11239 47
rect 11273 13 11311 47
rect 11345 13 11383 47
rect 11417 13 11455 47
rect 11489 13 11599 47
rect 11633 13 11671 47
rect 11705 13 11743 47
rect 11777 13 11815 47
rect 11849 13 11887 47
rect 11921 13 11959 47
rect 11993 13 12057 47
rect 12091 13 12129 47
rect 12163 13 12201 47
rect 12235 13 12273 47
rect 12307 13 12345 47
rect 12379 13 12417 47
rect 12451 13 12561 47
rect 12595 13 12633 47
rect 12667 13 12705 47
rect 12739 13 12777 47
rect 12811 13 12849 47
rect 12883 13 12921 47
rect 12955 13 13019 47
rect 13053 13 13091 47
rect 13125 13 13163 47
rect 13197 13 13235 47
rect 13269 13 13307 47
rect 13341 13 13379 47
rect 13413 13 13523 47
rect 13557 13 13595 47
rect 13629 13 13667 47
rect 13701 13 13739 47
rect 13773 13 13811 47
rect 13845 13 13883 47
rect 13917 13 13981 47
rect 14015 13 14053 47
rect 14087 13 14125 47
rect 14159 13 14197 47
rect 14231 13 14269 47
rect 14303 13 14341 47
rect 14375 13 14485 47
rect 14519 13 14557 47
rect 14591 13 14629 47
rect 14663 13 14701 47
rect 14735 13 14773 47
rect 14807 13 14845 47
rect 14879 13 14943 47
rect 14977 13 15015 47
rect 15049 13 15087 47
rect 15121 13 15159 47
rect 15193 13 15231 47
rect 15265 13 15303 47
rect 15337 13 15447 47
rect 15481 13 15519 47
rect 15553 13 15591 47
rect 15625 13 15663 47
rect 15697 13 15735 47
rect 15769 13 15807 47
rect 15841 13 15905 47
rect 15939 13 15977 47
rect 16011 13 16049 47
rect 16083 13 16121 47
rect 16155 13 16193 47
rect 16227 13 16265 47
rect 16299 13 16409 47
rect 16443 13 16481 47
rect 16515 13 16553 47
rect 16587 13 16625 47
rect 16659 13 16697 47
rect 16731 13 16769 47
rect 16803 13 16867 47
rect 16901 13 16939 47
rect 16973 13 17011 47
rect 17045 13 17083 47
rect 17117 13 17155 47
rect 17189 13 17227 47
rect 17261 13 17371 47
rect 17405 13 17443 47
rect 17477 13 17515 47
rect 17549 13 17587 47
rect 17621 13 17677 47
rect 17711 13 17749 47
rect 17783 13 17821 47
rect 17855 13 17893 47
rect 17927 13 18037 47
rect 18071 13 18109 47
rect 18143 13 18181 47
rect 18215 13 18253 47
rect 18287 13 18343 47
rect 18377 13 18415 47
rect 18449 13 18487 47
rect 18521 13 18559 47
rect 18593 13 18703 47
rect 18737 13 18775 47
rect 18809 13 18847 47
rect 18881 13 18919 47
rect 18953 13 19009 47
rect 19043 13 19081 47
rect 19115 13 19153 47
rect 19187 13 19225 47
rect 19259 13 19345 47
rect -31 0 19345 13
<< viali >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 343 1505 377 1539
rect 415 1505 449 1539
rect 513 1505 547 1539
rect 585 1505 619 1539
rect 657 1505 691 1539
rect 729 1505 763 1539
rect 801 1505 835 1539
rect 873 1505 907 1539
rect 1017 1505 1051 1539
rect 1089 1505 1123 1539
rect 1161 1505 1195 1539
rect 1233 1505 1267 1539
rect 1305 1505 1339 1539
rect 1377 1505 1411 1539
rect 1475 1505 1509 1539
rect 1547 1505 1581 1539
rect 1619 1505 1653 1539
rect 1691 1505 1725 1539
rect 1763 1505 1797 1539
rect 1835 1505 1869 1539
rect 1979 1505 2013 1539
rect 2051 1505 2085 1539
rect 2123 1505 2157 1539
rect 2195 1505 2229 1539
rect 2267 1505 2301 1539
rect 2339 1505 2373 1539
rect 2437 1505 2471 1539
rect 2509 1505 2543 1539
rect 2581 1505 2615 1539
rect 2653 1505 2687 1539
rect 2725 1505 2759 1539
rect 2797 1505 2831 1539
rect 2941 1505 2975 1539
rect 3013 1505 3047 1539
rect 3085 1505 3119 1539
rect 3157 1505 3191 1539
rect 3229 1505 3263 1539
rect 3301 1505 3335 1539
rect 3399 1505 3433 1539
rect 3471 1505 3505 1539
rect 3543 1505 3577 1539
rect 3615 1505 3649 1539
rect 3687 1505 3721 1539
rect 3759 1505 3793 1539
rect 3903 1505 3937 1539
rect 3975 1505 4009 1539
rect 4047 1505 4081 1539
rect 4119 1505 4153 1539
rect 4191 1505 4225 1539
rect 4263 1505 4297 1539
rect 4361 1505 4395 1539
rect 4433 1505 4467 1539
rect 4505 1505 4539 1539
rect 4577 1505 4611 1539
rect 4649 1505 4683 1539
rect 4721 1505 4755 1539
rect 4865 1505 4899 1539
rect 4937 1505 4971 1539
rect 5009 1505 5043 1539
rect 5081 1505 5115 1539
rect 5153 1505 5187 1539
rect 5225 1505 5259 1539
rect 5323 1505 5357 1539
rect 5395 1505 5429 1539
rect 5467 1505 5501 1539
rect 5539 1505 5573 1539
rect 5611 1505 5645 1539
rect 5683 1505 5717 1539
rect 5827 1505 5861 1539
rect 5899 1505 5933 1539
rect 5971 1505 6005 1539
rect 6043 1505 6077 1539
rect 6115 1505 6149 1539
rect 6187 1505 6221 1539
rect 6285 1505 6319 1539
rect 6357 1505 6391 1539
rect 6429 1505 6463 1539
rect 6501 1505 6535 1539
rect 6573 1505 6607 1539
rect 6645 1505 6679 1539
rect 6789 1505 6823 1539
rect 6861 1505 6895 1539
rect 6933 1505 6967 1539
rect 7005 1505 7039 1539
rect 7077 1505 7111 1539
rect 7149 1505 7183 1539
rect 7247 1505 7281 1539
rect 7319 1505 7353 1539
rect 7391 1505 7425 1539
rect 7463 1505 7497 1539
rect 7535 1505 7569 1539
rect 7607 1505 7641 1539
rect 7751 1505 7785 1539
rect 7823 1505 7857 1539
rect 7895 1505 7929 1539
rect 7967 1505 8001 1539
rect 8039 1505 8073 1539
rect 8111 1505 8145 1539
rect 8209 1505 8243 1539
rect 8281 1505 8315 1539
rect 8353 1505 8387 1539
rect 8425 1505 8459 1539
rect 8497 1505 8531 1539
rect 8569 1505 8603 1539
rect 8713 1505 8747 1539
rect 8785 1505 8819 1539
rect 8857 1505 8891 1539
rect 8929 1505 8963 1539
rect 9001 1505 9035 1539
rect 9073 1505 9107 1539
rect 9171 1505 9205 1539
rect 9243 1505 9277 1539
rect 9315 1505 9349 1539
rect 9387 1505 9421 1539
rect 9459 1505 9493 1539
rect 9531 1505 9565 1539
rect 9675 1505 9709 1539
rect 9747 1505 9781 1539
rect 9819 1505 9853 1539
rect 9891 1505 9925 1539
rect 9963 1505 9997 1539
rect 10035 1505 10069 1539
rect 10133 1505 10167 1539
rect 10205 1505 10239 1539
rect 10277 1505 10311 1539
rect 10349 1505 10383 1539
rect 10421 1505 10455 1539
rect 10493 1505 10527 1539
rect 10637 1505 10671 1539
rect 10709 1505 10743 1539
rect 10781 1505 10815 1539
rect 10853 1505 10887 1539
rect 10925 1505 10959 1539
rect 10997 1505 11031 1539
rect 11095 1505 11129 1539
rect 11167 1505 11201 1539
rect 11239 1505 11273 1539
rect 11311 1505 11345 1539
rect 11383 1505 11417 1539
rect 11455 1505 11489 1539
rect 11599 1505 11633 1539
rect 11671 1505 11705 1539
rect 11743 1505 11777 1539
rect 11815 1505 11849 1539
rect 11887 1505 11921 1539
rect 11959 1505 11993 1539
rect 12057 1505 12091 1539
rect 12129 1505 12163 1539
rect 12201 1505 12235 1539
rect 12273 1505 12307 1539
rect 12345 1505 12379 1539
rect 12417 1505 12451 1539
rect 12561 1505 12595 1539
rect 12633 1505 12667 1539
rect 12705 1505 12739 1539
rect 12777 1505 12811 1539
rect 12849 1505 12883 1539
rect 12921 1505 12955 1539
rect 13019 1505 13053 1539
rect 13091 1505 13125 1539
rect 13163 1505 13197 1539
rect 13235 1505 13269 1539
rect 13307 1505 13341 1539
rect 13379 1505 13413 1539
rect 13523 1505 13557 1539
rect 13595 1505 13629 1539
rect 13667 1505 13701 1539
rect 13739 1505 13773 1539
rect 13811 1505 13845 1539
rect 13883 1505 13917 1539
rect 13981 1505 14015 1539
rect 14053 1505 14087 1539
rect 14125 1505 14159 1539
rect 14197 1505 14231 1539
rect 14269 1505 14303 1539
rect 14341 1505 14375 1539
rect 14485 1505 14519 1539
rect 14557 1505 14591 1539
rect 14629 1505 14663 1539
rect 14701 1505 14735 1539
rect 14773 1505 14807 1539
rect 14845 1505 14879 1539
rect 14943 1505 14977 1539
rect 15015 1505 15049 1539
rect 15087 1505 15121 1539
rect 15159 1505 15193 1539
rect 15231 1505 15265 1539
rect 15303 1505 15337 1539
rect 15447 1505 15481 1539
rect 15519 1505 15553 1539
rect 15591 1505 15625 1539
rect 15663 1505 15697 1539
rect 15735 1505 15769 1539
rect 15807 1505 15841 1539
rect 15905 1505 15939 1539
rect 15977 1505 16011 1539
rect 16049 1505 16083 1539
rect 16121 1505 16155 1539
rect 16193 1505 16227 1539
rect 16265 1505 16299 1539
rect 16409 1505 16443 1539
rect 16481 1505 16515 1539
rect 16553 1505 16587 1539
rect 16625 1505 16659 1539
rect 16697 1505 16731 1539
rect 16769 1505 16803 1539
rect 16867 1505 16901 1539
rect 16939 1505 16973 1539
rect 17011 1505 17045 1539
rect 17083 1505 17117 1539
rect 17155 1505 17189 1539
rect 17227 1505 17261 1539
rect 17371 1505 17405 1539
rect 17443 1505 17477 1539
rect 17515 1505 17549 1539
rect 17587 1505 17621 1539
rect 17677 1505 17711 1539
rect 17749 1505 17783 1539
rect 17821 1505 17855 1539
rect 17893 1505 17927 1539
rect 18037 1505 18071 1539
rect 18109 1505 18143 1539
rect 18181 1505 18215 1539
rect 18253 1505 18287 1539
rect 18343 1505 18377 1539
rect 18415 1505 18449 1539
rect 18487 1505 18521 1539
rect 18559 1505 18593 1539
rect 18703 1505 18737 1539
rect 18775 1505 18809 1539
rect 18847 1505 18881 1539
rect 18919 1505 18953 1539
rect 19009 1505 19043 1539
rect 19081 1505 19115 1539
rect 19153 1505 19187 1539
rect 19225 1505 19259 1539
rect 205 871 239 905
rect 427 501 461 535
rect 649 723 683 757
rect 797 576 831 610
rect 1388 969 1389 979
rect 1389 969 1422 979
rect 1388 945 1422 969
rect 1167 576 1201 610
rect 1610 797 1644 831
rect 1759 723 1793 757
rect 2129 576 2163 610
rect 2351 461 2385 462
rect 2351 428 2385 461
rect 2573 797 2607 831
rect 2721 575 2755 609
rect 3091 575 3125 609
rect 3313 969 3347 979
rect 3313 945 3347 969
rect 3535 501 3569 535
rect 3683 797 3717 831
rect 4053 723 4087 757
rect 4275 501 4309 535
rect 4497 649 4531 683
rect 4645 723 4679 757
rect 5015 723 5049 757
rect 5237 427 5271 461
rect 5459 797 5493 831
rect 5977 871 6011 905
rect 5607 649 5641 683
rect 6199 501 6233 535
rect 6421 723 6455 757
rect 6569 576 6603 610
rect 7160 969 7161 979
rect 7161 969 7194 979
rect 7160 945 7194 969
rect 6939 576 6973 610
rect 7382 797 7416 831
rect 7531 723 7565 757
rect 7901 576 7935 610
rect 8123 461 8157 462
rect 8123 428 8157 461
rect 8345 797 8379 831
rect 8493 575 8527 609
rect 8863 575 8897 609
rect 9085 969 9119 979
rect 9085 945 9119 969
rect 9307 501 9341 535
rect 9455 797 9489 831
rect 9825 723 9859 757
rect 10047 501 10081 535
rect 10269 575 10303 609
rect 10417 723 10451 757
rect 10787 723 10821 757
rect 11009 427 11043 461
rect 11231 797 11265 831
rect 11749 871 11783 905
rect 11379 797 11413 831
rect 11379 575 11413 609
rect 11971 501 12005 535
rect 12193 723 12227 757
rect 12341 576 12375 610
rect 12932 969 12933 979
rect 12933 969 12966 979
rect 12932 945 12966 969
rect 12711 576 12745 610
rect 13154 797 13188 831
rect 13303 723 13337 757
rect 13673 576 13707 610
rect 13895 461 13929 462
rect 13895 428 13929 461
rect 14117 797 14151 831
rect 14265 575 14299 609
rect 14635 575 14669 609
rect 14857 969 14891 979
rect 14857 945 14891 969
rect 15079 501 15113 535
rect 15227 797 15261 831
rect 15597 723 15631 757
rect 15819 501 15853 535
rect 16041 575 16075 609
rect 16189 723 16223 757
rect 16559 723 16593 757
rect 16781 427 16815 461
rect 17003 797 17037 831
rect 17721 1071 17755 1105
rect 18121 1071 18155 1105
rect 18385 1071 18419 1105
rect 17447 970 17481 979
rect 17447 945 17481 970
rect 17151 797 17185 831
rect 17151 575 17185 609
rect 17447 797 17481 831
rect 18789 1071 18823 1105
rect 17669 871 17703 905
rect 18187 970 18221 979
rect 18187 945 18221 970
rect 18483 649 18517 683
rect 18483 427 18517 461
rect 17729 247 17763 281
rect 18779 427 18813 461
rect 19001 871 19035 905
rect 19149 797 19183 831
rect 18395 247 18429 281
rect 19061 247 19095 281
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 343 13 377 47
rect 415 13 449 47
rect 513 13 547 47
rect 585 13 619 47
rect 657 13 691 47
rect 729 13 763 47
rect 801 13 835 47
rect 873 13 907 47
rect 1017 13 1051 47
rect 1089 13 1123 47
rect 1161 13 1195 47
rect 1233 13 1267 47
rect 1305 13 1339 47
rect 1377 13 1411 47
rect 1475 13 1509 47
rect 1547 13 1581 47
rect 1619 13 1653 47
rect 1691 13 1725 47
rect 1763 13 1797 47
rect 1835 13 1869 47
rect 1979 13 2013 47
rect 2051 13 2085 47
rect 2123 13 2157 47
rect 2195 13 2229 47
rect 2267 13 2301 47
rect 2339 13 2373 47
rect 2437 13 2471 47
rect 2509 13 2543 47
rect 2581 13 2615 47
rect 2653 13 2687 47
rect 2725 13 2759 47
rect 2797 13 2831 47
rect 2941 13 2975 47
rect 3013 13 3047 47
rect 3085 13 3119 47
rect 3157 13 3191 47
rect 3229 13 3263 47
rect 3301 13 3335 47
rect 3399 13 3433 47
rect 3471 13 3505 47
rect 3543 13 3577 47
rect 3615 13 3649 47
rect 3687 13 3721 47
rect 3759 13 3793 47
rect 3903 13 3937 47
rect 3975 13 4009 47
rect 4047 13 4081 47
rect 4119 13 4153 47
rect 4191 13 4225 47
rect 4263 13 4297 47
rect 4361 13 4395 47
rect 4433 13 4467 47
rect 4505 13 4539 47
rect 4577 13 4611 47
rect 4649 13 4683 47
rect 4721 13 4755 47
rect 4865 13 4899 47
rect 4937 13 4971 47
rect 5009 13 5043 47
rect 5081 13 5115 47
rect 5153 13 5187 47
rect 5225 13 5259 47
rect 5323 13 5357 47
rect 5395 13 5429 47
rect 5467 13 5501 47
rect 5539 13 5573 47
rect 5611 13 5645 47
rect 5683 13 5717 47
rect 5827 13 5861 47
rect 5899 13 5933 47
rect 5971 13 6005 47
rect 6043 13 6077 47
rect 6115 13 6149 47
rect 6187 13 6221 47
rect 6285 13 6319 47
rect 6357 13 6391 47
rect 6429 13 6463 47
rect 6501 13 6535 47
rect 6573 13 6607 47
rect 6645 13 6679 47
rect 6789 13 6823 47
rect 6861 13 6895 47
rect 6933 13 6967 47
rect 7005 13 7039 47
rect 7077 13 7111 47
rect 7149 13 7183 47
rect 7247 13 7281 47
rect 7319 13 7353 47
rect 7391 13 7425 47
rect 7463 13 7497 47
rect 7535 13 7569 47
rect 7607 13 7641 47
rect 7751 13 7785 47
rect 7823 13 7857 47
rect 7895 13 7929 47
rect 7967 13 8001 47
rect 8039 13 8073 47
rect 8111 13 8145 47
rect 8209 13 8243 47
rect 8281 13 8315 47
rect 8353 13 8387 47
rect 8425 13 8459 47
rect 8497 13 8531 47
rect 8569 13 8603 47
rect 8713 13 8747 47
rect 8785 13 8819 47
rect 8857 13 8891 47
rect 8929 13 8963 47
rect 9001 13 9035 47
rect 9073 13 9107 47
rect 9171 13 9205 47
rect 9243 13 9277 47
rect 9315 13 9349 47
rect 9387 13 9421 47
rect 9459 13 9493 47
rect 9531 13 9565 47
rect 9675 13 9709 47
rect 9747 13 9781 47
rect 9819 13 9853 47
rect 9891 13 9925 47
rect 9963 13 9997 47
rect 10035 13 10069 47
rect 10133 13 10167 47
rect 10205 13 10239 47
rect 10277 13 10311 47
rect 10349 13 10383 47
rect 10421 13 10455 47
rect 10493 13 10527 47
rect 10637 13 10671 47
rect 10709 13 10743 47
rect 10781 13 10815 47
rect 10853 13 10887 47
rect 10925 13 10959 47
rect 10997 13 11031 47
rect 11095 13 11129 47
rect 11167 13 11201 47
rect 11239 13 11273 47
rect 11311 13 11345 47
rect 11383 13 11417 47
rect 11455 13 11489 47
rect 11599 13 11633 47
rect 11671 13 11705 47
rect 11743 13 11777 47
rect 11815 13 11849 47
rect 11887 13 11921 47
rect 11959 13 11993 47
rect 12057 13 12091 47
rect 12129 13 12163 47
rect 12201 13 12235 47
rect 12273 13 12307 47
rect 12345 13 12379 47
rect 12417 13 12451 47
rect 12561 13 12595 47
rect 12633 13 12667 47
rect 12705 13 12739 47
rect 12777 13 12811 47
rect 12849 13 12883 47
rect 12921 13 12955 47
rect 13019 13 13053 47
rect 13091 13 13125 47
rect 13163 13 13197 47
rect 13235 13 13269 47
rect 13307 13 13341 47
rect 13379 13 13413 47
rect 13523 13 13557 47
rect 13595 13 13629 47
rect 13667 13 13701 47
rect 13739 13 13773 47
rect 13811 13 13845 47
rect 13883 13 13917 47
rect 13981 13 14015 47
rect 14053 13 14087 47
rect 14125 13 14159 47
rect 14197 13 14231 47
rect 14269 13 14303 47
rect 14341 13 14375 47
rect 14485 13 14519 47
rect 14557 13 14591 47
rect 14629 13 14663 47
rect 14701 13 14735 47
rect 14773 13 14807 47
rect 14845 13 14879 47
rect 14943 13 14977 47
rect 15015 13 15049 47
rect 15087 13 15121 47
rect 15159 13 15193 47
rect 15231 13 15265 47
rect 15303 13 15337 47
rect 15447 13 15481 47
rect 15519 13 15553 47
rect 15591 13 15625 47
rect 15663 13 15697 47
rect 15735 13 15769 47
rect 15807 13 15841 47
rect 15905 13 15939 47
rect 15977 13 16011 47
rect 16049 13 16083 47
rect 16121 13 16155 47
rect 16193 13 16227 47
rect 16265 13 16299 47
rect 16409 13 16443 47
rect 16481 13 16515 47
rect 16553 13 16587 47
rect 16625 13 16659 47
rect 16697 13 16731 47
rect 16769 13 16803 47
rect 16867 13 16901 47
rect 16939 13 16973 47
rect 17011 13 17045 47
rect 17083 13 17117 47
rect 17155 13 17189 47
rect 17227 13 17261 47
rect 17371 13 17405 47
rect 17443 13 17477 47
rect 17515 13 17549 47
rect 17587 13 17621 47
rect 17677 13 17711 47
rect 17749 13 17783 47
rect 17821 13 17855 47
rect 17893 13 17927 47
rect 18037 13 18071 47
rect 18109 13 18143 47
rect 18181 13 18215 47
rect 18253 13 18287 47
rect 18343 13 18377 47
rect 18415 13 18449 47
rect 18487 13 18521 47
rect 18559 13 18593 47
rect 18703 13 18737 47
rect 18775 13 18809 47
rect 18847 13 18881 47
rect 18919 13 18953 47
rect 19009 13 19043 47
rect 19081 13 19115 47
rect 19153 13 19187 47
rect 19225 13 19259 47
<< metal1 >>
rect -31 1539 19345 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 343 1539
rect 377 1505 415 1539
rect 449 1505 513 1539
rect 547 1505 585 1539
rect 619 1505 657 1539
rect 691 1505 729 1539
rect 763 1505 801 1539
rect 835 1505 873 1539
rect 907 1505 1017 1539
rect 1051 1505 1089 1539
rect 1123 1505 1161 1539
rect 1195 1505 1233 1539
rect 1267 1505 1305 1539
rect 1339 1505 1377 1539
rect 1411 1505 1475 1539
rect 1509 1505 1547 1539
rect 1581 1505 1619 1539
rect 1653 1505 1691 1539
rect 1725 1505 1763 1539
rect 1797 1505 1835 1539
rect 1869 1505 1979 1539
rect 2013 1505 2051 1539
rect 2085 1505 2123 1539
rect 2157 1505 2195 1539
rect 2229 1505 2267 1539
rect 2301 1505 2339 1539
rect 2373 1505 2437 1539
rect 2471 1505 2509 1539
rect 2543 1505 2581 1539
rect 2615 1505 2653 1539
rect 2687 1505 2725 1539
rect 2759 1505 2797 1539
rect 2831 1505 2941 1539
rect 2975 1505 3013 1539
rect 3047 1505 3085 1539
rect 3119 1505 3157 1539
rect 3191 1505 3229 1539
rect 3263 1505 3301 1539
rect 3335 1505 3399 1539
rect 3433 1505 3471 1539
rect 3505 1505 3543 1539
rect 3577 1505 3615 1539
rect 3649 1505 3687 1539
rect 3721 1505 3759 1539
rect 3793 1505 3903 1539
rect 3937 1505 3975 1539
rect 4009 1505 4047 1539
rect 4081 1505 4119 1539
rect 4153 1505 4191 1539
rect 4225 1505 4263 1539
rect 4297 1505 4361 1539
rect 4395 1505 4433 1539
rect 4467 1505 4505 1539
rect 4539 1505 4577 1539
rect 4611 1505 4649 1539
rect 4683 1505 4721 1539
rect 4755 1505 4865 1539
rect 4899 1505 4937 1539
rect 4971 1505 5009 1539
rect 5043 1505 5081 1539
rect 5115 1505 5153 1539
rect 5187 1505 5225 1539
rect 5259 1505 5323 1539
rect 5357 1505 5395 1539
rect 5429 1505 5467 1539
rect 5501 1505 5539 1539
rect 5573 1505 5611 1539
rect 5645 1505 5683 1539
rect 5717 1505 5827 1539
rect 5861 1505 5899 1539
rect 5933 1505 5971 1539
rect 6005 1505 6043 1539
rect 6077 1505 6115 1539
rect 6149 1505 6187 1539
rect 6221 1505 6285 1539
rect 6319 1505 6357 1539
rect 6391 1505 6429 1539
rect 6463 1505 6501 1539
rect 6535 1505 6573 1539
rect 6607 1505 6645 1539
rect 6679 1505 6789 1539
rect 6823 1505 6861 1539
rect 6895 1505 6933 1539
rect 6967 1505 7005 1539
rect 7039 1505 7077 1539
rect 7111 1505 7149 1539
rect 7183 1505 7247 1539
rect 7281 1505 7319 1539
rect 7353 1505 7391 1539
rect 7425 1505 7463 1539
rect 7497 1505 7535 1539
rect 7569 1505 7607 1539
rect 7641 1505 7751 1539
rect 7785 1505 7823 1539
rect 7857 1505 7895 1539
rect 7929 1505 7967 1539
rect 8001 1505 8039 1539
rect 8073 1505 8111 1539
rect 8145 1505 8209 1539
rect 8243 1505 8281 1539
rect 8315 1505 8353 1539
rect 8387 1505 8425 1539
rect 8459 1505 8497 1539
rect 8531 1505 8569 1539
rect 8603 1505 8713 1539
rect 8747 1505 8785 1539
rect 8819 1505 8857 1539
rect 8891 1505 8929 1539
rect 8963 1505 9001 1539
rect 9035 1505 9073 1539
rect 9107 1505 9171 1539
rect 9205 1505 9243 1539
rect 9277 1505 9315 1539
rect 9349 1505 9387 1539
rect 9421 1505 9459 1539
rect 9493 1505 9531 1539
rect 9565 1505 9675 1539
rect 9709 1505 9747 1539
rect 9781 1505 9819 1539
rect 9853 1505 9891 1539
rect 9925 1505 9963 1539
rect 9997 1505 10035 1539
rect 10069 1505 10133 1539
rect 10167 1505 10205 1539
rect 10239 1505 10277 1539
rect 10311 1505 10349 1539
rect 10383 1505 10421 1539
rect 10455 1505 10493 1539
rect 10527 1505 10637 1539
rect 10671 1505 10709 1539
rect 10743 1505 10781 1539
rect 10815 1505 10853 1539
rect 10887 1505 10925 1539
rect 10959 1505 10997 1539
rect 11031 1505 11095 1539
rect 11129 1505 11167 1539
rect 11201 1505 11239 1539
rect 11273 1505 11311 1539
rect 11345 1505 11383 1539
rect 11417 1505 11455 1539
rect 11489 1505 11599 1539
rect 11633 1505 11671 1539
rect 11705 1505 11743 1539
rect 11777 1505 11815 1539
rect 11849 1505 11887 1539
rect 11921 1505 11959 1539
rect 11993 1505 12057 1539
rect 12091 1505 12129 1539
rect 12163 1505 12201 1539
rect 12235 1505 12273 1539
rect 12307 1505 12345 1539
rect 12379 1505 12417 1539
rect 12451 1505 12561 1539
rect 12595 1505 12633 1539
rect 12667 1505 12705 1539
rect 12739 1505 12777 1539
rect 12811 1505 12849 1539
rect 12883 1505 12921 1539
rect 12955 1505 13019 1539
rect 13053 1505 13091 1539
rect 13125 1505 13163 1539
rect 13197 1505 13235 1539
rect 13269 1505 13307 1539
rect 13341 1505 13379 1539
rect 13413 1505 13523 1539
rect 13557 1505 13595 1539
rect 13629 1505 13667 1539
rect 13701 1505 13739 1539
rect 13773 1505 13811 1539
rect 13845 1505 13883 1539
rect 13917 1505 13981 1539
rect 14015 1505 14053 1539
rect 14087 1505 14125 1539
rect 14159 1505 14197 1539
rect 14231 1505 14269 1539
rect 14303 1505 14341 1539
rect 14375 1505 14485 1539
rect 14519 1505 14557 1539
rect 14591 1505 14629 1539
rect 14663 1505 14701 1539
rect 14735 1505 14773 1539
rect 14807 1505 14845 1539
rect 14879 1505 14943 1539
rect 14977 1505 15015 1539
rect 15049 1505 15087 1539
rect 15121 1505 15159 1539
rect 15193 1505 15231 1539
rect 15265 1505 15303 1539
rect 15337 1505 15447 1539
rect 15481 1505 15519 1539
rect 15553 1505 15591 1539
rect 15625 1505 15663 1539
rect 15697 1505 15735 1539
rect 15769 1505 15807 1539
rect 15841 1505 15905 1539
rect 15939 1505 15977 1539
rect 16011 1505 16049 1539
rect 16083 1505 16121 1539
rect 16155 1505 16193 1539
rect 16227 1505 16265 1539
rect 16299 1505 16409 1539
rect 16443 1505 16481 1539
rect 16515 1505 16553 1539
rect 16587 1505 16625 1539
rect 16659 1505 16697 1539
rect 16731 1505 16769 1539
rect 16803 1505 16867 1539
rect 16901 1505 16939 1539
rect 16973 1505 17011 1539
rect 17045 1505 17083 1539
rect 17117 1505 17155 1539
rect 17189 1505 17227 1539
rect 17261 1505 17371 1539
rect 17405 1505 17443 1539
rect 17477 1505 17515 1539
rect 17549 1505 17587 1539
rect 17621 1505 17677 1539
rect 17711 1505 17749 1539
rect 17783 1505 17821 1539
rect 17855 1505 17893 1539
rect 17927 1505 18037 1539
rect 18071 1505 18109 1539
rect 18143 1505 18181 1539
rect 18215 1505 18253 1539
rect 18287 1505 18343 1539
rect 18377 1505 18415 1539
rect 18449 1505 18487 1539
rect 18521 1505 18559 1539
rect 18593 1505 18703 1539
rect 18737 1505 18775 1539
rect 18809 1505 18847 1539
rect 18881 1505 18919 1539
rect 18953 1505 19009 1539
rect 19043 1505 19081 1539
rect 19115 1505 19153 1539
rect 19187 1505 19225 1539
rect 19259 1505 19345 1539
rect -31 1492 19345 1505
rect 17715 1105 17761 1111
rect 18115 1105 18161 1111
rect 18379 1105 18425 1111
rect 18783 1105 18829 1111
rect 17709 1071 17721 1105
rect 17755 1071 18121 1105
rect 18155 1071 18167 1105
rect 18373 1071 18385 1105
rect 18419 1071 18789 1105
rect 18823 1071 18835 1105
rect 17715 1065 17761 1071
rect 18115 1065 18161 1071
rect 18379 1065 18425 1071
rect 18783 1065 18829 1071
rect 1382 979 1428 985
rect 3307 979 3353 985
rect 7154 979 7200 985
rect 9079 979 9125 985
rect 12926 979 12972 985
rect 14851 979 14897 985
rect 17441 979 17487 985
rect 18181 979 18227 985
rect 1376 945 1388 979
rect 1422 945 3313 979
rect 3347 945 7160 979
rect 7194 945 9085 979
rect 9119 945 12932 979
rect 12966 945 14857 979
rect 14891 945 14903 979
rect 17435 945 17447 979
rect 17481 945 18187 979
rect 18221 945 18233 979
rect 1382 939 1428 945
rect 3307 939 3353 945
rect 7154 939 7200 945
rect 9079 939 9125 945
rect 12926 939 12972 945
rect 14851 939 14897 945
rect 17441 939 17487 945
rect 18181 939 18227 945
rect 199 905 245 911
rect 5971 905 6017 911
rect 11743 905 11789 911
rect 17663 905 17709 911
rect 18995 905 19041 911
rect 169 871 205 905
rect 239 871 5977 905
rect 6011 871 11749 905
rect 11783 871 11819 905
rect 11971 871 17669 905
rect 17703 871 19001 905
rect 19035 871 19047 905
rect 199 865 245 871
rect 5971 865 6017 871
rect 11743 865 11789 871
rect 1604 831 1650 837
rect 2567 831 2613 837
rect 3677 831 3723 837
rect 5453 831 5499 837
rect 7376 831 7422 837
rect 8339 831 8385 837
rect 9449 831 9495 837
rect 11225 831 11271 837
rect 11373 831 11419 837
rect 11971 831 12005 871
rect 17663 865 17709 871
rect 18995 865 19041 871
rect 13148 831 13194 837
rect 14111 831 14157 837
rect 15221 831 15267 837
rect 16997 831 17043 837
rect 17145 831 17191 837
rect 17441 831 17487 837
rect 19143 831 19189 837
rect 1598 797 1610 831
rect 1644 797 2573 831
rect 2607 797 3683 831
rect 3717 797 5459 831
rect 5493 797 5505 831
rect 7370 797 7382 831
rect 7416 797 8345 831
rect 8379 797 9455 831
rect 9489 797 11231 831
rect 11265 797 11277 831
rect 11367 797 11379 831
rect 11413 797 12005 831
rect 13142 797 13154 831
rect 13188 797 14117 831
rect 14151 797 15227 831
rect 15261 797 17003 831
rect 17037 797 17049 831
rect 17139 797 17151 831
rect 17185 797 17447 831
rect 17481 797 17493 831
rect 19137 797 19149 831
rect 19183 797 19219 831
rect 1604 791 1650 797
rect 2567 791 2613 797
rect 3677 791 3723 797
rect 5453 791 5499 797
rect 7376 791 7422 797
rect 8339 791 8385 797
rect 9449 791 9495 797
rect 11225 791 11271 797
rect 11373 791 11419 797
rect 13148 791 13194 797
rect 14111 791 14157 797
rect 15221 791 15267 797
rect 16997 791 17043 797
rect 17145 791 17191 797
rect 17441 791 17487 797
rect 19143 791 19189 797
rect 643 757 689 763
rect 1753 757 1799 763
rect 4047 757 4093 763
rect 4639 757 4685 763
rect 5009 757 5055 763
rect 6415 757 6461 763
rect 7525 757 7571 763
rect 9819 757 9865 763
rect 10411 757 10457 763
rect 10781 757 10827 763
rect 12187 757 12233 763
rect 13297 757 13343 763
rect 15591 757 15637 763
rect 16183 757 16229 763
rect 16553 757 16599 763
rect 637 723 649 757
rect 683 723 1759 757
rect 1793 723 4053 757
rect 4087 723 4099 757
rect 4633 723 4645 757
rect 4679 723 5015 757
rect 5049 723 5061 757
rect 6409 723 6421 757
rect 6455 723 7531 757
rect 7565 723 9825 757
rect 9859 723 9871 757
rect 10405 723 10417 757
rect 10451 723 10787 757
rect 10821 723 10833 757
rect 12181 723 12193 757
rect 12227 723 13303 757
rect 13337 723 15597 757
rect 15631 723 15643 757
rect 16177 723 16189 757
rect 16223 723 16559 757
rect 16593 723 16605 757
rect 643 717 689 723
rect 1753 717 1799 723
rect 4047 717 4093 723
rect 4639 717 4685 723
rect 5009 717 5055 723
rect 6415 717 6461 723
rect 7525 717 7571 723
rect 9819 717 9865 723
rect 10411 717 10457 723
rect 10781 717 10827 723
rect 12187 717 12233 723
rect 13297 717 13343 723
rect 15591 717 15637 723
rect 16183 717 16229 723
rect 16553 717 16599 723
rect 4491 683 4537 689
rect 5601 683 5647 689
rect 18477 683 18523 689
rect 4485 649 4497 683
rect 4531 649 5607 683
rect 5641 649 18483 683
rect 18517 649 18529 683
rect 4491 643 4537 649
rect 5601 643 5647 649
rect 18477 643 18523 649
rect 791 610 837 616
rect 1161 610 1207 616
rect 2123 610 2169 616
rect 785 576 797 610
rect 831 576 1167 610
rect 1201 576 2129 610
rect 2163 576 2175 610
rect 2715 609 2761 615
rect 3085 609 3131 615
rect 6563 610 6609 616
rect 6933 610 6979 616
rect 7895 610 7941 616
rect 791 570 837 576
rect 1161 570 1207 576
rect 2123 570 2169 576
rect 2709 575 2721 609
rect 2755 575 3091 609
rect 3125 575 3137 609
rect 6557 576 6569 610
rect 6603 576 6939 610
rect 6973 576 7901 610
rect 7935 576 7947 610
rect 8487 609 8533 615
rect 8857 609 8903 615
rect 10263 609 10309 615
rect 11373 609 11419 615
rect 12335 610 12381 616
rect 12705 610 12751 616
rect 13667 610 13713 616
rect 2715 569 2761 575
rect 3085 569 3131 575
rect 6563 570 6609 576
rect 6933 570 6979 576
rect 7895 570 7941 576
rect 8481 575 8493 609
rect 8527 575 8863 609
rect 8897 575 8909 609
rect 10257 575 10269 609
rect 10303 575 11379 609
rect 11413 575 11425 609
rect 12329 576 12341 610
rect 12375 576 12711 610
rect 12745 576 13673 610
rect 13707 576 13719 610
rect 14259 609 14305 615
rect 14629 609 14675 615
rect 16035 609 16081 615
rect 17145 609 17191 615
rect 8487 569 8533 575
rect 8857 569 8903 575
rect 10263 569 10309 575
rect 11373 569 11419 575
rect 12335 570 12381 576
rect 12705 570 12751 576
rect 13667 570 13713 576
rect 14253 575 14265 609
rect 14299 575 14635 609
rect 14669 575 14681 609
rect 16029 575 16041 609
rect 16075 575 17151 609
rect 17185 575 17197 609
rect 14259 569 14305 575
rect 14629 569 14675 575
rect 16035 569 16081 575
rect 17145 569 17191 575
rect 421 535 467 541
rect 3529 535 3575 541
rect 4269 535 4315 541
rect 6193 535 6239 541
rect 9301 535 9347 541
rect 10041 535 10087 541
rect 11965 535 12011 541
rect 15073 535 15119 541
rect 15813 535 15859 541
rect 415 501 427 535
rect 461 501 3535 535
rect 3569 501 4275 535
rect 4309 501 6199 535
rect 6233 501 9307 535
rect 9341 501 10047 535
rect 10081 501 11971 535
rect 12005 501 15079 535
rect 15113 501 15819 535
rect 15853 501 15865 535
rect 421 495 467 501
rect 3529 495 3575 501
rect 4269 495 4315 501
rect 6193 495 6239 501
rect 9301 495 9347 501
rect 10041 495 10087 501
rect 11965 495 12011 501
rect 15073 495 15119 501
rect 15813 495 15859 501
rect 2345 462 2391 468
rect 2339 428 2351 462
rect 2385 461 2421 462
rect 5231 461 5277 467
rect 8117 462 8163 468
rect 8111 461 8123 462
rect 2385 428 5237 461
rect 2344 427 5237 428
rect 5271 428 8123 461
rect 8157 461 8193 462
rect 11003 461 11049 467
rect 13889 462 13935 468
rect 13883 461 13895 462
rect 8157 428 11009 461
rect 5271 427 11009 428
rect 11043 428 13895 461
rect 13929 461 13965 462
rect 16775 461 16821 467
rect 18477 461 18523 467
rect 18773 461 18819 467
rect 13929 428 16781 461
rect 11043 427 16781 428
rect 16815 427 16827 461
rect 18471 427 18483 461
rect 18517 427 18779 461
rect 18813 427 18825 461
rect 2345 422 2391 427
rect 5231 421 5277 427
rect 8117 422 8163 427
rect 11003 421 11049 427
rect 13889 422 13935 427
rect 16775 421 16821 427
rect 18477 421 18523 427
rect 18773 421 18819 427
rect 17723 281 17769 287
rect 18389 281 18435 287
rect 19055 281 19101 287
rect 17717 247 17729 281
rect 17763 247 18395 281
rect 18429 247 19061 281
rect 19095 247 19107 281
rect 17723 241 17769 247
rect 18389 241 18435 247
rect 19055 241 19101 247
rect -31 47 19345 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 343 47
rect 377 13 415 47
rect 449 13 513 47
rect 547 13 585 47
rect 619 13 657 47
rect 691 13 729 47
rect 763 13 801 47
rect 835 13 873 47
rect 907 13 1017 47
rect 1051 13 1089 47
rect 1123 13 1161 47
rect 1195 13 1233 47
rect 1267 13 1305 47
rect 1339 13 1377 47
rect 1411 13 1475 47
rect 1509 13 1547 47
rect 1581 13 1619 47
rect 1653 13 1691 47
rect 1725 13 1763 47
rect 1797 13 1835 47
rect 1869 13 1979 47
rect 2013 13 2051 47
rect 2085 13 2123 47
rect 2157 13 2195 47
rect 2229 13 2267 47
rect 2301 13 2339 47
rect 2373 13 2437 47
rect 2471 13 2509 47
rect 2543 13 2581 47
rect 2615 13 2653 47
rect 2687 13 2725 47
rect 2759 13 2797 47
rect 2831 13 2941 47
rect 2975 13 3013 47
rect 3047 13 3085 47
rect 3119 13 3157 47
rect 3191 13 3229 47
rect 3263 13 3301 47
rect 3335 13 3399 47
rect 3433 13 3471 47
rect 3505 13 3543 47
rect 3577 13 3615 47
rect 3649 13 3687 47
rect 3721 13 3759 47
rect 3793 13 3903 47
rect 3937 13 3975 47
rect 4009 13 4047 47
rect 4081 13 4119 47
rect 4153 13 4191 47
rect 4225 13 4263 47
rect 4297 13 4361 47
rect 4395 13 4433 47
rect 4467 13 4505 47
rect 4539 13 4577 47
rect 4611 13 4649 47
rect 4683 13 4721 47
rect 4755 13 4865 47
rect 4899 13 4937 47
rect 4971 13 5009 47
rect 5043 13 5081 47
rect 5115 13 5153 47
rect 5187 13 5225 47
rect 5259 13 5323 47
rect 5357 13 5395 47
rect 5429 13 5467 47
rect 5501 13 5539 47
rect 5573 13 5611 47
rect 5645 13 5683 47
rect 5717 13 5827 47
rect 5861 13 5899 47
rect 5933 13 5971 47
rect 6005 13 6043 47
rect 6077 13 6115 47
rect 6149 13 6187 47
rect 6221 13 6285 47
rect 6319 13 6357 47
rect 6391 13 6429 47
rect 6463 13 6501 47
rect 6535 13 6573 47
rect 6607 13 6645 47
rect 6679 13 6789 47
rect 6823 13 6861 47
rect 6895 13 6933 47
rect 6967 13 7005 47
rect 7039 13 7077 47
rect 7111 13 7149 47
rect 7183 13 7247 47
rect 7281 13 7319 47
rect 7353 13 7391 47
rect 7425 13 7463 47
rect 7497 13 7535 47
rect 7569 13 7607 47
rect 7641 13 7751 47
rect 7785 13 7823 47
rect 7857 13 7895 47
rect 7929 13 7967 47
rect 8001 13 8039 47
rect 8073 13 8111 47
rect 8145 13 8209 47
rect 8243 13 8281 47
rect 8315 13 8353 47
rect 8387 13 8425 47
rect 8459 13 8497 47
rect 8531 13 8569 47
rect 8603 13 8713 47
rect 8747 13 8785 47
rect 8819 13 8857 47
rect 8891 13 8929 47
rect 8963 13 9001 47
rect 9035 13 9073 47
rect 9107 13 9171 47
rect 9205 13 9243 47
rect 9277 13 9315 47
rect 9349 13 9387 47
rect 9421 13 9459 47
rect 9493 13 9531 47
rect 9565 13 9675 47
rect 9709 13 9747 47
rect 9781 13 9819 47
rect 9853 13 9891 47
rect 9925 13 9963 47
rect 9997 13 10035 47
rect 10069 13 10133 47
rect 10167 13 10205 47
rect 10239 13 10277 47
rect 10311 13 10349 47
rect 10383 13 10421 47
rect 10455 13 10493 47
rect 10527 13 10637 47
rect 10671 13 10709 47
rect 10743 13 10781 47
rect 10815 13 10853 47
rect 10887 13 10925 47
rect 10959 13 10997 47
rect 11031 13 11095 47
rect 11129 13 11167 47
rect 11201 13 11239 47
rect 11273 13 11311 47
rect 11345 13 11383 47
rect 11417 13 11455 47
rect 11489 13 11599 47
rect 11633 13 11671 47
rect 11705 13 11743 47
rect 11777 13 11815 47
rect 11849 13 11887 47
rect 11921 13 11959 47
rect 11993 13 12057 47
rect 12091 13 12129 47
rect 12163 13 12201 47
rect 12235 13 12273 47
rect 12307 13 12345 47
rect 12379 13 12417 47
rect 12451 13 12561 47
rect 12595 13 12633 47
rect 12667 13 12705 47
rect 12739 13 12777 47
rect 12811 13 12849 47
rect 12883 13 12921 47
rect 12955 13 13019 47
rect 13053 13 13091 47
rect 13125 13 13163 47
rect 13197 13 13235 47
rect 13269 13 13307 47
rect 13341 13 13379 47
rect 13413 13 13523 47
rect 13557 13 13595 47
rect 13629 13 13667 47
rect 13701 13 13739 47
rect 13773 13 13811 47
rect 13845 13 13883 47
rect 13917 13 13981 47
rect 14015 13 14053 47
rect 14087 13 14125 47
rect 14159 13 14197 47
rect 14231 13 14269 47
rect 14303 13 14341 47
rect 14375 13 14485 47
rect 14519 13 14557 47
rect 14591 13 14629 47
rect 14663 13 14701 47
rect 14735 13 14773 47
rect 14807 13 14845 47
rect 14879 13 14943 47
rect 14977 13 15015 47
rect 15049 13 15087 47
rect 15121 13 15159 47
rect 15193 13 15231 47
rect 15265 13 15303 47
rect 15337 13 15447 47
rect 15481 13 15519 47
rect 15553 13 15591 47
rect 15625 13 15663 47
rect 15697 13 15735 47
rect 15769 13 15807 47
rect 15841 13 15905 47
rect 15939 13 15977 47
rect 16011 13 16049 47
rect 16083 13 16121 47
rect 16155 13 16193 47
rect 16227 13 16265 47
rect 16299 13 16409 47
rect 16443 13 16481 47
rect 16515 13 16553 47
rect 16587 13 16625 47
rect 16659 13 16697 47
rect 16731 13 16769 47
rect 16803 13 16867 47
rect 16901 13 16939 47
rect 16973 13 17011 47
rect 17045 13 17083 47
rect 17117 13 17155 47
rect 17189 13 17227 47
rect 17261 13 17371 47
rect 17405 13 17443 47
rect 17477 13 17515 47
rect 17549 13 17587 47
rect 17621 13 17677 47
rect 17711 13 17749 47
rect 17783 13 17821 47
rect 17855 13 17893 47
rect 17927 13 18037 47
rect 18071 13 18109 47
rect 18143 13 18181 47
rect 18215 13 18253 47
rect 18287 13 18343 47
rect 18377 13 18415 47
rect 18449 13 18487 47
rect 18521 13 18559 47
rect 18593 13 18703 47
rect 18737 13 18775 47
rect 18809 13 18847 47
rect 18881 13 18919 47
rect 18953 13 19009 47
rect 19043 13 19081 47
rect 19115 13 19153 47
rect 19187 13 19225 47
rect 19259 13 19345 47
rect -31 0 19345 13
<< labels >>
rlabel metal1 19149 797 19183 831 1 QN
port 1 n
rlabel metal1 205 871 239 905 1 D
port 2 n
rlabel metal1 1388 945 1422 979 1 CLK
port 3 n
rlabel metal1 2351 427 2385 461 1 SN
port 4 n
rlabel metal1 427 501 461 535 1 RN
port 5 n
rlabel metal1 55 1505 89 1539 1 VDD
port 6 n
rlabel metal1 55 13 89 47 1 VSS
port 7 n
<< end >>
