* NGSPICE file created from 12T_ms_rhbd.ext - technology: sky130A

