magic
tech sky130A
magscale 1 2
timestamp 1645638419
<< nwell >>
rect -84 759 84 1353
<< psubdiff >>
rect -31 475 31 570
rect -31 441 -17 475
rect 17 441 31 475
rect -31 403 31 441
rect -31 369 -17 403
rect 17 369 31 403
rect -31 331 31 369
rect -31 297 -17 331
rect 17 297 31 331
rect -31 259 31 297
rect -31 225 -17 259
rect 17 225 31 259
rect -31 187 31 225
rect -31 153 -17 187
rect 17 153 31 187
rect -31 115 31 153
rect -31 81 -17 115
rect 17 81 31 115
rect -31 13 31 81
<< nsubdiff >>
rect -31 1249 31 1317
rect -31 1215 -17 1249
rect 17 1215 31 1249
rect -31 1177 31 1215
rect -31 1143 -17 1177
rect 17 1143 31 1177
rect -31 1105 31 1143
rect -31 1071 -17 1105
rect 17 1071 31 1105
rect -31 1033 31 1071
rect -31 999 -17 1033
rect 17 999 31 1033
rect -31 961 31 999
rect -31 927 -17 961
rect 17 927 31 961
rect -31 889 31 927
rect -31 855 -17 889
rect 17 855 31 889
rect -31 795 31 855
<< psubdiffcont >>
rect -17 441 17 475
rect -17 369 17 403
rect -17 297 17 331
rect -17 225 17 259
rect -17 153 17 187
rect -17 81 17 115
<< nsubdiffcont >>
rect -17 1215 17 1249
rect -17 1143 17 1177
rect -17 1071 17 1105
rect -17 999 17 1033
rect -17 927 17 961
rect -17 855 17 889
<< locali >>
rect -31 1249 31 1332
rect -31 1215 -17 1249
rect 17 1215 31 1249
rect -31 1177 31 1215
rect -31 1143 -17 1177
rect 17 1143 31 1177
rect -31 1105 31 1143
rect -31 1071 -17 1105
rect 17 1071 31 1105
rect -31 1033 31 1071
rect -31 999 -17 1033
rect 17 999 31 1033
rect -31 961 31 999
rect -31 927 -17 961
rect 17 927 31 961
rect -31 889 31 927
rect -31 855 -17 889
rect 17 855 31 889
rect -31 795 31 855
rect -31 475 31 570
rect -31 441 -17 475
rect 17 441 31 475
rect -31 403 31 441
rect -31 369 -17 403
rect 17 369 31 403
rect -31 331 31 369
rect -31 297 -17 331
rect 17 297 31 331
rect -31 259 31 297
rect -31 225 -17 259
rect 17 225 31 259
rect -31 187 31 225
rect -31 153 -17 187
rect 17 153 31 187
rect -31 115 31 153
rect -31 81 -17 115
rect 17 81 31 115
rect -31 0 31 81
<< viali >>
rect -17 1215 17 1249
rect -17 1143 17 1177
rect -17 1071 17 1105
rect -17 999 17 1033
rect -17 927 17 961
rect -17 855 17 889
rect -17 441 17 475
rect -17 369 17 403
rect -17 297 17 331
rect -17 225 17 259
rect -17 153 17 187
rect -17 81 17 115
<< metal1 >>
rect -31 1249 31 1332
rect -31 1215 -17 1249
rect 17 1215 31 1249
rect -31 1177 31 1215
rect -31 1143 -17 1177
rect 17 1143 31 1177
rect -31 1105 31 1143
rect -31 1071 -17 1105
rect 17 1071 31 1105
rect -31 1033 31 1071
rect -31 999 -17 1033
rect 17 999 31 1033
rect -31 961 31 999
rect -31 927 -17 961
rect 17 927 31 961
rect -31 889 31 927
rect -31 855 -17 889
rect 17 855 31 889
rect -31 795 31 855
rect -31 475 31 570
rect -31 441 -17 475
rect 17 441 31 475
rect -31 403 31 441
rect -31 369 -17 403
rect 17 369 31 403
rect -31 331 31 369
rect -31 297 -17 331
rect 17 297 31 331
rect -31 259 31 297
rect -31 225 -17 259
rect 17 225 31 259
rect -31 187 31 225
rect -31 153 -17 187
rect 17 153 31 187
rect -31 115 31 153
rect -31 81 -17 115
rect 17 81 31 115
rect -31 0 31 81
<< end >>
