* NGSPICE file created from DFFSNRNX1.ext - technology: sky130A

.subckt nmos_bottom a_86_101# a_56_85# a_0_0# VSUBS
X0 a_86_101# a_56_85# a_0_0# VSUBS sky130_fd_pr__nfet_01v8 ad=1.772p pd=1.56u as=1.152p ps=8.19u w=3u l=0.15u
.ends

.subckt nmos_top_trim1 a_56_92# a_86_108# a_0_0# VSUBS
X0 a_86_108# a_56_92# a_0_0# VSUBS sky130_fd_pr__nfet_01v8 ad=1.772p pd=1.56u as=1.15725p ps=8.12u w=3u l=0.15u
.ends

.subckt nmos_side_left a_87_107# a_57_91# a_0_0# VSUBS
X0 a_87_107# a_57_91# a_0_0# VSUBS sky130_fd_pr__nfet_01v8 ad=1.6345p pd=1.49u as=1.17945p ps=8.17u w=3u l=0.15u
.ends

.subckt pmos2 a_144_n460# a_262_n399# a_88_n399# w_52_n435# a_174_n399#
X0 a_174_n399# a_144_n460# a_88_n399# w_52_n435# sky130_fd_pr__pfet_01v8 ad=5.8p pd=4.58u as=5.6p ps=4.56u w=2u l=0.15u
X1 a_262_n399# a_144_n460# a_174_n399# w_52_n435# sky130_fd_pr__pfet_01v8 ad=5.4p pd=4.54u as=0p ps=0u w=2u l=0.15u
.ends

.subckt nand3x1_pcell VSS VDD a_289_1105# a_147_405# a_447_405# li_649_477# a_31_510#
Xnmos_bottom_0 VSS a_147_405# nmos_bottom_0/a_0_0# VSS nmos_bottom
Xnmos_top_trim1_0 li_649_477# a_289_1105# li_393_210# VSS nmos_top_trim1
Xnmos_side_left_0 li_393_210# a_447_405# nmos_bottom_0/a_0_0# VSS nmos_side_left
Xpmos2_0 a_147_405# VDD VDD VDD a_289_1105# pmos2
Xpmos2_1 a_447_405# VDD VDD VDD a_289_1105# pmos2
Xpmos2_2 li_649_477# VDD VDD VDD a_289_1105# pmos2
.ends

.subckt DFFSNRNX1 RN CLK SN Q QN D VDD VSS
Xnand3x1_pcell_0 VSS VDD m1_831_576# D m1_461_723# RN VSS nand3x1_pcell
Xnand3x1_pcell_1 VSS VDD m1_461_723# m1_1203_797# m1_831_576# CLK nand3x1_pcell_1/a_31_510#
+ nand3x1_pcell
Xnand3x1_pcell_2 VSS VDD m1_2757_575# m1_831_576# m1_1203_797# SN VSS nand3x1_pcell
Xnand3x1_pcell_3 VSS VDD m1_1203_797# RN CLK m1_2757_575# VSS nand3x1_pcell
Xnand3x1_pcell_4 VSS VDD QN RN m1_461_723# Q nand3x1_pcell_4/a_31_510# nand3x1_pcell
Xnand3x1_pcell_5 VSS VDD Q m1_1203_797# QN SN nand3x1_pcell_5/a_31_510# nand3x1_pcell
.ends

