magic
tech sky130A
magscale 1 2
timestamp 1647814117
<< nwell >>
rect 84 1554 582 1575
rect 31 1492 582 1554
rect 84 832 582 1492
rect 750 832 1248 1575
rect 1416 832 1914 1575
<< pdiffc >>
rect 141 1377 175 1411
rect 229 1377 263 1411
rect 317 1377 351 1411
rect 405 1377 439 1411
rect 493 1377 527 1411
rect 805 1377 839 1411
rect 981 1377 1015 1411
rect 1157 1377 1191 1411
rect 1473 1377 1507 1411
rect 1649 1377 1683 1411
rect 1825 1377 1859 1411
rect 141 1105 175 1139
rect 229 1105 263 1139
rect 493 1105 527 1139
rect 893 1105 927 1139
rect 1561 1105 1595 1139
rect 1737 1105 1771 1139
<< psubdiff >>
rect 31 510 635 572
rect 697 510 1301 572
rect 1363 510 1967 572
rect 31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 361 47
rect 395 13 433 47
rect 467 13 505 47
rect 539 13 577 47
rect 611 13 635 47
rect 697 13 721 47
rect 755 13 793 47
rect 827 13 865 47
rect 899 13 937 47
rect 971 13 1027 47
rect 1061 13 1099 47
rect 1133 13 1171 47
rect 1205 13 1243 47
rect 1277 13 1301 47
rect 1363 13 1387 47
rect 1421 13 1459 47
rect 1493 13 1531 47
rect 1565 13 1603 47
rect 1637 13 1693 47
rect 1727 13 1765 47
rect 1799 13 1837 47
rect 1871 13 1909 47
rect 1943 13 1967 47
<< nsubdiff >>
rect 31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 361 1539
rect 395 1505 433 1539
rect 467 1505 505 1539
rect 539 1505 577 1539
rect 611 1505 635 1539
rect 697 1505 721 1539
rect 755 1505 793 1539
rect 827 1505 865 1539
rect 899 1505 937 1539
rect 971 1505 1027 1539
rect 1061 1505 1099 1539
rect 1133 1505 1171 1539
rect 1205 1505 1243 1539
rect 1277 1505 1301 1539
rect 1363 1505 1387 1539
rect 1421 1505 1459 1539
rect 1493 1505 1531 1539
rect 1565 1505 1603 1539
rect 1637 1505 1693 1539
rect 1727 1505 1765 1539
rect 1799 1505 1837 1539
rect 1871 1505 1909 1539
rect 1943 1505 1967 1539
rect 31 868 635 930
rect 697 868 1301 930
rect 1363 868 1967 930
<< psubdiffcont >>
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 361 13 395 47
rect 433 13 467 47
rect 505 13 539 47
rect 577 13 611 47
rect 721 13 755 47
rect 793 13 827 47
rect 865 13 899 47
rect 937 13 971 47
rect 1027 13 1061 47
rect 1099 13 1133 47
rect 1171 13 1205 47
rect 1243 13 1277 47
rect 1387 13 1421 47
rect 1459 13 1493 47
rect 1531 13 1565 47
rect 1603 13 1637 47
rect 1693 13 1727 47
rect 1765 13 1799 47
rect 1837 13 1871 47
rect 1909 13 1943 47
<< nsubdiffcont >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 361 1505 395 1539
rect 433 1505 467 1539
rect 505 1505 539 1539
rect 577 1505 611 1539
rect 721 1505 755 1539
rect 793 1505 827 1539
rect 865 1505 899 1539
rect 937 1505 971 1539
rect 1027 1505 1061 1539
rect 1099 1505 1133 1539
rect 1171 1505 1205 1539
rect 1243 1505 1277 1539
rect 1387 1505 1421 1539
rect 1459 1505 1493 1539
rect 1531 1505 1565 1539
rect 1603 1505 1637 1539
rect 1693 1505 1727 1539
rect 1765 1505 1799 1539
rect 1837 1505 1871 1539
rect 1909 1505 1943 1539
<< poly >>
rect 175 990 187 1020
rect 1145 990 1157 1020
rect 1507 990 1519 1020
rect 168 403 198 441
rect 362 410 392 411
rect 834 403 864 441
rect 1134 410 1164 441
rect 1500 403 1530 441
rect 1694 410 1724 411
<< locali >>
rect 31 1539 635 1554
rect 31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 361 1539
rect 395 1505 433 1539
rect 467 1505 505 1539
rect 539 1505 577 1539
rect 611 1505 635 1539
rect 31 1492 635 1505
rect 697 1539 1301 1554
rect 697 1505 721 1539
rect 755 1505 793 1539
rect 827 1505 865 1539
rect 899 1505 937 1539
rect 971 1505 1027 1539
rect 1061 1505 1099 1539
rect 1133 1505 1171 1539
rect 1205 1505 1243 1539
rect 1277 1505 1301 1539
rect 697 1492 1301 1505
rect 1363 1539 1967 1554
rect 1363 1505 1387 1539
rect 1421 1505 1459 1539
rect 1493 1505 1531 1539
rect 1565 1505 1603 1539
rect 1637 1505 1693 1539
rect 1727 1505 1765 1539
rect 1799 1505 1837 1539
rect 1871 1505 1909 1539
rect 1943 1505 1967 1539
rect 1363 1492 1967 1505
rect 141 1411 175 1492
rect 141 1359 175 1377
rect 229 1411 265 1445
rect 317 1411 351 1492
rect 229 1359 263 1377
rect 317 1359 351 1377
rect 405 1411 439 1445
rect 405 1359 439 1377
rect 493 1411 527 1492
rect 493 1359 527 1377
rect 805 1411 1191 1445
rect 805 1359 839 1377
rect 981 1359 1015 1377
rect 1157 1359 1191 1377
rect 1473 1411 1859 1445
rect 1473 1359 1507 1377
rect 1649 1359 1683 1377
rect 1825 1359 1859 1377
rect 141 1139 175 1157
rect 141 1071 175 1105
rect 229 1139 263 1157
rect 405 1121 439 1157
rect 493 1139 527 1157
rect 805 1121 839 1173
rect 893 1139 927 1157
rect 229 1071 405 1105
rect 493 1071 527 1105
rect 1069 1121 1103 1157
rect 1157 1121 1191 1157
rect 1473 1121 1507 1157
rect 1561 1139 1595 1157
rect 1737 1139 1771 1173
rect 805 1069 839 1100
rect 893 1071 1103 1105
rect 1473 1071 1507 1084
rect 1561 1071 1867 1105
rect 131 461 165 988
rect 353 954 361 988
rect 353 847 387 954
rect 871 847 905 954
rect 1167 831 1201 988
rect 1463 847 1497 954
rect 353 469 387 501
rect 871 477 905 485
rect 353 461 357 469
rect 1167 461 1201 501
rect 1463 477 1497 486
rect 1685 461 1719 1020
rect 1833 374 1867 1071
rect 1745 340 1867 374
rect 1745 297 1779 340
rect 219 62 253 187
rect 885 62 919 187
rect 1551 62 1585 187
rect 31 47 635 62
rect 31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 361 47
rect 395 13 433 47
rect 467 13 505 47
rect 539 13 577 47
rect 611 13 635 47
rect 31 0 635 13
rect 697 47 1079 62
rect 1113 47 1301 62
rect 697 13 721 47
rect 755 13 793 47
rect 827 13 865 47
rect 899 13 937 47
rect 971 13 1027 47
rect 1061 13 1099 47
rect 1133 13 1171 47
rect 1205 13 1243 47
rect 1277 13 1301 47
rect 697 0 1301 13
rect 1363 47 1967 62
rect 1363 13 1387 47
rect 1421 13 1459 47
rect 1493 13 1531 47
rect 1565 13 1603 47
rect 1637 13 1693 47
rect 1727 13 1765 47
rect 1799 13 1837 47
rect 1871 13 1909 47
rect 1943 13 1967 47
rect 1363 0 1967 13
<< viali >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 361 1505 395 1539
rect 433 1505 467 1539
rect 505 1505 539 1539
rect 577 1505 611 1539
rect 721 1505 755 1539
rect 793 1505 827 1539
rect 865 1505 899 1539
rect 937 1505 971 1539
rect 1027 1505 1061 1539
rect 1099 1505 1133 1539
rect 1171 1505 1205 1539
rect 1243 1505 1277 1539
rect 1387 1505 1421 1539
rect 1459 1505 1493 1539
rect 1531 1505 1565 1539
rect 1603 1505 1637 1539
rect 1693 1505 1727 1539
rect 1765 1505 1799 1539
rect 1837 1505 1871 1539
rect 1909 1505 1943 1539
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 361 13 395 47
rect 433 13 467 47
rect 505 13 539 47
rect 577 13 611 47
rect 721 13 755 47
rect 793 13 827 47
rect 865 13 899 47
rect 937 13 971 47
rect 1027 13 1061 47
rect 1099 13 1133 47
rect 1171 13 1205 47
rect 1243 13 1277 47
rect 1387 13 1421 47
rect 1459 13 1493 47
rect 1531 13 1565 47
rect 1603 13 1637 47
rect 1693 13 1727 47
rect 1765 13 1799 47
rect 1837 13 1871 47
rect 1909 13 1943 47
<< metal1 >>
rect 31 1539 635 1554
rect 31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 361 1539
rect 395 1505 433 1539
rect 467 1505 505 1539
rect 539 1505 577 1539
rect 611 1505 635 1539
rect 31 1492 635 1505
rect 697 1539 1301 1554
rect 697 1505 721 1539
rect 755 1505 793 1539
rect 827 1505 865 1539
rect 899 1505 937 1539
rect 971 1505 1027 1539
rect 1061 1505 1099 1539
rect 1133 1505 1171 1539
rect 1205 1505 1243 1539
rect 1277 1505 1301 1539
rect 697 1492 1301 1505
rect 1363 1539 1967 1554
rect 1363 1505 1387 1539
rect 1421 1505 1459 1539
rect 1493 1505 1531 1539
rect 1565 1505 1603 1539
rect 1637 1505 1693 1539
rect 1727 1505 1765 1539
rect 1799 1505 1837 1539
rect 1871 1505 1909 1539
rect 1943 1505 1967 1539
rect 1363 1492 1967 1505
rect 475 1071 799 1105
rect 1135 1071 1466 1105
rect 166 871 1653 905
rect 389 797 839 831
rect 1201 797 1453 831
rect 387 501 844 535
rect 1201 501 1453 535
rect 449 247 1744 281
rect 31 47 635 62
rect 31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 361 47
rect 395 13 433 47
rect 467 13 505 47
rect 539 13 577 47
rect 611 13 635 47
rect 31 0 635 13
rect 697 47 1301 62
rect 697 13 721 47
rect 755 13 793 47
rect 827 13 865 47
rect 899 13 937 47
rect 971 13 1027 47
rect 1061 13 1099 47
rect 1133 13 1171 47
rect 1205 13 1243 47
rect 1277 13 1301 47
rect 697 0 1301 13
rect 1363 47 1967 62
rect 1363 13 1387 47
rect 1421 13 1459 47
rect 1493 13 1531 47
rect 1565 13 1603 47
rect 1637 13 1693 47
rect 1727 13 1765 47
rect 1799 13 1837 47
rect 1871 13 1909 47
rect 1943 13 1967 47
rect 1363 0 1967 13
use li1_M1_contact  li1_M1_contact_15
timestamp 1646004885
transform -1 0 148 0 1 888
box -53 -33 29 33
use diff_ring_side  diff_ring_side_1
timestamp 1646086970
transform 1 0 0 0 1 0
box -84 0 84 1575
use poly_li1_contact  poly_li1_contact_0
timestamp 1645652543
transform 0 1 148 -1 0 987
box -33 -27 33 27
use poly_li1_contact  poly_li1_contact_5
timestamp 1645652543
transform 0 1 148 -1 0 444
box -33 -27 33 27
use nmos_bottom  nmos_bottom_0
timestamp 1646007130
transform -1 0 360 0 1 101
box 0 0 248 302
use pmos2_1  pmos2_1_0
timestamp 1647326732
transform 1 0 43 0 1 1450
box 52 -460 352 37
use li1_M1_contact  li1_M1_contact_6
timestamp 1646004885
transform -1 0 370 0 1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_9
timestamp 1646004885
transform -1 0 370 0 1 518
box -53 -33 29 33
use nmos_top  nmos_top_0
timestamp 1645648650
transform -1 0 553 0 1 101
box -1 0 247 309
use pmos2_1  pmos2_1_1
timestamp 1647326732
transform 1 0 219 0 1 1450
box 52 -460 352 37
use li1_M1_contact  li1_M1_contact_3
timestamp 1646004885
transform -1 0 422 0 1 1088
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1646004885
transform -1 0 430 0 1 264
box -53 -33 29 33
use poly_li1_contact  poly_li1_contact_3
timestamp 1645652543
transform 0 1 378 -1 0 987
box -33 -27 33 27
use poly_li1_contact  poly_li1_contact_2
timestamp 1645652543
transform 0 -1 370 1 0 444
box -33 -27 33 27
use li1_M1_contact  li1_M1_contact_7
timestamp 1646004885
transform 1 0 822 0 -1 1088
box -53 -33 29 33
use pmos2_1  pmos2_1_3
timestamp 1647326732
transform -1 0 1113 0 1 1450
box 52 -460 352 37
use nmos_bottom  nmos_bottom_1
timestamp 1646007130
transform -1 0 1026 0 1 101
box 0 0 248 302
use diff_ring_side  diff_ring_side_2
timestamp 1646086970
transform 1 0 666 0 1 0
box -84 0 84 1575
use li1_M1_contact  li1_M1_contact_8
timestamp 1646004885
transform 1 0 888 0 1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_4
timestamp 1646004885
transform -1 0 1086 0 -1 1088
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_10
timestamp 1646004885
transform 1 0 888 0 1 518
box -53 -33 29 33
use poly_li1_contact  poly_li1_contact_7
timestamp 1645652543
transform 0 -1 888 -1 0 987
box -33 -27 33 27
use pmos2_1  pmos2_1_2
timestamp 1647326732
transform -1 0 1289 0 1 1450
box 52 -460 352 37
use poly_li1_contact  poly_li1_contact_4
timestamp 1645652543
transform 0 -1 888 -1 0 444
box -33 -27 33 27
use li1_M1_contact  li1_M1_contact_1
timestamp 1646004885
transform 1 0 1096 0 1 264
box -53 -33 29 33
use nmos_top_trim1  nmos_top_trim1_0
timestamp 1646008046
transform 1 0 972 0 1 101
box 0 0 248 309
use li1_M1_contact  li1_M1_contact_12
timestamp 1646004885
transform -1 0 1184 0 1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_11
timestamp 1646004885
transform -1 0 1184 0 1 518
box -53 -33 29 33
use poly_li1_contact  poly_li1_contact_6
timestamp 1645652543
transform 0 -1 1184 -1 0 987
box -33 -27 33 27
use poly_li1_contact  poly_li1_contact_1
timestamp 1645652543
transform 0 -1 1184 -1 0 444
box -33 -27 33 27
use diff_ring_side  diff_ring_side_3
timestamp 1646086970
transform 1 0 1332 0 1 0
box -84 0 84 1575
use li1_M1_contact  li1_M1_contact_14
timestamp 1646004885
transform 1 0 1480 0 1 518
box -53 -33 29 33
use poly_li1_contact  poly_li1_contact_10
timestamp 1645652543
transform 0 1 1480 -1 0 444
box -33 -27 33 27
use nmos_bottom  nmos_bottom_2
timestamp 1646007130
transform -1 0 1692 0 1 101
box 0 0 248 302
use poly_li1_contact  poly_li1_contact_11
timestamp 1645652543
transform 0 -1 1702 -1 0 444
box -33 -27 33 27
use nmos_top_trim2  nmos_top_trim2_2
timestamp 1647327697
transform -1 0 1886 0 1 101
box 0 0 248 309
use li1_M1_contact  li1_M1_contact_2
timestamp 1646004885
transform 1 0 1762 0 1 264
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_13
timestamp 1646004885
transform 1 0 1480 0 1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_16
timestamp 1646004885
transform 1 0 1702 0 1 888
box -53 -33 29 33
use poly_li1_contact  poly_li1_contact_8
timestamp 1645652543
transform 0 1 1480 -1 0 987
box -33 -27 33 27
use pmos2_1  pmos2_1_4
timestamp 1647326732
transform 1 0 1375 0 1 1450
box 52 -460 352 37
use poly_li1_contact  poly_li1_contact_9
timestamp 1645652543
transform 0 1 1707 -1 0 987
box -33 -27 33 27
use pmos2_1  pmos2_1_5
timestamp 1647326732
transform 1 0 1551 0 1 1450
box 52 -460 352 37
use li1_M1_contact  li1_M1_contact_5
timestamp 1646004885
transform 1 0 1490 0 1 1088
box -53 -33 29 33
use diff_ring_side  diff_ring_side_0
timestamp 1646086970
transform 1 0 1998 0 1 0
box -84 0 84 1575
<< end >>
