magic
tech sky130A
magscale 1 2
timestamp 1654886336
<< locali >>
rect 205 871 239 905
rect 427 871 461 905
rect 1389 871 1423 905
rect 3313 871 3347 905
rect 7161 871 7195 905
rect 9085 871 9119 905
rect 12933 871 12967 905
rect 14857 871 14891 905
rect 205 797 239 831
rect 5977 797 6011 831
rect 11749 797 11783 831
rect 11971 797 12005 831
rect 15079 797 15113 831
rect 205 723 239 757
rect 427 723 461 757
rect 1389 723 1423 757
rect 5977 723 6011 757
rect 6199 723 6233 757
rect 7161 723 7195 757
rect 205 649 239 683
rect 427 649 461 683
rect 4275 649 4309 683
rect 5977 649 6011 683
rect 6199 649 6233 683
rect 10047 649 10081 683
rect 11749 649 11783 683
rect 11971 649 12005 683
rect 15819 649 15853 683
rect 205 575 239 609
rect 427 575 461 609
rect 1389 575 1423 609
rect 2351 575 2385 609
rect 5237 575 5271 609
rect 8123 575 8157 609
rect 11009 575 11043 609
rect 13895 575 13929 609
rect 205 501 239 535
rect 427 501 461 535
rect 2351 501 2385 535
rect 3313 501 3347 535
rect 3535 501 3569 535
rect 4275 501 4309 535
rect 5237 501 5271 535
rect 5977 501 6011 535
rect 6199 501 6233 535
rect 8123 501 8157 535
rect 9085 501 9119 535
rect 9307 501 9341 535
rect 10047 501 10081 535
rect 11009 501 11043 535
rect 11749 501 11783 535
rect 11971 501 12005 535
rect 13895 501 13929 535
rect 14857 501 14891 535
rect 15079 501 15113 535
rect 15819 501 15853 535
rect 205 427 239 461
rect 427 427 461 461
rect 3535 427 3569 461
rect 4275 427 4309 461
rect 6199 427 6233 461
rect 9307 427 9341 461
rect 10047 427 10081 461
rect 11971 427 12005 461
rect 15079 427 15113 461
rect 15819 427 15853 461
<< metal1 >>
rect 5643 945 15039 979
rect 15005 905 15039 945
rect 1458 871 3277 905
rect 3359 871 7149 905
rect 7230 871 9049 905
rect 9131 871 12921 905
rect 13003 871 14822 905
rect 15005 873 17446 905
rect 15021 871 17446 873
rect 251 797 5965 831
rect 6047 797 11713 831
rect 13007 797 17701 831
rect 19593 797 19627 831
rect 13007 757 13041 797
rect 11449 723 13041 757
rect 4567 649 5645 683
rect 10339 649 11343 683
rect 2421 575 5201 609
rect 5283 575 8111 609
rect 8193 575 10973 609
rect 11055 575 13883 609
rect 4715 501 4979 535
rect 10487 501 10751 535
rect 16259 501 16523 535
rect 461 427 3523 461
rect 3605 427 4239 461
rect 4321 427 6187 461
rect 6269 427 9295 461
rect 9377 427 10011 461
rect 10093 427 11959 461
rect 12041 427 15067 461
rect 15149 427 15783 461
rect 16111 427 18523 461
use li1_M1_contact  li1_M1_contact_9 pcells
timestamp 1648061256
transform 1 0 5032 0 1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_8
timestamp 1648061256
transform -1 0 4662 0 -1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_6
timestamp 1648061256
transform 1 0 5624 0 1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_20
timestamp 1648061256
transform -1 0 5624 0 -1 962
box -53 -33 29 33
use dffsnrnx1_pcell  dffsnrnx1_pcell_0 pcells
timestamp 1654884202
transform 1 0 0 0 1 0
box -87 -34 5859 1550
use dffsnrnx1_pcell  dffsnrnx1_pcell_1
timestamp 1654884202
transform 1 0 5772 0 1 0
box -87 -34 5859 1550
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform 1 0 222 0 1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_15
timestamp 1648061256
transform -1 0 4514 0 -1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_17
timestamp 1648061256
transform 1 0 10804 0 1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_12
timestamp 1648061256
transform -1 0 10434 0 -1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_5
timestamp 1648061256
transform -1 0 10286 0 -1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_7
timestamp 1648061256
transform 1 0 11396 0 1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_3
timestamp 1648061256
transform -1 0 11396 0 -1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_2
timestamp 1648061256
transform 1 0 11766 0 1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform -1 0 5994 0 -1 814
box -53 -33 29 33
use dffsnrnx1_pcell  dffsnrnx1_pcell_2
timestamp 1654884202
transform 1 0 11544 0 1 0
box -87 -34 5859 1550
use li1_M1_contact  li1_M1_contact_14
timestamp 1648061256
transform 1 0 16576 0 1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_13
timestamp 1648061256
transform -1 0 16206 0 -1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_4
timestamp 1648061256
transform 1 0 17168 0 1 444
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_19
timestamp 1648061256
transform -1 0 16058 0 -1 444
box -53 -33 29 33
use voter3x1_pcell  voter3x1_pcell_0 pcells
timestamp 1652393968
transform 1 0 17316 0 1 0
box -87 -34 2529 1550
use li1_M1_contact  li1_M1_contact_16
timestamp 1648061256
transform -1 0 19610 0 -1 814
box -53 -33 29 33
use VOTER3X1  VOTER3X1_0
timestamp 1652394001
transform 1 0 17316 0 1 1703
box -87 -34 2529 1550
use DFFSNRNX1  DFFSNRNX1_2
timestamp 1652427256
transform 1 0 11544 0 1 1703
box -87 -34 5859 1550
use DFFSNRNX1  DFFSNRNX1_1
timestamp 1652427256
transform 1 0 5772 0 1 1703
box -87 -34 5859 1550
use DFFSNRNX1  DFFSNRNX1_0
timestamp 1652427256
transform 1 0 0 0 1 1703
box -87 -34 5859 1550
<< labels >>
rlabel metal1 19593 797 19627 831 1 Q
port 1 nsew signal output
rlabel locali 2351 575 2385 609 1 SN
port 4 nsew signal input
rlabel locali 427 427 461 461 1 RN
port 5 nsew signal input
rlabel locali 427 501 461 535 1 RN
port 5 nsew signal input
rlabel locali 427 575 461 609 1 RN
port 5 nsew signal input
rlabel locali 427 649 461 683 1 RN
port 5 nsew signal input
rlabel locali 427 723 461 757 1 RN
port 5 nsew signal input
rlabel locali 427 871 461 905 1 RN
port 5 nsew signal input
rlabel locali 205 797 239 831 1 D
port 2 nsew signal input
rlabel locali 205 723 239 757 1 D
port 2 nsew signal input
rlabel locali 205 649 239 683 1 D
port 2 nsew signal input
rlabel locali 205 575 239 609 1 D
port 2 nsew signal input
rlabel locali 205 501 239 535 1 D
port 2 nsew signal input
rlabel locali 205 427 239 461 1 D
port 2 nsew signal input
rlabel locali 205 871 239 905 1 D
port 2 nsew signal input
rlabel locali 2351 501 2385 535 1 SN
port 4 nsew signal input
rlabel locali 5977 797 6011 831 1 D
port 2 nsew signal input
rlabel locali 11749 797 11783 831 1 D
port 2 nsew signal input
rlabel locali 11749 501 11783 535 1 D
port 2 nsew signal input
rlabel locali 5977 723 6011 757 1 D
port 2 nsew signal input
rlabel locali 5977 501 6011 535 1 D
port 2 nsew signal input
rlabel locali 3535 427 3569 461 1 RN
port 5 nsew signal input
rlabel locali 4275 427 4309 461 1 RN
port 5 nsew signal input
rlabel locali 3535 501 3569 535 1 RN
port 5 nsew signal input
rlabel locali 4275 501 4309 535 1 RN
port 5 nsew signal input
rlabel locali 4275 649 4309 683 1 RN
port 5 nsew signal input
rlabel locali 6199 427 6233 461 1 RN
port 5 nsew signal input
rlabel locali 6199 501 6233 535 1 RN
port 5 nsew signal input
rlabel locali 6199 723 6233 757 1 RN
port 5 nsew signal input
rlabel locali 9307 427 9341 461 1 RN
port 5 nsew signal input
rlabel locali 9307 501 9341 535 1 RN
port 5 nsew signal input
rlabel locali 10047 427 10081 461 1 RN
port 5 nsew signal input
rlabel locali 10047 501 10081 535 1 RN
port 5 nsew signal input
rlabel locali 11971 427 12005 461 1 RN
port 5 nsew signal input
rlabel locali 11971 501 12005 535 1 RN
port 5 nsew signal input
rlabel locali 11971 797 12005 831 1 RN
port 5 nsew signal input
rlabel locali 15079 427 15113 461 1 RN
port 5 nsew signal input
rlabel locali 15819 427 15853 461 1 RN
port 5 nsew signal input
rlabel locali 15819 501 15853 535 1 RN
port 5 nsew signal input
rlabel locali 15079 501 15113 535 1 RN
port 5 nsew signal input
rlabel locali 9085 871 9119 905 1 CLK
port 3 nsew signal input
rlabel locali 7161 871 7195 905 1 CLK
port 3 nsew signal input
rlabel locali 3313 871 3347 905 1 CLK
port 3 nsew signal input
rlabel locali 1389 871 1423 905 1 CLK
port 3 nsew signal input
rlabel locali 1389 723 1423 757 1 CLK
port 3 nsew signal input
rlabel locali 1389 575 1423 609 1 CLK
port 3 nsew signal input
rlabel locali 3313 501 3347 535 1 CLK
port 3 nsew signal input
rlabel locali 7161 723 7195 757 1 CLK
port 3 nsew signal input
rlabel locali 12933 871 12967 905 1 CLK
port 3 nsew signal input
rlabel locali 14857 871 14891 905 1 CLK
port 3 nsew signal input
rlabel locali 14857 501 14891 535 1 CLK
port 3 nsew signal input
rlabel locali 5237 575 5271 609 1 SN
port 4 nsew signal input
rlabel locali 5237 501 5271 535 1 SN
port 4 nsew signal input
rlabel locali 8123 575 8157 609 1 SN
port 4 nsew signal input
rlabel locali 5977 649 6011 683 1 D
port 2 nsew signal input
rlabel locali 6199 649 6233 683 1 RN
port 5 nsew signal input
rlabel locali 8123 501 8157 535 1 SN
port 4 nsew signal input
rlabel locali 11009 575 11043 609 1 SN
port 4 nsew signal input
rlabel locali 11009 501 11043 535 1 SN
port 4 nsew signal input
rlabel locali 10047 649 10081 683 1 RN
port 5 nsew signal input
rlabel locali 13895 575 13929 609 1 SN
port 4 nsew signal input
rlabel locali 11971 649 12005 683 1 RN
port 5 nsew signal input
rlabel locali 11749 649 11783 683 1 D
port 2 nsew signal input
rlabel locali 15819 649 15853 683 1 RN
port 5 nsew signal input
rlabel locali 13895 501 13929 535 1 SN
port 4 nsew signal input
rlabel locali 9085 501 9119 535 1 CLK
port 3 nsew signal input
<< end >>
