* SPICE3 file created from VOTER3X1.ext - technology: sky130A

.subckt VOTER3X1 Y A B C VDD VSS
X0 Y a_392_209 VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8p pd=4.58u as=2.78p ps=2.278u w=2u l=0.15u M=2
X1 a_392_209 A a_881_1051 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X2 VDD B a_217_1051 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X3 a_881_1051 C a_217_1051 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X4 VSS B a_778_101 VSS sky130_fd_pr__nfet_01v8 ad=1.6781p pd=1.281u as=0p ps=0u w=3u l=0.15u
X5 VSS B a_112_101 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X6 VSS C a_1444_101 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X7 VDD A a_217_1051 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X8 a_881_1051 B a_217_1051 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X9 a_881_1051 C a_392_209 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X10 a_392_209 A a_1444_101 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X11 Y a_392_209 VSS VSS sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=0p ps=0u w=3u l=0.15u
X12 a_392_209 A a_112_101 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X13 a_392_209 C a_778_101 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
C0 VDD a_217_1051 3.12fF
C1 VDD VSS 4.82fF
.ends
