* SPICE3 file created from AO3X1.ext - technology: sky130A

.subckt AO3X1 Y A B C VDD VSS
X0 VDD B a_223_1051 VDD sky130_fd_pr__pfet_01v8 ad=2.78e+12p pd=2.278e+07u as=0p ps=0u w=2e+06u l=150000u M=2
X1 a_223_1051 C a_683_1051 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X2 a_223_1051 A a_108_101 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X3 Y a_223_1051 VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=150000u M=2
X4 a_223_1051 A VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X5 Y a_223_1051 VSS VSS sky130_fd_pr__nfet_01v8 ad=1.791e+11p pd=1.57e+06u as=1.499e+12p ps=1.124e+07u w=3e+06u l=150000u
X6 VSS B a_108_101 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X7 VSS C a_223_1051 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
C0 a_223_1051 VDD 2.81fF
C1 VDD VSS 2.67fF
.ends
