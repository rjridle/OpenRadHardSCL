magic
tech sky130A
magscale 1 2
timestamp 1642975841
<< nwell >>
rect -159 612 9 1353
<< psubdiff >>
rect -106 455 -44 549
rect -106 421 -91 455
rect -57 421 -44 455
rect -106 387 -44 421
rect -106 353 -91 387
rect -57 353 -44 387
rect -106 319 -44 353
rect -106 285 -91 319
rect -57 285 -44 319
rect -106 251 -44 285
rect -106 217 -91 251
rect -57 217 -44 251
rect -106 183 -44 217
rect -106 149 -91 183
rect -57 149 -44 183
rect -106 115 -44 149
rect -106 81 -92 115
rect -58 81 -44 115
rect -106 0 -44 81
<< nsubdiff >>
rect -106 1249 -44 1317
rect -106 1215 -92 1249
rect -57 1215 -44 1249
rect -106 1181 -44 1215
rect -106 1147 -92 1181
rect -57 1147 -44 1181
rect -106 1113 -44 1147
rect -106 1079 -92 1113
rect -57 1079 -44 1113
rect -106 1045 -44 1079
rect -106 1011 -92 1045
rect -57 1011 -44 1045
rect -106 977 -44 1011
rect -106 943 -92 977
rect -57 943 -44 977
rect -106 909 -44 943
rect -106 875 -92 909
rect -57 875 -44 909
rect -106 841 -44 875
rect -106 807 -92 841
rect -57 807 -44 841
rect -106 773 -44 807
rect -106 739 -92 773
rect -57 739 -44 773
rect -106 648 -44 739
<< psubdiffcont >>
rect -91 421 -57 455
rect -91 353 -57 387
rect -91 285 -57 319
rect -91 217 -57 251
rect -91 149 -57 183
rect -92 81 -58 115
<< nsubdiffcont >>
rect -92 1215 -57 1249
rect -92 1147 -57 1181
rect -92 1079 -57 1113
rect -92 1011 -57 1045
rect -92 943 -57 977
rect -92 875 -57 909
rect -92 807 -57 841
rect -92 739 -57 773
<< locali >>
rect -106 1249 -44 1332
rect -106 1215 -92 1249
rect -57 1215 -44 1249
rect -106 1181 -44 1215
rect -106 1147 -92 1181
rect -57 1147 -44 1181
rect -106 1113 -44 1147
rect -106 1079 -92 1113
rect -57 1079 -44 1113
rect -106 1045 -44 1079
rect -106 1011 -92 1045
rect -57 1011 -44 1045
rect -106 977 -44 1011
rect -106 943 -92 977
rect -57 943 -44 977
rect -106 909 -44 943
rect -106 875 -92 909
rect -57 875 -44 909
rect -106 841 -44 875
rect -106 807 -92 841
rect -57 807 -44 841
rect -106 773 -44 807
rect -106 739 -92 773
rect -57 739 -44 773
rect -106 648 -44 739
rect -106 455 -44 549
rect -106 421 -91 455
rect -57 421 -44 455
rect -106 387 -44 421
rect -106 353 -91 387
rect -57 353 -44 387
rect -106 319 -44 353
rect -106 285 -91 319
rect -57 285 -44 319
rect -106 251 -44 285
rect -106 217 -91 251
rect -57 217 -44 251
rect -106 183 -44 217
rect -106 149 -91 183
rect -57 149 -44 183
rect -106 115 -44 149
rect -106 81 -92 115
rect -58 81 -44 115
rect -106 0 -44 81
<< viali >>
rect -92 1215 -57 1249
rect -92 1147 -57 1181
rect -92 1079 -57 1113
rect -92 1011 -57 1045
rect -92 943 -57 977
rect -92 875 -57 909
rect -92 807 -57 841
rect -92 739 -57 773
rect -91 421 -57 455
rect -91 353 -57 387
rect -91 285 -57 319
rect -91 217 -57 251
rect -91 149 -57 183
rect -92 81 -58 115
<< metal1 >>
rect -106 1249 -44 1332
rect -106 1215 -92 1249
rect -57 1215 -44 1249
rect -106 1181 -44 1215
rect -106 1147 -92 1181
rect -57 1147 -44 1181
rect -106 1113 -44 1147
rect -106 1079 -92 1113
rect -57 1079 -44 1113
rect -106 1045 -44 1079
rect -106 1011 -92 1045
rect -57 1011 -44 1045
rect -106 977 -44 1011
rect -106 943 -92 977
rect -57 943 -44 977
rect -106 909 -44 943
rect -106 875 -92 909
rect -57 875 -44 909
rect -106 841 -44 875
rect -106 807 -92 841
rect -57 807 -44 841
rect -106 773 -44 807
rect -106 739 -92 773
rect -57 739 -44 773
rect -106 648 -44 739
rect -106 455 -44 549
rect -106 421 -91 455
rect -57 421 -44 455
rect -106 387 -44 421
rect -106 353 -91 387
rect -57 353 -44 387
rect -106 319 -44 353
rect -106 285 -91 319
rect -57 285 -44 319
rect -106 251 -44 285
rect -106 217 -91 251
rect -57 217 -44 251
rect -106 183 -44 217
rect -106 149 -91 183
rect -57 149 -44 183
rect -106 115 -44 149
rect -106 81 -92 115
rect -58 81 -44 115
rect -106 0 -44 81
<< end >>
