* SPICE3 file created from XOR2X1.ext - technology: sky130A

.subckt XOR2X1 Y A B VDD VSS
X0 a_807_990# B VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.36p ps=2.736u w=2u l=0.15u M=2
X1 a_185_209# A VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X2 VSS A a_556_101# VSS sky130_fd_pr__nfet_01v8 ad=2.6398p pd=1.934u as=0p ps=0u w=3u l=0.15u
X3 a_185_209# A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X4 a_575_1051# a_807_990# Y VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.16p ps=9.16u w=2u l=0.15u M=2
X5 Y a_185_209# a_1222_101# VSS sky130_fd_pr__nfet_01v8 ad=3.582p pd=3.14u as=0p ps=0u w=3u l=0.15u
X6 a_1241_1051# B VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X7 a_807_990# B VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X8 a_1241_1051# a_185_209# Y VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X9 Y B a_556_101# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X10 VDD A a_575_1051# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X11 VSS a_807_990# a_1222_101# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
C0 a_807_990# B 2.21fF
.ends
