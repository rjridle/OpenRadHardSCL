* SPICE3 file created from VOTERN3X1.ext - technology: sky130A

.subckt VOTERN3X1 YN A B C VDD GND
X0 YN C.t3 a_778_101.t0 GND sky130_fd_pr__nfet_01v8 ad=5.373p pd=4.72u as=0p ps=0u w=0u l=0u
X1 GND B.t1 a_778_101.t0 GND sky130_fd_pr__nfet_01v8 ad=5.373p pd=4.71u as=0p ps=0u w=0u l=0u
X2 GND B.t2 a_112_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X3 GND C.t1 a_1444_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X4 YN.t5 A.t0 a_881_1051.t6  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X5 VDD.t4 B.t0 a_217_1051.t5 VDD.t3 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X6 a_881_1051.t3 C.t0 a_217_1051.t1  sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X7 YN A.t2 a_1444_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X8 VDD.t12 A.t1 a_217_1051.t3  �M�	 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X9 a_881_1051.t5 B.t3 a_217_1051.t7 �M�	 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X10 a_881_1051.t0 C.t2 YN.t0  �M�	 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X11 YN A.t3 a_112_101.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X12 a_217_1051.t4 B.t4 VDD.t15 �M�	 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X13 a_217_1051.t6 B.t5 a_881_1051.t2  �M�	 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X14 a_217_1051.t2 A.t4 VDD.t10 �M�	 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X15 a_881_1051.t7 A.t5 YN.t4  �M�	 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X16 a_217_1051.t0 C.t4 a_881_1051.t1 �M�	 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X17 YN.t2 C.t5 a_881_1051.t4  �M�	 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
C0 YN VDD 0.73fF
C1 B A 0.96fF
C2 A C 0.26fF
C3 B C 0.15fF
C4 A VDD 1.95fF
C5 A YN 0.30fF
C6 B VDD 1.14fF
C7 C VDD 0.73fF
C8 B YN 0.05fF
C9 YN C 0.27fF
R0 A.n0 A.t5 475.572
R1 A.n2 A.t1 469.145
R2 A.n2 A.t4 384.527
R3 A.n0 A.t0 384.527
R4 A.n3 A.t3 370.613
R5 A.n1 A.t2 370.613
R6 A.n1 A.n0 128.028
R7 A.n3 A.n2 126.97
R8 A.n4 A.n1 9.501
R9 A.n4 A.n3 4.65
R10 A.n4 A 0.046
R11 a_881_1051.n4 a_881_1051.t7 179.895
R12 a_881_1051.n2 a_881_1051.n1 165.613
R13 a_881_1051.n2 a_881_1051.n0 142.653
R14 a_881_1051.n4 a_881_1051.n3 106.183
R15 a_881_1051.n5 a_881_1051.n4 99.358
R16 a_881_1051.n3 a_881_1051.n2 82.665
R17 a_881_1051.n3 a_881_1051.t4 73.712
R18 a_881_1051.n0 a_881_1051.t1 14.282
R19 a_881_1051.n0 a_881_1051.t3 14.282
R20 a_881_1051.n1 a_881_1051.t2 14.282
R21 a_881_1051.n1 a_881_1051.t5 14.282
R22 a_881_1051.n5 a_881_1051.t6 14.282
R23 a_881_1051.t0 a_881_1051.n5 14.282
R24 YN.n15 YN.n14 227.387
R25 YN.n2 YN.n1 165.613
R26 YN.n15 YN.n2 132.893
R27 YN.n10 YN.n5 126.225
R28 YN.n10 YN.n9 112.771
R29 YN.n14 YN.n13 106.052
R30 YN.n2 YN.n0 99.355
R31 YN.n13 YN.n11 80.526
R32 YN.n9 YN.n8 30
R33 YN.n13 YN.n12 30
R34 YN.n7 YN.n6 24.383
R35 YN.n9 YN.n7 23.684
R36 YN.n5 YN.n4 22.578
R37 YN.n0 YN.t4 14.282
R38 YN.n0 YN.t5 14.282
R39 YN.n1 YN.t0 14.282
R40 YN.n1 YN.t2 14.282
R41 YN.n5 YN.n3 8.58
R42 YN.n14 YN.n10 7.053
R43 YN.n16 YN.n15 4.65
R44 YN.n16 YN 0.046
R45 VDD.n75 VDD.n64 144.705
R46 VDD.n168 VDD.n157 144.705
R47 VDD.n113 VDD.t15 135.539
R48 VDD.n135 VDD.t12 135.539
R49 VDD.n127 VDD.n126 129.849
R50 VDD.n60 VDD.n59 92.5
R51 VDD.n58 VDD.n57 92.5
R52 VDD.n56 VDD.n55 92.5
R53 VDD.n54 VDD.n53 92.5
R54 VDD.n62 VDD.n61 92.5
R55 VDD.n153 VDD.n152 92.5
R56 VDD.n151 VDD.n150 92.5
R57 VDD.n149 VDD.n148 92.5
R58 VDD.n147 VDD.n146 92.5
R59 VDD.n155 VDD.n154 92.5
R60 VDD.n101 VDD.n100 92.5
R61 VDD.n99 VDD.n98 92.5
R62 VDD.n97 VDD.n96 92.5
R63 VDD.n95 VDD.n94 92.5
R64 VDD.n103 VDD.n102 92.5
R65 VDD.n14 VDD.n1 92.5
R66 VDD.n5 VDD.n4 92.5
R67 VDD.n7 VDD.n6 92.5
R68 VDD.n9 VDD.n8 92.5
R69 VDD.n11 VDD.n10 92.5
R70 VDD.n13 VDD.n12 92.5
R71 VDD.n21 VDD.n20 92.059
R72 VDD.n74 VDD.n73 92.059
R73 VDD.n167 VDD.n166 92.059
R74 VDD.n109 VDD.n108 92.059
R75 VDD.n20 VDD.n16 67.194
R76 VDD.n20 VDD.n17 67.194
R77 VDD.n20 VDD.n18 67.194
R78 VDD.n20 VDD.n19 67.194
R79 VDD.n93 VDD.n92 44.141
R80 VDD.n5 VDD.n3 44.141
R81 VDD.n92 VDD.n90 44.107
R82 VDD.n3 VDD.n2 44.107
R83 VDD.n20 VDD.n15 41.052
R84 VDD.n68 VDD.n66 39.742
R85 VDD.n68 VDD.n67 39.742
R86 VDD.n70 VDD.n69 39.742
R87 VDD.n105 VDD.n104 39.742
R88 VDD.n165 VDD.n162 39.742
R89 VDD.n165 VDD.n164 39.742
R90 VDD.n161 VDD.n160 39.742
R91 VDD.n92 VDD.n91 38
R92 VDD.n66 VDD.n65 36.774
R93 VDD.n164 VDD.n163 36.774
R94 VDD.n1 VDD.n0 30.923
R95 VDD.n73 VDD.n71 26.38
R96 VDD.n73 VDD.n70 26.38
R97 VDD.n73 VDD.n68 26.38
R98 VDD.n73 VDD.n72 26.38
R99 VDD.n108 VDD.n106 26.38
R100 VDD.n108 VDD.n105 26.38
R101 VDD.n108 VDD.n107 26.38
R102 VDD.n166 VDD.n165 26.38
R103 VDD.n166 VDD.n161 26.38
R104 VDD.n166 VDD.n159 26.38
R105 VDD.n166 VDD.n158 26.38
R106 VDD.n111 VDD.n103 22.915
R107 VDD.n23 VDD.n14 22.915
R108 VDD.n28  �M�	 20.457
R109 VDD.n175 �M�	 20.457
R110 VDD.n131  �M�	 20.457
R111 VDD.n39  �M�	 17.9
R112 VDD.n82 �M�	 17.9
R113 VDD.n118 �M�	 17.9
R114 VDD.n103 VDD.n101 14.864
R115 VDD.n101 VDD.n99 14.864
R116 VDD.n99 VDD.n97 14.864
R117 VDD.n97 VDD.n95 14.864
R118 VDD.n95 VDD.n93 14.864
R119 VDD.n62 VDD.n60 14.864
R120 VDD.n60 VDD.n58 14.864
R121 VDD.n58 VDD.n56 14.864
R122 VDD.n56 VDD.n54 14.864
R123 VDD.n54 VDD.n52 14.864
R124 VDD.n52 VDD.n51 14.864
R125 VDD.n155 VDD.n153 14.864
R126 VDD.n153 VDD.n151 14.864
R127 VDD.n151 VDD.n149 14.864
R128 VDD.n149 VDD.n147 14.864
R129 VDD.n147 VDD.n145 14.864
R130 VDD.n145 VDD.n144 14.864
R131 VDD.n14 VDD.n13 14.864
R132 VDD.n13 VDD.n11 14.864
R133 VDD.n11 VDD.n9 14.864
R134 VDD.n9 VDD.n7 14.864
R135 VDD.n7 VDD.n5 14.864
R136 VDD.n76 VDD.n63 14.864
R137 VDD.n169 VDD.n156 14.864
R138 VDD.n126 VDD.t10 14.282
R139 VDD.n126 VDD.t4 14.282
R140 VDD.n129 VDD.n127 9.083
R141 VDD.n23 VDD.n22 8.855
R142 VDD.n22 VDD.n21 8.855
R143 VDD.n26 VDD.n25 8.855
R144 VDD.n25 VDD.n24 8.855
R145 VDD.n30 VDD.n29 8.855
R146 VDD.n29 VDD.n28 8.855
R147 VDD.n33 VDD.n32 8.855
R148 VDD.n32 �ޞ�U 8.855
R149 VDD.n37 VDD.n36 8.855
R150 VDD.n36 VDD.n35 8.855
R151 VDD.n41 VDD.n40 8.855
R152 VDD.n40 VDD.n39 8.855
R153 VDD.n45 VDD.n44 8.855
R154 VDD.n44 VDD.n43 8.855
R155 VDD.n49 VDD.n48 8.855
R156 VDD.n48 VDD.n47 8.855
R157 VDD.n76 VDD.n75 8.855
R158 VDD.n75 VDD.n74 8.855
R159 VDD.n80 VDD.n79 8.855
R160 VDD.n79 VDD.n78 8.855
R161 VDD.n84 VDD.n83 8.855
R162 VDD.n83 VDD.n82 8.855
R163 VDD.n88 VDD.n87 8.855
R164 VDD.n87 VDD.n86 8.855
R165 VDD.n180 VDD.n179 8.855
R166 VDD.n179  �M�	 8.855
R167 VDD.n177 VDD.n176 8.855
R168 VDD.n176 VDD.n175 8.855
R169 VDD.n173 VDD.n172 8.855
R170 VDD.n172 VDD.n171 8.855
R171 VDD.n169 VDD.n168 8.855
R172 VDD.n168 VDD.n167 8.855
R173 VDD.n142 VDD.n141 8.855
R174 VDD.n141 VDD.n140 8.855
R175 VDD.n138 VDD.n137 8.855
R176 VDD.n137 VDD.n136 8.855
R177 VDD.n133 VDD.n132 8.855
R178 VDD.n132 VDD.n131 8.855
R179 VDD.n129 VDD.n128 8.855
R180 VDD.n128 �M�	 8.855
R181 VDD.n124 VDD.n123 8.855
R182 VDD.n123 VDD.n122 8.855
R183 VDD.n120 VDD.n119 8.855
R184 VDD.n119 VDD.n118 8.855
R185 VDD.n116 VDD.n115 8.855
R186 VDD.n115 VDD.n114 8.855
R187 VDD.n111 VDD.n110 8.855
R188 VDD.n110 VDD.n109 8.855
R189 VDD.n63 VDD.n62 8.051
R190 VDD.n156 VDD.n155 8.051
R191 VDD.n31 VDD.n30 4.65
R192 VDD.n34 VDD.n33 4.65
R193 VDD.n38 VDD.n37 4.65
R194 VDD.n42 VDD.n41 4.65
R195 VDD.n46 VDD.n45 4.65
R196 VDD.n50 VDD.n49 4.65
R197 VDD.n77 VDD.n76 4.65
R198 VDD.n81 VDD.n80 4.65
R199 VDD.n85 VDD.n84 4.65
R200 VDD.n89 VDD.n88 4.65
R201 VDD.n181 VDD.n180 4.65
R202 VDD.n178 VDD.n177 4.65
R203 VDD.n174 VDD.n173 4.65
R204 VDD.n170 VDD.n169 4.65
R205 VDD.n143 VDD.n142 4.65
R206 VDD.n139 VDD.n138 4.65
R207 VDD.n134 VDD.n133 4.65
R208 VDD.n130 VDD.n129 4.65
R209 VDD.n125 VDD.n124 4.65
R210 VDD.n121 VDD.n120 4.65
R211 VDD.n117 VDD.n116 4.65
R212 VDD.n112 VDD.n111 4.65
R213 VDD.n27 VDD.n23 2.933
R214 VDD.n116 VDD.n113 2.89
R215 VDD.n27 VDD.n26 2.844
R216 VDD.n35  �M�	 2.557
R217 VDD.n86  2.557
R218 VDD.n122 VDD.t3 2.557
R219 VDD.n138 VDD.n135 2.477
R220 VDD.n31 VDD.n27 1.063
R221 VDD.n77 VDD.n50 0.29
R222 VDD.n170 VDD.n143 0.29
R223 VDD.n112 VDD 0.207
R224 VDD.n38 VDD.n34 0.181
R225 VDD.n130 VDD.n125 0.181
R226 VDD.n34 VDD.n31 0.145
R227 VDD.n42 VDD.n38 0.145
R228 VDD.n46 VDD.n42 0.145
R229 VDD.n50 VDD.n46 0.145
R230 VDD.n81 VDD.n77 0.145
R231 VDD.n85 VDD.n81 0.145
R232 VDD.n89 VDD.n85 0.145
R233 VDD.n181 VDD.n178 0.145
R234 VDD.n178 VDD.n174 0.145
R235 VDD.n174 VDD.n170 0.145
R236 VDD.n143 VDD.n139 0.145
R237 VDD.n139 VDD.n134 0.145
R238 VDD.n134 VDD.n130 0.145
R239 VDD.n125 VDD.n121 0.145
R240 VDD.n121 VDD.n117 0.145
R241 VDD.n117 VDD.n112 0.145
R242 VDD VDD.n89 0.09
R243 VDD VDD.n181 0.09
R244 B.n2 B.t0 512.525
R245 B.n0 B.t5 477.179
R246 B.n1 B.t1 440.954
R247 B.n3 B.t2 434.527
R248 B.n0 B.t3 406.485
R249 B.n2 B.t4 371.139
R250 B.n3 B.n2 77.972
R251 B.n1 B.n0 21.4
R252 B.n4 B.n1 4.754
R253 B.n4 B.n3 2.079
R254 B.n4 B 0.046
R255 a_217_1051.n2 a_217_1051.t0 179.895
R256 a_217_1051.n4 a_217_1051.n0 157.021
R257 a_217_1051.n5 a_217_1051.n4 124.954
R258 a_217_1051.n3 a_217_1051.n2 106.183
R259 a_217_1051.n2 a_217_1051.n1 99.355
R260 a_217_1051.n4 a_217_1051.n3 82.65
R261 a_217_1051.n3 a_217_1051.t7 73.712
R262 a_217_1051.n1 a_217_1051.t1 14.282
R263 a_217_1051.n1 a_217_1051.t6 14.282
R264 a_217_1051.n0 a_217_1051.t5 14.282
R265 a_217_1051.n0 a_217_1051.t4 14.282
R266 a_217_1051.t3 a_217_1051.n5 14.282
R267 a_217_1051.n5 a_217_1051.t2 14.282
R268 C.n2 C.t0 512.525
R269 C.n0 C.t2 512.525
R270 C.n2 C.t4 371.139
R271 C.n0 C.t5 371.139
R272 C.n3 C.n2 343.521
R273 C.n1 C.n0 343.521
R274 C.n1 C.t1 172.106
R275 C.n3 C.t3 165.68
R276 C.n4 C.n1 5.693
R277 C.n4 C.n3 4.65
R278 C.n4 C 0.046
R279 a_778_101.t0 a_778_101.n0 93.333
R280 a_778_101.n3 a_778_101.n1 79.053
R281 a_778_101.n3 a_778_101.n2 2.109
R282 a_778_101.t0 a_778_101.n3 0.195
R283 GND.n31 GND.n30 237.558
R284 GND.n73 GND.n72 237.558
R285 GND.n28 GND.n27 210.82
R286 GND.n75 GND.n74 210.82
R287 GND.n83 GND.n82 172.612
R288 GND.n53 GND.n52 151.605
R289 GND.n17 GND.n16 151.605
R290 GND.n52 GND.n51 28.421
R291 GND.n16 GND.n15 28.421
R292 GND.n52 GND.n50 25.263
R293 GND.n16 GND.n14 25.263
R294 GND.n50 GND.n49 24.383
R295 GND.n14 GND.n13 24.383
R296 GND.n29 GND.n28 18.953
R297 GND.n76 GND.n75 18.953
R298 GND.n32 GND.n29 14.864
R299 GND.n77 GND.n76 14.864
R300 GND.n47 GND.n46 9.154
R301 GND.n55 GND.n54 9.154
R302 GND.n58 GND.n57 9.154
R303 GND.n61 GND.n60 9.154
R304 GND.n64 GND.n63 9.154
R305 GND.n67 GND.n66 9.154
R306 GND.n70 GND.n69 9.154
R307 GND.n77 GND.n73 9.154
R308 GND.n80 GND.n79 9.154
R309 GND.n85 GND.n84 9.154
R310 GND.n88 GND.n87 9.154
R311 GND.n41 GND.n40 9.154
R312 GND.n1 GND.n0 9.154
R313 GND.n5 GND.n4 9.154
R314 GND.n8 GND.n7 9.154
R315 GND.n11 GND.n10 9.154
R316 GND.n19 GND.n18 9.154
R317 GND.n22 GND.n21 9.154
R318 GND.n25 GND.n24 9.154
R319 GND.n32 GND.n31 9.154
R320 GND.n35 GND.n34 9.154
R321 GND.n38 GND.n37 9.154
R322 GND.n45 GND.n44 4.65
R323 GND.n42 GND.n41 4.65
R324 GND.n89 GND.n88 4.65
R325 GND.n86 GND.n85 4.65
R326 GND.n81 GND.n80 4.65
R327 GND.n78 GND.n77 4.65
R328 GND.n71 GND.n70 4.65
R329 GND.n68 GND.n67 4.65
R330 GND.n65 GND.n64 4.65
R331 GND.n62 GND.n61 4.65
R332 GND.n59 GND.n58 4.65
R333 GND.n56 GND.n55 4.65
R334 GND.n48 GND.n47 4.65
R335 GND.n6 GND.n5 4.65
R336 GND.n9 GND.n8 4.65
R337 GND.n12 GND.n11 4.65
R338 GND.n20 GND.n19 4.65
R339 GND.n23 GND.n22 4.65
R340 GND.n26 GND.n25 4.65
R341 GND.n33 GND.n32 4.65
R342 GND.n36 GND.n35 4.65
R343 GND.n39 GND.n38 4.65
R344 GND.n19 GND.n17 4.129
R345 GND.n85 GND.n83 4.129
R346 GND.n55 GND.n53 4.129
R347 GND.n3 GND.n2 3.408
R348 GND.n3 GND.n1 2.844
R349 GND.n6 GND.n3 1.063
R350 GND.n44 GND.n43 0.474
R351 GND.n33 GND.n26 0.29
R352 GND.n78 GND.n71 0.29
R353 GND.n45 GND 0.207
R354 GND.n12 GND.n9 0.181
R355 GND.n62 GND.n59 0.181
R356 GND.n9 GND.n6 0.145
R357 GND.n20 GND.n12 0.145
R358 GND.n23 GND.n20 0.145
R359 GND.n26 GND.n23 0.145
R360 GND.n36 GND.n33 0.145
R361 GND.n39 GND.n36 0.145
R362 GND.n42 GND.n39 0.145
R363 GND.n89 GND.n86 0.145
R364 GND.n86 GND.n81 0.145
R365 GND.n81 GND.n78 0.145
R366 GND.n71 GND.n68 0.145
R367 GND.n68 GND.n65 0.145
R368 GND.n65 GND.n62 0.145
R369 GND.n59 GND.n56 0.145
R370 GND.n56 GND.n48 0.145
R371 GND.n48 GND.n45 0.145
R372 GND GND.n42 0.09
R373 GND GND.n89 0.09
R374 a_112_101.n4 a_112_101.n2 41.528
R375 a_112_101.n1 a_112_101.n0 33.123
R376 a_112_101.t0 a_112_101.n1 10.642
R377 a_112_101.n6 a_112_101.n5 7.966
R378 a_112_101.n4 a_112_101.n3 3.644
R379 a_112_101.t0 a_112_101.n4 1.093
R380 a_112_101.t0 a_112_101.n6 0.088
R381 a_1444_101.n3 a_1444_101.n1 42.788
R382 a_1444_101.t0 a_1444_101.n0 8.137
R383 a_1444_101.n3 a_1444_101.n2 4.665
R384 a_1444_101.t0 a_1444_101.n3 0.06
C10 VDD GND 4.24fF
C11 a_1444_101.n0 GND 0.05fF
C12 a_1444_101.n1 GND 0.13fF
C13 a_1444_101.n2 GND 0.04fF
C14 a_1444_101.n3 GND 0.18fF
C15 a_112_101.n0 GND 0.09fF
C16 a_112_101.n1 GND 0.07fF
C17 a_112_101.n2 GND 0.10fF
C18 a_112_101.n3 GND 0.02fF
C19 a_112_101.n4 GND 0.02fF
C20 a_112_101.n5 GND 0.05fF
C21 a_112_101.n6 GND 0.20fF
C22 a_778_101.n0 GND 0.02fF
C23 a_778_101.n1 GND 0.13fF
C24 a_778_101.n2 GND 0.13fF
C25 a_778_101.n3 GND 0.15fF
C26 a_217_1051.n0 GND 0.42fF
C27 a_217_1051.n1 GND 0.32fF
C28 a_217_1051.n2 GND 0.52fF
C29 a_217_1051.n3 GND 0.30fF
C30 a_217_1051.n4 GND 0.79fF
C31 a_217_1051.n5 GND 0.36fF
C32 VDD.n1 GND 0.04fF
C33 VDD.n2 GND 0.15fF
C34 VDD.n3 GND 0.03fF
C35 VDD.n4 GND 0.02fF
C36 VDD.n5 GND 0.06fF
C37 VDD.n6 GND 0.02fF
C38 VDD.n7 GND 0.02fF
C39 VDD.n8 GND 0.02fF
C40 VDD.n9 GND 0.02fF
C41 VDD.n10 GND 0.02fF
C42 VDD.n11 GND 0.02fF
C43 VDD.n12 GND 0.02fF
C44 VDD.n13 GND 0.02fF
C45 VDD.n14 GND 0.04fF
C46 VDD.n15 GND 0.01fF
C47 VDD.n20 GND 0.50fF
C48 VDD.n21 GND 0.30fF
C49 VDD.n22 GND 0.02fF
C50 VDD.n23 GND 0.04fF
C51 VDD.n24 GND 0.27fF
C52 VDD.n25 GND 0.01fF
C53 VDD.n26 GND 0.02fF
C54 VDD.n27 GND 0.01fF
C55 VDD.n28 GND 0.18fF
C56 VDD.n29 GND 0.01fF
C57 VDD.n30 GND 0.02fF
C58 VDD.n31 GND 0.09fF
C59 VDD.n32 GND 0.02fF
C60 VDD.n33 GND 0.03fF
C61 VDD.n34 GND 0.03fF
C62 VDD.n35 GND 0.15fF
C63 VDD.n36 GND 0.02fF
C64 VDD.n37 GND 0.03fF
C65 VDD.n38 GND 0.03fF
C66 VDD.n39 GND 0.18fF
C67 VDD.n40 GND 0.01fF
C68 VDD.n41 GND 0.02fF
C69 VDD.n42 GND 0.02fF
C70 VDD.n43 GND 0.27fF
C71 VDD.n44 GND 0.01fF
C72 VDD.n45 GND 0.02fF
C73 VDD.n46 GND 0.02fF
C74 VDD.n47 GND 0.30fF
C75 VDD.n48 GND 0.01fF
C76 VDD.n49 GND 0.02fF
C77 VDD.n50 GND 0.04fF
C78 VDD.n51 GND 0.06fF
C79 VDD.n52 GND 0.02fF
C80 VDD.n53 GND 0.02fF
C81 VDD.n54 GND 0.02fF
C82 VDD.n55 GND 0.02fF
C83 VDD.n56 GND 0.02fF
C84 VDD.n57 GND 0.02fF
C85 VDD.n58 GND 0.02fF
C86 VDD.n59 GND 0.02fF
C87 VDD.n60 GND 0.02fF
C88 VDD.n61 GND 0.02fF
C89 VDD.n62 GND 0.02fF
C90 VDD.n63 GND 0.03fF
C91 VDD.n64 GND 0.03fF
C92 VDD.n65 GND 0.24fF
C93 VDD.n66 GND 0.02fF
C94 VDD.n67 GND 0.02fF
C95 VDD.n69 GND 0.02fF
C96 VDD.n73 GND 0.30fF
C97 VDD.n74 GND 0.30fF
C98 VDD.n75 GND 0.01fF
C99 VDD.n76 GND 0.02fF
C100 VDD.n77 GND 0.04fF
C101 VDD.n78 GND 0.27fF
C102 VDD.n79 GND 0.01fF
C103 VDD.n80 GND 0.02fF
C104 VDD.n81 GND 0.02fF
C105 VDD.n82 GND 0.18fF
C106 VDD.n83 GND 0.01fF
C107 VDD.n84 GND 0.02fF
C108 VDD.n85 GND 0.02fF
C109 VDD.n86 GND 0.15fF
C110 VDD.n87 GND 0.02fF
C111 VDD.n88 GND 0.03fF
C112 VDD.n89 GND 0.02fF
C113 VDD.n90 GND 0.15fF
C114 VDD.n91 GND 0.02fF
C115 VDD.n92 GND 0.02fF
C116 VDD.n93 GND 0.06fF
C117 VDD.n94 GND 0.02fF
C118 VDD.n95 GND 0.02fF
C119 VDD.n96 GND 0.02fF
C120 VDD.n97 GND 0.02fF
C121 VDD.n98 GND 0.02fF
C122 VDD.n99 GND 0.02fF
C123 VDD.n100 GND 0.02fF
C124 VDD.n101 GND 0.02fF
C125 VDD.n102 GND 0.04fF
C126 VDD.n103 GND 0.04fF
C127 VDD.n104 GND 0.02fF
C128 VDD.n108 GND 0.50fF
C129 VDD.n109 GND 0.30fF
C130 VDD.n110 GND 0.02fF
C131 VDD.n111 GND 0.04fF
C132 VDD.n112 GND 0.03fF
C133 VDD.n113 GND 0.07fF
C134 VDD.n114 GND 0.27fF
C135 VDD.n115 GND 0.01fF
C136 VDD.n116 GND 0.01fF
C137 VDD.n117 GND 0.02fF
C138 VDD.n118 GND 0.18fF
C139 VDD.n119 GND 0.01fF
C140 VDD.n120 GND 0.02fF
C141 VDD.n121 GND 0.02fF
C142 VDD.n122 GND 0.15fF
C143 VDD.n123 GND 0.02fF
C144 VDD.n124 GND 0.02fF
C145 VDD.n125 GND 0.03fF
C146 VDD.n126 GND 0.09fF
C147 VDD.n127 GND 0.06fF
C148 VDD.n128 GND 0.02fF
C149 VDD.n129 GND 0.02fF
C150 VDD.n130 GND 0.03fF
C151 VDD.n131 GND 0.18fF
C152 VDD.n132 GND 0.01fF
C153 VDD.n133 GND 0.02fF
C154 VDD.n134 GND 0.02fF
C155 VDD.n135 GND 0.07fF
C156 VDD.n136 GND 0.27fF
C157 VDD.n137 GND 0.01fF
C158 VDD.n138 GND 0.01fF
C159 VDD.n139 GND 0.02fF
C160 