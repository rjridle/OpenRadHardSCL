magic
tech sky130A
magscale 1 2
timestamp 1646086970
<< nwell >>
rect -84 832 84 1575
<< psubdiff >>
rect -31 547 31 572
rect -31 513 -17 547
rect 17 513 31 547
rect -31 475 31 513
rect -31 441 -17 475
rect 17 441 31 475
rect -31 403 31 441
rect -31 369 -17 403
rect 17 369 31 403
rect -31 331 31 369
rect -31 297 -17 331
rect 17 297 31 331
rect -31 259 31 297
rect -31 225 -17 259
rect 17 225 31 259
rect -31 187 31 225
rect -31 153 -17 187
rect 17 153 31 187
rect -31 115 31 153
rect -31 81 -17 115
rect 17 81 31 115
rect -31 13 31 81
<< nsubdiff >>
rect -31 1471 31 1539
rect -31 1437 -17 1471
rect 17 1437 31 1471
rect -31 1399 31 1437
rect -31 1365 -17 1399
rect 17 1365 31 1399
rect -31 1327 31 1365
rect -31 1293 -17 1327
rect 17 1293 31 1327
rect -31 1255 31 1293
rect -31 1221 -17 1255
rect 17 1221 31 1255
rect -31 1183 31 1221
rect -31 1149 -17 1183
rect 17 1149 31 1183
rect -31 1111 31 1149
rect -31 1077 -17 1111
rect 17 1077 31 1111
rect -31 1039 31 1077
rect -31 1005 -17 1039
rect 17 1005 31 1039
rect -31 967 31 1005
rect -31 933 -17 967
rect 17 933 31 967
rect -31 868 31 933
<< psubdiffcont >>
rect -17 513 17 547
rect -17 441 17 475
rect -17 369 17 403
rect -17 297 17 331
rect -17 225 17 259
rect -17 153 17 187
rect -17 81 17 115
<< nsubdiffcont >>
rect -17 1437 17 1471
rect -17 1365 17 1399
rect -17 1293 17 1327
rect -17 1221 17 1255
rect -17 1149 17 1183
rect -17 1077 17 1111
rect -17 1005 17 1039
rect -17 933 17 967
<< locali >>
rect -31 1471 31 1554
rect -31 1437 -17 1471
rect 17 1437 31 1471
rect -31 1399 31 1437
rect -31 1365 -17 1399
rect 17 1365 31 1399
rect -31 1327 31 1365
rect -31 1293 -17 1327
rect 17 1293 31 1327
rect -31 1255 31 1293
rect -31 1221 -17 1255
rect 17 1221 31 1255
rect -31 1183 31 1221
rect -31 1149 -17 1183
rect 17 1149 31 1183
rect -31 1111 31 1149
rect -31 1077 -17 1111
rect 17 1077 31 1111
rect -31 1039 31 1077
rect -31 1005 -17 1039
rect 17 1005 31 1039
rect -31 967 31 1005
rect -31 933 -17 967
rect 17 933 31 967
rect -31 868 31 933
rect -31 547 31 572
rect -31 513 -17 547
rect 17 513 31 547
rect -31 475 31 513
rect -31 441 -17 475
rect 17 441 31 475
rect -31 403 31 441
rect -31 369 -17 403
rect 17 369 31 403
rect -31 331 31 369
rect -31 297 -17 331
rect 17 297 31 331
rect -31 259 31 297
rect -31 225 -17 259
rect 17 225 31 259
rect -31 187 31 225
rect -31 153 -17 187
rect 17 153 31 187
rect -31 115 31 153
rect -31 81 -17 115
rect 17 81 31 115
rect -31 0 31 81
<< metal1 >>
rect -31 1492 31 1554
rect -31 0 31 62
<< end >>
