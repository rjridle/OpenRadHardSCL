* SPICE3 file created from TIEHI.ext - technology: sky130A

.subckt TIEHI Y VDD GND
X0 Y a_121_411# VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8p pd=4.58u as=1.1p ps=9.1u w=2u l=0.15u M=2
X1 a_121_411# a_121_411# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.1408p ps=8.1u w=3u l=0.15u
C0 a_121_411# Y 0.23fF
C1 a_121_411# VDD 0.39fF
C2 VDD Y 1.02fF
R0 Y.n1 Y.n0 205.342
R1 Y.n0 Y.t0 14.282
R2 Y.n0 Y.t1 14.282
R3 Y.n1 Y 0.046
R4 GND.n18 GND.n17 37.582
R5 GND.t0 GND.n15 32.601
R6 GND.n15 GND.n14 21.734
R7 GND.n24 GND.n22 20.705
R8 GND.n4 GND.n3 20.705
R9 GND.n19 GND.n18 20.705
R10 GND.n3 GND.n2 19.952
R11 GND.n17 GND.t0 15.644
R12 GND.n17 GND.n16 13.541
R13 GND.n20 GND.n11 9.154
R14 GND.n24 GND.n23 9.154
R15 GND.n6 GND.n5 9.154
R16 GND.n7 GND.n1 4.795
R17 GND.n10 GND.n9 4.65
R18 GND.n7 GND.n6 4.65
R19 GND.n25 GND.n24 4.65
R20 GND.n21 GND.n20 4.65
R21 GND.n13 GND.n12 4.504
R22 GND.n6 GND.n4 4.129
R23 GND.n20 GND.n19 3.716
R24 GND.t0 GND.n13 2.452
R25 GND.n1 GND.n0 0.474
R26 GND.n9 GND.n8 0.474
R27 GND.n10 GND 0.207
R28 GND.n25 GND.n7 0.157
R29 GND.n25 GND.n21 0.157
R30 GND.n21 GND.n10 0.145
C3 Y.t0 GND 0.15fF
C4 Y.t1 GND 0.15fF
C5 Y.n0 GND 0.61fF
C6 Y.n1 GND 0.31fF
.ends
